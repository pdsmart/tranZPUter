../../../../../cpu/zpu_uart_debug.vhd