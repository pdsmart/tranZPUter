-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"96",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"96",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"a1",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"c4",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"97",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"99",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"90",
           265 => x"0b",
           266 => x"04",
           267 => x"90",
           268 => x"0b",
           269 => x"04",
           270 => x"90",
           271 => x"0b",
           272 => x"04",
           273 => x"90",
           274 => x"0b",
           275 => x"04",
           276 => x"90",
           277 => x"0b",
           278 => x"04",
           279 => x"91",
           280 => x"0b",
           281 => x"04",
           282 => x"91",
           283 => x"0b",
           284 => x"04",
           285 => x"91",
           286 => x"0b",
           287 => x"04",
           288 => x"91",
           289 => x"0b",
           290 => x"04",
           291 => x"92",
           292 => x"0b",
           293 => x"04",
           294 => x"92",
           295 => x"0b",
           296 => x"04",
           297 => x"92",
           298 => x"0b",
           299 => x"04",
           300 => x"92",
           301 => x"0b",
           302 => x"04",
           303 => x"93",
           304 => x"0b",
           305 => x"04",
           306 => x"93",
           307 => x"0b",
           308 => x"04",
           309 => x"93",
           310 => x"0b",
           311 => x"04",
           312 => x"93",
           313 => x"0b",
           314 => x"04",
           315 => x"94",
           316 => x"0b",
           317 => x"04",
           318 => x"94",
           319 => x"0b",
           320 => x"04",
           321 => x"94",
           322 => x"0b",
           323 => x"04",
           324 => x"94",
           325 => x"0b",
           326 => x"04",
           327 => x"95",
           328 => x"0b",
           329 => x"04",
           330 => x"95",
           331 => x"0b",
           332 => x"04",
           333 => x"95",
           334 => x"0b",
           335 => x"04",
           336 => x"95",
           337 => x"0b",
           338 => x"04",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"00",
           386 => x"00",
           387 => x"00",
           388 => x"00",
           389 => x"00",
           390 => x"00",
           391 => x"00",
           392 => x"00",
           393 => x"00",
           394 => x"00",
           395 => x"00",
           396 => x"00",
           397 => x"00",
           398 => x"00",
           399 => x"00",
           400 => x"00",
           401 => x"00",
           402 => x"00",
           403 => x"00",
           404 => x"00",
           405 => x"00",
           406 => x"00",
           407 => x"00",
           408 => x"00",
           409 => x"00",
           410 => x"00",
           411 => x"00",
           412 => x"00",
           413 => x"00",
           414 => x"00",
           415 => x"00",
           416 => x"00",
           417 => x"00",
           418 => x"00",
           419 => x"00",
           420 => x"00",
           421 => x"00",
           422 => x"00",
           423 => x"00",
           424 => x"00",
           425 => x"00",
           426 => x"00",
           427 => x"00",
           428 => x"00",
           429 => x"00",
           430 => x"00",
           431 => x"00",
           432 => x"00",
           433 => x"00",
           434 => x"00",
           435 => x"00",
           436 => x"00",
           437 => x"00",
           438 => x"00",
           439 => x"00",
           440 => x"00",
           441 => x"00",
           442 => x"00",
           443 => x"00",
           444 => x"00",
           445 => x"00",
           446 => x"00",
           447 => x"00",
           448 => x"00",
           449 => x"00",
           450 => x"00",
           451 => x"00",
           452 => x"00",
           453 => x"00",
           454 => x"00",
           455 => x"00",
           456 => x"00",
           457 => x"00",
           458 => x"00",
           459 => x"00",
           460 => x"00",
           461 => x"00",
           462 => x"00",
           463 => x"00",
           464 => x"00",
           465 => x"00",
           466 => x"00",
           467 => x"00",
           468 => x"00",
           469 => x"00",
           470 => x"00",
           471 => x"00",
           472 => x"00",
           473 => x"00",
           474 => x"00",
           475 => x"00",
           476 => x"00",
           477 => x"00",
           478 => x"00",
           479 => x"00",
           480 => x"00",
           481 => x"00",
           482 => x"00",
           483 => x"00",
           484 => x"00",
           485 => x"00",
           486 => x"00",
           487 => x"00",
           488 => x"00",
           489 => x"00",
           490 => x"00",
           491 => x"00",
           492 => x"00",
           493 => x"00",
           494 => x"00",
           495 => x"00",
           496 => x"00",
           497 => x"00",
           498 => x"00",
           499 => x"00",
           500 => x"00",
           501 => x"00",
           502 => x"00",
           503 => x"00",
           504 => x"00",
           505 => x"00",
           506 => x"00",
           507 => x"00",
           508 => x"00",
           509 => x"00",
           510 => x"00",
           511 => x"00",
           512 => x"81",
           513 => x"d8",
           514 => x"2d",
           515 => x"08",
           516 => x"04",
           517 => x"0c",
           518 => x"81",
           519 => x"83",
           520 => x"81",
           521 => x"b1",
           522 => x"dc",
           523 => x"80",
           524 => x"dc",
           525 => x"80",
           526 => x"d8",
           527 => x"90",
           528 => x"d8",
           529 => x"2d",
           530 => x"08",
           531 => x"04",
           532 => x"0c",
           533 => x"81",
           534 => x"83",
           535 => x"81",
           536 => x"b2",
           537 => x"dc",
           538 => x"80",
           539 => x"dc",
           540 => x"d9",
           541 => x"d8",
           542 => x"90",
           543 => x"d8",
           544 => x"2d",
           545 => x"08",
           546 => x"04",
           547 => x"0c",
           548 => x"81",
           549 => x"83",
           550 => x"81",
           551 => x"b7",
           552 => x"dc",
           553 => x"80",
           554 => x"dc",
           555 => x"9e",
           556 => x"d8",
           557 => x"90",
           558 => x"d8",
           559 => x"2d",
           560 => x"08",
           561 => x"04",
           562 => x"0c",
           563 => x"81",
           564 => x"83",
           565 => x"81",
           566 => x"9f",
           567 => x"dc",
           568 => x"80",
           569 => x"dc",
           570 => x"df",
           571 => x"d8",
           572 => x"90",
           573 => x"d8",
           574 => x"2d",
           575 => x"08",
           576 => x"04",
           577 => x"0c",
           578 => x"2d",
           579 => x"08",
           580 => x"04",
           581 => x"0c",
           582 => x"2d",
           583 => x"08",
           584 => x"04",
           585 => x"0c",
           586 => x"2d",
           587 => x"08",
           588 => x"04",
           589 => x"0c",
           590 => x"2d",
           591 => x"08",
           592 => x"04",
           593 => x"0c",
           594 => x"2d",
           595 => x"08",
           596 => x"04",
           597 => x"0c",
           598 => x"2d",
           599 => x"08",
           600 => x"04",
           601 => x"0c",
           602 => x"2d",
           603 => x"08",
           604 => x"04",
           605 => x"0c",
           606 => x"2d",
           607 => x"08",
           608 => x"04",
           609 => x"0c",
           610 => x"2d",
           611 => x"08",
           612 => x"04",
           613 => x"0c",
           614 => x"2d",
           615 => x"08",
           616 => x"04",
           617 => x"0c",
           618 => x"2d",
           619 => x"08",
           620 => x"04",
           621 => x"0c",
           622 => x"2d",
           623 => x"08",
           624 => x"04",
           625 => x"0c",
           626 => x"2d",
           627 => x"08",
           628 => x"04",
           629 => x"0c",
           630 => x"2d",
           631 => x"08",
           632 => x"04",
           633 => x"0c",
           634 => x"2d",
           635 => x"08",
           636 => x"04",
           637 => x"0c",
           638 => x"2d",
           639 => x"08",
           640 => x"04",
           641 => x"0c",
           642 => x"2d",
           643 => x"08",
           644 => x"04",
           645 => x"0c",
           646 => x"2d",
           647 => x"08",
           648 => x"04",
           649 => x"0c",
           650 => x"2d",
           651 => x"08",
           652 => x"04",
           653 => x"0c",
           654 => x"2d",
           655 => x"08",
           656 => x"04",
           657 => x"0c",
           658 => x"2d",
           659 => x"08",
           660 => x"04",
           661 => x"0c",
           662 => x"2d",
           663 => x"08",
           664 => x"04",
           665 => x"0c",
           666 => x"2d",
           667 => x"08",
           668 => x"04",
           669 => x"0c",
           670 => x"2d",
           671 => x"08",
           672 => x"04",
           673 => x"0c",
           674 => x"2d",
           675 => x"08",
           676 => x"04",
           677 => x"0c",
           678 => x"81",
           679 => x"83",
           680 => x"81",
           681 => x"80",
           682 => x"81",
           683 => x"83",
           684 => x"81",
           685 => x"80",
           686 => x"81",
           687 => x"83",
           688 => x"81",
           689 => x"9f",
           690 => x"dc",
           691 => x"80",
           692 => x"dc",
           693 => x"b5",
           694 => x"d8",
           695 => x"90",
           696 => x"d8",
           697 => x"2d",
           698 => x"08",
           699 => x"04",
           700 => x"0c",
           701 => x"2d",
           702 => x"08",
           703 => x"04",
           704 => x"10",
           705 => x"10",
           706 => x"10",
           707 => x"10",
           708 => x"10",
           709 => x"10",
           710 => x"10",
           711 => x"10",
           712 => x"04",
           713 => x"81",
           714 => x"83",
           715 => x"05",
           716 => x"10",
           717 => x"72",
           718 => x"51",
           719 => x"72",
           720 => x"06",
           721 => x"72",
           722 => x"10",
           723 => x"10",
           724 => x"ed",
           725 => x"53",
           726 => x"dc",
           727 => x"f3",
           728 => x"38",
           729 => x"84",
           730 => x"0b",
           731 => x"dd",
           732 => x"51",
           733 => x"04",
           734 => x"d8",
           735 => x"dc",
           736 => x"3d",
           737 => x"81",
           738 => x"8c",
           739 => x"81",
           740 => x"88",
           741 => x"83",
           742 => x"dc",
           743 => x"81",
           744 => x"54",
           745 => x"81",
           746 => x"04",
           747 => x"08",
           748 => x"d8",
           749 => x"0d",
           750 => x"dc",
           751 => x"05",
           752 => x"dc",
           753 => x"05",
           754 => x"a1",
           755 => x"cc",
           756 => x"dc",
           757 => x"85",
           758 => x"dc",
           759 => x"81",
           760 => x"02",
           761 => x"0c",
           762 => x"80",
           763 => x"d8",
           764 => x"0c",
           765 => x"08",
           766 => x"80",
           767 => x"81",
           768 => x"88",
           769 => x"81",
           770 => x"88",
           771 => x"0b",
           772 => x"08",
           773 => x"81",
           774 => x"fc",
           775 => x"38",
           776 => x"dc",
           777 => x"05",
           778 => x"d8",
           779 => x"08",
           780 => x"08",
           781 => x"81",
           782 => x"8c",
           783 => x"25",
           784 => x"dc",
           785 => x"05",
           786 => x"dc",
           787 => x"05",
           788 => x"81",
           789 => x"f0",
           790 => x"dc",
           791 => x"05",
           792 => x"81",
           793 => x"d8",
           794 => x"0c",
           795 => x"08",
           796 => x"81",
           797 => x"fc",
           798 => x"53",
           799 => x"08",
           800 => x"52",
           801 => x"08",
           802 => x"51",
           803 => x"81",
           804 => x"70",
           805 => x"08",
           806 => x"54",
           807 => x"08",
           808 => x"80",
           809 => x"81",
           810 => x"f8",
           811 => x"81",
           812 => x"f8",
           813 => x"dc",
           814 => x"05",
           815 => x"dc",
           816 => x"89",
           817 => x"dc",
           818 => x"81",
           819 => x"02",
           820 => x"0c",
           821 => x"80",
           822 => x"d8",
           823 => x"0c",
           824 => x"08",
           825 => x"80",
           826 => x"81",
           827 => x"88",
           828 => x"81",
           829 => x"88",
           830 => x"0b",
           831 => x"08",
           832 => x"81",
           833 => x"8c",
           834 => x"25",
           835 => x"dc",
           836 => x"05",
           837 => x"dc",
           838 => x"05",
           839 => x"81",
           840 => x"8c",
           841 => x"81",
           842 => x"88",
           843 => x"bd",
           844 => x"cc",
           845 => x"dc",
           846 => x"05",
           847 => x"dc",
           848 => x"05",
           849 => x"90",
           850 => x"d8",
           851 => x"08",
           852 => x"d8",
           853 => x"0c",
           854 => x"08",
           855 => x"70",
           856 => x"0c",
           857 => x"0d",
           858 => x"0c",
           859 => x"d8",
           860 => x"dc",
           861 => x"3d",
           862 => x"81",
           863 => x"fc",
           864 => x"0b",
           865 => x"08",
           866 => x"81",
           867 => x"8c",
           868 => x"dc",
           869 => x"05",
           870 => x"38",
           871 => x"08",
           872 => x"80",
           873 => x"80",
           874 => x"d8",
           875 => x"08",
           876 => x"81",
           877 => x"8c",
           878 => x"81",
           879 => x"8c",
           880 => x"dc",
           881 => x"05",
           882 => x"dc",
           883 => x"05",
           884 => x"39",
           885 => x"08",
           886 => x"80",
           887 => x"38",
           888 => x"08",
           889 => x"81",
           890 => x"88",
           891 => x"ad",
           892 => x"d8",
           893 => x"08",
           894 => x"08",
           895 => x"31",
           896 => x"08",
           897 => x"81",
           898 => x"f8",
           899 => x"dc",
           900 => x"05",
           901 => x"dc",
           902 => x"05",
           903 => x"d8",
           904 => x"08",
           905 => x"dc",
           906 => x"05",
           907 => x"d8",
           908 => x"08",
           909 => x"dc",
           910 => x"05",
           911 => x"39",
           912 => x"08",
           913 => x"80",
           914 => x"81",
           915 => x"88",
           916 => x"81",
           917 => x"f4",
           918 => x"91",
           919 => x"d8",
           920 => x"08",
           921 => x"d8",
           922 => x"0c",
           923 => x"d8",
           924 => x"08",
           925 => x"0c",
           926 => x"81",
           927 => x"04",
           928 => x"76",
           929 => x"8c",
           930 => x"33",
           931 => x"55",
           932 => x"8a",
           933 => x"06",
           934 => x"2e",
           935 => x"12",
           936 => x"2e",
           937 => x"73",
           938 => x"55",
           939 => x"52",
           940 => x"09",
           941 => x"38",
           942 => x"cc",
           943 => x"0d",
           944 => x"88",
           945 => x"70",
           946 => x"07",
           947 => x"8f",
           948 => x"38",
           949 => x"84",
           950 => x"72",
           951 => x"05",
           952 => x"71",
           953 => x"53",
           954 => x"70",
           955 => x"0c",
           956 => x"71",
           957 => x"38",
           958 => x"90",
           959 => x"70",
           960 => x"0c",
           961 => x"71",
           962 => x"38",
           963 => x"8e",
           964 => x"0d",
           965 => x"72",
           966 => x"53",
           967 => x"93",
           968 => x"73",
           969 => x"54",
           970 => x"2e",
           971 => x"73",
           972 => x"71",
           973 => x"ff",
           974 => x"70",
           975 => x"38",
           976 => x"70",
           977 => x"81",
           978 => x"81",
           979 => x"71",
           980 => x"ff",
           981 => x"54",
           982 => x"38",
           983 => x"73",
           984 => x"75",
           985 => x"71",
           986 => x"dc",
           987 => x"52",
           988 => x"04",
           989 => x"f7",
           990 => x"14",
           991 => x"84",
           992 => x"06",
           993 => x"70",
           994 => x"14",
           995 => x"08",
           996 => x"71",
           997 => x"dc",
           998 => x"54",
           999 => x"39",
          1000 => x"dc",
          1001 => x"3d",
          1002 => x"3d",
          1003 => x"83",
          1004 => x"2b",
          1005 => x"3f",
          1006 => x"08",
          1007 => x"72",
          1008 => x"54",
          1009 => x"25",
          1010 => x"81",
          1011 => x"84",
          1012 => x"fb",
          1013 => x"70",
          1014 => x"53",
          1015 => x"2e",
          1016 => x"71",
          1017 => x"a0",
          1018 => x"06",
          1019 => x"12",
          1020 => x"71",
          1021 => x"81",
          1022 => x"73",
          1023 => x"ff",
          1024 => x"55",
          1025 => x"83",
          1026 => x"70",
          1027 => x"38",
          1028 => x"73",
          1029 => x"51",
          1030 => x"09",
          1031 => x"38",
          1032 => x"81",
          1033 => x"72",
          1034 => x"51",
          1035 => x"cc",
          1036 => x"0d",
          1037 => x"0d",
          1038 => x"08",
          1039 => x"38",
          1040 => x"05",
          1041 => x"9b",
          1042 => x"dc",
          1043 => x"38",
          1044 => x"39",
          1045 => x"81",
          1046 => x"86",
          1047 => x"fc",
          1048 => x"82",
          1049 => x"05",
          1050 => x"52",
          1051 => x"81",
          1052 => x"13",
          1053 => x"51",
          1054 => x"9e",
          1055 => x"38",
          1056 => x"51",
          1057 => x"97",
          1058 => x"38",
          1059 => x"51",
          1060 => x"bb",
          1061 => x"38",
          1062 => x"51",
          1063 => x"bb",
          1064 => x"38",
          1065 => x"55",
          1066 => x"87",
          1067 => x"d9",
          1068 => x"22",
          1069 => x"73",
          1070 => x"80",
          1071 => x"0b",
          1072 => x"9c",
          1073 => x"87",
          1074 => x"0c",
          1075 => x"87",
          1076 => x"0c",
          1077 => x"87",
          1078 => x"0c",
          1079 => x"87",
          1080 => x"0c",
          1081 => x"87",
          1082 => x"0c",
          1083 => x"87",
          1084 => x"0c",
          1085 => x"98",
          1086 => x"87",
          1087 => x"0c",
          1088 => x"c0",
          1089 => x"80",
          1090 => x"dc",
          1091 => x"3d",
          1092 => x"3d",
          1093 => x"87",
          1094 => x"5d",
          1095 => x"87",
          1096 => x"08",
          1097 => x"23",
          1098 => x"b8",
          1099 => x"82",
          1100 => x"c0",
          1101 => x"5a",
          1102 => x"34",
          1103 => x"b0",
          1104 => x"84",
          1105 => x"c0",
          1106 => x"5a",
          1107 => x"34",
          1108 => x"a8",
          1109 => x"86",
          1110 => x"c0",
          1111 => x"5c",
          1112 => x"23",
          1113 => x"a0",
          1114 => x"8a",
          1115 => x"7d",
          1116 => x"ff",
          1117 => x"7b",
          1118 => x"06",
          1119 => x"33",
          1120 => x"33",
          1121 => x"33",
          1122 => x"33",
          1123 => x"33",
          1124 => x"ff",
          1125 => x"81",
          1126 => x"94",
          1127 => x"3d",
          1128 => x"3d",
          1129 => x"05",
          1130 => x"70",
          1131 => x"52",
          1132 => x"0b",
          1133 => x"34",
          1134 => x"04",
          1135 => x"77",
          1136 => x"d8",
          1137 => x"81",
          1138 => x"55",
          1139 => x"94",
          1140 => x"80",
          1141 => x"87",
          1142 => x"51",
          1143 => x"96",
          1144 => x"06",
          1145 => x"70",
          1146 => x"38",
          1147 => x"70",
          1148 => x"51",
          1149 => x"72",
          1150 => x"81",
          1151 => x"70",
          1152 => x"38",
          1153 => x"70",
          1154 => x"51",
          1155 => x"38",
          1156 => x"06",
          1157 => x"94",
          1158 => x"80",
          1159 => x"87",
          1160 => x"52",
          1161 => x"75",
          1162 => x"0c",
          1163 => x"04",
          1164 => x"02",
          1165 => x"0b",
          1166 => x"f4",
          1167 => x"ff",
          1168 => x"56",
          1169 => x"84",
          1170 => x"2e",
          1171 => x"c0",
          1172 => x"70",
          1173 => x"2a",
          1174 => x"53",
          1175 => x"80",
          1176 => x"71",
          1177 => x"81",
          1178 => x"70",
          1179 => x"81",
          1180 => x"06",
          1181 => x"80",
          1182 => x"71",
          1183 => x"81",
          1184 => x"70",
          1185 => x"73",
          1186 => x"51",
          1187 => x"80",
          1188 => x"2e",
          1189 => x"c0",
          1190 => x"75",
          1191 => x"3d",
          1192 => x"3d",
          1193 => x"80",
          1194 => x"81",
          1195 => x"53",
          1196 => x"2e",
          1197 => x"71",
          1198 => x"81",
          1199 => x"81",
          1200 => x"70",
          1201 => x"59",
          1202 => x"87",
          1203 => x"51",
          1204 => x"86",
          1205 => x"94",
          1206 => x"08",
          1207 => x"70",
          1208 => x"54",
          1209 => x"2e",
          1210 => x"91",
          1211 => x"06",
          1212 => x"d7",
          1213 => x"32",
          1214 => x"51",
          1215 => x"2e",
          1216 => x"93",
          1217 => x"06",
          1218 => x"ff",
          1219 => x"81",
          1220 => x"87",
          1221 => x"52",
          1222 => x"86",
          1223 => x"94",
          1224 => x"72",
          1225 => x"74",
          1226 => x"ff",
          1227 => x"57",
          1228 => x"38",
          1229 => x"cc",
          1230 => x"0d",
          1231 => x"0d",
          1232 => x"d8",
          1233 => x"81",
          1234 => x"52",
          1235 => x"84",
          1236 => x"2e",
          1237 => x"c0",
          1238 => x"70",
          1239 => x"2a",
          1240 => x"51",
          1241 => x"80",
          1242 => x"71",
          1243 => x"51",
          1244 => x"80",
          1245 => x"2e",
          1246 => x"c0",
          1247 => x"71",
          1248 => x"ff",
          1249 => x"cc",
          1250 => x"3d",
          1251 => x"3d",
          1252 => x"81",
          1253 => x"70",
          1254 => x"52",
          1255 => x"94",
          1256 => x"80",
          1257 => x"87",
          1258 => x"52",
          1259 => x"82",
          1260 => x"06",
          1261 => x"ff",
          1262 => x"2e",
          1263 => x"81",
          1264 => x"87",
          1265 => x"52",
          1266 => x"86",
          1267 => x"94",
          1268 => x"08",
          1269 => x"70",
          1270 => x"53",
          1271 => x"dc",
          1272 => x"3d",
          1273 => x"3d",
          1274 => x"9e",
          1275 => x"9c",
          1276 => x"51",
          1277 => x"2e",
          1278 => x"87",
          1279 => x"08",
          1280 => x"0c",
          1281 => x"a8",
          1282 => x"fc",
          1283 => x"9e",
          1284 => x"d9",
          1285 => x"c0",
          1286 => x"81",
          1287 => x"87",
          1288 => x"08",
          1289 => x"0c",
          1290 => x"a0",
          1291 => x"8c",
          1292 => x"9e",
          1293 => x"d9",
          1294 => x"c0",
          1295 => x"81",
          1296 => x"87",
          1297 => x"08",
          1298 => x"0c",
          1299 => x"b8",
          1300 => x"9c",
          1301 => x"9e",
          1302 => x"d9",
          1303 => x"c0",
          1304 => x"81",
          1305 => x"87",
          1306 => x"08",
          1307 => x"0c",
          1308 => x"80",
          1309 => x"81",
          1310 => x"87",
          1311 => x"08",
          1312 => x"0c",
          1313 => x"88",
          1314 => x"b4",
          1315 => x"9e",
          1316 => x"d9",
          1317 => x"0b",
          1318 => x"34",
          1319 => x"c0",
          1320 => x"70",
          1321 => x"06",
          1322 => x"70",
          1323 => x"38",
          1324 => x"81",
          1325 => x"80",
          1326 => x"9e",
          1327 => x"88",
          1328 => x"51",
          1329 => x"80",
          1330 => x"81",
          1331 => x"d9",
          1332 => x"0b",
          1333 => x"90",
          1334 => x"80",
          1335 => x"52",
          1336 => x"2e",
          1337 => x"52",
          1338 => x"bf",
          1339 => x"87",
          1340 => x"08",
          1341 => x"80",
          1342 => x"52",
          1343 => x"83",
          1344 => x"71",
          1345 => x"34",
          1346 => x"c0",
          1347 => x"70",
          1348 => x"06",
          1349 => x"70",
          1350 => x"38",
          1351 => x"81",
          1352 => x"80",
          1353 => x"9e",
          1354 => x"90",
          1355 => x"51",
          1356 => x"80",
          1357 => x"81",
          1358 => x"d9",
          1359 => x"0b",
          1360 => x"90",
          1361 => x"80",
          1362 => x"52",
          1363 => x"2e",
          1364 => x"52",
          1365 => x"c3",
          1366 => x"87",
          1367 => x"08",
          1368 => x"80",
          1369 => x"52",
          1370 => x"83",
          1371 => x"71",
          1372 => x"34",
          1373 => x"c0",
          1374 => x"70",
          1375 => x"06",
          1376 => x"70",
          1377 => x"38",
          1378 => x"81",
          1379 => x"80",
          1380 => x"9e",
          1381 => x"80",
          1382 => x"51",
          1383 => x"80",
          1384 => x"81",
          1385 => x"d9",
          1386 => x"0b",
          1387 => x"90",
          1388 => x"80",
          1389 => x"52",
          1390 => x"83",
          1391 => x"71",
          1392 => x"34",
          1393 => x"90",
          1394 => x"80",
          1395 => x"2a",
          1396 => x"70",
          1397 => x"34",
          1398 => x"c0",
          1399 => x"70",
          1400 => x"51",
          1401 => x"80",
          1402 => x"81",
          1403 => x"d9",
          1404 => x"c0",
          1405 => x"70",
          1406 => x"70",
          1407 => x"51",
          1408 => x"d9",
          1409 => x"0b",
          1410 => x"90",
          1411 => x"06",
          1412 => x"70",
          1413 => x"38",
          1414 => x"81",
          1415 => x"87",
          1416 => x"08",
          1417 => x"51",
          1418 => x"d9",
          1419 => x"3d",
          1420 => x"3d",
          1421 => x"e4",
          1422 => x"3f",
          1423 => x"33",
          1424 => x"2e",
          1425 => x"c5",
          1426 => x"b4",
          1427 => x"8c",
          1428 => x"3f",
          1429 => x"33",
          1430 => x"2e",
          1431 => x"d9",
          1432 => x"d9",
          1433 => x"54",
          1434 => x"a4",
          1435 => x"3f",
          1436 => x"33",
          1437 => x"2e",
          1438 => x"d9",
          1439 => x"d9",
          1440 => x"54",
          1441 => x"c0",
          1442 => x"3f",
          1443 => x"33",
          1444 => x"2e",
          1445 => x"d8",
          1446 => x"d8",
          1447 => x"54",
          1448 => x"dc",
          1449 => x"3f",
          1450 => x"33",
          1451 => x"2e",
          1452 => x"d9",
          1453 => x"d9",
          1454 => x"54",
          1455 => x"f8",
          1456 => x"3f",
          1457 => x"33",
          1458 => x"2e",
          1459 => x"d9",
          1460 => x"d9",
          1461 => x"54",
          1462 => x"94",
          1463 => x"3f",
          1464 => x"33",
          1465 => x"2e",
          1466 => x"d9",
          1467 => x"81",
          1468 => x"89",
          1469 => x"d9",
          1470 => x"73",
          1471 => x"38",
          1472 => x"33",
          1473 => x"d0",
          1474 => x"3f",
          1475 => x"33",
          1476 => x"2e",
          1477 => x"d9",
          1478 => x"81",
          1479 => x"89",
          1480 => x"d9",
          1481 => x"73",
          1482 => x"38",
          1483 => x"51",
          1484 => x"81",
          1485 => x"54",
          1486 => x"88",
          1487 => x"a4",
          1488 => x"3f",
          1489 => x"33",
          1490 => x"2e",
          1491 => x"c8",
          1492 => x"ac",
          1493 => x"c5",
          1494 => x"80",
          1495 => x"81",
          1496 => x"83",
          1497 => x"d9",
          1498 => x"73",
          1499 => x"38",
          1500 => x"51",
          1501 => x"81",
          1502 => x"83",
          1503 => x"d9",
          1504 => x"81",
          1505 => x"88",
          1506 => x"d9",
          1507 => x"81",
          1508 => x"88",
          1509 => x"d9",
          1510 => x"81",
          1511 => x"88",
          1512 => x"c9",
          1513 => x"d8",
          1514 => x"ac",
          1515 => x"c9",
          1516 => x"b0",
          1517 => x"b0",
          1518 => x"84",
          1519 => x"51",
          1520 => x"81",
          1521 => x"bd",
          1522 => x"76",
          1523 => x"54",
          1524 => x"08",
          1525 => x"88",
          1526 => x"3f",
          1527 => x"33",
          1528 => x"2e",
          1529 => x"d9",
          1530 => x"bd",
          1531 => x"75",
          1532 => x"3f",
          1533 => x"08",
          1534 => x"29",
          1535 => x"54",
          1536 => x"cc",
          1537 => x"ca",
          1538 => x"d8",
          1539 => x"be",
          1540 => x"80",
          1541 => x"81",
          1542 => x"56",
          1543 => x"52",
          1544 => x"d5",
          1545 => x"cc",
          1546 => x"c0",
          1547 => x"31",
          1548 => x"dc",
          1549 => x"81",
          1550 => x"87",
          1551 => x"d6",
          1552 => x"bc",
          1553 => x"0d",
          1554 => x"0d",
          1555 => x"33",
          1556 => x"71",
          1557 => x"38",
          1558 => x"81",
          1559 => x"52",
          1560 => x"81",
          1561 => x"9d",
          1562 => x"94",
          1563 => x"81",
          1564 => x"91",
          1565 => x"a4",
          1566 => x"81",
          1567 => x"85",
          1568 => x"b0",
          1569 => x"3f",
          1570 => x"04",
          1571 => x"0c",
          1572 => x"87",
          1573 => x"0c",
          1574 => x"d0",
          1575 => x"96",
          1576 => x"fe",
          1577 => x"93",
          1578 => x"72",
          1579 => x"81",
          1580 => x"8d",
          1581 => x"81",
          1582 => x"52",
          1583 => x"90",
          1584 => x"34",
          1585 => x"08",
          1586 => x"dc",
          1587 => x"39",
          1588 => x"08",
          1589 => x"2e",
          1590 => x"51",
          1591 => x"3d",
          1592 => x"3d",
          1593 => x"05",
          1594 => x"dc",
          1595 => x"dc",
          1596 => x"51",
          1597 => x"72",
          1598 => x"0c",
          1599 => x"04",
          1600 => x"75",
          1601 => x"70",
          1602 => x"53",
          1603 => x"2e",
          1604 => x"81",
          1605 => x"81",
          1606 => x"87",
          1607 => x"85",
          1608 => x"fc",
          1609 => x"81",
          1610 => x"78",
          1611 => x"0c",
          1612 => x"33",
          1613 => x"06",
          1614 => x"80",
          1615 => x"72",
          1616 => x"51",
          1617 => x"fe",
          1618 => x"39",
          1619 => x"dc",
          1620 => x"0d",
          1621 => x"0d",
          1622 => x"59",
          1623 => x"05",
          1624 => x"75",
          1625 => x"f8",
          1626 => x"2e",
          1627 => x"82",
          1628 => x"70",
          1629 => x"05",
          1630 => x"5b",
          1631 => x"2e",
          1632 => x"85",
          1633 => x"8b",
          1634 => x"2e",
          1635 => x"8a",
          1636 => x"78",
          1637 => x"5a",
          1638 => x"aa",
          1639 => x"06",
          1640 => x"84",
          1641 => x"7b",
          1642 => x"5d",
          1643 => x"59",
          1644 => x"d0",
          1645 => x"89",
          1646 => x"7a",
          1647 => x"10",
          1648 => x"d0",
          1649 => x"81",
          1650 => x"57",
          1651 => x"75",
          1652 => x"70",
          1653 => x"07",
          1654 => x"80",
          1655 => x"30",
          1656 => x"80",
          1657 => x"53",
          1658 => x"55",
          1659 => x"2e",
          1660 => x"84",
          1661 => x"81",
          1662 => x"57",
          1663 => x"2e",
          1664 => x"75",
          1665 => x"76",
          1666 => x"e0",
          1667 => x"ff",
          1668 => x"73",
          1669 => x"81",
          1670 => x"80",
          1671 => x"38",
          1672 => x"2e",
          1673 => x"73",
          1674 => x"8b",
          1675 => x"c2",
          1676 => x"38",
          1677 => x"73",
          1678 => x"81",
          1679 => x"8f",
          1680 => x"d5",
          1681 => x"38",
          1682 => x"24",
          1683 => x"80",
          1684 => x"38",
          1685 => x"73",
          1686 => x"80",
          1687 => x"ef",
          1688 => x"19",
          1689 => x"59",
          1690 => x"33",
          1691 => x"75",
          1692 => x"81",
          1693 => x"70",
          1694 => x"55",
          1695 => x"79",
          1696 => x"90",
          1697 => x"16",
          1698 => x"7b",
          1699 => x"a0",
          1700 => x"3f",
          1701 => x"53",
          1702 => x"e9",
          1703 => x"fc",
          1704 => x"81",
          1705 => x"72",
          1706 => x"b0",
          1707 => x"fb",
          1708 => x"39",
          1709 => x"83",
          1710 => x"59",
          1711 => x"82",
          1712 => x"88",
          1713 => x"8a",
          1714 => x"90",
          1715 => x"75",
          1716 => x"3f",
          1717 => x"79",
          1718 => x"81",
          1719 => x"72",
          1720 => x"38",
          1721 => x"59",
          1722 => x"84",
          1723 => x"58",
          1724 => x"80",
          1725 => x"30",
          1726 => x"80",
          1727 => x"55",
          1728 => x"25",
          1729 => x"80",
          1730 => x"74",
          1731 => x"07",
          1732 => x"0b",
          1733 => x"57",
          1734 => x"51",
          1735 => x"81",
          1736 => x"81",
          1737 => x"53",
          1738 => x"e0",
          1739 => x"dc",
          1740 => x"89",
          1741 => x"38",
          1742 => x"75",
          1743 => x"84",
          1744 => x"53",
          1745 => x"06",
          1746 => x"53",
          1747 => x"81",
          1748 => x"81",
          1749 => x"70",
          1750 => x"2a",
          1751 => x"76",
          1752 => x"38",
          1753 => x"38",
          1754 => x"70",
          1755 => x"53",
          1756 => x"8e",
          1757 => x"77",
          1758 => x"53",
          1759 => x"81",
          1760 => x"7a",
          1761 => x"55",
          1762 => x"83",
          1763 => x"79",
          1764 => x"81",
          1765 => x"72",
          1766 => x"17",
          1767 => x"27",
          1768 => x"51",
          1769 => x"75",
          1770 => x"72",
          1771 => x"81",
          1772 => x"7a",
          1773 => x"38",
          1774 => x"05",
          1775 => x"ff",
          1776 => x"70",
          1777 => x"57",
          1778 => x"76",
          1779 => x"81",
          1780 => x"72",
          1781 => x"84",
          1782 => x"f9",
          1783 => x"39",
          1784 => x"04",
          1785 => x"86",
          1786 => x"84",
          1787 => x"55",
          1788 => x"fa",
          1789 => x"3d",
          1790 => x"3d",
          1791 => x"dc",
          1792 => x"3d",
          1793 => x"75",
          1794 => x"3f",
          1795 => x"08",
          1796 => x"34",
          1797 => x"dc",
          1798 => x"3d",
          1799 => x"3d",
          1800 => x"dc",
          1801 => x"dc",
          1802 => x"3d",
          1803 => x"77",
          1804 => x"a1",
          1805 => x"dc",
          1806 => x"3d",
          1807 => x"3d",
          1808 => x"81",
          1809 => x"70",
          1810 => x"55",
          1811 => x"80",
          1812 => x"38",
          1813 => x"08",
          1814 => x"81",
          1815 => x"81",
          1816 => x"72",
          1817 => x"cb",
          1818 => x"2e",
          1819 => x"88",
          1820 => x"70",
          1821 => x"51",
          1822 => x"2e",
          1823 => x"80",
          1824 => x"ff",
          1825 => x"39",
          1826 => x"c8",
          1827 => x"52",
          1828 => x"c0",
          1829 => x"52",
          1830 => x"81",
          1831 => x"51",
          1832 => x"ff",
          1833 => x"15",
          1834 => x"34",
          1835 => x"f3",
          1836 => x"72",
          1837 => x"0c",
          1838 => x"04",
          1839 => x"81",
          1840 => x"75",
          1841 => x"0c",
          1842 => x"52",
          1843 => x"3f",
          1844 => x"e0",
          1845 => x"0d",
          1846 => x"0d",
          1847 => x"56",
          1848 => x"0c",
          1849 => x"70",
          1850 => x"73",
          1851 => x"81",
          1852 => x"81",
          1853 => x"ed",
          1854 => x"2e",
          1855 => x"8e",
          1856 => x"08",
          1857 => x"76",
          1858 => x"56",
          1859 => x"b0",
          1860 => x"06",
          1861 => x"75",
          1862 => x"76",
          1863 => x"70",
          1864 => x"73",
          1865 => x"8b",
          1866 => x"73",
          1867 => x"85",
          1868 => x"82",
          1869 => x"76",
          1870 => x"70",
          1871 => x"ac",
          1872 => x"a0",
          1873 => x"fa",
          1874 => x"53",
          1875 => x"57",
          1876 => x"98",
          1877 => x"39",
          1878 => x"80",
          1879 => x"26",
          1880 => x"86",
          1881 => x"80",
          1882 => x"57",
          1883 => x"74",
          1884 => x"38",
          1885 => x"27",
          1886 => x"14",
          1887 => x"06",
          1888 => x"14",
          1889 => x"06",
          1890 => x"74",
          1891 => x"f9",
          1892 => x"ff",
          1893 => x"89",
          1894 => x"38",
          1895 => x"c5",
          1896 => x"29",
          1897 => x"81",
          1898 => x"76",
          1899 => x"56",
          1900 => x"ba",
          1901 => x"2e",
          1902 => x"30",
          1903 => x"0c",
          1904 => x"81",
          1905 => x"8a",
          1906 => x"f8",
          1907 => x"7c",
          1908 => x"70",
          1909 => x"75",
          1910 => x"55",
          1911 => x"2e",
          1912 => x"87",
          1913 => x"76",
          1914 => x"73",
          1915 => x"81",
          1916 => x"81",
          1917 => x"77",
          1918 => x"70",
          1919 => x"58",
          1920 => x"09",
          1921 => x"c2",
          1922 => x"81",
          1923 => x"75",
          1924 => x"55",
          1925 => x"e2",
          1926 => x"90",
          1927 => x"f8",
          1928 => x"8f",
          1929 => x"81",
          1930 => x"75",
          1931 => x"55",
          1932 => x"81",
          1933 => x"27",
          1934 => x"d0",
          1935 => x"55",
          1936 => x"73",
          1937 => x"80",
          1938 => x"14",
          1939 => x"72",
          1940 => x"e0",
          1941 => x"80",
          1942 => x"39",
          1943 => x"55",
          1944 => x"80",
          1945 => x"e0",
          1946 => x"38",
          1947 => x"81",
          1948 => x"53",
          1949 => x"81",
          1950 => x"53",
          1951 => x"8e",
          1952 => x"70",
          1953 => x"55",
          1954 => x"27",
          1955 => x"77",
          1956 => x"74",
          1957 => x"76",
          1958 => x"77",
          1959 => x"70",
          1960 => x"55",
          1961 => x"77",
          1962 => x"38",
          1963 => x"74",
          1964 => x"55",
          1965 => x"cc",
          1966 => x"0d",
          1967 => x"0d",
          1968 => x"33",
          1969 => x"70",
          1970 => x"38",
          1971 => x"11",
          1972 => x"81",
          1973 => x"83",
          1974 => x"fc",
          1975 => x"9b",
          1976 => x"84",
          1977 => x"33",
          1978 => x"51",
          1979 => x"80",
          1980 => x"84",
          1981 => x"92",
          1982 => x"51",
          1983 => x"80",
          1984 => x"81",
          1985 => x"72",
          1986 => x"92",
          1987 => x"81",
          1988 => x"0b",
          1989 => x"8c",
          1990 => x"71",
          1991 => x"06",
          1992 => x"80",
          1993 => x"87",
          1994 => x"08",
          1995 => x"38",
          1996 => x"80",
          1997 => x"71",
          1998 => x"c0",
          1999 => x"51",
          2000 => x"87",
          2001 => x"d9",
          2002 => x"81",
          2003 => x"33",
          2004 => x"dc",
          2005 => x"3d",
          2006 => x"3d",
          2007 => x"64",
          2008 => x"bf",
          2009 => x"40",
          2010 => x"74",
          2011 => x"cd",
          2012 => x"cc",
          2013 => x"7a",
          2014 => x"81",
          2015 => x"72",
          2016 => x"87",
          2017 => x"11",
          2018 => x"8c",
          2019 => x"92",
          2020 => x"5a",
          2021 => x"58",
          2022 => x"c0",
          2023 => x"76",
          2024 => x"76",
          2025 => x"70",
          2026 => x"81",
          2027 => x"54",
          2028 => x"8e",
          2029 => x"52",
          2030 => x"81",
          2031 => x"81",
          2032 => x"74",
          2033 => x"53",
          2034 => x"83",
          2035 => x"78",
          2036 => x"8f",
          2037 => x"2e",
          2038 => x"c0",
          2039 => x"52",
          2040 => x"87",
          2041 => x"08",
          2042 => x"2e",
          2043 => x"84",
          2044 => x"38",
          2045 => x"87",
          2046 => x"15",
          2047 => x"70",
          2048 => x"52",
          2049 => x"ff",
          2050 => x"39",
          2051 => x"81",
          2052 => x"ff",
          2053 => x"57",
          2054 => x"90",
          2055 => x"80",
          2056 => x"71",
          2057 => x"78",
          2058 => x"38",
          2059 => x"80",
          2060 => x"80",
          2061 => x"81",
          2062 => x"72",
          2063 => x"0c",
          2064 => x"04",
          2065 => x"60",
          2066 => x"8c",
          2067 => x"33",
          2068 => x"5b",
          2069 => x"74",
          2070 => x"e1",
          2071 => x"cc",
          2072 => x"79",
          2073 => x"78",
          2074 => x"06",
          2075 => x"77",
          2076 => x"87",
          2077 => x"11",
          2078 => x"8c",
          2079 => x"92",
          2080 => x"59",
          2081 => x"85",
          2082 => x"98",
          2083 => x"7d",
          2084 => x"0c",
          2085 => x"08",
          2086 => x"70",
          2087 => x"53",
          2088 => x"2e",
          2089 => x"70",
          2090 => x"33",
          2091 => x"18",
          2092 => x"2a",
          2093 => x"51",
          2094 => x"2e",
          2095 => x"c0",
          2096 => x"52",
          2097 => x"87",
          2098 => x"08",
          2099 => x"2e",
          2100 => x"84",
          2101 => x"38",
          2102 => x"87",
          2103 => x"15",
          2104 => x"70",
          2105 => x"52",
          2106 => x"ff",
          2107 => x"39",
          2108 => x"81",
          2109 => x"80",
          2110 => x"52",
          2111 => x"90",
          2112 => x"80",
          2113 => x"71",
          2114 => x"7a",
          2115 => x"38",
          2116 => x"80",
          2117 => x"80",
          2118 => x"81",
          2119 => x"72",
          2120 => x"0c",
          2121 => x"04",
          2122 => x"7a",
          2123 => x"a3",
          2124 => x"88",
          2125 => x"33",
          2126 => x"56",
          2127 => x"3f",
          2128 => x"08",
          2129 => x"83",
          2130 => x"fe",
          2131 => x"87",
          2132 => x"0c",
          2133 => x"76",
          2134 => x"38",
          2135 => x"93",
          2136 => x"2b",
          2137 => x"8c",
          2138 => x"71",
          2139 => x"38",
          2140 => x"71",
          2141 => x"c6",
          2142 => x"39",
          2143 => x"81",
          2144 => x"06",
          2145 => x"71",
          2146 => x"38",
          2147 => x"8c",
          2148 => x"e8",
          2149 => x"98",
          2150 => x"71",
          2151 => x"73",
          2152 => x"92",
          2153 => x"72",
          2154 => x"06",
          2155 => x"f7",
          2156 => x"80",
          2157 => x"88",
          2158 => x"0c",
          2159 => x"80",
          2160 => x"56",
          2161 => x"56",
          2162 => x"81",
          2163 => x"88",
          2164 => x"fe",
          2165 => x"81",
          2166 => x"33",
          2167 => x"07",
          2168 => x"0c",
          2169 => x"3d",
          2170 => x"3d",
          2171 => x"11",
          2172 => x"33",
          2173 => x"71",
          2174 => x"81",
          2175 => x"72",
          2176 => x"75",
          2177 => x"81",
          2178 => x"52",
          2179 => x"54",
          2180 => x"0d",
          2181 => x"0d",
          2182 => x"05",
          2183 => x"52",
          2184 => x"70",
          2185 => x"34",
          2186 => x"51",
          2187 => x"83",
          2188 => x"ff",
          2189 => x"75",
          2190 => x"72",
          2191 => x"54",
          2192 => x"2a",
          2193 => x"70",
          2194 => x"34",
          2195 => x"51",
          2196 => x"81",
          2197 => x"70",
          2198 => x"70",
          2199 => x"3d",
          2200 => x"3d",
          2201 => x"77",
          2202 => x"70",
          2203 => x"38",
          2204 => x"05",
          2205 => x"70",
          2206 => x"34",
          2207 => x"eb",
          2208 => x"0d",
          2209 => x"0d",
          2210 => x"54",
          2211 => x"72",
          2212 => x"54",
          2213 => x"51",
          2214 => x"84",
          2215 => x"fc",
          2216 => x"77",
          2217 => x"53",
          2218 => x"05",
          2219 => x"70",
          2220 => x"33",
          2221 => x"ff",
          2222 => x"52",
          2223 => x"2e",
          2224 => x"80",
          2225 => x"71",
          2226 => x"0c",
          2227 => x"04",
          2228 => x"74",
          2229 => x"89",
          2230 => x"2e",
          2231 => x"11",
          2232 => x"52",
          2233 => x"70",
          2234 => x"cc",
          2235 => x"0d",
          2236 => x"81",
          2237 => x"04",
          2238 => x"dc",
          2239 => x"f7",
          2240 => x"56",
          2241 => x"17",
          2242 => x"74",
          2243 => x"d6",
          2244 => x"b0",
          2245 => x"b4",
          2246 => x"81",
          2247 => x"59",
          2248 => x"81",
          2249 => x"7a",
          2250 => x"06",
          2251 => x"dc",
          2252 => x"17",
          2253 => x"08",
          2254 => x"08",
          2255 => x"08",
          2256 => x"74",
          2257 => x"38",
          2258 => x"55",
          2259 => x"09",
          2260 => x"38",
          2261 => x"18",
          2262 => x"81",
          2263 => x"f9",
          2264 => x"39",
          2265 => x"81",
          2266 => x"8b",
          2267 => x"fa",
          2268 => x"7a",
          2269 => x"57",
          2270 => x"08",
          2271 => x"75",
          2272 => x"3f",
          2273 => x"08",
          2274 => x"cc",
          2275 => x"81",
          2276 => x"b4",
          2277 => x"16",
          2278 => x"be",
          2279 => x"cc",
          2280 => x"85",
          2281 => x"81",
          2282 => x"17",
          2283 => x"dc",
          2284 => x"3d",
          2285 => x"3d",
          2286 => x"52",
          2287 => x"3f",
          2288 => x"08",
          2289 => x"cc",
          2290 => x"38",
          2291 => x"74",
          2292 => x"81",
          2293 => x"38",
          2294 => x"59",
          2295 => x"09",
          2296 => x"e3",
          2297 => x"53",
          2298 => x"08",
          2299 => x"70",
          2300 => x"91",
          2301 => x"d5",
          2302 => x"17",
          2303 => x"3f",
          2304 => x"a4",
          2305 => x"51",
          2306 => x"86",
          2307 => x"f2",
          2308 => x"17",
          2309 => x"3f",
          2310 => x"52",
          2311 => x"51",
          2312 => x"8c",
          2313 => x"84",
          2314 => x"fc",
          2315 => x"17",
          2316 => x"70",
          2317 => x"79",
          2318 => x"52",
          2319 => x"51",
          2320 => x"77",
          2321 => x"80",
          2322 => x"81",
          2323 => x"f9",
          2324 => x"dc",
          2325 => x"2e",
          2326 => x"58",
          2327 => x"cc",
          2328 => x"0d",
          2329 => x"0d",
          2330 => x"98",
          2331 => x"05",
          2332 => x"80",
          2333 => x"27",
          2334 => x"14",
          2335 => x"29",
          2336 => x"05",
          2337 => x"81",
          2338 => x"87",
          2339 => x"f9",
          2340 => x"7a",
          2341 => x"54",
          2342 => x"27",
          2343 => x"76",
          2344 => x"27",
          2345 => x"ff",
          2346 => x"58",
          2347 => x"80",
          2348 => x"82",
          2349 => x"72",
          2350 => x"38",
          2351 => x"72",
          2352 => x"8e",
          2353 => x"39",
          2354 => x"17",
          2355 => x"a4",
          2356 => x"53",
          2357 => x"fd",
          2358 => x"dc",
          2359 => x"9f",
          2360 => x"ff",
          2361 => x"11",
          2362 => x"70",
          2363 => x"18",
          2364 => x"76",
          2365 => x"53",
          2366 => x"81",
          2367 => x"80",
          2368 => x"83",
          2369 => x"b4",
          2370 => x"88",
          2371 => x"79",
          2372 => x"84",
          2373 => x"58",
          2374 => x"80",
          2375 => x"9f",
          2376 => x"80",
          2377 => x"88",
          2378 => x"08",
          2379 => x"51",
          2380 => x"81",
          2381 => x"80",
          2382 => x"10",
          2383 => x"74",
          2384 => x"51",
          2385 => x"81",
          2386 => x"83",
          2387 => x"58",
          2388 => x"87",
          2389 => x"08",
          2390 => x"51",
          2391 => x"81",
          2392 => x"9b",
          2393 => x"2b",
          2394 => x"74",
          2395 => x"51",
          2396 => x"81",
          2397 => x"f0",
          2398 => x"83",
          2399 => x"77",
          2400 => x"0c",
          2401 => x"04",
          2402 => x"7a",
          2403 => x"58",
          2404 => x"81",
          2405 => x"9e",
          2406 => x"17",
          2407 => x"96",
          2408 => x"53",
          2409 => x"81",
          2410 => x"79",
          2411 => x"72",
          2412 => x"38",
          2413 => x"72",
          2414 => x"b8",
          2415 => x"39",
          2416 => x"17",
          2417 => x"a4",
          2418 => x"53",
          2419 => x"fb",
          2420 => x"dc",
          2421 => x"81",
          2422 => x"81",
          2423 => x"83",
          2424 => x"b4",
          2425 => x"78",
          2426 => x"56",
          2427 => x"76",
          2428 => x"38",
          2429 => x"9f",
          2430 => x"33",
          2431 => x"07",
          2432 => x"74",
          2433 => x"83",
          2434 => x"89",
          2435 => x"08",
          2436 => x"51",
          2437 => x"81",
          2438 => x"59",
          2439 => x"08",
          2440 => x"74",
          2441 => x"16",
          2442 => x"84",
          2443 => x"76",
          2444 => x"88",
          2445 => x"81",
          2446 => x"8f",
          2447 => x"53",
          2448 => x"80",
          2449 => x"88",
          2450 => x"08",
          2451 => x"51",
          2452 => x"81",
          2453 => x"59",
          2454 => x"08",
          2455 => x"77",
          2456 => x"06",
          2457 => x"83",
          2458 => x"05",
          2459 => x"f7",
          2460 => x"39",
          2461 => x"a4",
          2462 => x"52",
          2463 => x"ef",
          2464 => x"cc",
          2465 => x"dc",
          2466 => x"38",
          2467 => x"06",
          2468 => x"83",
          2469 => x"18",
          2470 => x"54",
          2471 => x"f6",
          2472 => x"dc",
          2473 => x"0a",
          2474 => x"52",
          2475 => x"83",
          2476 => x"83",
          2477 => x"81",
          2478 => x"8a",
          2479 => x"f8",
          2480 => x"7c",
          2481 => x"59",
          2482 => x"81",
          2483 => x"38",
          2484 => x"08",
          2485 => x"73",
          2486 => x"38",
          2487 => x"52",
          2488 => x"a4",
          2489 => x"cc",
          2490 => x"dc",
          2491 => x"f2",
          2492 => x"82",
          2493 => x"39",
          2494 => x"e6",
          2495 => x"cc",
          2496 => x"de",
          2497 => x"78",
          2498 => x"3f",
          2499 => x"08",
          2500 => x"cc",
          2501 => x"80",
          2502 => x"dc",
          2503 => x"2e",
          2504 => x"dc",
          2505 => x"2e",
          2506 => x"53",
          2507 => x"51",
          2508 => x"81",
          2509 => x"c5",
          2510 => x"08",
          2511 => x"18",
          2512 => x"57",
          2513 => x"90",
          2514 => x"90",
          2515 => x"16",
          2516 => x"54",
          2517 => x"34",
          2518 => x"78",
          2519 => x"38",
          2520 => x"81",
          2521 => x"8a",
          2522 => x"f6",
          2523 => x"7e",
          2524 => x"5b",
          2525 => x"38",
          2526 => x"58",
          2527 => x"88",
          2528 => x"08",
          2529 => x"38",
          2530 => x"39",
          2531 => x"51",
          2532 => x"81",
          2533 => x"dc",
          2534 => x"82",
          2535 => x"dc",
          2536 => x"81",
          2537 => x"ff",
          2538 => x"38",
          2539 => x"81",
          2540 => x"26",
          2541 => x"79",
          2542 => x"08",
          2543 => x"73",
          2544 => x"b9",
          2545 => x"2e",
          2546 => x"80",
          2547 => x"1a",
          2548 => x"08",
          2549 => x"38",
          2550 => x"52",
          2551 => x"af",
          2552 => x"81",
          2553 => x"81",
          2554 => x"06",
          2555 => x"dc",
          2556 => x"81",
          2557 => x"09",
          2558 => x"72",
          2559 => x"70",
          2560 => x"dc",
          2561 => x"51",
          2562 => x"73",
          2563 => x"81",
          2564 => x"80",
          2565 => x"8c",
          2566 => x"81",
          2567 => x"38",
          2568 => x"08",
          2569 => x"73",
          2570 => x"75",
          2571 => x"77",
          2572 => x"56",
          2573 => x"76",
          2574 => x"82",
          2575 => x"26",
          2576 => x"75",
          2577 => x"f8",
          2578 => x"dc",
          2579 => x"2e",
          2580 => x"59",
          2581 => x"08",
          2582 => x"81",
          2583 => x"81",
          2584 => x"59",
          2585 => x"08",
          2586 => x"70",
          2587 => x"25",
          2588 => x"51",
          2589 => x"73",
          2590 => x"75",
          2591 => x"81",
          2592 => x"38",
          2593 => x"f5",
          2594 => x"75",
          2595 => x"f9",
          2596 => x"dc",
          2597 => x"dc",
          2598 => x"70",
          2599 => x"08",
          2600 => x"51",
          2601 => x"80",
          2602 => x"73",
          2603 => x"38",
          2604 => x"52",
          2605 => x"d0",
          2606 => x"cc",
          2607 => x"a5",
          2608 => x"18",
          2609 => x"08",
          2610 => x"18",
          2611 => x"74",
          2612 => x"38",
          2613 => x"18",
          2614 => x"33",
          2615 => x"73",
          2616 => x"97",
          2617 => x"74",
          2618 => x"38",
          2619 => x"55",
          2620 => x"dc",
          2621 => x"85",
          2622 => x"75",
          2623 => x"dc",
          2624 => x"3d",
          2625 => x"3d",
          2626 => x"52",
          2627 => x"3f",
          2628 => x"08",
          2629 => x"81",
          2630 => x"80",
          2631 => x"52",
          2632 => x"c1",
          2633 => x"cc",
          2634 => x"cc",
          2635 => x"0c",
          2636 => x"53",
          2637 => x"15",
          2638 => x"f2",
          2639 => x"56",
          2640 => x"16",
          2641 => x"22",
          2642 => x"27",
          2643 => x"54",
          2644 => x"76",
          2645 => x"33",
          2646 => x"3f",
          2647 => x"08",
          2648 => x"38",
          2649 => x"76",
          2650 => x"70",
          2651 => x"9f",
          2652 => x"56",
          2653 => x"dc",
          2654 => x"3d",
          2655 => x"3d",
          2656 => x"71",
          2657 => x"57",
          2658 => x"0a",
          2659 => x"38",
          2660 => x"53",
          2661 => x"38",
          2662 => x"0c",
          2663 => x"54",
          2664 => x"75",
          2665 => x"73",
          2666 => x"a8",
          2667 => x"73",
          2668 => x"85",
          2669 => x"0b",
          2670 => x"5a",
          2671 => x"27",
          2672 => x"a8",
          2673 => x"18",
          2674 => x"39",
          2675 => x"70",
          2676 => x"58",
          2677 => x"b2",
          2678 => x"76",
          2679 => x"3f",
          2680 => x"08",
          2681 => x"cc",
          2682 => x"bd",
          2683 => x"81",
          2684 => x"27",
          2685 => x"16",
          2686 => x"cc",
          2687 => x"38",
          2688 => x"39",
          2689 => x"55",
          2690 => x"52",
          2691 => x"d5",
          2692 => x"cc",
          2693 => x"0c",
          2694 => x"0c",
          2695 => x"53",
          2696 => x"80",
          2697 => x"85",
          2698 => x"94",
          2699 => x"2a",
          2700 => x"0c",
          2701 => x"06",
          2702 => x"9c",
          2703 => x"58",
          2704 => x"cc",
          2705 => x"0d",
          2706 => x"0d",
          2707 => x"90",
          2708 => x"05",
          2709 => x"f0",
          2710 => x"27",
          2711 => x"0b",
          2712 => x"98",
          2713 => x"84",
          2714 => x"2e",
          2715 => x"76",
          2716 => x"58",
          2717 => x"38",
          2718 => x"15",
          2719 => x"08",
          2720 => x"38",
          2721 => x"88",
          2722 => x"53",
          2723 => x"81",
          2724 => x"c0",
          2725 => x"22",
          2726 => x"89",
          2727 => x"72",
          2728 => x"74",
          2729 => x"f3",
          2730 => x"dc",
          2731 => x"82",
          2732 => x"81",
          2733 => x"27",
          2734 => x"81",
          2735 => x"cc",
          2736 => x"80",
          2737 => x"16",
          2738 => x"cc",
          2739 => x"ca",
          2740 => x"38",
          2741 => x"0c",
          2742 => x"dd",
          2743 => x"08",
          2744 => x"f9",
          2745 => x"dc",
          2746 => x"87",
          2747 => x"cc",
          2748 => x"80",
          2749 => x"55",
          2750 => x"08",
          2751 => x"38",
          2752 => x"dc",
          2753 => x"2e",
          2754 => x"dc",
          2755 => x"75",
          2756 => x"3f",
          2757 => x"08",
          2758 => x"94",
          2759 => x"52",
          2760 => x"c1",
          2761 => x"cc",
          2762 => x"0c",
          2763 => x"0c",
          2764 => x"05",
          2765 => x"80",
          2766 => x"dc",
          2767 => x"3d",
          2768 => x"3d",
          2769 => x"71",
          2770 => x"57",
          2771 => x"51",
          2772 => x"81",
          2773 => x"54",
          2774 => x"08",
          2775 => x"81",
          2776 => x"56",
          2777 => x"52",
          2778 => x"83",
          2779 => x"cc",
          2780 => x"dc",
          2781 => x"d2",
          2782 => x"cc",
          2783 => x"08",
          2784 => x"54",
          2785 => x"e5",
          2786 => x"06",
          2787 => x"58",
          2788 => x"08",
          2789 => x"38",
          2790 => x"75",
          2791 => x"80",
          2792 => x"81",
          2793 => x"7a",
          2794 => x"06",
          2795 => x"39",
          2796 => x"08",
          2797 => x"76",
          2798 => x"3f",
          2799 => x"08",
          2800 => x"cc",
          2801 => x"ff",
          2802 => x"84",
          2803 => x"06",
          2804 => x"54",
          2805 => x"cc",
          2806 => x"0d",
          2807 => x"0d",
          2808 => x"52",
          2809 => x"3f",
          2810 => x"08",
          2811 => x"06",
          2812 => x"51",
          2813 => x"83",
          2814 => x"06",
          2815 => x"14",
          2816 => x"3f",
          2817 => x"08",
          2818 => x"07",
          2819 => x"dc",
          2820 => x"3d",
          2821 => x"3d",
          2822 => x"70",
          2823 => x"06",
          2824 => x"53",
          2825 => x"ed",
          2826 => x"33",
          2827 => x"83",
          2828 => x"06",
          2829 => x"90",
          2830 => x"15",
          2831 => x"3f",
          2832 => x"04",
          2833 => x"7b",
          2834 => x"84",
          2835 => x"58",
          2836 => x"80",
          2837 => x"38",
          2838 => x"52",
          2839 => x"8f",
          2840 => x"cc",
          2841 => x"dc",
          2842 => x"f5",
          2843 => x"08",
          2844 => x"53",
          2845 => x"84",
          2846 => x"39",
          2847 => x"70",
          2848 => x"81",
          2849 => x"51",
          2850 => x"16",
          2851 => x"cc",
          2852 => x"81",
          2853 => x"38",
          2854 => x"ae",
          2855 => x"81",
          2856 => x"54",
          2857 => x"2e",
          2858 => x"8f",
          2859 => x"81",
          2860 => x"76",
          2861 => x"54",
          2862 => x"09",
          2863 => x"38",
          2864 => x"7a",
          2865 => x"80",
          2866 => x"fa",
          2867 => x"dc",
          2868 => x"81",
          2869 => x"89",
          2870 => x"08",
          2871 => x"86",
          2872 => x"98",
          2873 => x"81",
          2874 => x"8b",
          2875 => x"fb",
          2876 => x"70",
          2877 => x"81",
          2878 => x"fc",
          2879 => x"dc",
          2880 => x"81",
          2881 => x"b4",
          2882 => x"08",
          2883 => x"ec",
          2884 => x"dc",
          2885 => x"81",
          2886 => x"a0",
          2887 => x"81",
          2888 => x"52",
          2889 => x"51",
          2890 => x"8b",
          2891 => x"52",
          2892 => x"51",
          2893 => x"81",
          2894 => x"34",
          2895 => x"cc",
          2896 => x"0d",
          2897 => x"0d",
          2898 => x"98",
          2899 => x"70",
          2900 => x"ec",
          2901 => x"dc",
          2902 => x"38",
          2903 => x"53",
          2904 => x"81",
          2905 => x"34",
          2906 => x"04",
          2907 => x"78",
          2908 => x"80",
          2909 => x"34",
          2910 => x"80",
          2911 => x"38",
          2912 => x"18",
          2913 => x"9c",
          2914 => x"70",
          2915 => x"56",
          2916 => x"a0",
          2917 => x"71",
          2918 => x"81",
          2919 => x"81",
          2920 => x"89",
          2921 => x"06",
          2922 => x"73",
          2923 => x"55",
          2924 => x"55",
          2925 => x"81",
          2926 => x"81",
          2927 => x"74",
          2928 => x"75",
          2929 => x"52",
          2930 => x"13",
          2931 => x"08",
          2932 => x"33",
          2933 => x"9c",
          2934 => x"11",
          2935 => x"8a",
          2936 => x"cc",
          2937 => x"96",
          2938 => x"e7",
          2939 => x"cc",
          2940 => x"23",
          2941 => x"e7",
          2942 => x"dc",
          2943 => x"17",
          2944 => x"0d",
          2945 => x"0d",
          2946 => x"5e",
          2947 => x"70",
          2948 => x"55",
          2949 => x"83",
          2950 => x"73",
          2951 => x"91",
          2952 => x"2e",
          2953 => x"1d",
          2954 => x"0c",
          2955 => x"15",
          2956 => x"70",
          2957 => x"56",
          2958 => x"09",
          2959 => x"38",
          2960 => x"80",
          2961 => x"30",
          2962 => x"78",
          2963 => x"54",
          2964 => x"73",
          2965 => x"60",
          2966 => x"54",
          2967 => x"96",
          2968 => x"0b",
          2969 => x"80",
          2970 => x"f6",
          2971 => x"dc",
          2972 => x"85",
          2973 => x"3d",
          2974 => x"5c",
          2975 => x"53",
          2976 => x"51",
          2977 => x"80",
          2978 => x"88",
          2979 => x"5c",
          2980 => x"09",
          2981 => x"d4",
          2982 => x"70",
          2983 => x"71",
          2984 => x"30",
          2985 => x"73",
          2986 => x"51",
          2987 => x"57",
          2988 => x"38",
          2989 => x"75",
          2990 => x"17",
          2991 => x"75",
          2992 => x"30",
          2993 => x"51",
          2994 => x"80",
          2995 => x"38",
          2996 => x"87",
          2997 => x"26",
          2998 => x"77",
          2999 => x"a4",
          3000 => x"27",
          3001 => x"a0",
          3002 => x"39",
          3003 => x"33",
          3004 => x"57",
          3005 => x"27",
          3006 => x"75",
          3007 => x"30",
          3008 => x"32",
          3009 => x"80",
          3010 => x"25",
          3011 => x"56",
          3012 => x"80",
          3013 => x"84",
          3014 => x"58",
          3015 => x"70",
          3016 => x"55",
          3017 => x"09",
          3018 => x"38",
          3019 => x"80",
          3020 => x"30",
          3021 => x"77",
          3022 => x"54",
          3023 => x"81",
          3024 => x"ae",
          3025 => x"06",
          3026 => x"54",
          3027 => x"74",
          3028 => x"80",
          3029 => x"7b",
          3030 => x"30",
          3031 => x"70",
          3032 => x"25",
          3033 => x"07",
          3034 => x"51",
          3035 => x"a7",
          3036 => x"8b",
          3037 => x"39",
          3038 => x"54",
          3039 => x"8c",
          3040 => x"ff",
          3041 => x"9c",
          3042 => x"54",
          3043 => x"e1",
          3044 => x"cc",
          3045 => x"b2",
          3046 => x"70",
          3047 => x"71",
          3048 => x"54",
          3049 => x"81",
          3050 => x"80",
          3051 => x"38",
          3052 => x"76",
          3053 => x"df",
          3054 => x"54",
          3055 => x"81",
          3056 => x"55",
          3057 => x"34",
          3058 => x"52",
          3059 => x"51",
          3060 => x"81",
          3061 => x"bf",
          3062 => x"16",
          3063 => x"26",
          3064 => x"16",
          3065 => x"06",
          3066 => x"17",
          3067 => x"34",
          3068 => x"fd",
          3069 => x"19",
          3070 => x"80",
          3071 => x"79",
          3072 => x"81",
          3073 => x"81",
          3074 => x"85",
          3075 => x"54",
          3076 => x"8f",
          3077 => x"86",
          3078 => x"39",
          3079 => x"f3",
          3080 => x"73",
          3081 => x"80",
          3082 => x"52",
          3083 => x"ce",
          3084 => x"cc",
          3085 => x"dc",
          3086 => x"d7",
          3087 => x"08",
          3088 => x"e6",
          3089 => x"dc",
          3090 => x"81",
          3091 => x"80",
          3092 => x"1b",
          3093 => x"55",
          3094 => x"2e",
          3095 => x"8b",
          3096 => x"06",
          3097 => x"1c",
          3098 => x"33",
          3099 => x"70",
          3100 => x"55",
          3101 => x"38",
          3102 => x"52",
          3103 => x"9f",
          3104 => x"cc",
          3105 => x"8b",
          3106 => x"7a",
          3107 => x"3f",
          3108 => x"75",
          3109 => x"57",
          3110 => x"2e",
          3111 => x"84",
          3112 => x"06",
          3113 => x"75",
          3114 => x"81",
          3115 => x"2a",
          3116 => x"73",
          3117 => x"38",
          3118 => x"54",
          3119 => x"fb",
          3120 => x"80",
          3121 => x"34",
          3122 => x"c1",
          3123 => x"06",
          3124 => x"38",
          3125 => x"39",
          3126 => x"70",
          3127 => x"54",
          3128 => x"86",
          3129 => x"84",
          3130 => x"06",
          3131 => x"73",
          3132 => x"38",
          3133 => x"83",
          3134 => x"b4",
          3135 => x"51",
          3136 => x"81",
          3137 => x"88",
          3138 => x"ea",
          3139 => x"dc",
          3140 => x"3d",
          3141 => x"3d",
          3142 => x"ff",
          3143 => x"71",
          3144 => x"5c",
          3145 => x"80",
          3146 => x"38",
          3147 => x"05",
          3148 => x"a0",
          3149 => x"71",
          3150 => x"38",
          3151 => x"71",
          3152 => x"81",
          3153 => x"38",
          3154 => x"11",
          3155 => x"06",
          3156 => x"70",
          3157 => x"38",
          3158 => x"81",
          3159 => x"05",
          3160 => x"76",
          3161 => x"38",
          3162 => x"cc",
          3163 => x"77",
          3164 => x"57",
          3165 => x"05",
          3166 => x"70",
          3167 => x"33",
          3168 => x"53",
          3169 => x"99",
          3170 => x"e0",
          3171 => x"ff",
          3172 => x"ff",
          3173 => x"70",
          3174 => x"38",
          3175 => x"81",
          3176 => x"51",
          3177 => x"9f",
          3178 => x"72",
          3179 => x"81",
          3180 => x"70",
          3181 => x"72",
          3182 => x"32",
          3183 => x"72",
          3184 => x"73",
          3185 => x"53",
          3186 => x"70",
          3187 => x"38",
          3188 => x"19",
          3189 => x"75",
          3190 => x"38",
          3191 => x"83",
          3192 => x"74",
          3193 => x"59",
          3194 => x"39",
          3195 => x"33",
          3196 => x"dc",
          3197 => x"3d",
          3198 => x"3d",
          3199 => x"80",
          3200 => x"34",
          3201 => x"17",
          3202 => x"75",
          3203 => x"3f",
          3204 => x"dc",
          3205 => x"80",
          3206 => x"16",
          3207 => x"3f",
          3208 => x"08",
          3209 => x"06",
          3210 => x"73",
          3211 => x"2e",
          3212 => x"80",
          3213 => x"0b",
          3214 => x"56",
          3215 => x"e9",
          3216 => x"06",
          3217 => x"57",
          3218 => x"32",
          3219 => x"80",
          3220 => x"51",
          3221 => x"8a",
          3222 => x"e8",
          3223 => x"06",
          3224 => x"53",
          3225 => x"52",
          3226 => x"51",
          3227 => x"81",
          3228 => x"55",
          3229 => x"08",
          3230 => x"38",
          3231 => x"cb",
          3232 => x"86",
          3233 => x"97",
          3234 => x"cc",
          3235 => x"dc",
          3236 => x"2e",
          3237 => x"55",
          3238 => x"cc",
          3239 => x"0d",
          3240 => x"0d",
          3241 => x"05",
          3242 => x"33",
          3243 => x"75",
          3244 => x"fc",
          3245 => x"dc",
          3246 => x"8b",
          3247 => x"81",
          3248 => x"24",
          3249 => x"81",
          3250 => x"84",
          3251 => x"e8",
          3252 => x"55",
          3253 => x"73",
          3254 => x"e6",
          3255 => x"0c",
          3256 => x"06",
          3257 => x"57",
          3258 => x"ae",
          3259 => x"33",
          3260 => x"3f",
          3261 => x"08",
          3262 => x"70",
          3263 => x"55",
          3264 => x"76",
          3265 => x"b8",
          3266 => x"2a",
          3267 => x"51",
          3268 => x"72",
          3269 => x"86",
          3270 => x"74",
          3271 => x"15",
          3272 => x"81",
          3273 => x"d7",
          3274 => x"dc",
          3275 => x"ff",
          3276 => x"06",
          3277 => x"56",
          3278 => x"38",
          3279 => x"8f",
          3280 => x"2a",
          3281 => x"51",
          3282 => x"72",
          3283 => x"80",
          3284 => x"52",
          3285 => x"3f",
          3286 => x"08",
          3287 => x"57",
          3288 => x"09",
          3289 => x"e2",
          3290 => x"74",
          3291 => x"56",
          3292 => x"33",
          3293 => x"72",
          3294 => x"38",
          3295 => x"51",
          3296 => x"81",
          3297 => x"57",
          3298 => x"84",
          3299 => x"ff",
          3300 => x"56",
          3301 => x"25",
          3302 => x"0b",
          3303 => x"56",
          3304 => x"05",
          3305 => x"83",
          3306 => x"2e",
          3307 => x"52",
          3308 => x"c6",
          3309 => x"cc",
          3310 => x"06",
          3311 => x"27",
          3312 => x"16",
          3313 => x"27",
          3314 => x"56",
          3315 => x"84",
          3316 => x"56",
          3317 => x"84",
          3318 => x"14",
          3319 => x"3f",
          3320 => x"08",
          3321 => x"06",
          3322 => x"80",
          3323 => x"06",
          3324 => x"80",
          3325 => x"db",
          3326 => x"dc",
          3327 => x"ff",
          3328 => x"77",
          3329 => x"d8",
          3330 => x"de",
          3331 => x"cc",
          3332 => x"9c",
          3333 => x"c4",
          3334 => x"15",
          3335 => x"14",
          3336 => x"70",
          3337 => x"51",
          3338 => x"56",
          3339 => x"84",
          3340 => x"81",
          3341 => x"71",
          3342 => x"16",
          3343 => x"53",
          3344 => x"23",
          3345 => x"8b",
          3346 => x"73",
          3347 => x"80",
          3348 => x"8d",
          3349 => x"39",
          3350 => x"51",
          3351 => x"81",
          3352 => x"53",
          3353 => x"08",
          3354 => x"72",
          3355 => x"8d",
          3356 => x"ce",
          3357 => x"14",
          3358 => x"3f",
          3359 => x"08",
          3360 => x"06",
          3361 => x"38",
          3362 => x"51",
          3363 => x"81",
          3364 => x"55",
          3365 => x"51",
          3366 => x"81",
          3367 => x"83",
          3368 => x"53",
          3369 => x"80",
          3370 => x"38",
          3371 => x"78",
          3372 => x"2a",
          3373 => x"78",
          3374 => x"86",
          3375 => x"22",
          3376 => x"31",
          3377 => x"b1",
          3378 => x"cc",
          3379 => x"dc",
          3380 => x"2e",
          3381 => x"81",
          3382 => x"80",
          3383 => x"f5",
          3384 => x"83",
          3385 => x"ff",
          3386 => x"38",
          3387 => x"9f",
          3388 => x"38",
          3389 => x"39",
          3390 => x"80",
          3391 => x"38",
          3392 => x"98",
          3393 => x"a0",
          3394 => x"1c",
          3395 => x"0c",
          3396 => x"17",
          3397 => x"76",
          3398 => x"81",
          3399 => x"80",
          3400 => x"d9",
          3401 => x"dc",
          3402 => x"ff",
          3403 => x"8d",
          3404 => x"8e",
          3405 => x"8a",
          3406 => x"14",
          3407 => x"3f",
          3408 => x"08",
          3409 => x"74",
          3410 => x"a2",
          3411 => x"79",
          3412 => x"ee",
          3413 => x"a8",
          3414 => x"15",
          3415 => x"2e",
          3416 => x"10",
          3417 => x"2a",
          3418 => x"05",
          3419 => x"ff",
          3420 => x"53",
          3421 => x"9c",
          3422 => x"81",
          3423 => x"0b",
          3424 => x"ff",
          3425 => x"0c",
          3426 => x"84",
          3427 => x"83",
          3428 => x"06",
          3429 => x"80",
          3430 => x"d8",
          3431 => x"dc",
          3432 => x"ff",
          3433 => x"72",
          3434 => x"81",
          3435 => x"38",
          3436 => x"73",
          3437 => x"3f",
          3438 => x"08",
          3439 => x"81",
          3440 => x"84",
          3441 => x"b2",
          3442 => x"87",
          3443 => x"cc",
          3444 => x"ff",
          3445 => x"82",
          3446 => x"09",
          3447 => x"c8",
          3448 => x"51",
          3449 => x"81",
          3450 => x"84",
          3451 => x"d2",
          3452 => x"06",
          3453 => x"98",
          3454 => x"ee",
          3455 => x"cc",
          3456 => x"85",
          3457 => x"09",
          3458 => x"38",
          3459 => x"51",
          3460 => x"81",
          3461 => x"90",
          3462 => x"a0",
          3463 => x"ca",
          3464 => x"cc",
          3465 => x"0c",
          3466 => x"81",
          3467 => x"81",
          3468 => x"81",
          3469 => x"72",
          3470 => x"80",
          3471 => x"0c",
          3472 => x"81",
          3473 => x"90",
          3474 => x"fb",
          3475 => x"54",
          3476 => x"80",
          3477 => x"73",
          3478 => x"80",
          3479 => x"72",
          3480 => x"80",
          3481 => x"86",
          3482 => x"15",
          3483 => x"71",
          3484 => x"81",
          3485 => x"81",
          3486 => x"d0",
          3487 => x"dc",
          3488 => x"06",
          3489 => x"38",
          3490 => x"54",
          3491 => x"80",
          3492 => x"71",
          3493 => x"81",
          3494 => x"87",
          3495 => x"fa",
          3496 => x"ab",
          3497 => x"58",
          3498 => x"05",
          3499 => x"e6",
          3500 => x"80",
          3501 => x"cc",
          3502 => x"38",
          3503 => x"08",
          3504 => x"dc",
          3505 => x"08",
          3506 => x"80",
          3507 => x"80",
          3508 => x"54",
          3509 => x"84",
          3510 => x"34",
          3511 => x"75",
          3512 => x"2e",
          3513 => x"53",
          3514 => x"53",
          3515 => x"f7",
          3516 => x"dc",
          3517 => x"73",
          3518 => x"0c",
          3519 => x"04",
          3520 => x"67",
          3521 => x"80",
          3522 => x"59",
          3523 => x"78",
          3524 => x"c8",
          3525 => x"06",
          3526 => x"3d",
          3527 => x"99",
          3528 => x"52",
          3529 => x"3f",
          3530 => x"08",
          3531 => x"cc",
          3532 => x"38",
          3533 => x"52",
          3534 => x"52",
          3535 => x"3f",
          3536 => x"08",
          3537 => x"cc",
          3538 => x"02",
          3539 => x"33",
          3540 => x"55",
          3541 => x"25",
          3542 => x"55",
          3543 => x"54",
          3544 => x"81",
          3545 => x"80",
          3546 => x"74",
          3547 => x"81",
          3548 => x"75",
          3549 => x"3f",
          3550 => x"08",
          3551 => x"02",
          3552 => x"91",
          3553 => x"81",
          3554 => x"82",
          3555 => x"06",
          3556 => x"80",
          3557 => x"88",
          3558 => x"39",
          3559 => x"58",
          3560 => x"38",
          3561 => x"70",
          3562 => x"54",
          3563 => x"81",
          3564 => x"52",
          3565 => x"a5",
          3566 => x"cc",
          3567 => x"88",
          3568 => x"62",
          3569 => x"d4",
          3570 => x"54",
          3571 => x"15",
          3572 => x"62",
          3573 => x"e8",
          3574 => x"52",
          3575 => x"51",
          3576 => x"7a",
          3577 => x"83",
          3578 => x"80",
          3579 => x"38",
          3580 => x"08",
          3581 => x"53",
          3582 => x"3d",
          3583 => x"dd",
          3584 => x"dc",
          3585 => x"81",
          3586 => x"82",
          3587 => x"39",
          3588 => x"38",
          3589 => x"33",
          3590 => x"70",
          3591 => x"55",
          3592 => x"2e",
          3593 => x"55",
          3594 => x"77",
          3595 => x"81",
          3596 => x"73",
          3597 => x"38",
          3598 => x"54",
          3599 => x"a0",
          3600 => x"82",
          3601 => x"52",
          3602 => x"a3",
          3603 => x"cc",
          3604 => x"18",
          3605 => x"55",
          3606 => x"cc",
          3607 => x"38",
          3608 => x"70",
          3609 => x"54",
          3610 => x"86",
          3611 => x"c0",
          3612 => x"b0",
          3613 => x"1b",
          3614 => x"1b",
          3615 => x"70",
          3616 => x"d9",
          3617 => x"cc",
          3618 => x"cc",
          3619 => x"0c",
          3620 => x"52",
          3621 => x"3f",
          3622 => x"08",
          3623 => x"08",
          3624 => x"77",
          3625 => x"86",
          3626 => x"1a",
          3627 => x"1a",
          3628 => x"91",
          3629 => x"0b",
          3630 => x"80",
          3631 => x"0c",
          3632 => x"70",
          3633 => x"54",
          3634 => x"81",
          3635 => x"dc",
          3636 => x"2e",
          3637 => x"81",
          3638 => x"94",
          3639 => x"17",
          3640 => x"2b",
          3641 => x"57",
          3642 => x"52",
          3643 => x"9f",
          3644 => x"cc",
          3645 => x"dc",
          3646 => x"26",
          3647 => x"55",
          3648 => x"08",
          3649 => x"81",
          3650 => x"79",
          3651 => x"31",
          3652 => x"70",
          3653 => x"25",
          3654 => x"76",
          3655 => x"81",
          3656 => x"55",
          3657 => x"38",
          3658 => x"0c",
          3659 => x"75",
          3660 => x"54",
          3661 => x"a2",
          3662 => x"7a",
          3663 => x"3f",
          3664 => x"08",
          3665 => x"55",
          3666 => x"89",
          3667 => x"cc",
          3668 => x"1a",
          3669 => x"80",
          3670 => x"54",
          3671 => x"cc",
          3672 => x"0d",
          3673 => x"0d",
          3674 => x"64",
          3675 => x"59",
          3676 => x"90",
          3677 => x"52",
          3678 => x"cf",
          3679 => x"cc",
          3680 => x"dc",
          3681 => x"38",
          3682 => x"55",
          3683 => x"86",
          3684 => x"82",
          3685 => x"19",
          3686 => x"55",
          3687 => x"80",
          3688 => x"38",
          3689 => x"0b",
          3690 => x"82",
          3691 => x"39",
          3692 => x"1a",
          3693 => x"82",
          3694 => x"19",
          3695 => x"08",
          3696 => x"7c",
          3697 => x"74",
          3698 => x"2e",
          3699 => x"94",
          3700 => x"83",
          3701 => x"56",
          3702 => x"38",
          3703 => x"22",
          3704 => x"89",
          3705 => x"55",
          3706 => x"75",
          3707 => x"19",
          3708 => x"39",
          3709 => x"52",
          3710 => x"93",
          3711 => x"cc",
          3712 => x"75",
          3713 => x"38",
          3714 => x"ff",
          3715 => x"98",
          3716 => x"19",
          3717 => x"51",
          3718 => x"81",
          3719 => x"80",
          3720 => x"38",
          3721 => x"08",
          3722 => x"2a",
          3723 => x"80",
          3724 => x"38",
          3725 => x"8a",
          3726 => x"5c",
          3727 => x"27",
          3728 => x"7a",
          3729 => x"54",
          3730 => x"52",
          3731 => x"51",
          3732 => x"81",
          3733 => x"fe",
          3734 => x"83",
          3735 => x"56",
          3736 => x"9f",
          3737 => x"08",
          3738 => x"74",
          3739 => x"38",
          3740 => x"b4",
          3741 => x"16",
          3742 => x"89",
          3743 => x"51",
          3744 => x"77",
          3745 => x"b9",
          3746 => x"1a",
          3747 => x"08",
          3748 => x"84",
          3749 => x"57",
          3750 => x"27",
          3751 => x"56",
          3752 => x"52",
          3753 => x"c7",
          3754 => x"cc",
          3755 => x"38",
          3756 => x"19",
          3757 => x"06",
          3758 => x"52",
          3759 => x"a2",
          3760 => x"31",
          3761 => x"7f",
          3762 => x"94",
          3763 => x"94",
          3764 => x"5c",
          3765 => x"80",
          3766 => x"dc",
          3767 => x"3d",
          3768 => x"3d",
          3769 => x"65",
          3770 => x"5d",
          3771 => x"0c",
          3772 => x"05",
          3773 => x"f6",
          3774 => x"dc",
          3775 => x"81",
          3776 => x"8a",
          3777 => x"33",
          3778 => x"2e",
          3779 => x"56",
          3780 => x"90",
          3781 => x"81",
          3782 => x"06",
          3783 => x"87",
          3784 => x"2e",
          3785 => x"95",
          3786 => x"91",
          3787 => x"56",
          3788 => x"81",
          3789 => x"34",
          3790 => x"8e",
          3791 => x"08",
          3792 => x"56",
          3793 => x"84",
          3794 => x"5c",
          3795 => x"82",
          3796 => x"18",
          3797 => x"ff",
          3798 => x"74",
          3799 => x"7e",
          3800 => x"ff",
          3801 => x"2a",
          3802 => x"7a",
          3803 => x"8c",
          3804 => x"08",
          3805 => x"38",
          3806 => x"39",
          3807 => x"52",
          3808 => x"e7",
          3809 => x"cc",
          3810 => x"dc",
          3811 => x"2e",
          3812 => x"74",
          3813 => x"91",
          3814 => x"2e",
          3815 => x"74",
          3816 => x"88",
          3817 => x"38",
          3818 => x"0c",
          3819 => x"15",
          3820 => x"08",
          3821 => x"06",
          3822 => x"51",
          3823 => x"81",
          3824 => x"fe",
          3825 => x"18",
          3826 => x"51",
          3827 => x"81",
          3828 => x"80",
          3829 => x"38",
          3830 => x"08",
          3831 => x"2a",
          3832 => x"80",
          3833 => x"38",
          3834 => x"8a",
          3835 => x"5b",
          3836 => x"27",
          3837 => x"7b",
          3838 => x"54",
          3839 => x"52",
          3840 => x"51",
          3841 => x"81",
          3842 => x"fe",
          3843 => x"b0",
          3844 => x"31",
          3845 => x"79",
          3846 => x"84",
          3847 => x"16",
          3848 => x"89",
          3849 => x"52",
          3850 => x"cc",
          3851 => x"55",
          3852 => x"16",
          3853 => x"2b",
          3854 => x"39",
          3855 => x"94",
          3856 => x"93",
          3857 => x"cd",
          3858 => x"dc",
          3859 => x"e3",
          3860 => x"b0",
          3861 => x"76",
          3862 => x"94",
          3863 => x"ff",
          3864 => x"71",
          3865 => x"7b",
          3866 => x"38",
          3867 => x"18",
          3868 => x"51",
          3869 => x"81",
          3870 => x"fd",
          3871 => x"53",
          3872 => x"18",
          3873 => x"06",
          3874 => x"51",
          3875 => x"7e",
          3876 => x"83",
          3877 => x"76",
          3878 => x"17",
          3879 => x"1e",
          3880 => x"18",
          3881 => x"0c",
          3882 => x"58",
          3883 => x"74",
          3884 => x"38",
          3885 => x"8c",
          3886 => x"90",
          3887 => x"33",
          3888 => x"55",
          3889 => x"34",
          3890 => x"81",
          3891 => x"90",
          3892 => x"f8",
          3893 => x"8b",
          3894 => x"53",
          3895 => x"f2",
          3896 => x"dc",
          3897 => x"81",
          3898 => x"80",
          3899 => x"16",
          3900 => x"2a",
          3901 => x"51",
          3902 => x"80",
          3903 => x"38",
          3904 => x"52",
          3905 => x"e7",
          3906 => x"cc",
          3907 => x"dc",
          3908 => x"d4",
          3909 => x"08",
          3910 => x"a0",
          3911 => x"73",
          3912 => x"88",
          3913 => x"74",
          3914 => x"51",
          3915 => x"8c",
          3916 => x"9c",
          3917 => x"fb",
          3918 => x"b2",
          3919 => x"15",
          3920 => x"3f",
          3921 => x"15",
          3922 => x"3f",
          3923 => x"0b",
          3924 => x"78",
          3925 => x"3f",
          3926 => x"08",
          3927 => x"81",
          3928 => x"57",
          3929 => x"34",
          3930 => x"cc",
          3931 => x"0d",
          3932 => x"0d",
          3933 => x"54",
          3934 => x"81",
          3935 => x"53",
          3936 => x"08",
          3937 => x"3d",
          3938 => x"73",
          3939 => x"3f",
          3940 => x"08",
          3941 => x"cc",
          3942 => x"81",
          3943 => x"74",
          3944 => x"dc",
          3945 => x"3d",
          3946 => x"3d",
          3947 => x"51",
          3948 => x"8b",
          3949 => x"81",
          3950 => x"24",
          3951 => x"dc",
          3952 => x"dc",
          3953 => x"52",
          3954 => x"cc",
          3955 => x"0d",
          3956 => x"0d",
          3957 => x"3d",
          3958 => x"94",
          3959 => x"c1",
          3960 => x"cc",
          3961 => x"dc",
          3962 => x"e0",
          3963 => x"63",
          3964 => x"d4",
          3965 => x"8d",
          3966 => x"cc",
          3967 => x"dc",
          3968 => x"38",
          3969 => x"05",
          3970 => x"2b",
          3971 => x"80",
          3972 => x"76",
          3973 => x"0c",
          3974 => x"02",
          3975 => x"70",
          3976 => x"81",
          3977 => x"56",
          3978 => x"9e",
          3979 => x"53",
          3980 => x"db",
          3981 => x"dc",
          3982 => x"15",
          3983 => x"81",
          3984 => x"84",
          3985 => x"06",
          3986 => x"55",
          3987 => x"cc",
          3988 => x"0d",
          3989 => x"0d",
          3990 => x"5b",
          3991 => x"80",
          3992 => x"ff",
          3993 => x"9f",
          3994 => x"b5",
          3995 => x"cc",
          3996 => x"dc",
          3997 => x"fc",
          3998 => x"7a",
          3999 => x"08",
          4000 => x"64",
          4001 => x"2e",
          4002 => x"a0",
          4003 => x"70",
          4004 => x"ea",
          4005 => x"cc",
          4006 => x"dc",
          4007 => x"d4",
          4008 => x"7b",
          4009 => x"3f",
          4010 => x"08",
          4011 => x"cc",
          4012 => x"38",
          4013 => x"51",
          4014 => x"81",
          4015 => x"45",
          4016 => x"51",
          4017 => x"81",
          4018 => x"57",
          4019 => x"08",
          4020 => x"80",
          4021 => x"da",
          4022 => x"dc",
          4023 => x"81",
          4024 => x"a4",
          4025 => x"7b",
          4026 => x"3f",
          4027 => x"cc",
          4028 => x"38",
          4029 => x"51",
          4030 => x"81",
          4031 => x"57",
          4032 => x"08",
          4033 => x"38",
          4034 => x"09",
          4035 => x"38",
          4036 => x"e0",
          4037 => x"dc",
          4038 => x"ff",
          4039 => x"74",
          4040 => x"3f",
          4041 => x"78",
          4042 => x"33",
          4043 => x"56",
          4044 => x"91",
          4045 => x"05",
          4046 => x"81",
          4047 => x"56",
          4048 => x"f5",
          4049 => x"54",
          4050 => x"81",
          4051 => x"80",
          4052 => x"78",
          4053 => x"55",
          4054 => x"11",
          4055 => x"18",
          4056 => x"58",
          4057 => x"34",
          4058 => x"ff",
          4059 => x"55",
          4060 => x"34",
          4061 => x"77",
          4062 => x"81",
          4063 => x"ff",
          4064 => x"55",
          4065 => x"34",
          4066 => x"dc",
          4067 => x"84",
          4068 => x"8c",
          4069 => x"70",
          4070 => x"56",
          4071 => x"76",
          4072 => x"81",
          4073 => x"70",
          4074 => x"56",
          4075 => x"82",
          4076 => x"78",
          4077 => x"80",
          4078 => x"27",
          4079 => x"19",
          4080 => x"7a",
          4081 => x"5c",
          4082 => x"55",
          4083 => x"7a",
          4084 => x"5c",
          4085 => x"2e",
          4086 => x"85",
          4087 => x"94",
          4088 => x"81",
          4089 => x"73",
          4090 => x"81",
          4091 => x"7a",
          4092 => x"38",
          4093 => x"76",
          4094 => x"0c",
          4095 => x"04",
          4096 => x"7b",
          4097 => x"fc",
          4098 => x"53",
          4099 => x"bb",
          4100 => x"cc",
          4101 => x"dc",
          4102 => x"fa",
          4103 => x"33",
          4104 => x"f2",
          4105 => x"08",
          4106 => x"27",
          4107 => x"15",
          4108 => x"2a",
          4109 => x"51",
          4110 => x"83",
          4111 => x"94",
          4112 => x"80",
          4113 => x"0c",
          4114 => x"2e",
          4115 => x"79",
          4116 => x"70",
          4117 => x"51",
          4118 => x"2e",
          4119 => x"52",
          4120 => x"ff",
          4121 => x"81",
          4122 => x"ff",
          4123 => x"70",
          4124 => x"ff",
          4125 => x"81",
          4126 => x"73",
          4127 => x"76",
          4128 => x"06",
          4129 => x"0c",
          4130 => x"98",
          4131 => x"58",
          4132 => x"39",
          4133 => x"54",
          4134 => x"73",
          4135 => x"cd",
          4136 => x"dc",
          4137 => x"81",
          4138 => x"81",
          4139 => x"38",
          4140 => x"08",
          4141 => x"9b",
          4142 => x"cc",
          4143 => x"0c",
          4144 => x"0c",
          4145 => x"81",
          4146 => x"76",
          4147 => x"38",
          4148 => x"94",
          4149 => x"94",
          4150 => x"16",
          4151 => x"2a",
          4152 => x"51",
          4153 => x"72",
          4154 => x"38",
          4155 => x"51",
          4156 => x"81",
          4157 => x"54",
          4158 => x"08",
          4159 => x"dc",
          4160 => x"a7",
          4161 => x"74",
          4162 => x"3f",
          4163 => x"08",
          4164 => x"2e",
          4165 => x"74",
          4166 => x"79",
          4167 => x"14",
          4168 => x"38",
          4169 => x"0c",
          4170 => x"94",
          4171 => x"94",
          4172 => x"83",
          4173 => x"72",
          4174 => x"38",
          4175 => x"51",
          4176 => x"81",
          4177 => x"94",
          4178 => x"91",
          4179 => x"53",
          4180 => x"81",
          4181 => x"34",
          4182 => x"39",
          4183 => x"81",
          4184 => x"05",
          4185 => x"08",
          4186 => x"08",
          4187 => x"38",
          4188 => x"0c",
          4189 => x"80",
          4190 => x"72",
          4191 => x"73",
          4192 => x"53",
          4193 => x"8c",
          4194 => x"16",
          4195 => x"38",
          4196 => x"0c",
          4197 => x"81",
          4198 => x"8b",
          4199 => x"f9",
          4200 => x"56",
          4201 => x"80",
          4202 => x"38",
          4203 => x"3d",
          4204 => x"8a",
          4205 => x"51",
          4206 => x"81",
          4207 => x"55",
          4208 => x"08",
          4209 => x"77",
          4210 => x"52",
          4211 => x"b5",
          4212 => x"cc",
          4213 => x"dc",
          4214 => x"c3",
          4215 => x"33",
          4216 => x"55",
          4217 => x"24",
          4218 => x"16",
          4219 => x"2a",
          4220 => x"51",
          4221 => x"80",
          4222 => x"9c",
          4223 => x"77",
          4224 => x"3f",
          4225 => x"08",
          4226 => x"77",
          4227 => x"22",
          4228 => x"74",
          4229 => x"ce",
          4230 => x"dc",
          4231 => x"74",
          4232 => x"81",
          4233 => x"85",
          4234 => x"74",
          4235 => x"38",
          4236 => x"74",
          4237 => x"dc",
          4238 => x"3d",
          4239 => x"3d",
          4240 => x"3d",
          4241 => x"70",
          4242 => x"ff",
          4243 => x"cc",
          4244 => x"81",
          4245 => x"73",
          4246 => x"0d",
          4247 => x"0d",
          4248 => x"3d",
          4249 => x"71",
          4250 => x"e7",
          4251 => x"dc",
          4252 => x"81",
          4253 => x"80",
          4254 => x"93",
          4255 => x"cc",
          4256 => x"51",
          4257 => x"81",
          4258 => x"53",
          4259 => x"81",
          4260 => x"52",
          4261 => x"ac",
          4262 => x"cc",
          4263 => x"dc",
          4264 => x"2e",
          4265 => x"85",
          4266 => x"87",
          4267 => x"cc",
          4268 => x"74",
          4269 => x"d5",
          4270 => x"52",
          4271 => x"89",
          4272 => x"cc",
          4273 => x"70",
          4274 => x"07",
          4275 => x"81",
          4276 => x"06",
          4277 => x"54",
          4278 => x"cc",
          4279 => x"0d",
          4280 => x"0d",
          4281 => x"53",
          4282 => x"53",
          4283 => x"56",
          4284 => x"81",
          4285 => x"55",
          4286 => x"08",
          4287 => x"52",
          4288 => x"81",
          4289 => x"cc",
          4290 => x"dc",
          4291 => x"38",
          4292 => x"05",
          4293 => x"2b",
          4294 => x"80",
          4295 => x"86",
          4296 => x"76",
          4297 => x"38",
          4298 => x"51",
          4299 => x"74",
          4300 => x"0c",
          4301 => x"04",
          4302 => x"63",
          4303 => x"80",
          4304 => x"ec",
          4305 => x"3d",
          4306 => x"3f",
          4307 => x"08",
          4308 => x"cc",
          4309 => x"38",
          4310 => x"73",
          4311 => x"08",
          4312 => x"13",
          4313 => x"58",
          4314 => x"26",
          4315 => x"7c",
          4316 => x"39",
          4317 => x"cc",
          4318 => x"81",
          4319 => x"dc",
          4320 => x"33",
          4321 => x"81",
          4322 => x"06",
          4323 => x"75",
          4324 => x"52",
          4325 => x"05",
          4326 => x"3f",
          4327 => x"08",
          4328 => x"38",
          4329 => x"08",
          4330 => x"38",
          4331 => x"08",
          4332 => x"dc",
          4333 => x"80",
          4334 => x"81",
          4335 => x"59",
          4336 => x"14",
          4337 => x"ca",
          4338 => x"39",
          4339 => x"81",
          4340 => x"57",
          4341 => x"38",
          4342 => x"18",
          4343 => x"ff",
          4344 => x"81",
          4345 => x"5b",
          4346 => x"08",
          4347 => x"7c",
          4348 => x"12",
          4349 => x"52",
          4350 => x"82",
          4351 => x"06",
          4352 => x"14",
          4353 => x"cb",
          4354 => x"cc",
          4355 => x"ff",
          4356 => x"70",
          4357 => x"82",
          4358 => x"51",
          4359 => x"b4",
          4360 => x"bb",
          4361 => x"dc",
          4362 => x"0a",
          4363 => x"70",
          4364 => x"84",
          4365 => x"51",
          4366 => x"ff",
          4367 => x"56",
          4368 => x"38",
          4369 => x"7c",
          4370 => x"0c",
          4371 => x"81",
          4372 => x"74",
          4373 => x"7a",
          4374 => x"0c",
          4375 => x"04",
          4376 => x"79",
          4377 => x"05",
          4378 => x"57",
          4379 => x"81",
          4380 => x"56",
          4381 => x"08",
          4382 => x"91",
          4383 => x"75",
          4384 => x"90",
          4385 => x"81",
          4386 => x"06",
          4387 => x"87",
          4388 => x"2e",
          4389 => x"94",
          4390 => x"73",
          4391 => x"27",
          4392 => x"73",
          4393 => x"dc",
          4394 => x"88",
          4395 => x"76",
          4396 => x"3f",
          4397 => x"08",
          4398 => x"0c",
          4399 => x"39",
          4400 => x"52",
          4401 => x"bf",
          4402 => x"dc",
          4403 => x"2e",
          4404 => x"83",
          4405 => x"81",
          4406 => x"81",
          4407 => x"06",
          4408 => x"56",
          4409 => x"a0",
          4410 => x"81",
          4411 => x"98",
          4412 => x"94",
          4413 => x"08",
          4414 => x"cc",
          4415 => x"51",
          4416 => x"81",
          4417 => x"56",
          4418 => x"8c",
          4419 => x"17",
          4420 => x"07",
          4421 => x"18",
          4422 => x"2e",
          4423 => x"91",
          4424 => x"55",
          4425 => x"cc",
          4426 => x"0d",
          4427 => x"0d",
          4428 => x"3d",
          4429 => x"52",
          4430 => x"da",
          4431 => x"dc",
          4432 => x"81",
          4433 => x"81",
          4434 => x"45",
          4435 => x"52",
          4436 => x"52",
          4437 => x"3f",
          4438 => x"08",
          4439 => x"cc",
          4440 => x"38",
          4441 => x"05",
          4442 => x"2a",
          4443 => x"51",
          4444 => x"55",
          4445 => x"38",
          4446 => x"54",
          4447 => x"81",
          4448 => x"80",
          4449 => x"70",
          4450 => x"54",
          4451 => x"81",
          4452 => x"52",
          4453 => x"c5",
          4454 => x"cc",
          4455 => x"2a",
          4456 => x"51",
          4457 => x"80",
          4458 => x"38",
          4459 => x"dc",
          4460 => x"15",
          4461 => x"86",
          4462 => x"81",
          4463 => x"5c",
          4464 => x"3d",
          4465 => x"c7",
          4466 => x"dc",
          4467 => x"81",
          4468 => x"80",
          4469 => x"dc",
          4470 => x"73",
          4471 => x"3f",
          4472 => x"08",
          4473 => x"cc",
          4474 => x"87",
          4475 => x"39",
          4476 => x"08",
          4477 => x"38",
          4478 => x"08",
          4479 => x"77",
          4480 => x"3f",
          4481 => x"08",
          4482 => x"08",
          4483 => x"dc",
          4484 => x"80",
          4485 => x"55",
          4486 => x"94",
          4487 => x"2e",
          4488 => x"53",
          4489 => x"51",
          4490 => x"81",
          4491 => x"55",
          4492 => x"78",
          4493 => x"fe",
          4494 => x"cc",
          4495 => x"81",
          4496 => x"a0",
          4497 => x"e9",
          4498 => x"53",
          4499 => x"05",
          4500 => x"51",
          4501 => x"81",
          4502 => x"54",
          4503 => x"08",
          4504 => x"78",
          4505 => x"8e",
          4506 => x"58",
          4507 => x"81",
          4508 => x"54",
          4509 => x"08",
          4510 => x"54",
          4511 => x"81",
          4512 => x"84",
          4513 => x"06",
          4514 => x"02",
          4515 => x"33",
          4516 => x"81",
          4517 => x"86",
          4518 => x"f6",
          4519 => x"74",
          4520 => x"70",
          4521 => x"c3",
          4522 => x"cc",
          4523 => x"56",
          4524 => x"08",
          4525 => x"54",
          4526 => x"08",
          4527 => x"81",
          4528 => x"82",
          4529 => x"cc",
          4530 => x"09",
          4531 => x"38",
          4532 => x"b4",
          4533 => x"b0",
          4534 => x"cc",
          4535 => x"51",
          4536 => x"81",
          4537 => x"54",
          4538 => x"08",
          4539 => x"8b",
          4540 => x"b4",
          4541 => x"b7",
          4542 => x"54",
          4543 => x"15",
          4544 => x"90",
          4545 => x"34",
          4546 => x"0a",
          4547 => x"19",
          4548 => x"9f",
          4549 => x"78",
          4550 => x"51",
          4551 => x"a0",
          4552 => x"11",
          4553 => x"05",
          4554 => x"b6",
          4555 => x"ae",
          4556 => x"15",
          4557 => x"78",
          4558 => x"53",
          4559 => x"3f",
          4560 => x"0b",
          4561 => x"77",
          4562 => x"3f",
          4563 => x"08",
          4564 => x"cc",
          4565 => x"82",
          4566 => x"52",
          4567 => x"51",
          4568 => x"3f",
          4569 => x"52",
          4570 => x"aa",
          4571 => x"90",
          4572 => x"34",
          4573 => x"0b",
          4574 => x"78",
          4575 => x"b6",
          4576 => x"cc",
          4577 => x"39",
          4578 => x"52",
          4579 => x"be",
          4580 => x"81",
          4581 => x"99",
          4582 => x"da",
          4583 => x"3d",
          4584 => x"d2",
          4585 => x"53",
          4586 => x"84",
          4587 => x"3d",
          4588 => x"3f",
          4589 => x"08",
          4590 => x"cc",
          4591 => x"38",
          4592 => x"3d",
          4593 => x"3d",
          4594 => x"cc",
          4595 => x"dc",
          4596 => x"81",
          4597 => x"82",
          4598 => x"81",
          4599 => x"81",
          4600 => x"86",
          4601 => x"aa",
          4602 => x"a4",
          4603 => x"a8",
          4604 => x"05",
          4605 => x"ea",
          4606 => x"77",
          4607 => x"70",
          4608 => x"b4",
          4609 => x"3d",
          4610 => x"51",
          4611 => x"81",
          4612 => x"55",
          4613 => x"08",
          4614 => x"6f",
          4615 => x"06",
          4616 => x"a2",
          4617 => x"92",
          4618 => x"81",
          4619 => x"dc",
          4620 => x"2e",
          4621 => x"81",
          4622 => x"51",
          4623 => x"81",
          4624 => x"55",
          4625 => x"08",
          4626 => x"68",
          4627 => x"a8",
          4628 => x"05",
          4629 => x"51",
          4630 => x"3f",
          4631 => x"33",
          4632 => x"8b",
          4633 => x"84",
          4634 => x"06",
          4635 => x"73",
          4636 => x"a0",
          4637 => x"8b",
          4638 => x"54",
          4639 => x"15",
          4640 => x"33",
          4641 => x"70",
          4642 => x"55",
          4643 => x"2e",
          4644 => x"6e",
          4645 => x"df",
          4646 => x"78",
          4647 => x"3f",
          4648 => x"08",
          4649 => x"ff",
          4650 => x"82",
          4651 => x"cc",
          4652 => x"80",
          4653 => x"dc",
          4654 => x"78",
          4655 => x"af",
          4656 => x"cc",
          4657 => x"d4",
          4658 => x"55",
          4659 => x"08",
          4660 => x"81",
          4661 => x"73",
          4662 => x"81",
          4663 => x"63",
          4664 => x"76",
          4665 => x"3f",
          4666 => x"0b",
          4667 => x"87",
          4668 => x"cc",
          4669 => x"77",
          4670 => x"3f",
          4671 => x"08",
          4672 => x"cc",
          4673 => x"78",
          4674 => x"aa",
          4675 => x"cc",
          4676 => x"81",
          4677 => x"a8",
          4678 => x"ed",
          4679 => x"80",
          4680 => x"02",
          4681 => x"df",
          4682 => x"57",
          4683 => x"3d",
          4684 => x"96",
          4685 => x"e9",
          4686 => x"cc",
          4687 => x"dc",
          4688 => x"cf",
          4689 => x"65",
          4690 => x"d4",
          4691 => x"b5",
          4692 => x"cc",
          4693 => x"dc",
          4694 => x"38",
          4695 => x"05",
          4696 => x"06",
          4697 => x"73",
          4698 => x"a7",
          4699 => x"09",
          4700 => x"71",
          4701 => x"06",
          4702 => x"55",
          4703 => x"15",
          4704 => x"81",
          4705 => x"34",
          4706 => x"b4",
          4707 => x"dc",
          4708 => x"74",
          4709 => x"0c",
          4710 => x"04",
          4711 => x"64",
          4712 => x"93",
          4713 => x"52",
          4714 => x"d1",
          4715 => x"dc",
          4716 => x"81",
          4717 => x"80",
          4718 => x"58",
          4719 => x"3d",
          4720 => x"c8",
          4721 => x"dc",
          4722 => x"81",
          4723 => x"b4",
          4724 => x"c7",
          4725 => x"a0",
          4726 => x"55",
          4727 => x"84",
          4728 => x"17",
          4729 => x"2b",
          4730 => x"96",
          4731 => x"b0",
          4732 => x"54",
          4733 => x"15",
          4734 => x"ff",
          4735 => x"81",
          4736 => x"55",
          4737 => x"cc",
          4738 => x"0d",
          4739 => x"0d",
          4740 => x"5a",
          4741 => x"3d",
          4742 => x"99",
          4743 => x"81",
          4744 => x"cc",
          4745 => x"cc",
          4746 => x"81",
          4747 => x"07",
          4748 => x"55",
          4749 => x"2e",
          4750 => x"81",
          4751 => x"55",
          4752 => x"2e",
          4753 => x"7b",
          4754 => x"80",
          4755 => x"70",
          4756 => x"be",
          4757 => x"dc",
          4758 => x"81",
          4759 => x"80",
          4760 => x"52",
          4761 => x"dc",
          4762 => x"cc",
          4763 => x"dc",
          4764 => x"38",
          4765 => x"08",
          4766 => x"08",
          4767 => x"56",
          4768 => x"19",
          4769 => x"59",
          4770 => x"74",
          4771 => x"56",
          4772 => x"ec",
          4773 => x"75",
          4774 => x"74",
          4775 => x"2e",
          4776 => x"16",
          4777 => x"33",
          4778 => x"73",
          4779 => x"38",
          4780 => x"84",
          4781 => x"06",
          4782 => x"7a",
          4783 => x"76",
          4784 => x"07",
          4785 => x"54",
          4786 => x"80",
          4787 => x"80",
          4788 => x"7b",
          4789 => x"53",
          4790 => x"93",
          4791 => x"cc",
          4792 => x"dc",
          4793 => x"38",
          4794 => x"55",
          4795 => x"56",
          4796 => x"8b",
          4797 => x"56",
          4798 => x"83",
          4799 => x"75",
          4800 => x"51",
          4801 => x"3f",
          4802 => x"08",
          4803 => x"81",
          4804 => x"98",
          4805 => x"e6",
          4806 => x"53",
          4807 => x"b8",
          4808 => x"3d",
          4809 => x"3f",
          4810 => x"08",
          4811 => x"08",
          4812 => x"dc",
          4813 => x"98",
          4814 => x"a0",
          4815 => x"70",
          4816 => x"ae",
          4817 => x"6d",
          4818 => x"81",
          4819 => x"57",
          4820 => x"74",
          4821 => x"38",
          4822 => x"81",
          4823 => x"81",
          4824 => x"52",
          4825 => x"89",
          4826 => x"cc",
          4827 => x"a5",
          4828 => x"33",
          4829 => x"54",
          4830 => x"3f",
          4831 => x"08",
          4832 => x"38",
          4833 => x"76",
          4834 => x"05",
          4835 => x"39",
          4836 => x"08",
          4837 => x"15",
          4838 => x"ff",
          4839 => x"73",
          4840 => x"38",
          4841 => x"83",
          4842 => x"56",
          4843 => x"75",
          4844 => x"81",
          4845 => x"33",
          4846 => x"2e",
          4847 => x"52",
          4848 => x"51",
          4849 => x"3f",
          4850 => x"08",
          4851 => x"ff",
          4852 => x"38",
          4853 => x"88",
          4854 => x"8a",
          4855 => x"38",
          4856 => x"ec",
          4857 => x"75",
          4858 => x"74",
          4859 => x"73",
          4860 => x"05",
          4861 => x"17",
          4862 => x"70",
          4863 => x"34",
          4864 => x"70",
          4865 => x"ff",
          4866 => x"55",
          4867 => x"26",
          4868 => x"8b",
          4869 => x"86",
          4870 => x"e5",
          4871 => x"38",
          4872 => x"99",
          4873 => x"05",
          4874 => x"70",
          4875 => x"73",
          4876 => x"81",
          4877 => x"ff",
          4878 => x"ed",
          4879 => x"80",
          4880 => x"91",
          4881 => x"55",
          4882 => x"3f",
          4883 => x"08",
          4884 => x"cc",
          4885 => x"38",
          4886 => x"51",
          4887 => x"3f",
          4888 => x"08",
          4889 => x"cc",
          4890 => x"76",
          4891 => x"67",
          4892 => x"34",
          4893 => x"81",
          4894 => x"84",
          4895 => x"06",
          4896 => x"80",
          4897 => x"2e",
          4898 => x"81",
          4899 => x"ff",
          4900 => x"81",
          4901 => x"54",
          4902 => x"08",
          4903 => x"53",
          4904 => x"08",
          4905 => x"ff",
          4906 => x"67",
          4907 => x"8b",
          4908 => x"53",
          4909 => x"51",
          4910 => x"3f",
          4911 => x"0b",
          4912 => x"79",
          4913 => x"ee",
          4914 => x"cc",
          4915 => x"55",
          4916 => x"cc",
          4917 => x"0d",
          4918 => x"0d",
          4919 => x"88",
          4920 => x"05",
          4921 => x"fc",
          4922 => x"54",
          4923 => x"d2",
          4924 => x"dc",
          4925 => x"81",
          4926 => x"82",
          4927 => x"1a",
          4928 => x"82",
          4929 => x"80",
          4930 => x"8c",
          4931 => x"78",
          4932 => x"1a",
          4933 => x"2a",
          4934 => x"51",
          4935 => x"90",
          4936 => x"82",
          4937 => x"58",
          4938 => x"81",
          4939 => x"39",
          4940 => x"22",
          4941 => x"70",
          4942 => x"56",
          4943 => x"fc",
          4944 => x"14",
          4945 => x"30",
          4946 => x"9f",
          4947 => x"cc",
          4948 => x"19",
          4949 => x"5a",
          4950 => x"81",
          4951 => x"38",
          4952 => x"77",
          4953 => x"82",
          4954 => x"56",
          4955 => x"74",
          4956 => x"ff",
          4957 => x"81",
          4958 => x"55",
          4959 => x"75",
          4960 => x"82",
          4961 => x"cc",
          4962 => x"ff",
          4963 => x"dc",
          4964 => x"2e",
          4965 => x"81",
          4966 => x"8e",
          4967 => x"56",
          4968 => x"09",
          4969 => x"38",
          4970 => x"59",
          4971 => x"77",
          4972 => x"06",
          4973 => x"87",
          4974 => x"39",
          4975 => x"ba",
          4976 => x"55",
          4977 => x"2e",
          4978 => x"15",
          4979 => x"2e",
          4980 => x"83",
          4981 => x"75",
          4982 => x"7e",
          4983 => x"a8",
          4984 => x"cc",
          4985 => x"dc",
          4986 => x"ce",
          4987 => x"16",
          4988 => x"56",
          4989 => x"38",
          4990 => x"19",
          4991 => x"8c",
          4992 => x"7d",
          4993 => x"38",
          4994 => x"0c",
          4995 => x"0c",
          4996 => x"80",
          4997 => x"73",
          4998 => x"98",
          4999 => x"05",
          5000 => x"57",
          5001 => x"26",
          5002 => x"7b",
          5003 => x"0c",
          5004 => x"81",
          5005 => x"84",
          5006 => x"54",
          5007 => x"cc",
          5008 => x"0d",
          5009 => x"0d",
          5010 => x"88",
          5011 => x"05",
          5012 => x"54",
          5013 => x"c5",
          5014 => x"56",
          5015 => x"dc",
          5016 => x"8b",
          5017 => x"dc",
          5018 => x"29",
          5019 => x"05",
          5020 => x"55",
          5021 => x"84",
          5022 => x"34",
          5023 => x"08",
          5024 => x"5f",
          5025 => x"51",
          5026 => x"3f",
          5027 => x"08",
          5028 => x"70",
          5029 => x"57",
          5030 => x"8b",
          5031 => x"82",
          5032 => x"06",
          5033 => x"56",
          5034 => x"38",
          5035 => x"05",
          5036 => x"7e",
          5037 => x"f0",
          5038 => x"cc",
          5039 => x"67",
          5040 => x"2e",
          5041 => x"82",
          5042 => x"8b",
          5043 => x"75",
          5044 => x"80",
          5045 => x"81",
          5046 => x"2e",
          5047 => x"80",
          5048 => x"38",
          5049 => x"0a",
          5050 => x"ff",
          5051 => x"55",
          5052 => x"86",
          5053 => x"8a",
          5054 => x"89",
          5055 => x"2a",
          5056 => x"77",
          5057 => x"59",
          5058 => x"81",
          5059 => x"70",
          5060 => x"07",
          5061 => x"56",
          5062 => x"38",
          5063 => x"05",
          5064 => x"7e",
          5065 => x"80",
          5066 => x"81",
          5067 => x"8a",
          5068 => x"83",
          5069 => x"06",
          5070 => x"08",
          5071 => x"74",
          5072 => x"41",
          5073 => x"56",
          5074 => x"8a",
          5075 => x"61",
          5076 => x"55",
          5077 => x"27",
          5078 => x"93",
          5079 => x"80",
          5080 => x"38",
          5081 => x"70",
          5082 => x"43",
          5083 => x"95",
          5084 => x"06",
          5085 => x"2e",
          5086 => x"77",
          5087 => x"74",
          5088 => x"83",
          5089 => x"06",
          5090 => x"82",
          5091 => x"2e",
          5092 => x"78",
          5093 => x"2e",
          5094 => x"80",
          5095 => x"ae",
          5096 => x"2a",
          5097 => x"81",
          5098 => x"56",
          5099 => x"2e",
          5100 => x"77",
          5101 => x"81",
          5102 => x"79",
          5103 => x"70",
          5104 => x"5a",
          5105 => x"86",
          5106 => x"27",
          5107 => x"52",
          5108 => x"f7",
          5109 => x"dc",
          5110 => x"29",
          5111 => x"70",
          5112 => x"55",
          5113 => x"0b",
          5114 => x"08",
          5115 => x"05",
          5116 => x"ff",
          5117 => x"27",
          5118 => x"88",
          5119 => x"ae",
          5120 => x"2a",
          5121 => x"81",
          5122 => x"56",
          5123 => x"2e",
          5124 => x"77",
          5125 => x"81",
          5126 => x"79",
          5127 => x"70",
          5128 => x"5a",
          5129 => x"86",
          5130 => x"27",
          5131 => x"52",
          5132 => x"f6",
          5133 => x"dc",
          5134 => x"84",
          5135 => x"dc",
          5136 => x"f5",
          5137 => x"81",
          5138 => x"cc",
          5139 => x"dc",
          5140 => x"71",
          5141 => x"83",
          5142 => x"5e",
          5143 => x"89",
          5144 => x"5c",
          5145 => x"1c",
          5146 => x"05",
          5147 => x"ff",
          5148 => x"70",
          5149 => x"31",
          5150 => x"57",
          5151 => x"83",
          5152 => x"06",
          5153 => x"1c",
          5154 => x"5c",
          5155 => x"1d",
          5156 => x"29",
          5157 => x"31",
          5158 => x"55",
          5159 => x"87",
          5160 => x"7c",
          5161 => x"7a",
          5162 => x"31",
          5163 => x"f5",
          5164 => x"dc",
          5165 => x"7d",
          5166 => x"81",
          5167 => x"81",
          5168 => x"83",
          5169 => x"80",
          5170 => x"87",
          5171 => x"81",
          5172 => x"fd",
          5173 => x"f8",
          5174 => x"2e",
          5175 => x"80",
          5176 => x"ff",
          5177 => x"dc",
          5178 => x"a0",
          5179 => x"38",
          5180 => x"74",
          5181 => x"86",
          5182 => x"fd",
          5183 => x"81",
          5184 => x"80",
          5185 => x"83",
          5186 => x"39",
          5187 => x"08",
          5188 => x"92",
          5189 => x"b8",
          5190 => x"59",
          5191 => x"27",
          5192 => x"86",
          5193 => x"55",
          5194 => x"09",
          5195 => x"38",
          5196 => x"f5",
          5197 => x"38",
          5198 => x"55",
          5199 => x"86",
          5200 => x"80",
          5201 => x"7a",
          5202 => x"b9",
          5203 => x"81",
          5204 => x"7a",
          5205 => x"8a",
          5206 => x"52",
          5207 => x"ff",
          5208 => x"79",
          5209 => x"7b",
          5210 => x"06",
          5211 => x"51",
          5212 => x"3f",
          5213 => x"1c",
          5214 => x"32",
          5215 => x"96",
          5216 => x"06",
          5217 => x"91",
          5218 => x"a1",
          5219 => x"55",
          5220 => x"ff",
          5221 => x"74",
          5222 => x"06",
          5223 => x"51",
          5224 => x"3f",
          5225 => x"52",
          5226 => x"ff",
          5227 => x"f8",
          5228 => x"34",
          5229 => x"1b",
          5230 => x"d9",
          5231 => x"52",
          5232 => x"ff",
          5233 => x"60",
          5234 => x"51",
          5235 => x"3f",
          5236 => x"09",
          5237 => x"cb",
          5238 => x"b2",
          5239 => x"c3",
          5240 => x"a0",
          5241 => x"52",
          5242 => x"ff",
          5243 => x"82",
          5244 => x"51",
          5245 => x"3f",
          5246 => x"1b",
          5247 => x"95",
          5248 => x"b2",
          5249 => x"a0",
          5250 => x"80",
          5251 => x"1c",
          5252 => x"80",
          5253 => x"93",
          5254 => x"e4",
          5255 => x"1b",
          5256 => x"82",
          5257 => x"52",
          5258 => x"ff",
          5259 => x"7c",
          5260 => x"06",
          5261 => x"51",
          5262 => x"3f",
          5263 => x"a4",
          5264 => x"0b",
          5265 => x"93",
          5266 => x"f8",
          5267 => x"51",
          5268 => x"3f",
          5269 => x"52",
          5270 => x"70",
          5271 => x"9f",
          5272 => x"54",
          5273 => x"52",
          5274 => x"9b",
          5275 => x"56",
          5276 => x"08",
          5277 => x"7d",
          5278 => x"81",
          5279 => x"38",
          5280 => x"86",
          5281 => x"52",
          5282 => x"9b",
          5283 => x"80",
          5284 => x"7a",
          5285 => x"ed",
          5286 => x"85",
          5287 => x"7a",
          5288 => x"8f",
          5289 => x"85",
          5290 => x"83",
          5291 => x"ff",
          5292 => x"ff",
          5293 => x"e8",
          5294 => x"9e",
          5295 => x"52",
          5296 => x"51",
          5297 => x"3f",
          5298 => x"52",
          5299 => x"9e",
          5300 => x"54",
          5301 => x"53",
          5302 => x"51",
          5303 => x"3f",
          5304 => x"16",
          5305 => x"7e",
          5306 => x"d8",
          5307 => x"80",
          5308 => x"ff",
          5309 => x"7f",
          5310 => x"7d",
          5311 => x"81",
          5312 => x"f8",
          5313 => x"ff",
          5314 => x"ff",
          5315 => x"51",
          5316 => x"3f",
          5317 => x"88",
          5318 => x"39",
          5319 => x"f8",
          5320 => x"2e",
          5321 => x"55",
          5322 => x"51",
          5323 => x"3f",
          5324 => x"57",
          5325 => x"83",
          5326 => x"76",
          5327 => x"7a",
          5328 => x"ff",
          5329 => x"81",
          5330 => x"82",
          5331 => x"80",
          5332 => x"cc",
          5333 => x"51",
          5334 => x"3f",
          5335 => x"78",
          5336 => x"74",
          5337 => x"18",
          5338 => x"2e",
          5339 => x"79",
          5340 => x"2e",
          5341 => x"55",
          5342 => x"62",
          5343 => x"74",
          5344 => x"75",
          5345 => x"7e",
          5346 => x"b8",
          5347 => x"cc",
          5348 => x"38",
          5349 => x"78",
          5350 => x"74",
          5351 => x"56",
          5352 => x"93",
          5353 => x"66",
          5354 => x"26",
          5355 => x"56",
          5356 => x"83",
          5357 => x"64",
          5358 => x"77",
          5359 => x"84",
          5360 => x"52",
          5361 => x"9d",
          5362 => x"d4",
          5363 => x"51",
          5364 => x"3f",
          5365 => x"55",
          5366 => x"81",
          5367 => x"34",
          5368 => x"16",
          5369 => x"16",
          5370 => x"16",
          5371 => x"05",
          5372 => x"c1",
          5373 => x"fe",
          5374 => x"fe",
          5375 => x"34",
          5376 => x"08",
          5377 => x"07",
          5378 => x"16",
          5379 => x"cc",
          5380 => x"34",
          5381 => x"c6",
          5382 => x"9c",
          5383 => x"52",
          5384 => x"51",
          5385 => x"3f",
          5386 => x"53",
          5387 => x"51",
          5388 => x"3f",
          5389 => x"dc",
          5390 => x"38",
          5391 => x"52",
          5392 => x"99",
          5393 => x"56",
          5394 => x"08",
          5395 => x"39",
          5396 => x"39",
          5397 => x"39",
          5398 => x"08",
          5399 => x"dc",
          5400 => x"3d",
          5401 => x"3d",
          5402 => x"5b",
          5403 => x"60",
          5404 => x"57",
          5405 => x"25",
          5406 => x"3d",
          5407 => x"55",
          5408 => x"15",
          5409 => x"c9",
          5410 => x"81",
          5411 => x"06",
          5412 => x"3d",
          5413 => x"8d",
          5414 => x"74",
          5415 => x"05",
          5416 => x"17",
          5417 => x"2e",
          5418 => x"c9",
          5419 => x"34",
          5420 => x"83",
          5421 => x"74",
          5422 => x"0c",
          5423 => x"04",
          5424 => x"78",
          5425 => x"55",
          5426 => x"80",
          5427 => x"38",
          5428 => x"77",
          5429 => x"33",
          5430 => x"39",
          5431 => x"80",
          5432 => x"56",
          5433 => x"83",
          5434 => x"73",
          5435 => x"2a",
          5436 => x"53",
          5437 => x"73",
          5438 => x"81",
          5439 => x"72",
          5440 => x"05",
          5441 => x"56",
          5442 => x"81",
          5443 => x"77",
          5444 => x"08",
          5445 => x"f3",
          5446 => x"dc",
          5447 => x"38",
          5448 => x"53",
          5449 => x"ff",
          5450 => x"16",
          5451 => x"06",
          5452 => x"76",
          5453 => x"ff",
          5454 => x"dc",
          5455 => x"3d",
          5456 => x"3d",
          5457 => x"71",
          5458 => x"8e",
          5459 => x"29",
          5460 => x"05",
          5461 => x"04",
          5462 => x"51",
          5463 => x"81",
          5464 => x"80",
          5465 => x"cf",
          5466 => x"f2",
          5467 => x"9c",
          5468 => x"39",
          5469 => x"51",
          5470 => x"81",
          5471 => x"80",
          5472 => x"cf",
          5473 => x"d6",
          5474 => x"e0",
          5475 => x"39",
          5476 => x"51",
          5477 => x"81",
          5478 => x"80",
          5479 => x"d0",
          5480 => x"39",
          5481 => x"51",
          5482 => x"d0",
          5483 => x"39",
          5484 => x"51",
          5485 => x"d1",
          5486 => x"39",
          5487 => x"51",
          5488 => x"d1",
          5489 => x"39",
          5490 => x"51",
          5491 => x"d1",
          5492 => x"39",
          5493 => x"51",
          5494 => x"d2",
          5495 => x"86",
          5496 => x"3d",
          5497 => x"3d",
          5498 => x"56",
          5499 => x"e7",
          5500 => x"74",
          5501 => x"e8",
          5502 => x"39",
          5503 => x"74",
          5504 => x"f5",
          5505 => x"cc",
          5506 => x"51",
          5507 => x"3f",
          5508 => x"08",
          5509 => x"75",
          5510 => x"b0",
          5511 => x"c4",
          5512 => x"0d",
          5513 => x"0d",
          5514 => x"05",
          5515 => x"33",
          5516 => x"68",
          5517 => x"7a",
          5518 => x"51",
          5519 => x"78",
          5520 => x"ff",
          5521 => x"81",
          5522 => x"07",
          5523 => x"06",
          5524 => x"56",
          5525 => x"38",
          5526 => x"52",
          5527 => x"52",
          5528 => x"3f",
          5529 => x"08",
          5530 => x"cc",
          5531 => x"81",
          5532 => x"87",
          5533 => x"0c",
          5534 => x"08",
          5535 => x"d4",
          5536 => x"80",
          5537 => x"75",
          5538 => x"3f",
          5539 => x"08",
          5540 => x"cc",
          5541 => x"7a",
          5542 => x"2e",
          5543 => x"19",
          5544 => x"59",
          5545 => x"3d",
          5546 => x"cd",
          5547 => x"30",
          5548 => x"80",
          5549 => x"70",
          5550 => x"06",
          5551 => x"56",
          5552 => x"90",
          5553 => x"d4",
          5554 => x"98",
          5555 => x"78",
          5556 => x"3f",
          5557 => x"81",
          5558 => x"96",
          5559 => x"f9",
          5560 => x"02",
          5561 => x"05",
          5562 => x"ff",
          5563 => x"7a",
          5564 => x"fe",
          5565 => x"dc",
          5566 => x"38",
          5567 => x"88",
          5568 => x"2e",
          5569 => x"39",
          5570 => x"54",
          5571 => x"53",
          5572 => x"51",
          5573 => x"dc",
          5574 => x"83",
          5575 => x"76",
          5576 => x"0c",
          5577 => x"04",
          5578 => x"7f",
          5579 => x"8c",
          5580 => x"05",
          5581 => x"15",
          5582 => x"5c",
          5583 => x"5e",
          5584 => x"d2",
          5585 => x"89",
          5586 => x"d2",
          5587 => x"83",
          5588 => x"55",
          5589 => x"80",
          5590 => x"90",
          5591 => x"7b",
          5592 => x"38",
          5593 => x"74",
          5594 => x"7a",
          5595 => x"72",
          5596 => x"d2",
          5597 => x"88",
          5598 => x"39",
          5599 => x"51",
          5600 => x"3f",
          5601 => x"80",
          5602 => x"18",
          5603 => x"27",
          5604 => x"08",
          5605 => x"dc",
          5606 => x"c8",
          5607 => x"81",
          5608 => x"ff",
          5609 => x"84",
          5610 => x"39",
          5611 => x"72",
          5612 => x"38",
          5613 => x"81",
          5614 => x"ff",
          5615 => x"89",
          5616 => x"84",
          5617 => x"b8",
          5618 => x"55",
          5619 => x"81",
          5620 => x"80",
          5621 => x"88",
          5622 => x"a4",
          5623 => x"74",
          5624 => x"38",
          5625 => x"33",
          5626 => x"56",
          5627 => x"83",
          5628 => x"80",
          5629 => x"27",
          5630 => x"53",
          5631 => x"70",
          5632 => x"51",
          5633 => x"2e",
          5634 => x"80",
          5635 => x"38",
          5636 => x"39",
          5637 => x"81",
          5638 => x"15",
          5639 => x"81",
          5640 => x"ff",
          5641 => x"78",
          5642 => x"5c",
          5643 => x"de",
          5644 => x"cc",
          5645 => x"70",
          5646 => x"57",
          5647 => x"09",
          5648 => x"38",
          5649 => x"3f",
          5650 => x"08",
          5651 => x"98",
          5652 => x"32",
          5653 => x"9b",
          5654 => x"70",
          5655 => x"75",
          5656 => x"58",
          5657 => x"51",
          5658 => x"24",
          5659 => x"9b",
          5660 => x"06",
          5661 => x"53",
          5662 => x"1e",
          5663 => x"26",
          5664 => x"ff",
          5665 => x"dc",
          5666 => x"3d",
          5667 => x"3d",
          5668 => x"05",
          5669 => x"90",
          5670 => x"94",
          5671 => x"86",
          5672 => x"d9",
          5673 => x"fe",
          5674 => x"81",
          5675 => x"81",
          5676 => x"81",
          5677 => x"52",
          5678 => x"51",
          5679 => x"3f",
          5680 => x"85",
          5681 => x"ea",
          5682 => x"0d",
          5683 => x"0d",
          5684 => x"80",
          5685 => x"ff",
          5686 => x"51",
          5687 => x"3f",
          5688 => x"51",
          5689 => x"3f",
          5690 => x"f1",
          5691 => x"81",
          5692 => x"06",
          5693 => x"80",
          5694 => x"81",
          5695 => x"a2",
          5696 => x"e8",
          5697 => x"9a",
          5698 => x"fe",
          5699 => x"72",
          5700 => x"81",
          5701 => x"71",
          5702 => x"38",
          5703 => x"f1",
          5704 => x"d3",
          5705 => x"f2",
          5706 => x"51",
          5707 => x"3f",
          5708 => x"70",
          5709 => x"52",
          5710 => x"95",
          5711 => x"fe",
          5712 => x"81",
          5713 => x"fe",
          5714 => x"80",
          5715 => x"d2",
          5716 => x"2a",
          5717 => x"51",
          5718 => x"2e",
          5719 => x"51",
          5720 => x"3f",
          5721 => x"51",
          5722 => x"3f",
          5723 => x"f0",
          5724 => x"85",
          5725 => x"06",
          5726 => x"80",
          5727 => x"81",
          5728 => x"9e",
          5729 => x"b4",
          5730 => x"96",
          5731 => x"fe",
          5732 => x"72",
          5733 => x"81",
          5734 => x"71",
          5735 => x"38",
          5736 => x"ef",
          5737 => x"d4",
          5738 => x"f1",
          5739 => x"51",
          5740 => x"3f",
          5741 => x"70",
          5742 => x"52",
          5743 => x"95",
          5744 => x"fe",
          5745 => x"81",
          5746 => x"fe",
          5747 => x"80",
          5748 => x"ce",
          5749 => x"2a",
          5750 => x"51",
          5751 => x"2e",
          5752 => x"51",
          5753 => x"3f",
          5754 => x"51",
          5755 => x"3f",
          5756 => x"ef",
          5757 => x"fd",
          5758 => x"3d",
          5759 => x"3d",
          5760 => x"70",
          5761 => x"80",
          5762 => x"fe",
          5763 => x"81",
          5764 => x"54",
          5765 => x"81",
          5766 => x"b0",
          5767 => x"d0",
          5768 => x"dc",
          5769 => x"cc",
          5770 => x"81",
          5771 => x"07",
          5772 => x"71",
          5773 => x"54",
          5774 => x"d8",
          5775 => x"d8",
          5776 => x"81",
          5777 => x"06",
          5778 => x"f3",
          5779 => x"52",
          5780 => x"92",
          5781 => x"cc",
          5782 => x"8c",
          5783 => x"cc",
          5784 => x"fd",
          5785 => x"39",
          5786 => x"51",
          5787 => x"82",
          5788 => x"d8",
          5789 => x"d8",
          5790 => x"82",
          5791 => x"06",
          5792 => x"52",
          5793 => x"83",
          5794 => x"0b",
          5795 => x"0c",
          5796 => x"04",
          5797 => x"80",
          5798 => x"f3",
          5799 => x"5d",
          5800 => x"51",
          5801 => x"3f",
          5802 => x"08",
          5803 => x"59",
          5804 => x"09",
          5805 => x"38",
          5806 => x"52",
          5807 => x"52",
          5808 => x"b6",
          5809 => x"78",
          5810 => x"fc",
          5811 => x"cf",
          5812 => x"cc",
          5813 => x"88",
          5814 => x"c4",
          5815 => x"39",
          5816 => x"5d",
          5817 => x"51",
          5818 => x"3f",
          5819 => x"46",
          5820 => x"52",
          5821 => x"86",
          5822 => x"ff",
          5823 => x"f3",
          5824 => x"dc",
          5825 => x"2b",
          5826 => x"51",
          5827 => x"c2",
          5828 => x"38",
          5829 => x"24",
          5830 => x"bd",
          5831 => x"38",
          5832 => x"90",
          5833 => x"2e",
          5834 => x"78",
          5835 => x"da",
          5836 => x"39",
          5837 => x"2e",
          5838 => x"78",
          5839 => x"85",
          5840 => x"bf",
          5841 => x"38",
          5842 => x"78",
          5843 => x"89",
          5844 => x"80",
          5845 => x"38",
          5846 => x"2e",
          5847 => x"78",
          5848 => x"89",
          5849 => x"b4",
          5850 => x"83",
          5851 => x"38",
          5852 => x"24",
          5853 => x"81",
          5854 => x"fd",
          5855 => x"39",
          5856 => x"2e",
          5857 => x"8a",
          5858 => x"3d",
          5859 => x"53",
          5860 => x"51",
          5861 => x"3f",
          5862 => x"08",
          5863 => x"c4",
          5864 => x"fe",
          5865 => x"ff",
          5866 => x"ff",
          5867 => x"81",
          5868 => x"80",
          5869 => x"38",
          5870 => x"f8",
          5871 => x"84",
          5872 => x"82",
          5873 => x"dc",
          5874 => x"38",
          5875 => x"08",
          5876 => x"80",
          5877 => x"a8",
          5878 => x"5c",
          5879 => x"27",
          5880 => x"61",
          5881 => x"70",
          5882 => x"0c",
          5883 => x"f5",
          5884 => x"39",
          5885 => x"80",
          5886 => x"84",
          5887 => x"81",
          5888 => x"dc",
          5889 => x"2e",
          5890 => x"b4",
          5891 => x"11",
          5892 => x"05",
          5893 => x"c1",
          5894 => x"cc",
          5895 => x"fd",
          5896 => x"3d",
          5897 => x"53",
          5898 => x"51",
          5899 => x"3f",
          5900 => x"08",
          5901 => x"ac",
          5902 => x"90",
          5903 => x"c0",
          5904 => x"79",
          5905 => x"8c",
          5906 => x"79",
          5907 => x"5b",
          5908 => x"61",
          5909 => x"eb",
          5910 => x"ff",
          5911 => x"ff",
          5912 => x"ff",
          5913 => x"81",
          5914 => x"80",
          5915 => x"38",
          5916 => x"fc",
          5917 => x"84",
          5918 => x"80",
          5919 => x"dc",
          5920 => x"2e",
          5921 => x"b4",
          5922 => x"11",
          5923 => x"05",
          5924 => x"c5",
          5925 => x"cc",
          5926 => x"fc",
          5927 => x"d6",
          5928 => x"f8",
          5929 => x"5a",
          5930 => x"a8",
          5931 => x"33",
          5932 => x"5a",
          5933 => x"2e",
          5934 => x"55",
          5935 => x"33",
          5936 => x"81",
          5937 => x"fe",
          5938 => x"81",
          5939 => x"05",
          5940 => x"39",
          5941 => x"51",
          5942 => x"b4",
          5943 => x"11",
          5944 => x"05",
          5945 => x"f1",
          5946 => x"cc",
          5947 => x"38",
          5948 => x"33",
          5949 => x"2e",
          5950 => x"d8",
          5951 => x"80",
          5952 => x"d9",
          5953 => x"78",
          5954 => x"38",
          5955 => x"08",
          5956 => x"81",
          5957 => x"59",
          5958 => x"88",
          5959 => x"88",
          5960 => x"39",
          5961 => x"33",
          5962 => x"2e",
          5963 => x"d9",
          5964 => x"9a",
          5965 => x"be",
          5966 => x"80",
          5967 => x"81",
          5968 => x"44",
          5969 => x"d9",
          5970 => x"80",
          5971 => x"3d",
          5972 => x"53",
          5973 => x"51",
          5974 => x"3f",
          5975 => x"08",
          5976 => x"81",
          5977 => x"59",
          5978 => x"89",
          5979 => x"fc",
          5980 => x"cc",
          5981 => x"c1",
          5982 => x"80",
          5983 => x"81",
          5984 => x"43",
          5985 => x"d9",
          5986 => x"78",
          5987 => x"38",
          5988 => x"08",
          5989 => x"81",
          5990 => x"59",
          5991 => x"88",
          5992 => x"94",
          5993 => x"39",
          5994 => x"33",
          5995 => x"2e",
          5996 => x"d9",
          5997 => x"88",
          5998 => x"a8",
          5999 => x"43",
          6000 => x"f8",
          6001 => x"84",
          6002 => x"fe",
          6003 => x"dc",
          6004 => x"2e",
          6005 => x"62",
          6006 => x"88",
          6007 => x"81",
          6008 => x"32",
          6009 => x"72",
          6010 => x"70",
          6011 => x"51",
          6012 => x"80",
          6013 => x"7a",
          6014 => x"38",
          6015 => x"d6",
          6016 => x"f5",
          6017 => x"55",
          6018 => x"53",
          6019 => x"51",
          6020 => x"81",
          6021 => x"fe",
          6022 => x"f9",
          6023 => x"3d",
          6024 => x"53",
          6025 => x"51",
          6026 => x"3f",
          6027 => x"08",
          6028 => x"b0",
          6029 => x"fe",
          6030 => x"ff",
          6031 => x"fe",
          6032 => x"81",
          6033 => x"80",
          6034 => x"63",
          6035 => x"cb",
          6036 => x"34",
          6037 => x"44",
          6038 => x"fc",
          6039 => x"84",
          6040 => x"fc",
          6041 => x"dc",
          6042 => x"38",
          6043 => x"63",
          6044 => x"52",
          6045 => x"51",
          6046 => x"3f",
          6047 => x"79",
          6048 => x"ba",
          6049 => x"79",
          6050 => x"ae",
          6051 => x"38",
          6052 => x"a0",
          6053 => x"fe",
          6054 => x"ff",
          6055 => x"fe",
          6056 => x"81",
          6057 => x"80",
          6058 => x"63",
          6059 => x"cb",
          6060 => x"34",
          6061 => x"44",
          6062 => x"81",
          6063 => x"fe",
          6064 => x"ff",
          6065 => x"3d",
          6066 => x"53",
          6067 => x"51",
          6068 => x"3f",
          6069 => x"08",
          6070 => x"88",
          6071 => x"fe",
          6072 => x"ff",
          6073 => x"fe",
          6074 => x"81",
          6075 => x"80",
          6076 => x"60",
          6077 => x"05",
          6078 => x"82",
          6079 => x"78",
          6080 => x"fe",
          6081 => x"ff",
          6082 => x"fe",
          6083 => x"81",
          6084 => x"df",
          6085 => x"39",
          6086 => x"54",
          6087 => x"f8",
          6088 => x"c0",
          6089 => x"52",
          6090 => x"fa",
          6091 => x"45",
          6092 => x"78",
          6093 => x"ac",
          6094 => x"26",
          6095 => x"82",
          6096 => x"39",
          6097 => x"f0",
          6098 => x"84",
          6099 => x"fc",
          6100 => x"dc",
          6101 => x"2e",
          6102 => x"59",
          6103 => x"22",
          6104 => x"05",
          6105 => x"41",
          6106 => x"81",
          6107 => x"fe",
          6108 => x"ff",
          6109 => x"3d",
          6110 => x"53",
          6111 => x"51",
          6112 => x"3f",
          6113 => x"08",
          6114 => x"d8",
          6115 => x"fe",
          6116 => x"ff",
          6117 => x"fe",
          6118 => x"81",
          6119 => x"80",
          6120 => x"60",
          6121 => x"59",
          6122 => x"41",
          6123 => x"f0",
          6124 => x"84",
          6125 => x"fc",
          6126 => x"dc",
          6127 => x"38",
          6128 => x"60",
          6129 => x"52",
          6130 => x"51",
          6131 => x"3f",
          6132 => x"79",
          6133 => x"e6",
          6134 => x"79",
          6135 => x"ae",
          6136 => x"38",
          6137 => x"9c",
          6138 => x"fe",
          6139 => x"ff",
          6140 => x"fe",
          6141 => x"81",
          6142 => x"80",
          6143 => x"60",
          6144 => x"59",
          6145 => x"41",
          6146 => x"81",
          6147 => x"fe",
          6148 => x"ff",
          6149 => x"3d",
          6150 => x"53",
          6151 => x"51",
          6152 => x"3f",
          6153 => x"08",
          6154 => x"b8",
          6155 => x"81",
          6156 => x"fe",
          6157 => x"63",
          6158 => x"b4",
          6159 => x"11",
          6160 => x"05",
          6161 => x"91",
          6162 => x"cc",
          6163 => x"f5",
          6164 => x"52",
          6165 => x"51",
          6166 => x"3f",
          6167 => x"2d",
          6168 => x"08",
          6169 => x"fc",
          6170 => x"cc",
          6171 => x"d7",
          6172 => x"f6",
          6173 => x"ec",
          6174 => x"e4",
          6175 => x"80",
          6176 => x"d6",
          6177 => x"39",
          6178 => x"51",
          6179 => x"3f",
          6180 => x"a5",
          6181 => x"9a",
          6182 => x"39",
          6183 => x"51",
          6184 => x"2e",
          6185 => x"7d",
          6186 => x"78",
          6187 => x"d8",
          6188 => x"ff",
          6189 => x"fe",
          6190 => x"81",
          6191 => x"5c",
          6192 => x"82",
          6193 => x"7a",
          6194 => x"38",
          6195 => x"8c",
          6196 => x"39",
          6197 => x"b0",
          6198 => x"39",
          6199 => x"56",
          6200 => x"d8",
          6201 => x"53",
          6202 => x"52",
          6203 => x"b0",
          6204 => x"f6",
          6205 => x"39",
          6206 => x"52",
          6207 => x"b0",
          6208 => x"f5",
          6209 => x"39",
          6210 => x"d8",
          6211 => x"53",
          6212 => x"52",
          6213 => x"b0",
          6214 => x"f5",
          6215 => x"39",
          6216 => x"53",
          6217 => x"52",
          6218 => x"b0",
          6219 => x"f5",
          6220 => x"d8",
          6221 => x"dd",
          6222 => x"56",
          6223 => x"46",
          6224 => x"80",
          6225 => x"80",
          6226 => x"80",
          6227 => x"ff",
          6228 => x"eb",
          6229 => x"dc",
          6230 => x"dc",
          6231 => x"70",
          6232 => x"07",
          6233 => x"5b",
          6234 => x"5a",
          6235 => x"83",
          6236 => x"78",
          6237 => x"78",
          6238 => x"38",
          6239 => x"81",
          6240 => x"59",
          6241 => x"38",
          6242 => x"7d",
          6243 => x"59",
          6244 => x"7e",
          6245 => x"81",
          6246 => x"38",
          6247 => x"51",
          6248 => x"3f",
          6249 => x"fc",
          6250 => x"0b",
          6251 => x"34",
          6252 => x"8c",
          6253 => x"55",
          6254 => x"52",
          6255 => x"d3",
          6256 => x"dc",
          6257 => x"2b",
          6258 => x"53",
          6259 => x"52",
          6260 => x"d3",
          6261 => x"81",
          6262 => x"07",
          6263 => x"c0",
          6264 => x"08",
          6265 => x"84",
          6266 => x"51",
          6267 => x"3f",
          6268 => x"08",
          6269 => x"08",
          6270 => x"84",
          6271 => x"51",
          6272 => x"3f",
          6273 => x"cc",
          6274 => x"0c",
          6275 => x"0b",
          6276 => x"84",
          6277 => x"83",
          6278 => x"94",
          6279 => x"bc",
          6280 => x"dc",
          6281 => x"0b",
          6282 => x"0c",
          6283 => x"3f",
          6284 => x"3f",
          6285 => x"51",
          6286 => x"3f",
          6287 => x"51",
          6288 => x"3f",
          6289 => x"51",
          6290 => x"3f",
          6291 => x"be",
          6292 => x"3f",
          6293 => x"00",
          6294 => x"ff",
          6295 => x"ff",
          6296 => x"ff",
          6297 => x"00",
          6298 => x"63",
          6299 => x"69",
          6300 => x"6f",
          6301 => x"75",
          6302 => x"7b",
          6303 => x"d4",
          6304 => x"58",
          6305 => x"5f",
          6306 => x"66",
          6307 => x"6d",
          6308 => x"74",
          6309 => x"7b",
          6310 => x"82",
          6311 => x"89",
          6312 => x"90",
          6313 => x"97",
          6314 => x"9e",
          6315 => x"a4",
          6316 => x"aa",
          6317 => x"b0",
          6318 => x"b6",
          6319 => x"bc",
          6320 => x"c2",
          6321 => x"c8",
          6322 => x"ce",
          6323 => x"25",
          6324 => x"64",
          6325 => x"3a",
          6326 => x"25",
          6327 => x"64",
          6328 => x"00",
          6329 => x"20",
          6330 => x"66",
          6331 => x"72",
          6332 => x"6f",
          6333 => x"00",
          6334 => x"72",
          6335 => x"53",
          6336 => x"63",
          6337 => x"69",
          6338 => x"00",
          6339 => x"65",
          6340 => x"65",
          6341 => x"6d",
          6342 => x"6d",
          6343 => x"65",
          6344 => x"00",
          6345 => x"20",
          6346 => x"53",
          6347 => x"4d",
          6348 => x"25",
          6349 => x"3a",
          6350 => x"58",
          6351 => x"00",
          6352 => x"20",
          6353 => x"41",
          6354 => x"20",
          6355 => x"25",
          6356 => x"3a",
          6357 => x"58",
          6358 => x"00",
          6359 => x"20",
          6360 => x"4e",
          6361 => x"41",
          6362 => x"25",
          6363 => x"3a",
          6364 => x"58",
          6365 => x"00",
          6366 => x"20",
          6367 => x"4d",
          6368 => x"20",
          6369 => x"25",
          6370 => x"3a",
          6371 => x"58",
          6372 => x"00",
          6373 => x"20",
          6374 => x"20",
          6375 => x"20",
          6376 => x"25",
          6377 => x"3a",
          6378 => x"58",
          6379 => x"00",
          6380 => x"20",
          6381 => x"43",
          6382 => x"20",
          6383 => x"44",
          6384 => x"63",
          6385 => x"3d",
          6386 => x"64",
          6387 => x"00",
          6388 => x"20",
          6389 => x"45",
          6390 => x"20",
          6391 => x"54",
          6392 => x"72",
          6393 => x"3d",
          6394 => x"64",
          6395 => x"00",
          6396 => x"20",
          6397 => x"52",
          6398 => x"52",
          6399 => x"43",
          6400 => x"6e",
          6401 => x"3d",
          6402 => x"64",
          6403 => x"00",
          6404 => x"20",
          6405 => x"48",
          6406 => x"45",
          6407 => x"53",
          6408 => x"00",
          6409 => x"20",
          6410 => x"49",
          6411 => x"00",
          6412 => x"20",
          6413 => x"54",
          6414 => x"00",
          6415 => x"20",
          6416 => x"0a",
          6417 => x"00",
          6418 => x"20",
          6419 => x"0a",
          6420 => x"00",
          6421 => x"72",
          6422 => x"65",
          6423 => x"00",
          6424 => x"20",
          6425 => x"20",
          6426 => x"65",
          6427 => x"65",
          6428 => x"72",
          6429 => x"64",
          6430 => x"73",
          6431 => x"25",
          6432 => x"0a",
          6433 => x"00",
          6434 => x"20",
          6435 => x"20",
          6436 => x"6f",
          6437 => x"53",
          6438 => x"74",
          6439 => x"64",
          6440 => x"73",
          6441 => x"25",
          6442 => x"0a",
          6443 => x"00",
          6444 => x"20",
          6445 => x"63",
          6446 => x"74",
          6447 => x"20",
          6448 => x"72",
          6449 => x"20",
          6450 => x"20",
          6451 => x"25",
          6452 => x"0a",
          6453 => x"00",
          6454 => x"63",
          6455 => x"00",
          6456 => x"20",
          6457 => x"20",
          6458 => x"20",
          6459 => x"20",
          6460 => x"20",
          6461 => x"20",
          6462 => x"20",
          6463 => x"25",
          6464 => x"0a",
          6465 => x"00",
          6466 => x"20",
          6467 => x"74",
          6468 => x"43",
          6469 => x"6b",
          6470 => x"65",
          6471 => x"20",
          6472 => x"20",
          6473 => x"25",
          6474 => x"30",
          6475 => x"48",
          6476 => x"00",
          6477 => x"20",
          6478 => x"41",
          6479 => x"6c",
          6480 => x"20",
          6481 => x"71",
          6482 => x"20",
          6483 => x"20",
          6484 => x"25",
          6485 => x"30",
          6486 => x"48",
          6487 => x"00",
          6488 => x"20",
          6489 => x"68",
          6490 => x"65",
          6491 => x"52",
          6492 => x"43",
          6493 => x"6b",
          6494 => x"65",
          6495 => x"25",
          6496 => x"30",
          6497 => x"48",
          6498 => x"00",
          6499 => x"6c",
          6500 => x"00",
          6501 => x"69",
          6502 => x"00",
          6503 => x"78",
          6504 => x"00",
          6505 => x"00",
          6506 => x"6d",
          6507 => x"00",
          6508 => x"6e",
          6509 => x"00",
          6510 => x"00",
          6511 => x"2c",
          6512 => x"3d",
          6513 => x"5d",
          6514 => x"00",
          6515 => x"00",
          6516 => x"33",
          6517 => x"00",
          6518 => x"4d",
          6519 => x"53",
          6520 => x"00",
          6521 => x"4e",
          6522 => x"20",
          6523 => x"46",
          6524 => x"32",
          6525 => x"00",
          6526 => x"4e",
          6527 => x"20",
          6528 => x"46",
          6529 => x"20",
          6530 => x"00",
          6531 => x"b8",
          6532 => x"00",
          6533 => x"00",
          6534 => x"00",
          6535 => x"41",
          6536 => x"80",
          6537 => x"49",
          6538 => x"8f",
          6539 => x"4f",
          6540 => x"55",
          6541 => x"9b",
          6542 => x"9f",
          6543 => x"55",
          6544 => x"a7",
          6545 => x"ab",
          6546 => x"af",
          6547 => x"b3",
          6548 => x"b7",
          6549 => x"bb",
          6550 => x"bf",
          6551 => x"c3",
          6552 => x"c7",
          6553 => x"cb",
          6554 => x"cf",
          6555 => x"d3",
          6556 => x"d7",
          6557 => x"db",
          6558 => x"df",
          6559 => x"e3",
          6560 => x"e7",
          6561 => x"eb",
          6562 => x"ef",
          6563 => x"f3",
          6564 => x"f7",
          6565 => x"fb",
          6566 => x"ff",
          6567 => x"3b",
          6568 => x"2f",
          6569 => x"3a",
          6570 => x"7c",
          6571 => x"00",
          6572 => x"04",
          6573 => x"40",
          6574 => x"00",
          6575 => x"00",
          6576 => x"02",
          6577 => x"08",
          6578 => x"20",
          6579 => x"00",
          6580 => x"69",
          6581 => x"00",
          6582 => x"63",
          6583 => x"00",
          6584 => x"69",
          6585 => x"00",
          6586 => x"61",
          6587 => x"00",
          6588 => x"65",
          6589 => x"00",
          6590 => x"65",
          6591 => x"00",
          6592 => x"70",
          6593 => x"00",
          6594 => x"66",
          6595 => x"00",
          6596 => x"6d",
          6597 => x"00",
          6598 => x"00",
          6599 => x"00",
          6600 => x"00",
          6601 => x"00",
          6602 => x"00",
          6603 => x"00",
          6604 => x"00",
          6605 => x"6c",
          6606 => x"00",
          6607 => x"00",
          6608 => x"74",
          6609 => x"00",
          6610 => x"65",
          6611 => x"00",
          6612 => x"6f",
          6613 => x"00",
          6614 => x"74",
          6615 => x"00",
          6616 => x"73",
          6617 => x"00",
          6618 => x"6b",
          6619 => x"72",
          6620 => x"00",
          6621 => x"65",
          6622 => x"6c",
          6623 => x"72",
          6624 => x"0a",
          6625 => x"00",
          6626 => x"6b",
          6627 => x"74",
          6628 => x"61",
          6629 => x"0a",
          6630 => x"00",
          6631 => x"66",
          6632 => x"20",
          6633 => x"6e",
          6634 => x"00",
          6635 => x"70",
          6636 => x"20",
          6637 => x"6e",
          6638 => x"00",
          6639 => x"61",
          6640 => x"20",
          6641 => x"65",
          6642 => x"65",
          6643 => x"00",
          6644 => x"65",
          6645 => x"64",
          6646 => x"65",
          6647 => x"00",
          6648 => x"65",
          6649 => x"72",
          6650 => x"79",
          6651 => x"69",
          6652 => x"2e",
          6653 => x"00",
          6654 => x"65",
          6655 => x"6e",
          6656 => x"20",
          6657 => x"61",
          6658 => x"2e",
          6659 => x"00",
          6660 => x"69",
          6661 => x"72",
          6662 => x"20",
          6663 => x"74",
          6664 => x"65",
          6665 => x"00",
          6666 => x"76",
          6667 => x"75",
          6668 => x"72",
          6669 => x"20",
          6670 => x"61",
          6671 => x"2e",
          6672 => x"00",
          6673 => x"6b",
          6674 => x"74",
          6675 => x"61",
          6676 => x"64",
          6677 => x"00",
          6678 => x"63",
          6679 => x"61",
          6680 => x"6c",
          6681 => x"69",
          6682 => x"79",
          6683 => x"6d",
          6684 => x"75",
          6685 => x"6f",
          6686 => x"69",
          6687 => x"0a",
          6688 => x"00",
          6689 => x"6d",
          6690 => x"61",
          6691 => x"74",
          6692 => x"0a",
          6693 => x"00",
          6694 => x"65",
          6695 => x"2c",
          6696 => x"65",
          6697 => x"69",
          6698 => x"63",
          6699 => x"65",
          6700 => x"64",
          6701 => x"00",
          6702 => x"65",
          6703 => x"20",
          6704 => x"6b",
          6705 => x"0a",
          6706 => x"00",
          6707 => x"75",
          6708 => x"63",
          6709 => x"74",
          6710 => x"6d",
          6711 => x"2e",
          6712 => x"00",
          6713 => x"20",
          6714 => x"79",
          6715 => x"65",
          6716 => x"69",
          6717 => x"2e",
          6718 => x"00",
          6719 => x"61",
          6720 => x"65",
          6721 => x"69",
          6722 => x"72",
          6723 => x"74",
          6724 => x"00",
          6725 => x"63",
          6726 => x"2e",
          6727 => x"00",
          6728 => x"6e",
          6729 => x"20",
          6730 => x"6f",
          6731 => x"00",
          6732 => x"75",
          6733 => x"74",
          6734 => x"25",
          6735 => x"74",
          6736 => x"75",
          6737 => x"74",
          6738 => x"73",
          6739 => x"0a",
          6740 => x"00",
          6741 => x"64",
          6742 => x"00",
          6743 => x"58",
          6744 => x"00",
          6745 => x"00",
          6746 => x"58",
          6747 => x"00",
          6748 => x"20",
          6749 => x"20",
          6750 => x"00",
          6751 => x"58",
          6752 => x"00",
          6753 => x"00",
          6754 => x"00",
          6755 => x"00",
          6756 => x"00",
          6757 => x"20",
          6758 => x"28",
          6759 => x"00",
          6760 => x"30",
          6761 => x"30",
          6762 => x"00",
          6763 => x"30",
          6764 => x"00",
          6765 => x"55",
          6766 => x"65",
          6767 => x"30",
          6768 => x"20",
          6769 => x"25",
          6770 => x"2a",
          6771 => x"00",
          6772 => x"20",
          6773 => x"65",
          6774 => x"70",
          6775 => x"61",
          6776 => x"65",
          6777 => x"00",
          6778 => x"65",
          6779 => x"6e",
          6780 => x"72",
          6781 => x"0a",
          6782 => x"00",
          6783 => x"20",
          6784 => x"65",
          6785 => x"70",
          6786 => x"00",
          6787 => x"54",
          6788 => x"44",
          6789 => x"74",
          6790 => x"75",
          6791 => x"00",
          6792 => x"54",
          6793 => x"52",
          6794 => x"74",
          6795 => x"75",
          6796 => x"00",
          6797 => x"54",
          6798 => x"58",
          6799 => x"74",
          6800 => x"75",
          6801 => x"00",
          6802 => x"54",
          6803 => x"58",
          6804 => x"74",
          6805 => x"75",
          6806 => x"00",
          6807 => x"54",
          6808 => x"58",
          6809 => x"74",
          6810 => x"75",
          6811 => x"00",
          6812 => x"54",
          6813 => x"58",
          6814 => x"74",
          6815 => x"75",
          6816 => x"00",
          6817 => x"74",
          6818 => x"20",
          6819 => x"74",
          6820 => x"72",
          6821 => x"0a",
          6822 => x"00",
          6823 => x"62",
          6824 => x"67",
          6825 => x"6d",
          6826 => x"2e",
          6827 => x"00",
          6828 => x"6f",
          6829 => x"63",
          6830 => x"74",
          6831 => x"00",
          6832 => x"00",
          6833 => x"6c",
          6834 => x"74",
          6835 => x"6e",
          6836 => x"61",
          6837 => x"65",
          6838 => x"20",
          6839 => x"64",
          6840 => x"20",
          6841 => x"61",
          6842 => x"69",
          6843 => x"20",
          6844 => x"75",
          6845 => x"79",
          6846 => x"00",
          6847 => x"00",
          6848 => x"61",
          6849 => x"67",
          6850 => x"2e",
          6851 => x"00",
          6852 => x"79",
          6853 => x"2e",
          6854 => x"00",
          6855 => x"70",
          6856 => x"6e",
          6857 => x"2e",
          6858 => x"00",
          6859 => x"6c",
          6860 => x"30",
          6861 => x"2d",
          6862 => x"38",
          6863 => x"25",
          6864 => x"29",
          6865 => x"00",
          6866 => x"70",
          6867 => x"6d",
          6868 => x"0a",
          6869 => x"00",
          6870 => x"6d",
          6871 => x"74",
          6872 => x"00",
          6873 => x"58",
          6874 => x"32",
          6875 => x"00",
          6876 => x"0a",
          6877 => x"00",
          6878 => x"58",
          6879 => x"34",
          6880 => x"00",
          6881 => x"58",
          6882 => x"38",
          6883 => x"00",
          6884 => x"63",
          6885 => x"6e",
          6886 => x"6f",
          6887 => x"40",
          6888 => x"38",
          6889 => x"2e",
          6890 => x"00",
          6891 => x"6c",
          6892 => x"20",
          6893 => x"65",
          6894 => x"25",
          6895 => x"20",
          6896 => x"0a",
          6897 => x"00",
          6898 => x"6c",
          6899 => x"74",
          6900 => x"65",
          6901 => x"6f",
          6902 => x"28",
          6903 => x"2e",
          6904 => x"00",
          6905 => x"74",
          6906 => x"69",
          6907 => x"61",
          6908 => x"69",
          6909 => x"69",
          6910 => x"2e",
          6911 => x"00",
          6912 => x"64",
          6913 => x"62",
          6914 => x"69",
          6915 => x"2e",
          6916 => x"00",
          6917 => x"00",
          6918 => x"00",
          6919 => x"5c",
          6920 => x"25",
          6921 => x"73",
          6922 => x"00",
          6923 => x"5c",
          6924 => x"25",
          6925 => x"00",
          6926 => x"5c",
          6927 => x"00",
          6928 => x"20",
          6929 => x"6d",
          6930 => x"2e",
          6931 => x"00",
          6932 => x"6e",
          6933 => x"2e",
          6934 => x"00",
          6935 => x"62",
          6936 => x"67",
          6937 => x"74",
          6938 => x"75",
          6939 => x"2e",
          6940 => x"00",
          6941 => x"00",
          6942 => x"00",
          6943 => x"ff",
          6944 => x"00",
          6945 => x"ff",
          6946 => x"00",
          6947 => x"ff",
          6948 => x"00",
          6949 => x"00",
          6950 => x"00",
          6951 => x"ff",
          6952 => x"00",
          6953 => x"00",
          6954 => x"00",
          6955 => x"00",
          6956 => x"00",
          6957 => x"00",
          6958 => x"00",
          6959 => x"00",
          6960 => x"01",
          6961 => x"01",
          6962 => x"01",
          6963 => x"00",
          6964 => x"00",
          6965 => x"00",
          6966 => x"00",
          6967 => x"d0",
          6968 => x"00",
          6969 => x"00",
          6970 => x"00",
          6971 => x"d8",
          6972 => x"00",
          6973 => x"00",
          6974 => x"00",
          6975 => x"e0",
          6976 => x"00",
          6977 => x"00",
          6978 => x"00",
          6979 => x"e8",
          6980 => x"00",
          6981 => x"00",
          6982 => x"00",
          6983 => x"f0",
          6984 => x"00",
          6985 => x"00",
          6986 => x"00",
          6987 => x"f8",
          6988 => x"00",
          6989 => x"00",
          6990 => x"00",
          6991 => x"00",
          6992 => x"00",
          6993 => x"00",
          6994 => x"00",
          6995 => x"08",
          6996 => x"00",
          6997 => x"00",
          6998 => x"00",
          6999 => x"10",
          7000 => x"00",
          7001 => x"00",
          7002 => x"00",
          7003 => x"18",
          7004 => x"00",
          7005 => x"00",
          7006 => x"00",
          7007 => x"1c",
          7008 => x"00",
          7009 => x"00",
          7010 => x"00",
          7011 => x"20",
          7012 => x"00",
          7013 => x"00",
          7014 => x"00",
          7015 => x"24",
          7016 => x"00",
          7017 => x"00",
          7018 => x"00",
          7019 => x"28",
          7020 => x"00",
          7021 => x"00",
          7022 => x"00",
          7023 => x"2c",
          7024 => x"00",
          7025 => x"00",
          7026 => x"00",
          7027 => x"30",
          7028 => x"00",
          7029 => x"00",
          7030 => x"00",
          7031 => x"34",
          7032 => x"00",
          7033 => x"00",
          7034 => x"00",
          7035 => x"3c",
          7036 => x"00",
          7037 => x"00",
          7038 => x"00",
          7039 => x"40",
          7040 => x"00",
          7041 => x"00",
          7042 => x"00",
          7043 => x"48",
          7044 => x"00",
          7045 => x"00",
          7046 => x"00",
          7047 => x"50",
          7048 => x"00",
          7049 => x"00",
          7050 => x"00",
          7051 => x"58",
          7052 => x"00",
          7053 => x"00",
          7054 => x"00",
          7055 => x"60",
          7056 => x"00",
          7057 => x"00",
          7058 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"96",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"81",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"08",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a3",
           270 => x"0b",
           271 => x"0b",
           272 => x"c1",
           273 => x"0b",
           274 => x"0b",
           275 => x"df",
           276 => x"0b",
           277 => x"0b",
           278 => x"fd",
           279 => x"0b",
           280 => x"0b",
           281 => x"9b",
           282 => x"0b",
           283 => x"0b",
           284 => x"b9",
           285 => x"0b",
           286 => x"0b",
           287 => x"d7",
           288 => x"0b",
           289 => x"0b",
           290 => x"f5",
           291 => x"0b",
           292 => x"0b",
           293 => x"94",
           294 => x"0b",
           295 => x"0b",
           296 => x"b4",
           297 => x"0b",
           298 => x"0b",
           299 => x"d4",
           300 => x"0b",
           301 => x"0b",
           302 => x"f4",
           303 => x"0b",
           304 => x"0b",
           305 => x"94",
           306 => x"0b",
           307 => x"0b",
           308 => x"b4",
           309 => x"0b",
           310 => x"0b",
           311 => x"d4",
           312 => x"0b",
           313 => x"0b",
           314 => x"f4",
           315 => x"0b",
           316 => x"0b",
           317 => x"94",
           318 => x"0b",
           319 => x"0b",
           320 => x"b4",
           321 => x"0b",
           322 => x"0b",
           323 => x"d4",
           324 => x"0b",
           325 => x"0b",
           326 => x"f4",
           327 => x"0b",
           328 => x"0b",
           329 => x"94",
           330 => x"0b",
           331 => x"0b",
           332 => x"b3",
           333 => x"0b",
           334 => x"0b",
           335 => x"d2",
           336 => x"0b",
           337 => x"0b",
           338 => x"f0",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"00",
           386 => x"00",
           387 => x"00",
           388 => x"00",
           389 => x"00",
           390 => x"00",
           391 => x"00",
           392 => x"00",
           393 => x"00",
           394 => x"00",
           395 => x"00",
           396 => x"00",
           397 => x"00",
           398 => x"00",
           399 => x"00",
           400 => x"00",
           401 => x"00",
           402 => x"00",
           403 => x"00",
           404 => x"00",
           405 => x"00",
           406 => x"00",
           407 => x"00",
           408 => x"00",
           409 => x"00",
           410 => x"00",
           411 => x"00",
           412 => x"00",
           413 => x"00",
           414 => x"00",
           415 => x"00",
           416 => x"00",
           417 => x"00",
           418 => x"00",
           419 => x"00",
           420 => x"00",
           421 => x"00",
           422 => x"00",
           423 => x"00",
           424 => x"00",
           425 => x"00",
           426 => x"00",
           427 => x"00",
           428 => x"00",
           429 => x"00",
           430 => x"00",
           431 => x"00",
           432 => x"00",
           433 => x"00",
           434 => x"00",
           435 => x"00",
           436 => x"00",
           437 => x"00",
           438 => x"00",
           439 => x"00",
           440 => x"00",
           441 => x"00",
           442 => x"00",
           443 => x"00",
           444 => x"00",
           445 => x"00",
           446 => x"00",
           447 => x"00",
           448 => x"00",
           449 => x"00",
           450 => x"00",
           451 => x"00",
           452 => x"00",
           453 => x"00",
           454 => x"00",
           455 => x"00",
           456 => x"00",
           457 => x"00",
           458 => x"00",
           459 => x"00",
           460 => x"00",
           461 => x"00",
           462 => x"00",
           463 => x"00",
           464 => x"00",
           465 => x"00",
           466 => x"00",
           467 => x"00",
           468 => x"00",
           469 => x"00",
           470 => x"00",
           471 => x"00",
           472 => x"00",
           473 => x"00",
           474 => x"00",
           475 => x"00",
           476 => x"00",
           477 => x"00",
           478 => x"00",
           479 => x"00",
           480 => x"00",
           481 => x"00",
           482 => x"00",
           483 => x"00",
           484 => x"00",
           485 => x"00",
           486 => x"00",
           487 => x"00",
           488 => x"00",
           489 => x"00",
           490 => x"00",
           491 => x"00",
           492 => x"00",
           493 => x"00",
           494 => x"00",
           495 => x"00",
           496 => x"00",
           497 => x"00",
           498 => x"00",
           499 => x"00",
           500 => x"00",
           501 => x"00",
           502 => x"00",
           503 => x"00",
           504 => x"00",
           505 => x"00",
           506 => x"00",
           507 => x"00",
           508 => x"00",
           509 => x"00",
           510 => x"00",
           511 => x"00",
           512 => x"90",
           513 => x"dc",
           514 => x"b0",
           515 => x"d8",
           516 => x"90",
           517 => x"d8",
           518 => x"2d",
           519 => x"08",
           520 => x"04",
           521 => x"0c",
           522 => x"81",
           523 => x"83",
           524 => x"81",
           525 => x"b2",
           526 => x"dc",
           527 => x"80",
           528 => x"dc",
           529 => x"be",
           530 => x"d8",
           531 => x"90",
           532 => x"d8",
           533 => x"2d",
           534 => x"08",
           535 => x"04",
           536 => x"0c",
           537 => x"81",
           538 => x"83",
           539 => x"81",
           540 => x"b9",
           541 => x"dc",
           542 => x"80",
           543 => x"dc",
           544 => x"cb",
           545 => x"d8",
           546 => x"90",
           547 => x"d8",
           548 => x"2d",
           549 => x"08",
           550 => x"04",
           551 => x"0c",
           552 => x"81",
           553 => x"83",
           554 => x"81",
           555 => x"b8",
           556 => x"dc",
           557 => x"80",
           558 => x"dc",
           559 => x"bd",
           560 => x"d8",
           561 => x"90",
           562 => x"d8",
           563 => x"2d",
           564 => x"08",
           565 => x"04",
           566 => x"0c",
           567 => x"81",
           568 => x"83",
           569 => x"81",
           570 => x"a0",
           571 => x"dc",
           572 => x"80",
           573 => x"dc",
           574 => x"92",
           575 => x"d8",
           576 => x"90",
           577 => x"d8",
           578 => x"80",
           579 => x"d8",
           580 => x"90",
           581 => x"d8",
           582 => x"f1",
           583 => x"d8",
           584 => x"90",
           585 => x"d8",
           586 => x"e5",
           587 => x"d8",
           588 => x"90",
           589 => x"d8",
           590 => x"e2",
           591 => x"d8",
           592 => x"90",
           593 => x"d8",
           594 => x"80",
           595 => x"d8",
           596 => x"90",
           597 => x"d8",
           598 => x"e0",
           599 => x"d8",
           600 => x"90",
           601 => x"d8",
           602 => x"d3",
           603 => x"d8",
           604 => x"90",
           605 => x"d8",
           606 => x"9f",
           607 => x"d8",
           608 => x"90",
           609 => x"d8",
           610 => x"be",
           611 => x"d8",
           612 => x"90",
           613 => x"d8",
           614 => x"dd",
           615 => x"d8",
           616 => x"90",
           617 => x"d8",
           618 => x"c7",
           619 => x"d8",
           620 => x"90",
           621 => x"d8",
           622 => x"ad",
           623 => x"d8",
           624 => x"90",
           625 => x"d8",
           626 => x"9b",
           627 => x"d8",
           628 => x"90",
           629 => x"d8",
           630 => x"e1",
           631 => x"d8",
           632 => x"90",
           633 => x"d8",
           634 => x"9b",
           635 => x"d8",
           636 => x"90",
           637 => x"d8",
           638 => x"9c",
           639 => x"d8",
           640 => x"90",
           641 => x"d8",
           642 => x"d1",
           643 => x"d8",
           644 => x"90",
           645 => x"d8",
           646 => x"aa",
           647 => x"d8",
           648 => x"90",
           649 => x"d8",
           650 => x"d5",
           651 => x"d8",
           652 => x"90",
           653 => x"d8",
           654 => x"b8",
           655 => x"d8",
           656 => x"90",
           657 => x"d8",
           658 => x"8d",
           659 => x"d8",
           660 => x"90",
           661 => x"d8",
           662 => x"97",
           663 => x"d8",
           664 => x"90",
           665 => x"d8",
           666 => x"d9",
           667 => x"d8",
           668 => x"90",
           669 => x"d8",
           670 => x"9f",
           671 => x"d8",
           672 => x"90",
           673 => x"d8",
           674 => x"c5",
           675 => x"d8",
           676 => x"90",
           677 => x"d8",
           678 => x"2d",
           679 => x"08",
           680 => x"04",
           681 => x"0c",
           682 => x"2d",
           683 => x"08",
           684 => x"04",
           685 => x"0c",
           686 => x"2d",
           687 => x"08",
           688 => x"04",
           689 => x"0c",
           690 => x"81",
           691 => x"83",
           692 => x"81",
           693 => x"a0",
           694 => x"dc",
           695 => x"80",
           696 => x"dc",
           697 => x"a2",
           698 => x"d8",
           699 => x"90",
           700 => x"d8",
           701 => x"c2",
           702 => x"d8",
           703 => x"90",
           704 => x"10",
           705 => x"10",
           706 => x"10",
           707 => x"10",
           708 => x"10",
           709 => x"10",
           710 => x"10",
           711 => x"10",
           712 => x"51",
           713 => x"73",
           714 => x"73",
           715 => x"81",
           716 => x"10",
           717 => x"07",
           718 => x"0c",
           719 => x"72",
           720 => x"81",
           721 => x"09",
           722 => x"71",
           723 => x"0a",
           724 => x"72",
           725 => x"51",
           726 => x"81",
           727 => x"81",
           728 => x"8e",
           729 => x"70",
           730 => x"0c",
           731 => x"96",
           732 => x"81",
           733 => x"a7",
           734 => x"dc",
           735 => x"81",
           736 => x"fd",
           737 => x"53",
           738 => x"08",
           739 => x"52",
           740 => x"08",
           741 => x"51",
           742 => x"81",
           743 => x"70",
           744 => x"0c",
           745 => x"0d",
           746 => x"0c",
           747 => x"d8",
           748 => x"dc",
           749 => x"3d",
           750 => x"81",
           751 => x"8c",
           752 => x"81",
           753 => x"88",
           754 => x"83",
           755 => x"dc",
           756 => x"81",
           757 => x"54",
           758 => x"81",
           759 => x"04",
           760 => x"08",
           761 => x"d8",
           762 => x"0d",
           763 => x"dc",
           764 => x"05",
           765 => x"d8",
           766 => x"08",
           767 => x"38",
           768 => x"08",
           769 => x"30",
           770 => x"08",
           771 => x"80",
           772 => x"d8",
           773 => x"0c",
           774 => x"08",
           775 => x"8a",
           776 => x"81",
           777 => x"f4",
           778 => x"dc",
           779 => x"05",
           780 => x"d8",
           781 => x"0c",
           782 => x"08",
           783 => x"80",
           784 => x"81",
           785 => x"8c",
           786 => x"81",
           787 => x"8c",
           788 => x"0b",
           789 => x"08",
           790 => x"81",
           791 => x"fc",
           792 => x"38",
           793 => x"dc",
           794 => x"05",
           795 => x"d8",
           796 => x"08",
           797 => x"08",
           798 => x"80",
           799 => x"d8",
           800 => x"08",
           801 => x"d8",
           802 => x"08",
           803 => x"3f",
           804 => x"08",
           805 => x"d8",
           806 => x"0c",
           807 => x"d8",
           808 => x"08",
           809 => x"38",
           810 => x"08",
           811 => x"30",
           812 => x"08",
           813 => x"81",
           814 => x"f8",
           815 => x"81",
           816 => x"54",
           817 => x"81",
           818 => x"04",
           819 => x"08",
           820 => x"d8",
           821 => x"0d",
           822 => x"dc",
           823 => x"05",
           824 => x"d8",
           825 => x"08",
           826 => x"38",
           827 => x"08",
           828 => x"30",
           829 => x"08",
           830 => x"81",
           831 => x"d8",
           832 => x"0c",
           833 => x"08",
           834 => x"80",
           835 => x"81",
           836 => x"8c",
           837 => x"81",
           838 => x"8c",
           839 => x"53",
           840 => x"08",
           841 => x"52",
           842 => x"08",
           843 => x"51",
           844 => x"dc",
           845 => x"81",
           846 => x"f8",
           847 => x"81",
           848 => x"fc",
           849 => x"2e",
           850 => x"dc",
           851 => x"05",
           852 => x"dc",
           853 => x"05",
           854 => x"d8",
           855 => x"08",
           856 => x"cc",
           857 => x"3d",
           858 => x"d8",
           859 => x"dc",
           860 => x"81",
           861 => x"fd",
           862 => x"0b",
           863 => x"08",
           864 => x"80",
           865 => x"d8",
           866 => x"0c",
           867 => x"08",
           868 => x"81",
           869 => x"88",
           870 => x"b9",
           871 => x"d8",
           872 => x"08",
           873 => x"38",
           874 => x"dc",
           875 => x"05",
           876 => x"38",
           877 => x"08",
           878 => x"10",
           879 => x"08",
           880 => x"81",
           881 => x"fc",
           882 => x"81",
           883 => x"fc",
           884 => x"b8",
           885 => x"d8",
           886 => x"08",
           887 => x"e1",
           888 => x"d8",
           889 => x"08",
           890 => x"08",
           891 => x"26",
           892 => x"dc",
           893 => x"05",
           894 => x"d8",
           895 => x"08",
           896 => x"d8",
           897 => x"0c",
           898 => x"08",
           899 => x"81",
           900 => x"fc",
           901 => x"81",
           902 => x"f8",
           903 => x"dc",
           904 => x"05",
           905 => x"81",
           906 => x"fc",
           907 => x"dc",
           908 => x"05",
           909 => x"81",
           910 => x"8c",
           911 => x"95",
           912 => x"d8",
           913 => x"08",
           914 => x"38",
           915 => x"08",
           916 => x"70",
           917 => x"08",
           918 => x"51",
           919 => x"dc",
           920 => x"05",
           921 => x"dc",
           922 => x"05",
           923 => x"dc",
           924 => x"05",
           925 => x"cc",
           926 => x"0d",
           927 => x"0c",
           928 => x"0d",
           929 => x"02",
           930 => x"05",
           931 => x"53",
           932 => x"27",
           933 => x"83",
           934 => x"80",
           935 => x"ff",
           936 => x"ff",
           937 => x"73",
           938 => x"05",
           939 => x"12",
           940 => x"2e",
           941 => x"ef",
           942 => x"dc",
           943 => x"3d",
           944 => x"74",
           945 => x"07",
           946 => x"2b",
           947 => x"51",
           948 => x"a5",
           949 => x"70",
           950 => x"0c",
           951 => x"84",
           952 => x"72",
           953 => x"05",
           954 => x"71",
           955 => x"53",
           956 => x"52",
           957 => x"dd",
           958 => x"27",
           959 => x"71",
           960 => x"53",
           961 => x"52",
           962 => x"f2",
           963 => x"ff",
           964 => x"3d",
           965 => x"70",
           966 => x"06",
           967 => x"70",
           968 => x"73",
           969 => x"56",
           970 => x"08",
           971 => x"38",
           972 => x"52",
           973 => x"81",
           974 => x"54",
           975 => x"9d",
           976 => x"55",
           977 => x"09",
           978 => x"38",
           979 => x"14",
           980 => x"81",
           981 => x"56",
           982 => x"e5",
           983 => x"55",
           984 => x"06",
           985 => x"06",
           986 => x"81",
           987 => x"52",
           988 => x"0d",
           989 => x"70",
           990 => x"ff",
           991 => x"f8",
           992 => x"80",
           993 => x"51",
           994 => x"84",
           995 => x"71",
           996 => x"54",
           997 => x"2e",
           998 => x"75",
           999 => x"94",
          1000 => x"81",
          1001 => x"87",
          1002 => x"fe",
          1003 => x"52",
          1004 => x"88",
          1005 => x"86",
          1006 => x"cc",
          1007 => x"06",
          1008 => x"14",
          1009 => x"80",
          1010 => x"71",
          1011 => x"0c",
          1012 => x"04",
          1013 => x"77",
          1014 => x"53",
          1015 => x"80",
          1016 => x"38",
          1017 => x"70",
          1018 => x"81",
          1019 => x"81",
          1020 => x"39",
          1021 => x"39",
          1022 => x"80",
          1023 => x"81",
          1024 => x"55",
          1025 => x"2e",
          1026 => x"55",
          1027 => x"84",
          1028 => x"38",
          1029 => x"06",
          1030 => x"2e",
          1031 => x"88",
          1032 => x"70",
          1033 => x"34",
          1034 => x"71",
          1035 => x"dc",
          1036 => x"3d",
          1037 => x"3d",
          1038 => x"72",
          1039 => x"91",
          1040 => x"fc",
          1041 => x"51",
          1042 => x"81",
          1043 => x"85",
          1044 => x"83",
          1045 => x"72",
          1046 => x"0c",
          1047 => x"04",
          1048 => x"76",
          1049 => x"ff",
          1050 => x"81",
          1051 => x"26",
          1052 => x"83",
          1053 => x"05",
          1054 => x"70",
          1055 => x"8a",
          1056 => x"33",
          1057 => x"70",
          1058 => x"fe",
          1059 => x"33",
          1060 => x"70",
          1061 => x"f2",
          1062 => x"33",
          1063 => x"70",
          1064 => x"e6",
          1065 => x"22",
          1066 => x"74",
          1067 => x"80",
          1068 => x"13",
          1069 => x"52",
          1070 => x"26",
          1071 => x"81",
          1072 => x"98",
          1073 => x"22",
          1074 => x"bc",
          1075 => x"33",
          1076 => x"b8",
          1077 => x"33",
          1078 => x"b4",
          1079 => x"33",
          1080 => x"b0",
          1081 => x"33",
          1082 => x"ac",
          1083 => x"33",
          1084 => x"a8",
          1085 => x"c0",
          1086 => x"73",
          1087 => x"a0",
          1088 => x"87",
          1089 => x"0c",
          1090 => x"81",
          1091 => x"86",
          1092 => x"f3",
          1093 => x"5b",
          1094 => x"9c",
          1095 => x"0c",
          1096 => x"bc",
          1097 => x"7b",
          1098 => x"98",
          1099 => x"79",
          1100 => x"87",
          1101 => x"08",
          1102 => x"1c",
          1103 => x"98",
          1104 => x"79",
          1105 => x"87",
          1106 => x"08",
          1107 => x"1c",
          1108 => x"98",
          1109 => x"79",
          1110 => x"87",
          1111 => x"08",
          1112 => x"1c",
          1113 => x"98",
          1114 => x"79",
          1115 => x"80",
          1116 => x"83",
          1117 => x"59",
          1118 => x"ff",
          1119 => x"1b",
          1120 => x"1b",
          1121 => x"1b",
          1122 => x"1b",
          1123 => x"1b",
          1124 => x"83",
          1125 => x"52",
          1126 => x"51",
          1127 => x"8f",
          1128 => x"ff",
          1129 => x"8f",
          1130 => x"30",
          1131 => x"51",
          1132 => x"0b",
          1133 => x"f4",
          1134 => x"0d",
          1135 => x"0d",
          1136 => x"81",
          1137 => x"70",
          1138 => x"57",
          1139 => x"c0",
          1140 => x"74",
          1141 => x"38",
          1142 => x"94",
          1143 => x"70",
          1144 => x"81",
          1145 => x"52",
          1146 => x"8c",
          1147 => x"2a",
          1148 => x"51",
          1149 => x"38",
          1150 => x"70",
          1151 => x"51",
          1152 => x"8d",
          1153 => x"2a",
          1154 => x"51",
          1155 => x"be",
          1156 => x"ff",
          1157 => x"c0",
          1158 => x"70",
          1159 => x"38",
          1160 => x"90",
          1161 => x"0c",
          1162 => x"cc",
          1163 => x"0d",
          1164 => x"0d",
          1165 => x"33",
          1166 => x"d8",
          1167 => x"81",
          1168 => x"55",
          1169 => x"94",
          1170 => x"80",
          1171 => x"87",
          1172 => x"51",
          1173 => x"96",
          1174 => x"06",
          1175 => x"70",
          1176 => x"38",
          1177 => x"70",
          1178 => x"51",
          1179 => x"72",
          1180 => x"81",
          1181 => x"70",
          1182 => x"38",
          1183 => x"70",
          1184 => x"51",
          1185 => x"38",
          1186 => x"06",
          1187 => x"94",
          1188 => x"80",
          1189 => x"87",
          1190 => x"52",
          1191 => x"87",
          1192 => x"f9",
          1193 => x"54",
          1194 => x"70",
          1195 => x"53",
          1196 => x"77",
          1197 => x"38",
          1198 => x"06",
          1199 => x"0b",
          1200 => x"33",
          1201 => x"06",
          1202 => x"58",
          1203 => x"84",
          1204 => x"2e",
          1205 => x"c0",
          1206 => x"70",
          1207 => x"2a",
          1208 => x"53",
          1209 => x"80",
          1210 => x"71",
          1211 => x"81",
          1212 => x"70",
          1213 => x"81",
          1214 => x"06",
          1215 => x"80",
          1216 => x"71",
          1217 => x"81",
          1218 => x"70",
          1219 => x"74",
          1220 => x"51",
          1221 => x"80",
          1222 => x"2e",
          1223 => x"c0",
          1224 => x"77",
          1225 => x"17",
          1226 => x"81",
          1227 => x"53",
          1228 => x"84",
          1229 => x"dc",
          1230 => x"3d",
          1231 => x"3d",
          1232 => x"81",
          1233 => x"70",
          1234 => x"54",
          1235 => x"94",
          1236 => x"80",
          1237 => x"87",
          1238 => x"51",
          1239 => x"82",
          1240 => x"06",
          1241 => x"70",
          1242 => x"38",
          1243 => x"06",
          1244 => x"94",
          1245 => x"80",
          1246 => x"87",
          1247 => x"52",
          1248 => x"81",
          1249 => x"dc",
          1250 => x"84",
          1251 => x"fe",
          1252 => x"0b",
          1253 => x"33",
          1254 => x"06",
          1255 => x"c0",
          1256 => x"70",
          1257 => x"38",
          1258 => x"94",
          1259 => x"70",
          1260 => x"81",
          1261 => x"51",
          1262 => x"80",
          1263 => x"72",
          1264 => x"51",
          1265 => x"80",
          1266 => x"2e",
          1267 => x"c0",
          1268 => x"71",
          1269 => x"2b",
          1270 => x"51",
          1271 => x"81",
          1272 => x"84",
          1273 => x"ff",
          1274 => x"c0",
          1275 => x"70",
          1276 => x"06",
          1277 => x"80",
          1278 => x"38",
          1279 => x"a4",
          1280 => x"f8",
          1281 => x"9e",
          1282 => x"d8",
          1283 => x"c0",
          1284 => x"81",
          1285 => x"87",
          1286 => x"08",
          1287 => x"0c",
          1288 => x"9c",
          1289 => x"88",
          1290 => x"9e",
          1291 => x"d9",
          1292 => x"c0",
          1293 => x"81",
          1294 => x"87",
          1295 => x"08",
          1296 => x"0c",
          1297 => x"b4",
          1298 => x"98",
          1299 => x"9e",
          1300 => x"d9",
          1301 => x"c0",
          1302 => x"81",
          1303 => x"87",
          1304 => x"08",
          1305 => x"0c",
          1306 => x"c4",
          1307 => x"a8",
          1308 => x"9e",
          1309 => x"70",
          1310 => x"23",
          1311 => x"84",
          1312 => x"b0",
          1313 => x"9e",
          1314 => x"d9",
          1315 => x"c0",
          1316 => x"81",
          1317 => x"81",
          1318 => x"bc",
          1319 => x"87",
          1320 => x"08",
          1321 => x"0a",
          1322 => x"52",
          1323 => x"83",
          1324 => x"71",
          1325 => x"34",
          1326 => x"c0",
          1327 => x"70",
          1328 => x"06",
          1329 => x"70",
          1330 => x"38",
          1331 => x"81",
          1332 => x"80",
          1333 => x"9e",
          1334 => x"90",
          1335 => x"51",
          1336 => x"80",
          1337 => x"81",
          1338 => x"d9",
          1339 => x"0b",
          1340 => x"90",
          1341 => x"80",
          1342 => x"52",
          1343 => x"2e",
          1344 => x"52",
          1345 => x"c0",
          1346 => x"87",
          1347 => x"08",
          1348 => x"80",
          1349 => x"52",
          1350 => x"83",
          1351 => x"71",
          1352 => x"34",
          1353 => x"c0",
          1354 => x"70",
          1355 => x"06",
          1356 => x"70",
          1357 => x"38",
          1358 => x"81",
          1359 => x"80",
          1360 => x"9e",
          1361 => x"84",
          1362 => x"51",
          1363 => x"80",
          1364 => x"81",
          1365 => x"d9",
          1366 => x"0b",
          1367 => x"90",
          1368 => x"80",
          1369 => x"52",
          1370 => x"2e",
          1371 => x"52",
          1372 => x"c4",
          1373 => x"87",
          1374 => x"08",
          1375 => x"80",
          1376 => x"52",
          1377 => x"83",
          1378 => x"71",
          1379 => x"34",
          1380 => x"c0",
          1381 => x"70",
          1382 => x"06",
          1383 => x"70",
          1384 => x"38",
          1385 => x"81",
          1386 => x"80",
          1387 => x"9e",
          1388 => x"a0",
          1389 => x"52",
          1390 => x"2e",
          1391 => x"52",
          1392 => x"c7",
          1393 => x"9e",
          1394 => x"98",
          1395 => x"8a",
          1396 => x"51",
          1397 => x"c8",
          1398 => x"87",
          1399 => x"08",
          1400 => x"06",
          1401 => x"70",
          1402 => x"38",
          1403 => x"81",
          1404 => x"87",
          1405 => x"08",
          1406 => x"06",
          1407 => x"51",
          1408 => x"81",
          1409 => x"80",
          1410 => x"9e",
          1411 => x"88",
          1412 => x"52",
          1413 => x"83",
          1414 => x"71",
          1415 => x"34",
          1416 => x"90",
          1417 => x"06",
          1418 => x"81",
          1419 => x"83",
          1420 => x"fb",
          1421 => x"c5",
          1422 => x"c5",
          1423 => x"bc",
          1424 => x"80",
          1425 => x"81",
          1426 => x"85",
          1427 => x"c6",
          1428 => x"ad",
          1429 => x"be",
          1430 => x"80",
          1431 => x"81",
          1432 => x"81",
          1433 => x"11",
          1434 => x"c6",
          1435 => x"f5",
          1436 => x"c3",
          1437 => x"80",
          1438 => x"81",
          1439 => x"81",
          1440 => x"11",
          1441 => x"c6",
          1442 => x"d9",
          1443 => x"c0",
          1444 => x"80",
          1445 => x"81",
          1446 => x"81",
          1447 => x"11",
          1448 => x"c6",
          1449 => x"bd",
          1450 => x"c1",
          1451 => x"80",
          1452 => x"81",
          1453 => x"81",
          1454 => x"11",
          1455 => x"c6",
          1456 => x"a1",
          1457 => x"c2",
          1458 => x"80",
          1459 => x"81",
          1460 => x"81",
          1461 => x"11",
          1462 => x"c7",
          1463 => x"85",
          1464 => x"c7",
          1465 => x"80",
          1466 => x"81",
          1467 => x"52",
          1468 => x"51",
          1469 => x"81",
          1470 => x"54",
          1471 => x"8d",
          1472 => x"cc",
          1473 => x"c7",
          1474 => x"d9",
          1475 => x"c9",
          1476 => x"80",
          1477 => x"81",
          1478 => x"52",
          1479 => x"51",
          1480 => x"81",
          1481 => x"54",
          1482 => x"88",
          1483 => x"90",
          1484 => x"3f",
          1485 => x"33",
          1486 => x"2e",
          1487 => x"c8",
          1488 => x"bd",
          1489 => x"c4",
          1490 => x"80",
          1491 => x"81",
          1492 => x"83",
          1493 => x"d9",
          1494 => x"73",
          1495 => x"38",
          1496 => x"51",
          1497 => x"81",
          1498 => x"54",
          1499 => x"88",
          1500 => x"c8",
          1501 => x"3f",
          1502 => x"51",
          1503 => x"81",
          1504 => x"52",
          1505 => x"51",
          1506 => x"81",
          1507 => x"52",
          1508 => x"51",
          1509 => x"81",
          1510 => x"52",
          1511 => x"51",
          1512 => x"81",
          1513 => x"82",
          1514 => x"d9",
          1515 => x"81",
          1516 => x"88",
          1517 => x"d9",
          1518 => x"bd",
          1519 => x"75",
          1520 => x"3f",
          1521 => x"08",
          1522 => x"29",
          1523 => x"54",
          1524 => x"cc",
          1525 => x"ca",
          1526 => x"89",
          1527 => x"c3",
          1528 => x"80",
          1529 => x"81",
          1530 => x"56",
          1531 => x"52",
          1532 => x"86",
          1533 => x"cc",
          1534 => x"c0",
          1535 => x"31",
          1536 => x"dc",
          1537 => x"81",
          1538 => x"87",
          1539 => x"d9",
          1540 => x"73",
          1541 => x"38",
          1542 => x"08",
          1543 => x"c0",
          1544 => x"e6",
          1545 => x"dc",
          1546 => x"84",
          1547 => x"71",
          1548 => x"81",
          1549 => x"52",
          1550 => x"51",
          1551 => x"81",
          1552 => x"81",
          1553 => x"3d",
          1554 => x"3d",
          1555 => x"05",
          1556 => x"52",
          1557 => x"aa",
          1558 => x"29",
          1559 => x"05",
          1560 => x"04",
          1561 => x"51",
          1562 => x"cb",
          1563 => x"39",
          1564 => x"51",
          1565 => x"cb",
          1566 => x"39",
          1567 => x"51",
          1568 => x"cb",
          1569 => x"f9",
          1570 => x"0d",
          1571 => x"80",
          1572 => x"0b",
          1573 => x"84",
          1574 => x"d9",
          1575 => x"c0",
          1576 => x"04",
          1577 => x"02",
          1578 => x"53",
          1579 => x"09",
          1580 => x"38",
          1581 => x"3f",
          1582 => x"08",
          1583 => x"2e",
          1584 => x"72",
          1585 => x"e4",
          1586 => x"81",
          1587 => x"8f",
          1588 => x"dc",
          1589 => x"80",
          1590 => x"72",
          1591 => x"84",
          1592 => x"fe",
          1593 => x"97",
          1594 => x"dc",
          1595 => x"81",
          1596 => x"54",
          1597 => x"3f",
          1598 => x"dc",
          1599 => x"0d",
          1600 => x"0d",
          1601 => x"33",
          1602 => x"06",
          1603 => x"80",
          1604 => x"72",
          1605 => x"51",
          1606 => x"ff",
          1607 => x"39",
          1608 => x"04",
          1609 => x"77",
          1610 => x"08",
          1611 => x"dc",
          1612 => x"73",
          1613 => x"ff",
          1614 => x"71",
          1615 => x"38",
          1616 => x"06",
          1617 => x"54",
          1618 => x"e7",
          1619 => x"dc",
          1620 => x"3d",
          1621 => x"3d",
          1622 => x"59",
          1623 => x"81",
          1624 => x"56",
          1625 => x"84",
          1626 => x"a5",
          1627 => x"06",
          1628 => x"80",
          1629 => x"81",
          1630 => x"58",
          1631 => x"b0",
          1632 => x"06",
          1633 => x"5a",
          1634 => x"ad",
          1635 => x"06",
          1636 => x"5a",
          1637 => x"05",
          1638 => x"75",
          1639 => x"81",
          1640 => x"77",
          1641 => x"08",
          1642 => x"05",
          1643 => x"5d",
          1644 => x"39",
          1645 => x"72",
          1646 => x"38",
          1647 => x"7b",
          1648 => x"05",
          1649 => x"70",
          1650 => x"33",
          1651 => x"39",
          1652 => x"32",
          1653 => x"72",
          1654 => x"78",
          1655 => x"70",
          1656 => x"07",
          1657 => x"07",
          1658 => x"51",
          1659 => x"80",
          1660 => x"79",
          1661 => x"70",
          1662 => x"33",
          1663 => x"80",
          1664 => x"38",
          1665 => x"e0",
          1666 => x"38",
          1667 => x"81",
          1668 => x"53",
          1669 => x"2e",
          1670 => x"73",
          1671 => x"a2",
          1672 => x"c3",
          1673 => x"38",
          1674 => x"24",
          1675 => x"80",
          1676 => x"8c",
          1677 => x"39",
          1678 => x"2e",
          1679 => x"81",
          1680 => x"80",
          1681 => x"80",
          1682 => x"d5",
          1683 => x"73",
          1684 => x"8e",
          1685 => x"39",
          1686 => x"2e",
          1687 => x"80",
          1688 => x"84",
          1689 => x"56",
          1690 => x"74",
          1691 => x"72",
          1692 => x"38",
          1693 => x"15",
          1694 => x"54",
          1695 => x"38",
          1696 => x"56",
          1697 => x"81",
          1698 => x"72",
          1699 => x"38",
          1700 => x"90",
          1701 => x"06",
          1702 => x"2e",
          1703 => x"51",
          1704 => x"74",
          1705 => x"53",
          1706 => x"fd",
          1707 => x"51",
          1708 => x"ef",
          1709 => x"19",
          1710 => x"53",
          1711 => x"39",
          1712 => x"39",
          1713 => x"39",
          1714 => x"39",
          1715 => x"39",
          1716 => x"d0",
          1717 => x"39",
          1718 => x"70",
          1719 => x"53",
          1720 => x"88",
          1721 => x"19",
          1722 => x"39",
          1723 => x"54",
          1724 => x"74",
          1725 => x"70",
          1726 => x"07",
          1727 => x"55",
          1728 => x"80",
          1729 => x"72",
          1730 => x"38",
          1731 => x"90",
          1732 => x"80",
          1733 => x"5e",
          1734 => x"74",
          1735 => x"3f",
          1736 => x"08",
          1737 => x"7c",
          1738 => x"54",
          1739 => x"81",
          1740 => x"55",
          1741 => x"92",
          1742 => x"53",
          1743 => x"2e",
          1744 => x"14",
          1745 => x"ff",
          1746 => x"14",
          1747 => x"70",
          1748 => x"34",
          1749 => x"30",
          1750 => x"9f",
          1751 => x"57",
          1752 => x"85",
          1753 => x"b1",
          1754 => x"2a",
          1755 => x"51",
          1756 => x"2e",
          1757 => x"3d",
          1758 => x"05",
          1759 => x"34",
          1760 => x"76",
          1761 => x"54",
          1762 => x"72",
          1763 => x"54",
          1764 => x"70",
          1765 => x"56",
          1766 => x"81",
          1767 => x"7b",
          1768 => x"73",
          1769 => x"3f",
          1770 => x"53",
          1771 => x"74",
          1772 => x"53",
          1773 => x"eb",
          1774 => x"77",
          1775 => x"53",
          1776 => x"14",
          1777 => x"54",
          1778 => x"3f",
          1779 => x"74",
          1780 => x"53",
          1781 => x"fb",
          1782 => x"51",
          1783 => x"ef",
          1784 => x"0d",
          1785 => x"0d",
          1786 => x"70",
          1787 => x"08",
          1788 => x"51",
          1789 => x"85",
          1790 => x"fe",
          1791 => x"81",
          1792 => x"85",
          1793 => x"52",
          1794 => x"ca",
          1795 => x"e4",
          1796 => x"73",
          1797 => x"81",
          1798 => x"84",
          1799 => x"fd",
          1800 => x"dc",
          1801 => x"81",
          1802 => x"87",
          1803 => x"53",
          1804 => x"fa",
          1805 => x"81",
          1806 => x"85",
          1807 => x"fb",
          1808 => x"79",
          1809 => x"08",
          1810 => x"57",
          1811 => x"71",
          1812 => x"e0",
          1813 => x"e0",
          1814 => x"2d",
          1815 => x"08",
          1816 => x"53",
          1817 => x"80",
          1818 => x"8d",
          1819 => x"72",
          1820 => x"30",
          1821 => x"51",
          1822 => x"80",
          1823 => x"71",
          1824 => x"38",
          1825 => x"97",
          1826 => x"25",
          1827 => x"16",
          1828 => x"25",
          1829 => x"14",
          1830 => x"34",
          1831 => x"72",
          1832 => x"3f",
          1833 => x"73",
          1834 => x"72",
          1835 => x"f7",
          1836 => x"53",
          1837 => x"cc",
          1838 => x"0d",
          1839 => x"0d",
          1840 => x"08",
          1841 => x"e0",
          1842 => x"76",
          1843 => x"ef",
          1844 => x"dc",
          1845 => x"3d",
          1846 => x"3d",
          1847 => x"5a",
          1848 => x"7a",
          1849 => x"08",
          1850 => x"53",
          1851 => x"09",
          1852 => x"38",
          1853 => x"0c",
          1854 => x"ad",
          1855 => x"06",
          1856 => x"76",
          1857 => x"0c",
          1858 => x"33",
          1859 => x"73",
          1860 => x"81",
          1861 => x"38",
          1862 => x"05",
          1863 => x"08",
          1864 => x"53",
          1865 => x"2e",
          1866 => x"57",
          1867 => x"2e",
          1868 => x"39",
          1869 => x"13",
          1870 => x"08",
          1871 => x"53",
          1872 => x"55",
          1873 => x"80",
          1874 => x"14",
          1875 => x"88",
          1876 => x"27",
          1877 => x"eb",
          1878 => x"53",
          1879 => x"89",
          1880 => x"38",
          1881 => x"55",
          1882 => x"8a",
          1883 => x"a0",
          1884 => x"c2",
          1885 => x"74",
          1886 => x"e0",
          1887 => x"ff",
          1888 => x"d0",
          1889 => x"ff",
          1890 => x"90",
          1891 => x"38",
          1892 => x"81",
          1893 => x"53",
          1894 => x"ca",
          1895 => x"27",
          1896 => x"77",
          1897 => x"08",
          1898 => x"0c",
          1899 => x"33",
          1900 => x"ff",
          1901 => x"80",
          1902 => x"74",
          1903 => x"79",
          1904 => x"74",
          1905 => x"0c",
          1906 => x"04",
          1907 => x"7a",
          1908 => x"80",
          1909 => x"58",
          1910 => x"33",
          1911 => x"a0",
          1912 => x"06",
          1913 => x"13",
          1914 => x"39",
          1915 => x"09",
          1916 => x"38",
          1917 => x"11",
          1918 => x"08",
          1919 => x"54",
          1920 => x"2e",
          1921 => x"80",
          1922 => x"08",
          1923 => x"0c",
          1924 => x"33",
          1925 => x"80",
          1926 => x"38",
          1927 => x"80",
          1928 => x"38",
          1929 => x"57",
          1930 => x"0c",
          1931 => x"33",
          1932 => x"39",
          1933 => x"74",
          1934 => x"38",
          1935 => x"80",
          1936 => x"89",
          1937 => x"38",
          1938 => x"d0",
          1939 => x"55",
          1940 => x"80",
          1941 => x"39",
          1942 => x"d9",
          1943 => x"80",
          1944 => x"27",
          1945 => x"80",
          1946 => x"89",
          1947 => x"70",
          1948 => x"55",
          1949 => x"70",
          1950 => x"55",
          1951 => x"27",
          1952 => x"14",
          1953 => x"06",
          1954 => x"74",
          1955 => x"73",
          1956 => x"38",
          1957 => x"14",
          1958 => x"05",
          1959 => x"08",
          1960 => x"54",
          1961 => x"39",
          1962 => x"84",
          1963 => x"55",
          1964 => x"81",
          1965 => x"dc",
          1966 => x"3d",
          1967 => x"3d",
          1968 => x"05",
          1969 => x"52",
          1970 => x"87",
          1971 => x"d4",
          1972 => x"71",
          1973 => x"0c",
          1974 => x"04",
          1975 => x"02",
          1976 => x"02",
          1977 => x"05",
          1978 => x"83",
          1979 => x"26",
          1980 => x"72",
          1981 => x"c0",
          1982 => x"53",
          1983 => x"74",
          1984 => x"38",
          1985 => x"73",
          1986 => x"c0",
          1987 => x"51",
          1988 => x"85",
          1989 => x"98",
          1990 => x"52",
          1991 => x"82",
          1992 => x"70",
          1993 => x"38",
          1994 => x"8c",
          1995 => x"ec",
          1996 => x"fc",
          1997 => x"52",
          1998 => x"87",
          1999 => x"08",
          2000 => x"2e",
          2001 => x"81",
          2002 => x"34",
          2003 => x"13",
          2004 => x"81",
          2005 => x"86",
          2006 => x"f3",
          2007 => x"62",
          2008 => x"05",
          2009 => x"57",
          2010 => x"83",
          2011 => x"fe",
          2012 => x"dc",
          2013 => x"06",
          2014 => x"71",
          2015 => x"71",
          2016 => x"2b",
          2017 => x"80",
          2018 => x"92",
          2019 => x"c0",
          2020 => x"41",
          2021 => x"5a",
          2022 => x"87",
          2023 => x"0c",
          2024 => x"84",
          2025 => x"08",
          2026 => x"70",
          2027 => x"53",
          2028 => x"2e",
          2029 => x"08",
          2030 => x"70",
          2031 => x"34",
          2032 => x"80",
          2033 => x"53",
          2034 => x"2e",
          2035 => x"53",
          2036 => x"26",
          2037 => x"80",
          2038 => x"87",
          2039 => x"08",
          2040 => x"38",
          2041 => x"8c",
          2042 => x"80",
          2043 => x"78",
          2044 => x"99",
          2045 => x"0c",
          2046 => x"8c",
          2047 => x"08",
          2048 => x"51",
          2049 => x"38",
          2050 => x"8d",
          2051 => x"17",
          2052 => x"81",
          2053 => x"53",
          2054 => x"2e",
          2055 => x"fc",
          2056 => x"52",
          2057 => x"7d",
          2058 => x"ed",
          2059 => x"80",
          2060 => x"71",
          2061 => x"38",
          2062 => x"53",
          2063 => x"cc",
          2064 => x"0d",
          2065 => x"0d",
          2066 => x"02",
          2067 => x"05",
          2068 => x"58",
          2069 => x"80",
          2070 => x"fc",
          2071 => x"dc",
          2072 => x"06",
          2073 => x"71",
          2074 => x"81",
          2075 => x"38",
          2076 => x"2b",
          2077 => x"80",
          2078 => x"92",
          2079 => x"c0",
          2080 => x"40",
          2081 => x"5a",
          2082 => x"c0",
          2083 => x"76",
          2084 => x"76",
          2085 => x"75",
          2086 => x"2a",
          2087 => x"51",
          2088 => x"80",
          2089 => x"7a",
          2090 => x"5c",
          2091 => x"81",
          2092 => x"81",
          2093 => x"06",
          2094 => x"80",
          2095 => x"87",
          2096 => x"08",
          2097 => x"38",
          2098 => x"8c",
          2099 => x"80",
          2100 => x"77",
          2101 => x"99",
          2102 => x"0c",
          2103 => x"8c",
          2104 => x"08",
          2105 => x"51",
          2106 => x"38",
          2107 => x"8d",
          2108 => x"70",
          2109 => x"84",
          2110 => x"5b",
          2111 => x"2e",
          2112 => x"fc",
          2113 => x"52",
          2114 => x"7d",
          2115 => x"f8",
          2116 => x"80",
          2117 => x"71",
          2118 => x"38",
          2119 => x"53",
          2120 => x"cc",
          2121 => x"0d",
          2122 => x"0d",
          2123 => x"05",
          2124 => x"02",
          2125 => x"05",
          2126 => x"54",
          2127 => x"fe",
          2128 => x"cc",
          2129 => x"53",
          2130 => x"80",
          2131 => x"0b",
          2132 => x"8c",
          2133 => x"71",
          2134 => x"dc",
          2135 => x"24",
          2136 => x"84",
          2137 => x"92",
          2138 => x"54",
          2139 => x"8d",
          2140 => x"39",
          2141 => x"80",
          2142 => x"cb",
          2143 => x"70",
          2144 => x"81",
          2145 => x"52",
          2146 => x"8a",
          2147 => x"98",
          2148 => x"71",
          2149 => x"c0",
          2150 => x"52",
          2151 => x"81",
          2152 => x"c0",
          2153 => x"53",
          2154 => x"82",
          2155 => x"71",
          2156 => x"39",
          2157 => x"39",
          2158 => x"77",
          2159 => x"81",
          2160 => x"72",
          2161 => x"84",
          2162 => x"73",
          2163 => x"0c",
          2164 => x"04",
          2165 => x"74",
          2166 => x"71",
          2167 => x"2b",
          2168 => x"cc",
          2169 => x"84",
          2170 => x"fd",
          2171 => x"83",
          2172 => x"12",
          2173 => x"2b",
          2174 => x"07",
          2175 => x"70",
          2176 => x"2b",
          2177 => x"07",
          2178 => x"0c",
          2179 => x"56",
          2180 => x"3d",
          2181 => x"3d",
          2182 => x"84",
          2183 => x"22",
          2184 => x"72",
          2185 => x"54",
          2186 => x"2a",
          2187 => x"34",
          2188 => x"04",
          2189 => x"73",
          2190 => x"70",
          2191 => x"05",
          2192 => x"88",
          2193 => x"72",
          2194 => x"54",
          2195 => x"2a",
          2196 => x"70",
          2197 => x"34",
          2198 => x"51",
          2199 => x"83",
          2200 => x"fe",
          2201 => x"75",
          2202 => x"51",
          2203 => x"92",
          2204 => x"81",
          2205 => x"73",
          2206 => x"55",
          2207 => x"51",
          2208 => x"3d",
          2209 => x"3d",
          2210 => x"76",
          2211 => x"72",
          2212 => x"05",
          2213 => x"11",
          2214 => x"38",
          2215 => x"04",
          2216 => x"78",
          2217 => x"56",
          2218 => x"81",
          2219 => x"74",
          2220 => x"56",
          2221 => x"31",
          2222 => x"52",
          2223 => x"80",
          2224 => x"71",
          2225 => x"38",
          2226 => x"cc",
          2227 => x"0d",
          2228 => x"0d",
          2229 => x"51",
          2230 => x"73",
          2231 => x"81",
          2232 => x"33",
          2233 => x"38",
          2234 => x"dc",
          2235 => x"3d",
          2236 => x"0b",
          2237 => x"0c",
          2238 => x"81",
          2239 => x"04",
          2240 => x"7b",
          2241 => x"83",
          2242 => x"5a",
          2243 => x"80",
          2244 => x"54",
          2245 => x"53",
          2246 => x"53",
          2247 => x"52",
          2248 => x"3f",
          2249 => x"08",
          2250 => x"81",
          2251 => x"81",
          2252 => x"83",
          2253 => x"16",
          2254 => x"18",
          2255 => x"18",
          2256 => x"58",
          2257 => x"9f",
          2258 => x"33",
          2259 => x"2e",
          2260 => x"93",
          2261 => x"76",
          2262 => x"52",
          2263 => x"51",
          2264 => x"83",
          2265 => x"79",
          2266 => x"0c",
          2267 => x"04",
          2268 => x"78",
          2269 => x"80",
          2270 => x"17",
          2271 => x"38",
          2272 => x"fc",
          2273 => x"cc",
          2274 => x"dc",
          2275 => x"38",
          2276 => x"53",
          2277 => x"81",
          2278 => x"f7",
          2279 => x"dc",
          2280 => x"2e",
          2281 => x"55",
          2282 => x"b0",
          2283 => x"81",
          2284 => x"88",
          2285 => x"f8",
          2286 => x"70",
          2287 => x"c0",
          2288 => x"cc",
          2289 => x"dc",
          2290 => x"91",
          2291 => x"55",
          2292 => x"09",
          2293 => x"f0",
          2294 => x"33",
          2295 => x"2e",
          2296 => x"80",
          2297 => x"80",
          2298 => x"cc",
          2299 => x"17",
          2300 => x"fd",
          2301 => x"d4",
          2302 => x"b2",
          2303 => x"96",
          2304 => x"85",
          2305 => x"75",
          2306 => x"3f",
          2307 => x"e4",
          2308 => x"98",
          2309 => x"9c",
          2310 => x"08",
          2311 => x"17",
          2312 => x"3f",
          2313 => x"52",
          2314 => x"51",
          2315 => x"a0",
          2316 => x"05",
          2317 => x"0c",
          2318 => x"75",
          2319 => x"33",
          2320 => x"3f",
          2321 => x"34",
          2322 => x"52",
          2323 => x"51",
          2324 => x"81",
          2325 => x"80",
          2326 => x"81",
          2327 => x"dc",
          2328 => x"3d",
          2329 => x"3d",
          2330 => x"1a",
          2331 => x"fe",
          2332 => x"54",
          2333 => x"73",
          2334 => x"8a",
          2335 => x"71",
          2336 => x"08",
          2337 => x"75",
          2338 => x"0c",
          2339 => x"04",
          2340 => x"7a",
          2341 => x"56",
          2342 => x"77",
          2343 => x"38",
          2344 => x"08",
          2345 => x"38",
          2346 => x"54",
          2347 => x"2e",
          2348 => x"72",
          2349 => x"38",
          2350 => x"8d",
          2351 => x"39",
          2352 => x"81",
          2353 => x"b6",
          2354 => x"2a",
          2355 => x"2a",
          2356 => x"05",
          2357 => x"55",
          2358 => x"81",
          2359 => x"81",
          2360 => x"83",
          2361 => x"b4",
          2362 => x"17",
          2363 => x"a4",
          2364 => x"55",
          2365 => x"57",
          2366 => x"3f",
          2367 => x"08",
          2368 => x"74",
          2369 => x"14",
          2370 => x"70",
          2371 => x"07",
          2372 => x"71",
          2373 => x"52",
          2374 => x"72",
          2375 => x"75",
          2376 => x"58",
          2377 => x"76",
          2378 => x"15",
          2379 => x"73",
          2380 => x"3f",
          2381 => x"08",
          2382 => x"76",
          2383 => x"06",
          2384 => x"05",
          2385 => x"3f",
          2386 => x"08",
          2387 => x"06",
          2388 => x"76",
          2389 => x"15",
          2390 => x"73",
          2391 => x"3f",
          2392 => x"08",
          2393 => x"82",
          2394 => x"06",
          2395 => x"05",
          2396 => x"3f",
          2397 => x"08",
          2398 => x"58",
          2399 => x"58",
          2400 => x"cc",
          2401 => x"0d",
          2402 => x"0d",
          2403 => x"5a",
          2404 => x"59",
          2405 => x"82",
          2406 => x"98",
          2407 => x"82",
          2408 => x"33",
          2409 => x"2e",
          2410 => x"72",
          2411 => x"38",
          2412 => x"8d",
          2413 => x"39",
          2414 => x"81",
          2415 => x"f7",
          2416 => x"2a",
          2417 => x"2a",
          2418 => x"05",
          2419 => x"55",
          2420 => x"81",
          2421 => x"59",
          2422 => x"08",
          2423 => x"74",
          2424 => x"16",
          2425 => x"16",
          2426 => x"59",
          2427 => x"53",
          2428 => x"8f",
          2429 => x"2b",
          2430 => x"74",
          2431 => x"71",
          2432 => x"72",
          2433 => x"0b",
          2434 => x"74",
          2435 => x"17",
          2436 => x"75",
          2437 => x"3f",
          2438 => x"08",
          2439 => x"cc",
          2440 => x"38",
          2441 => x"06",
          2442 => x"78",
          2443 => x"54",
          2444 => x"77",
          2445 => x"33",
          2446 => x"71",
          2447 => x"51",
          2448 => x"34",
          2449 => x"76",
          2450 => x"17",
          2451 => x"75",
          2452 => x"3f",
          2453 => x"08",
          2454 => x"cc",
          2455 => x"38",
          2456 => x"ff",
          2457 => x"10",
          2458 => x"76",
          2459 => x"51",
          2460 => x"be",
          2461 => x"2a",
          2462 => x"05",
          2463 => x"f9",
          2464 => x"dc",
          2465 => x"81",
          2466 => x"ab",
          2467 => x"0a",
          2468 => x"2b",
          2469 => x"70",
          2470 => x"70",
          2471 => x"54",
          2472 => x"81",
          2473 => x"8f",
          2474 => x"07",
          2475 => x"f7",
          2476 => x"0b",
          2477 => x"78",
          2478 => x"0c",
          2479 => x"04",
          2480 => x"7a",
          2481 => x"08",
          2482 => x"59",
          2483 => x"a4",
          2484 => x"17",
          2485 => x"38",
          2486 => x"aa",
          2487 => x"73",
          2488 => x"fd",
          2489 => x"dc",
          2490 => x"81",
          2491 => x"80",
          2492 => x"39",
          2493 => x"eb",
          2494 => x"80",
          2495 => x"dc",
          2496 => x"80",
          2497 => x"52",
          2498 => x"84",
          2499 => x"cc",
          2500 => x"dc",
          2501 => x"2e",
          2502 => x"81",
          2503 => x"81",
          2504 => x"81",
          2505 => x"ff",
          2506 => x"80",
          2507 => x"75",
          2508 => x"3f",
          2509 => x"08",
          2510 => x"16",
          2511 => x"90",
          2512 => x"55",
          2513 => x"27",
          2514 => x"15",
          2515 => x"84",
          2516 => x"07",
          2517 => x"17",
          2518 => x"76",
          2519 => x"a6",
          2520 => x"73",
          2521 => x"0c",
          2522 => x"04",
          2523 => x"7c",
          2524 => x"59",
          2525 => x"95",
          2526 => x"08",
          2527 => x"2e",
          2528 => x"17",
          2529 => x"b2",
          2530 => x"ae",
          2531 => x"7a",
          2532 => x"3f",
          2533 => x"81",
          2534 => x"27",
          2535 => x"81",
          2536 => x"55",
          2537 => x"08",
          2538 => x"d2",
          2539 => x"08",
          2540 => x"08",
          2541 => x"38",
          2542 => x"17",
          2543 => x"54",
          2544 => x"82",
          2545 => x"7a",
          2546 => x"06",
          2547 => x"81",
          2548 => x"17",
          2549 => x"83",
          2550 => x"75",
          2551 => x"f9",
          2552 => x"59",
          2553 => x"08",
          2554 => x"81",
          2555 => x"81",
          2556 => x"59",
          2557 => x"08",
          2558 => x"70",
          2559 => x"25",
          2560 => x"81",
          2561 => x"54",
          2562 => x"55",
          2563 => x"38",
          2564 => x"08",
          2565 => x"38",
          2566 => x"54",
          2567 => x"90",
          2568 => x"18",
          2569 => x"38",
          2570 => x"39",
          2571 => x"38",
          2572 => x"16",
          2573 => x"08",
          2574 => x"38",
          2575 => x"78",
          2576 => x"38",
          2577 => x"51",
          2578 => x"81",
          2579 => x"80",
          2580 => x"80",
          2581 => x"cc",
          2582 => x"09",
          2583 => x"38",
          2584 => x"08",
          2585 => x"cc",
          2586 => x"30",
          2587 => x"80",
          2588 => x"07",
          2589 => x"55",
          2590 => x"38",
          2591 => x"09",
          2592 => x"ae",
          2593 => x"80",
          2594 => x"53",
          2595 => x"51",
          2596 => x"81",
          2597 => x"81",
          2598 => x"30",
          2599 => x"cc",
          2600 => x"25",
          2601 => x"79",
          2602 => x"38",
          2603 => x"8f",
          2604 => x"79",
          2605 => x"f9",
          2606 => x"dc",
          2607 => x"74",
          2608 => x"8c",
          2609 => x"17",
          2610 => x"90",
          2611 => x"54",
          2612 => x"86",
          2613 => x"90",
          2614 => x"17",
          2615 => x"54",
          2616 => x"34",
          2617 => x"56",
          2618 => x"90",
          2619 => x"80",
          2620 => x"81",
          2621 => x"55",
          2622 => x"56",
          2623 => x"81",
          2624 => x"8c",
          2625 => x"f8",
          2626 => x"70",
          2627 => x"f0",
          2628 => x"cc",
          2629 => x"56",
          2630 => x"08",
          2631 => x"7b",
          2632 => x"f6",
          2633 => x"dc",
          2634 => x"dc",
          2635 => x"17",
          2636 => x"80",
          2637 => x"b4",
          2638 => x"57",
          2639 => x"77",
          2640 => x"81",
          2641 => x"15",
          2642 => x"78",
          2643 => x"81",
          2644 => x"53",
          2645 => x"15",
          2646 => x"e9",
          2647 => x"cc",
          2648 => x"df",
          2649 => x"22",
          2650 => x"30",
          2651 => x"70",
          2652 => x"51",
          2653 => x"81",
          2654 => x"8a",
          2655 => x"f8",
          2656 => x"7c",
          2657 => x"56",
          2658 => x"80",
          2659 => x"f1",
          2660 => x"06",
          2661 => x"e9",
          2662 => x"18",
          2663 => x"08",
          2664 => x"38",
          2665 => x"82",
          2666 => x"38",
          2667 => x"54",
          2668 => x"74",
          2669 => x"82",
          2670 => x"22",
          2671 => x"79",
          2672 => x"38",
          2673 => x"98",
          2674 => x"cd",
          2675 => x"22",
          2676 => x"54",
          2677 => x"26",
          2678 => x"52",
          2679 => x"b0",
          2680 => x"cc",
          2681 => x"dc",
          2682 => x"2e",
          2683 => x"0b",
          2684 => x"08",
          2685 => x"98",
          2686 => x"dc",
          2687 => x"85",
          2688 => x"bd",
          2689 => x"31",
          2690 => x"73",
          2691 => x"f4",
          2692 => x"dc",
          2693 => x"18",
          2694 => x"18",
          2695 => x"08",
          2696 => x"72",
          2697 => x"38",
          2698 => x"58",
          2699 => x"89",
          2700 => x"18",
          2701 => x"ff",
          2702 => x"05",
          2703 => x"80",
          2704 => x"dc",
          2705 => x"3d",
          2706 => x"3d",
          2707 => x"08",
          2708 => x"a0",
          2709 => x"54",
          2710 => x"77",
          2711 => x"80",
          2712 => x"0c",
          2713 => x"53",
          2714 => x"80",
          2715 => x"38",
          2716 => x"06",
          2717 => x"b5",
          2718 => x"98",
          2719 => x"14",
          2720 => x"92",
          2721 => x"2a",
          2722 => x"56",
          2723 => x"26",
          2724 => x"80",
          2725 => x"16",
          2726 => x"77",
          2727 => x"53",
          2728 => x"38",
          2729 => x"51",
          2730 => x"81",
          2731 => x"53",
          2732 => x"0b",
          2733 => x"08",
          2734 => x"38",
          2735 => x"dc",
          2736 => x"2e",
          2737 => x"98",
          2738 => x"dc",
          2739 => x"80",
          2740 => x"8a",
          2741 => x"15",
          2742 => x"80",
          2743 => x"14",
          2744 => x"51",
          2745 => x"81",
          2746 => x"53",
          2747 => x"dc",
          2748 => x"2e",
          2749 => x"82",
          2750 => x"cc",
          2751 => x"ba",
          2752 => x"81",
          2753 => x"ff",
          2754 => x"81",
          2755 => x"52",
          2756 => x"f3",
          2757 => x"cc",
          2758 => x"72",
          2759 => x"72",
          2760 => x"f2",
          2761 => x"dc",
          2762 => x"15",
          2763 => x"15",
          2764 => x"b4",
          2765 => x"0c",
          2766 => x"81",
          2767 => x"8a",
          2768 => x"f7",
          2769 => x"7d",
          2770 => x"5b",
          2771 => x"76",
          2772 => x"3f",
          2773 => x"08",
          2774 => x"cc",
          2775 => x"38",
          2776 => x"08",
          2777 => x"08",
          2778 => x"f0",
          2779 => x"dc",
          2780 => x"81",
          2781 => x"80",
          2782 => x"dc",
          2783 => x"18",
          2784 => x"51",
          2785 => x"81",
          2786 => x"81",
          2787 => x"81",
          2788 => x"cc",
          2789 => x"83",
          2790 => x"77",
          2791 => x"72",
          2792 => x"38",
          2793 => x"75",
          2794 => x"81",
          2795 => x"a5",
          2796 => x"cc",
          2797 => x"52",
          2798 => x"8e",
          2799 => x"cc",
          2800 => x"dc",
          2801 => x"2e",
          2802 => x"73",
          2803 => x"81",
          2804 => x"87",
          2805 => x"dc",
          2806 => x"3d",
          2807 => x"3d",
          2808 => x"11",
          2809 => x"ec",
          2810 => x"cc",
          2811 => x"ff",
          2812 => x"33",
          2813 => x"71",
          2814 => x"81",
          2815 => x"94",
          2816 => x"d0",
          2817 => x"cc",
          2818 => x"73",
          2819 => x"81",
          2820 => x"85",
          2821 => x"fc",
          2822 => x"79",
          2823 => x"ff",
          2824 => x"12",
          2825 => x"eb",
          2826 => x"70",
          2827 => x"72",
          2828 => x"81",
          2829 => x"73",
          2830 => x"94",
          2831 => x"d6",
          2832 => x"0d",
          2833 => x"0d",
          2834 => x"55",
          2835 => x"5a",
          2836 => x"08",
          2837 => x"8a",
          2838 => x"08",
          2839 => x"ee",
          2840 => x"dc",
          2841 => x"81",
          2842 => x"80",
          2843 => x"15",
          2844 => x"55",
          2845 => x"38",
          2846 => x"e6",
          2847 => x"33",
          2848 => x"70",
          2849 => x"58",
          2850 => x"86",
          2851 => x"dc",
          2852 => x"73",
          2853 => x"83",
          2854 => x"73",
          2855 => x"38",
          2856 => x"06",
          2857 => x"80",
          2858 => x"75",
          2859 => x"38",
          2860 => x"08",
          2861 => x"54",
          2862 => x"2e",
          2863 => x"83",
          2864 => x"73",
          2865 => x"38",
          2866 => x"51",
          2867 => x"81",
          2868 => x"58",
          2869 => x"08",
          2870 => x"15",
          2871 => x"38",
          2872 => x"0b",
          2873 => x"77",
          2874 => x"0c",
          2875 => x"04",
          2876 => x"77",
          2877 => x"54",
          2878 => x"51",
          2879 => x"81",
          2880 => x"55",
          2881 => x"08",
          2882 => x"14",
          2883 => x"51",
          2884 => x"81",
          2885 => x"55",
          2886 => x"08",
          2887 => x"53",
          2888 => x"08",
          2889 => x"08",
          2890 => x"3f",
          2891 => x"14",
          2892 => x"08",
          2893 => x"3f",
          2894 => x"17",
          2895 => x"dc",
          2896 => x"3d",
          2897 => x"3d",
          2898 => x"08",
          2899 => x"54",
          2900 => x"53",
          2901 => x"81",
          2902 => x"8d",
          2903 => x"08",
          2904 => x"34",
          2905 => x"15",
          2906 => x"0d",
          2907 => x"0d",
          2908 => x"57",
          2909 => x"17",
          2910 => x"08",
          2911 => x"82",
          2912 => x"89",
          2913 => x"55",
          2914 => x"14",
          2915 => x"16",
          2916 => x"71",
          2917 => x"38",
          2918 => x"09",
          2919 => x"38",
          2920 => x"73",
          2921 => x"81",
          2922 => x"ae",
          2923 => x"05",
          2924 => x"15",
          2925 => x"70",
          2926 => x"34",
          2927 => x"8a",
          2928 => x"38",
          2929 => x"05",
          2930 => x"81",
          2931 => x"17",
          2932 => x"12",
          2933 => x"34",
          2934 => x"9c",
          2935 => x"e8",
          2936 => x"dc",
          2937 => x"0c",
          2938 => x"e7",
          2939 => x"dc",
          2940 => x"17",
          2941 => x"51",
          2942 => x"81",
          2943 => x"84",
          2944 => x"3d",
          2945 => x"3d",
          2946 => x"08",
          2947 => x"61",
          2948 => x"55",
          2949 => x"2e",
          2950 => x"55",
          2951 => x"2e",
          2952 => x"80",
          2953 => x"94",
          2954 => x"1c",
          2955 => x"81",
          2956 => x"61",
          2957 => x"56",
          2958 => x"2e",
          2959 => x"83",
          2960 => x"73",
          2961 => x"70",
          2962 => x"25",
          2963 => x"51",
          2964 => x"38",
          2965 => x"0c",
          2966 => x"51",
          2967 => x"26",
          2968 => x"80",
          2969 => x"34",
          2970 => x"51",
          2971 => x"81",
          2972 => x"55",
          2973 => x"91",
          2974 => x"1d",
          2975 => x"8b",
          2976 => x"79",
          2977 => x"3f",
          2978 => x"57",
          2979 => x"55",
          2980 => x"2e",
          2981 => x"80",
          2982 => x"18",
          2983 => x"1a",
          2984 => x"70",
          2985 => x"2a",
          2986 => x"07",
          2987 => x"5a",
          2988 => x"8c",
          2989 => x"54",
          2990 => x"81",
          2991 => x"39",
          2992 => x"70",
          2993 => x"2a",
          2994 => x"75",
          2995 => x"8c",
          2996 => x"2e",
          2997 => x"a0",
          2998 => x"38",
          2999 => x"0c",
          3000 => x"76",
          3001 => x"38",
          3002 => x"b8",
          3003 => x"70",
          3004 => x"5a",
          3005 => x"76",
          3006 => x"38",
          3007 => x"70",
          3008 => x"dc",
          3009 => x"72",
          3010 => x"80",
          3011 => x"51",
          3012 => x"73",
          3013 => x"38",
          3014 => x"18",
          3015 => x"1a",
          3016 => x"55",
          3017 => x"2e",
          3018 => x"83",
          3019 => x"73",
          3020 => x"70",
          3021 => x"25",
          3022 => x"51",
          3023 => x"38",
          3024 => x"75",
          3025 => x"81",
          3026 => x"81",
          3027 => x"27",
          3028 => x"73",
          3029 => x"38",
          3030 => x"70",
          3031 => x"32",
          3032 => x"80",
          3033 => x"2a",
          3034 => x"56",
          3035 => x"81",
          3036 => x"57",
          3037 => x"f5",
          3038 => x"2b",
          3039 => x"25",
          3040 => x"80",
          3041 => x"cc",
          3042 => x"57",
          3043 => x"e6",
          3044 => x"dc",
          3045 => x"2e",
          3046 => x"18",
          3047 => x"1a",
          3048 => x"56",
          3049 => x"3f",
          3050 => x"08",
          3051 => x"e8",
          3052 => x"54",
          3053 => x"80",
          3054 => x"17",
          3055 => x"34",
          3056 => x"11",
          3057 => x"74",
          3058 => x"75",
          3059 => x"bc",
          3060 => x"3f",
          3061 => x"08",
          3062 => x"9f",
          3063 => x"99",
          3064 => x"e0",
          3065 => x"ff",
          3066 => x"79",
          3067 => x"74",
          3068 => x"57",
          3069 => x"77",
          3070 => x"76",
          3071 => x"38",
          3072 => x"73",
          3073 => x"09",
          3074 => x"38",
          3075 => x"84",
          3076 => x"27",
          3077 => x"39",
          3078 => x"f2",
          3079 => x"80",
          3080 => x"54",
          3081 => x"34",
          3082 => x"58",
          3083 => x"f2",
          3084 => x"dc",
          3085 => x"81",
          3086 => x"80",
          3087 => x"1b",
          3088 => x"51",
          3089 => x"81",
          3090 => x"56",
          3091 => x"08",
          3092 => x"9c",
          3093 => x"33",
          3094 => x"80",
          3095 => x"38",
          3096 => x"bf",
          3097 => x"86",
          3098 => x"15",
          3099 => x"2a",
          3100 => x"51",
          3101 => x"92",
          3102 => x"79",
          3103 => x"e4",
          3104 => x"dc",
          3105 => x"2e",
          3106 => x"52",
          3107 => x"ba",
          3108 => x"39",
          3109 => x"33",
          3110 => x"80",
          3111 => x"74",
          3112 => x"81",
          3113 => x"38",
          3114 => x"70",
          3115 => x"82",
          3116 => x"54",
          3117 => x"96",
          3118 => x"06",
          3119 => x"2e",
          3120 => x"ff",
          3121 => x"1c",
          3122 => x"80",
          3123 => x"81",
          3124 => x"ba",
          3125 => x"b6",
          3126 => x"2a",
          3127 => x"51",
          3128 => x"38",
          3129 => x"70",
          3130 => x"81",
          3131 => x"55",
          3132 => x"e1",
          3133 => x"08",
          3134 => x"1d",
          3135 => x"7c",
          3136 => x"3f",
          3137 => x"08",
          3138 => x"fa",
          3139 => x"81",
          3140 => x"8f",
          3141 => x"f6",
          3142 => x"5b",
          3143 => x"70",
          3144 => x"59",
          3145 => x"73",
          3146 => x"c6",
          3147 => x"81",
          3148 => x"70",
          3149 => x"52",
          3150 => x"8d",
          3151 => x"38",
          3152 => x"09",
          3153 => x"a5",
          3154 => x"d0",
          3155 => x"ff",
          3156 => x"53",
          3157 => x"91",
          3158 => x"73",
          3159 => x"d0",
          3160 => x"71",
          3161 => x"f7",
          3162 => x"81",
          3163 => x"55",
          3164 => x"55",
          3165 => x"81",
          3166 => x"74",
          3167 => x"56",
          3168 => x"12",
          3169 => x"70",
          3170 => x"38",
          3171 => x"81",
          3172 => x"51",
          3173 => x"51",
          3174 => x"89",
          3175 => x"70",
          3176 => x"53",
          3177 => x"70",
          3178 => x"51",
          3179 => x"09",
          3180 => x"38",
          3181 => x"38",
          3182 => x"77",
          3183 => x"70",
          3184 => x"2a",
          3185 => x"07",
          3186 => x"51",
          3187 => x"8f",
          3188 => x"84",
          3189 => x"83",
          3190 => x"94",
          3191 => x"74",
          3192 => x"38",
          3193 => x"0c",
          3194 => x"86",
          3195 => x"fc",
          3196 => x"81",
          3197 => x"8c",
          3198 => x"fa",
          3199 => x"56",
          3200 => x"17",
          3201 => x"b0",
          3202 => x"52",
          3203 => x"e0",
          3204 => x"81",
          3205 => x"81",
          3206 => x"b2",
          3207 => x"b4",
          3208 => x"cc",
          3209 => x"ff",
          3210 => x"55",
          3211 => x"d5",
          3212 => x"06",
          3213 => x"80",
          3214 => x"33",
          3215 => x"81",
          3216 => x"81",
          3217 => x"81",
          3218 => x"eb",
          3219 => x"70",
          3220 => x"07",
          3221 => x"73",
          3222 => x"81",
          3223 => x"81",
          3224 => x"83",
          3225 => x"cc",
          3226 => x"16",
          3227 => x"3f",
          3228 => x"08",
          3229 => x"cc",
          3230 => x"9d",
          3231 => x"81",
          3232 => x"81",
          3233 => x"e0",
          3234 => x"dc",
          3235 => x"81",
          3236 => x"80",
          3237 => x"82",
          3238 => x"dc",
          3239 => x"3d",
          3240 => x"3d",
          3241 => x"84",
          3242 => x"05",
          3243 => x"80",
          3244 => x"51",
          3245 => x"81",
          3246 => x"58",
          3247 => x"0b",
          3248 => x"08",
          3249 => x"38",
          3250 => x"08",
          3251 => x"dc",
          3252 => x"08",
          3253 => x"56",
          3254 => x"86",
          3255 => x"75",
          3256 => x"fe",
          3257 => x"54",
          3258 => x"2e",
          3259 => x"14",
          3260 => x"ca",
          3261 => x"cc",
          3262 => x"06",
          3263 => x"54",
          3264 => x"38",
          3265 => x"86",
          3266 => x"82",
          3267 => x"06",
          3268 => x"56",
          3269 => x"38",
          3270 => x"80",
          3271 => x"81",
          3272 => x"52",
          3273 => x"51",
          3274 => x"81",
          3275 => x"81",
          3276 => x"81",
          3277 => x"83",
          3278 => x"87",
          3279 => x"2e",
          3280 => x"82",
          3281 => x"06",
          3282 => x"56",
          3283 => x"38",
          3284 => x"74",
          3285 => x"a3",
          3286 => x"cc",
          3287 => x"06",
          3288 => x"2e",
          3289 => x"80",
          3290 => x"3d",
          3291 => x"83",
          3292 => x"15",
          3293 => x"53",
          3294 => x"8d",
          3295 => x"15",
          3296 => x"3f",
          3297 => x"08",
          3298 => x"70",
          3299 => x"0c",
          3300 => x"16",
          3301 => x"80",
          3302 => x"80",
          3303 => x"54",
          3304 => x"84",
          3305 => x"5b",
          3306 => x"80",
          3307 => x"7a",
          3308 => x"fc",
          3309 => x"dc",
          3310 => x"ff",
          3311 => x"77",
          3312 => x"81",
          3313 => x"76",
          3314 => x"81",
          3315 => x"2e",
          3316 => x"8d",
          3317 => x"26",
          3318 => x"bf",
          3319 => x"f4",
          3320 => x"cc",
          3321 => x"ff",
          3322 => x"84",
          3323 => x"81",
          3324 => x"38",
          3325 => x"51",
          3326 => x"81",
          3327 => x"83",
          3328 => x"58",
          3329 => x"80",
          3330 => x"db",
          3331 => x"dc",
          3332 => x"77",
          3333 => x"80",
          3334 => x"82",
          3335 => x"c4",
          3336 => x"11",
          3337 => x"06",
          3338 => x"8d",
          3339 => x"26",
          3340 => x"74",
          3341 => x"78",
          3342 => x"c1",
          3343 => x"59",
          3344 => x"15",
          3345 => x"2e",
          3346 => x"13",
          3347 => x"72",
          3348 => x"38",
          3349 => x"eb",
          3350 => x"14",
          3351 => x"3f",
          3352 => x"08",
          3353 => x"cc",
          3354 => x"23",
          3355 => x"57",
          3356 => x"83",
          3357 => x"c7",
          3358 => x"d8",
          3359 => x"cc",
          3360 => x"ff",
          3361 => x"8d",
          3362 => x"14",
          3363 => x"3f",
          3364 => x"08",
          3365 => x"14",
          3366 => x"3f",
          3367 => x"08",
          3368 => x"06",
          3369 => x"72",
          3370 => x"97",
          3371 => x"22",
          3372 => x"84",
          3373 => x"5a",
          3374 => x"83",
          3375 => x"14",
          3376 => x"79",
          3377 => x"ad",
          3378 => x"dc",
          3379 => x"81",
          3380 => x"80",
          3381 => x"38",
          3382 => x"08",
          3383 => x"ff",
          3384 => x"38",
          3385 => x"83",
          3386 => x"83",
          3387 => x"74",
          3388 => x"85",
          3389 => x"89",
          3390 => x"76",
          3391 => x"c3",
          3392 => x"70",
          3393 => x"7b",
          3394 => x"73",
          3395 => x"17",
          3396 => x"ac",
          3397 => x"55",
          3398 => x"09",
          3399 => x"38",
          3400 => x"51",
          3401 => x"81",
          3402 => x"83",
          3403 => x"53",
          3404 => x"82",
          3405 => x"82",
          3406 => x"e0",
          3407 => x"ab",
          3408 => x"cc",
          3409 => x"0c",
          3410 => x"53",
          3411 => x"56",
          3412 => x"81",
          3413 => x"13",
          3414 => x"74",
          3415 => x"82",
          3416 => x"74",
          3417 => x"81",
          3418 => x"06",
          3419 => x"83",
          3420 => x"2a",
          3421 => x"72",
          3422 => x"26",
          3423 => x"ff",
          3424 => x"0c",
          3425 => x"15",
          3426 => x"0b",
          3427 => x"76",
          3428 => x"81",
          3429 => x"38",
          3430 => x"51",
          3431 => x"81",
          3432 => x"83",
          3433 => x"53",
          3434 => x"09",
          3435 => x"f9",
          3436 => x"52",
          3437 => x"b8",
          3438 => x"cc",
          3439 => x"38",
          3440 => x"08",
          3441 => x"84",
          3442 => x"d8",
          3443 => x"dc",
          3444 => x"ff",
          3445 => x"72",
          3446 => x"2e",
          3447 => x"80",
          3448 => x"14",
          3449 => x"3f",
          3450 => x"08",
          3451 => x"a4",
          3452 => x"81",
          3453 => x"84",
          3454 => x"d7",
          3455 => x"dc",
          3456 => x"8a",
          3457 => x"2e",
          3458 => x"9d",
          3459 => x"14",
          3460 => x"3f",
          3461 => x"08",
          3462 => x"84",
          3463 => x"d7",
          3464 => x"dc",
          3465 => x"15",
          3466 => x"34",
          3467 => x"22",
          3468 => x"72",
          3469 => x"23",
          3470 => x"23",
          3471 => x"15",
          3472 => x"75",
          3473 => x"0c",
          3474 => x"04",
          3475 => x"77",
          3476 => x"73",
          3477 => x"38",
          3478 => x"72",
          3479 => x"38",
          3480 => x"71",
          3481 => x"38",
          3482 => x"84",
          3483 => x"52",
          3484 => x"09",
          3485 => x"38",
          3486 => x"51",
          3487 => x"81",
          3488 => x"81",
          3489 => x"88",
          3490 => x"08",
          3491 => x"39",
          3492 => x"73",
          3493 => x"74",
          3494 => x"0c",
          3495 => x"04",
          3496 => x"02",
          3497 => x"7a",
          3498 => x"fc",
          3499 => x"f4",
          3500 => x"54",
          3501 => x"dc",
          3502 => x"bc",
          3503 => x"cc",
          3504 => x"81",
          3505 => x"70",
          3506 => x"73",
          3507 => x"38",
          3508 => x"78",
          3509 => x"2e",
          3510 => x"74",
          3511 => x"0c",
          3512 => x"80",
          3513 => x"80",
          3514 => x"70",
          3515 => x"51",
          3516 => x"81",
          3517 => x"54",
          3518 => x"cc",
          3519 => x"0d",
          3520 => x"0d",
          3521 => x"05",
          3522 => x"33",
          3523 => x"54",
          3524 => x"84",
          3525 => x"bf",
          3526 => x"98",
          3527 => x"53",
          3528 => x"05",
          3529 => x"fa",
          3530 => x"cc",
          3531 => x"dc",
          3532 => x"a4",
          3533 => x"68",
          3534 => x"70",
          3535 => x"c6",
          3536 => x"cc",
          3537 => x"dc",
          3538 => x"38",
          3539 => x"05",
          3540 => x"2b",
          3541 => x"80",
          3542 => x"86",
          3543 => x"06",
          3544 => x"2e",
          3545 => x"74",
          3546 => x"38",
          3547 => x"09",
          3548 => x"38",
          3549 => x"f8",
          3550 => x"cc",
          3551 => x"39",
          3552 => x"33",
          3553 => x"73",
          3554 => x"77",
          3555 => x"81",
          3556 => x"73",
          3557 => x"38",
          3558 => x"bc",
          3559 => x"07",
          3560 => x"b4",
          3561 => x"2a",
          3562 => x"51",
          3563 => x"2e",
          3564 => x"62",
          3565 => x"e8",
          3566 => x"dc",
          3567 => x"82",
          3568 => x"52",
          3569 => x"51",
          3570 => x"62",
          3571 => x"8b",
          3572 => x"53",
          3573 => x"51",
          3574 => x"80",
          3575 => x"05",
          3576 => x"3f",
          3577 => x"0b",
          3578 => x"75",
          3579 => x"f1",
          3580 => x"11",
          3581 => x"80",
          3582 => x"97",
          3583 => x"51",
          3584 => x"81",
          3585 => x"55",
          3586 => x"08",
          3587 => x"b7",
          3588 => x"c4",
          3589 => x"05",
          3590 => x"2a",
          3591 => x"51",
          3592 => x"80",
          3593 => x"84",
          3594 => x"39",
          3595 => x"70",
          3596 => x"54",
          3597 => x"a9",
          3598 => x"06",
          3599 => x"2e",
          3600 => x"55",
          3601 => x"73",
          3602 => x"d6",
          3603 => x"dc",
          3604 => x"ff",
          3605 => x"0c",
          3606 => x"dc",
          3607 => x"f8",
          3608 => x"2a",
          3609 => x"51",
          3610 => x"2e",
          3611 => x"80",
          3612 => x"7a",
          3613 => x"a0",
          3614 => x"a4",
          3615 => x"53",
          3616 => x"e6",
          3617 => x"dc",
          3618 => x"dc",
          3619 => x"1b",
          3620 => x"05",
          3621 => x"d3",
          3622 => x"cc",
          3623 => x"cc",
          3624 => x"0c",
          3625 => x"56",
          3626 => x"84",
          3627 => x"90",
          3628 => x"0b",
          3629 => x"80",
          3630 => x"0c",
          3631 => x"1a",
          3632 => x"2a",
          3633 => x"51",
          3634 => x"2e",
          3635 => x"81",
          3636 => x"80",
          3637 => x"38",
          3638 => x"08",
          3639 => x"8a",
          3640 => x"89",
          3641 => x"59",
          3642 => x"76",
          3643 => x"d7",
          3644 => x"dc",
          3645 => x"81",
          3646 => x"81",
          3647 => x"82",
          3648 => x"cc",
          3649 => x"09",
          3650 => x"38",
          3651 => x"78",
          3652 => x"30",
          3653 => x"80",
          3654 => x"77",
          3655 => x"38",
          3656 => x"06",
          3657 => x"c3",
          3658 => x"1a",
          3659 => x"38",
          3660 => x"06",
          3661 => x"2e",
          3662 => x"52",
          3663 => x"a6",
          3664 => x"cc",
          3665 => x"82",
          3666 => x"75",
          3667 => x"dc",
          3668 => x"9c",
          3669 => x"39",
          3670 => x"74",
          3671 => x"dc",
          3672 => x"3d",
          3673 => x"3d",
          3674 => x"65",
          3675 => x"5d",
          3676 => x"0c",
          3677 => x"05",
          3678 => x"f9",
          3679 => x"dc",
          3680 => x"81",
          3681 => x"8a",
          3682 => x"33",
          3683 => x"2e",
          3684 => x"56",
          3685 => x"90",
          3686 => x"06",
          3687 => x"74",
          3688 => x"b6",
          3689 => x"82",
          3690 => x"34",
          3691 => x"aa",
          3692 => x"91",
          3693 => x"56",
          3694 => x"8c",
          3695 => x"1a",
          3696 => x"74",
          3697 => x"38",
          3698 => x"80",
          3699 => x"38",
          3700 => x"70",
          3701 => x"56",
          3702 => x"b2",
          3703 => x"11",
          3704 => x"77",
          3705 => x"5b",
          3706 => x"38",
          3707 => x"88",
          3708 => x"8f",
          3709 => x"08",
          3710 => x"d5",
          3711 => x"dc",
          3712 => x"81",
          3713 => x"9f",
          3714 => x"2e",
          3715 => x"74",
          3716 => x"98",
          3717 => x"7e",
          3718 => x"3f",
          3719 => x"08",
          3720 => x"83",
          3721 => x"cc",
          3722 => x"89",
          3723 => x"77",
          3724 => x"d6",
          3725 => x"7f",
          3726 => x"58",
          3727 => x"75",
          3728 => x"75",
          3729 => x"77",
          3730 => x"7c",
          3731 => x"33",
          3732 => x"3f",
          3733 => x"08",
          3734 => x"7e",
          3735 => x"56",
          3736 => x"2e",
          3737 => x"16",
          3738 => x"55",
          3739 => x"94",
          3740 => x"53",
          3741 => x"b0",
          3742 => x"31",
          3743 => x"05",
          3744 => x"3f",
          3745 => x"56",
          3746 => x"9c",
          3747 => x"19",
          3748 => x"06",
          3749 => x"31",
          3750 => x"76",
          3751 => x"7b",
          3752 => x"08",
          3753 => x"d1",
          3754 => x"dc",
          3755 => x"81",
          3756 => x"94",
          3757 => x"ff",
          3758 => x"05",
          3759 => x"cf",
          3760 => x"76",
          3761 => x"17",
          3762 => x"1e",
          3763 => x"18",
          3764 => x"5e",
          3765 => x"39",
          3766 => x"81",
          3767 => x"90",
          3768 => x"f2",
          3769 => x"63",
          3770 => x"40",
          3771 => x"7e",
          3772 => x"fc",
          3773 => x"51",
          3774 => x"81",
          3775 => x"55",
          3776 => x"08",
          3777 => x"18",
          3778 => x"80",
          3779 => x"74",
          3780 => x"39",
          3781 => x"70",
          3782 => x"81",
          3783 => x"56",
          3784 => x"80",
          3785 => x"38",
          3786 => x"0b",
          3787 => x"82",
          3788 => x"39",
          3789 => x"19",
          3790 => x"83",
          3791 => x"18",
          3792 => x"56",
          3793 => x"27",
          3794 => x"09",
          3795 => x"2e",
          3796 => x"94",
          3797 => x"83",
          3798 => x"56",
          3799 => x"38",
          3800 => x"22",
          3801 => x"89",
          3802 => x"55",
          3803 => x"75",
          3804 => x"18",
          3805 => x"9c",
          3806 => x"85",
          3807 => x"08",
          3808 => x"d7",
          3809 => x"dc",
          3810 => x"81",
          3811 => x"80",
          3812 => x"38",
          3813 => x"ff",
          3814 => x"ff",
          3815 => x"38",
          3816 => x"0c",
          3817 => x"85",
          3818 => x"19",
          3819 => x"b0",
          3820 => x"19",
          3821 => x"81",
          3822 => x"74",
          3823 => x"3f",
          3824 => x"08",
          3825 => x"98",
          3826 => x"7e",
          3827 => x"3f",
          3828 => x"08",
          3829 => x"d2",
          3830 => x"cc",
          3831 => x"89",
          3832 => x"78",
          3833 => x"d5",
          3834 => x"7f",
          3835 => x"58",
          3836 => x"75",
          3837 => x"75",
          3838 => x"78",
          3839 => x"7c",
          3840 => x"33",
          3841 => x"3f",
          3842 => x"08",
          3843 => x"7e",
          3844 => x"78",
          3845 => x"74",
          3846 => x"38",
          3847 => x"b0",
          3848 => x"31",
          3849 => x"05",
          3850 => x"51",
          3851 => x"7e",
          3852 => x"83",
          3853 => x"89",
          3854 => x"db",
          3855 => x"08",
          3856 => x"26",
          3857 => x"51",
          3858 => x"81",
          3859 => x"fd",
          3860 => x"77",
          3861 => x"55",
          3862 => x"0c",
          3863 => x"83",
          3864 => x"80",
          3865 => x"55",
          3866 => x"83",
          3867 => x"9c",
          3868 => x"7e",
          3869 => x"3f",
          3870 => x"08",
          3871 => x"75",
          3872 => x"94",
          3873 => x"ff",
          3874 => x"05",
          3875 => x"3f",
          3876 => x"0b",
          3877 => x"7b",
          3878 => x"08",
          3879 => x"76",
          3880 => x"08",
          3881 => x"1c",
          3882 => x"08",
          3883 => x"5c",
          3884 => x"83",
          3885 => x"74",
          3886 => x"fd",
          3887 => x"18",
          3888 => x"07",
          3889 => x"19",
          3890 => x"75",
          3891 => x"0c",
          3892 => x"04",
          3893 => x"7a",
          3894 => x"05",
          3895 => x"56",
          3896 => x"81",
          3897 => x"57",
          3898 => x"08",
          3899 => x"90",
          3900 => x"86",
          3901 => x"06",
          3902 => x"73",
          3903 => x"e9",
          3904 => x"08",
          3905 => x"cc",
          3906 => x"dc",
          3907 => x"81",
          3908 => x"80",
          3909 => x"16",
          3910 => x"33",
          3911 => x"55",
          3912 => x"34",
          3913 => x"53",
          3914 => x"08",
          3915 => x"3f",
          3916 => x"52",
          3917 => x"c9",
          3918 => x"88",
          3919 => x"96",
          3920 => x"f0",
          3921 => x"92",
          3922 => x"ca",
          3923 => x"81",
          3924 => x"34",
          3925 => x"df",
          3926 => x"cc",
          3927 => x"33",
          3928 => x"55",
          3929 => x"17",
          3930 => x"dc",
          3931 => x"3d",
          3932 => x"3d",
          3933 => x"52",
          3934 => x"3f",
          3935 => x"08",
          3936 => x"cc",
          3937 => x"86",
          3938 => x"52",
          3939 => x"bc",
          3940 => x"cc",
          3941 => x"dc",
          3942 => x"38",
          3943 => x"08",
          3944 => x"81",
          3945 => x"86",
          3946 => x"ff",
          3947 => x"3d",
          3948 => x"3f",
          3949 => x"0b",
          3950 => x"08",
          3951 => x"81",
          3952 => x"81",
          3953 => x"80",
          3954 => x"dc",
          3955 => x"3d",
          3956 => x"3d",
          3957 => x"93",
          3958 => x"52",
          3959 => x"e9",
          3960 => x"dc",
          3961 => x"81",
          3962 => x"80",
          3963 => x"58",
          3964 => x"3d",
          3965 => x"e0",
          3966 => x"dc",
          3967 => x"81",
          3968 => x"bc",
          3969 => x"c7",
          3970 => x"98",
          3971 => x"73",
          3972 => x"38",
          3973 => x"12",
          3974 => x"39",
          3975 => x"33",
          3976 => x"70",
          3977 => x"55",
          3978 => x"2e",
          3979 => x"7f",
          3980 => x"54",
          3981 => x"81",
          3982 => x"94",
          3983 => x"39",
          3984 => x"08",
          3985 => x"81",
          3986 => x"85",
          3987 => x"dc",
          3988 => x"3d",
          3989 => x"3d",
          3990 => x"5b",
          3991 => x"34",
          3992 => x"3d",
          3993 => x"52",
          3994 => x"e8",
          3995 => x"dc",
          3996 => x"81",
          3997 => x"82",
          3998 => x"43",
          3999 => x"11",
          4000 => x"58",
          4001 => x"80",
          4002 => x"38",
          4003 => x"3d",
          4004 => x"d5",
          4005 => x"dc",
          4006 => x"81",
          4007 => x"82",
          4008 => x"52",
          4009 => x"c8",
          4010 => x"cc",
          4011 => x"dc",
          4012 => x"c1",
          4013 => x"7b",
          4014 => x"3f",
          4015 => x"08",
          4016 => x"74",
          4017 => x"3f",
          4018 => x"08",
          4019 => x"cc",
          4020 => x"38",
          4021 => x"51",
          4022 => x"81",
          4023 => x"57",
          4024 => x"08",
          4025 => x"52",
          4026 => x"f2",
          4027 => x"dc",
          4028 => x"a6",
          4029 => x"74",
          4030 => x"3f",
          4031 => x"08",
          4032 => x"cc",
          4033 => x"cc",
          4034 => x"2e",
          4035 => x"86",
          4036 => x"81",
          4037 => x"81",
          4038 => x"3d",
          4039 => x"52",
          4040 => x"c9",
          4041 => x"3d",
          4042 => x"11",
          4043 => x"5a",
          4044 => x"2e",
          4045 => x"b9",
          4046 => x"16",
          4047 => x"33",
          4048 => x"73",
          4049 => x"16",
          4050 => x"26",
          4051 => x"75",
          4052 => x"38",
          4053 => x"05",
          4054 => x"6f",
          4055 => x"ff",
          4056 => x"55",
          4057 => x"74",
          4058 => x"38",
          4059 => x"11",
          4060 => x"74",
          4061 => x"39",
          4062 => x"09",
          4063 => x"38",
          4064 => x"11",
          4065 => x"74",
          4066 => x"81",
          4067 => x"70",
          4068 => x"cc",
          4069 => x"08",
          4070 => x"5c",
          4071 => x"73",
          4072 => x"38",
          4073 => x"1a",
          4074 => x"55",
          4075 => x"38",
          4076 => x"73",
          4077 => x"38",
          4078 => x"76",
          4079 => x"74",
          4080 => x"33",
          4081 => x"05",
          4082 => x"15",
          4083 => x"ba",
          4084 => x"05",
          4085 => x"ff",
          4086 => x"06",
          4087 => x"57",
          4088 => x"18",
          4089 => x"54",
          4090 => x"70",
          4091 => x"34",
          4092 => x"ee",
          4093 => x"34",
          4094 => x"cc",
          4095 => x"0d",
          4096 => x"0d",
          4097 => x"3d",
          4098 => x"71",
          4099 => x"ec",
          4100 => x"dc",
          4101 => x"81",
          4102 => x"82",
          4103 => x"15",
          4104 => x"82",
          4105 => x"15",
          4106 => x"76",
          4107 => x"90",
          4108 => x"81",
          4109 => x"06",
          4110 => x"72",
          4111 => x"56",
          4112 => x"54",
          4113 => x"17",
          4114 => x"78",
          4115 => x"38",
          4116 => x"22",
          4117 => x"59",
          4118 => x"78",
          4119 => x"76",
          4120 => x"51",
          4121 => x"3f",
          4122 => x"08",
          4123 => x"54",
          4124 => x"53",
          4125 => x"3f",
          4126 => x"08",
          4127 => x"38",
          4128 => x"75",
          4129 => x"18",
          4130 => x"31",
          4131 => x"57",
          4132 => x"b1",
          4133 => x"08",
          4134 => x"38",
          4135 => x"51",
          4136 => x"81",
          4137 => x"54",
          4138 => x"08",
          4139 => x"9a",
          4140 => x"cc",
          4141 => x"81",
          4142 => x"dc",
          4143 => x"16",
          4144 => x"16",
          4145 => x"2e",
          4146 => x"76",
          4147 => x"dc",
          4148 => x"31",
          4149 => x"18",
          4150 => x"90",
          4151 => x"81",
          4152 => x"06",
          4153 => x"56",
          4154 => x"9a",
          4155 => x"74",
          4156 => x"3f",
          4157 => x"08",
          4158 => x"cc",
          4159 => x"81",
          4160 => x"56",
          4161 => x"52",
          4162 => x"84",
          4163 => x"cc",
          4164 => x"ff",
          4165 => x"81",
          4166 => x"38",
          4167 => x"98",
          4168 => x"a6",
          4169 => x"16",
          4170 => x"39",
          4171 => x"16",
          4172 => x"75",
          4173 => x"53",
          4174 => x"aa",
          4175 => x"79",
          4176 => x"3f",
          4177 => x"08",
          4178 => x"0b",
          4179 => x"82",
          4180 => x"39",
          4181 => x"16",
          4182 => x"bb",
          4183 => x"2a",
          4184 => x"08",
          4185 => x"15",
          4186 => x"15",
          4187 => x"90",
          4188 => x"16",
          4189 => x"33",
          4190 => x"53",
          4191 => x"34",
          4192 => x"06",
          4193 => x"2e",
          4194 => x"9c",
          4195 => x"85",
          4196 => x"16",
          4197 => x"72",
          4198 => x"0c",
          4199 => x"04",
          4200 => x"79",
          4201 => x"75",
          4202 => x"8a",
          4203 => x"89",
          4204 => x"52",
          4205 => x"05",
          4206 => x"3f",
          4207 => x"08",
          4208 => x"cc",
          4209 => x"38",
          4210 => x"7a",
          4211 => x"d8",
          4212 => x"dc",
          4213 => x"81",
          4214 => x"80",
          4215 => x"16",
          4216 => x"2b",
          4217 => x"74",
          4218 => x"86",
          4219 => x"84",
          4220 => x"06",
          4221 => x"73",
          4222 => x"38",
          4223 => x"52",
          4224 => x"da",
          4225 => x"cc",
          4226 => x"0c",
          4227 => x"14",
          4228 => x"23",
          4229 => x"51",
          4230 => x"81",
          4231 => x"55",
          4232 => x"09",
          4233 => x"38",
          4234 => x"39",
          4235 => x"84",
          4236 => x"0c",
          4237 => x"81",
          4238 => x"89",
          4239 => x"fc",
          4240 => x"87",
          4241 => x"53",
          4242 => x"e7",
          4243 => x"dc",
          4244 => x"38",
          4245 => x"08",
          4246 => x"3d",
          4247 => x"3d",
          4248 => x"89",
          4249 => x"54",
          4250 => x"54",
          4251 => x"81",
          4252 => x"53",
          4253 => x"08",
          4254 => x"74",
          4255 => x"dc",
          4256 => x"73",
          4257 => x"3f",
          4258 => x"08",
          4259 => x"39",
          4260 => x"08",
          4261 => x"d3",
          4262 => x"dc",
          4263 => x"81",
          4264 => x"84",
          4265 => x"06",
          4266 => x"53",
          4267 => x"dc",
          4268 => x"38",
          4269 => x"51",
          4270 => x"72",
          4271 => x"cf",
          4272 => x"dc",
          4273 => x"32",
          4274 => x"72",
          4275 => x"70",
          4276 => x"08",
          4277 => x"54",
          4278 => x"dc",
          4279 => x"3d",
          4280 => x"3d",
          4281 => x"80",
          4282 => x"70",
          4283 => x"52",
          4284 => x"3f",
          4285 => x"08",
          4286 => x"cc",
          4287 => x"64",
          4288 => x"d6",
          4289 => x"dc",
          4290 => x"81",
          4291 => x"a0",
          4292 => x"cb",
          4293 => x"98",
          4294 => x"73",
          4295 => x"38",
          4296 => x"39",
          4297 => x"88",
          4298 => x"75",
          4299 => x"3f",
          4300 => x"cc",
          4301 => x"0d",
          4302 => x"0d",
          4303 => x"5c",
          4304 => x"3d",
          4305 => x"93",
          4306 => x"d6",
          4307 => x"cc",
          4308 => x"dc",
          4309 => x"80",
          4310 => x"0c",
          4311 => x"11",
          4312 => x"90",
          4313 => x"56",
          4314 => x"74",
          4315 => x"75",
          4316 => x"e4",
          4317 => x"81",
          4318 => x"5b",
          4319 => x"81",
          4320 => x"75",
          4321 => x"73",
          4322 => x"81",
          4323 => x"82",
          4324 => x"76",
          4325 => x"f0",
          4326 => x"f4",
          4327 => x"cc",
          4328 => x"d1",
          4329 => x"cc",
          4330 => x"ce",
          4331 => x"cc",
          4332 => x"81",
          4333 => x"07",
          4334 => x"05",
          4335 => x"53",
          4336 => x"98",
          4337 => x"26",
          4338 => x"f9",
          4339 => x"08",
          4340 => x"08",
          4341 => x"98",
          4342 => x"81",
          4343 => x"58",
          4344 => x"3f",
          4345 => x"08",
          4346 => x"cc",
          4347 => x"38",
          4348 => x"77",
          4349 => x"5d",
          4350 => x"74",
          4351 => x"81",
          4352 => x"b4",
          4353 => x"bb",
          4354 => x"dc",
          4355 => x"ff",
          4356 => x"30",
          4357 => x"1b",
          4358 => x"5b",
          4359 => x"39",
          4360 => x"ff",
          4361 => x"81",
          4362 => x"f0",
          4363 => x"30",
          4364 => x"1b",
          4365 => x"5b",
          4366 => x"83",
          4367 => x"58",
          4368 => x"92",
          4369 => x"0c",
          4370 => x"12",
          4371 => x"33",
          4372 => x"54",
          4373 => x"34",
          4374 => x"cc",
          4375 => x"0d",
          4376 => x"0d",
          4377 => x"fc",
          4378 => x"52",
          4379 => x"3f",
          4380 => x"08",
          4381 => x"cc",
          4382 => x"38",
          4383 => x"56",
          4384 => x"38",
          4385 => x"70",
          4386 => x"81",
          4387 => x"55",
          4388 => x"80",
          4389 => x"38",
          4390 => x"54",
          4391 => x"08",
          4392 => x"38",
          4393 => x"81",
          4394 => x"53",
          4395 => x"52",
          4396 => x"8c",
          4397 => x"cc",
          4398 => x"19",
          4399 => x"c9",
          4400 => x"08",
          4401 => x"ff",
          4402 => x"81",
          4403 => x"ff",
          4404 => x"06",
          4405 => x"56",
          4406 => x"08",
          4407 => x"81",
          4408 => x"82",
          4409 => x"75",
          4410 => x"54",
          4411 => x"08",
          4412 => x"27",
          4413 => x"17",
          4414 => x"dc",
          4415 => x"76",
          4416 => x"3f",
          4417 => x"08",
          4418 => x"08",
          4419 => x"90",
          4420 => x"c0",
          4421 => x"90",
          4422 => x"80",
          4423 => x"75",
          4424 => x"75",
          4425 => x"dc",
          4426 => x"3d",
          4427 => x"3d",
          4428 => x"a0",
          4429 => x"05",
          4430 => x"51",
          4431 => x"81",
          4432 => x"55",
          4433 => x"08",
          4434 => x"78",
          4435 => x"08",
          4436 => x"70",
          4437 => x"ae",
          4438 => x"cc",
          4439 => x"dc",
          4440 => x"db",
          4441 => x"fb",
          4442 => x"85",
          4443 => x"06",
          4444 => x"86",
          4445 => x"c7",
          4446 => x"2b",
          4447 => x"24",
          4448 => x"02",
          4449 => x"33",
          4450 => x"58",
          4451 => x"76",
          4452 => x"6b",
          4453 => x"cc",
          4454 => x"dc",
          4455 => x"84",
          4456 => x"06",
          4457 => x"73",
          4458 => x"d4",
          4459 => x"81",
          4460 => x"94",
          4461 => x"81",
          4462 => x"5a",
          4463 => x"08",
          4464 => x"8a",
          4465 => x"54",
          4466 => x"81",
          4467 => x"55",
          4468 => x"08",
          4469 => x"81",
          4470 => x"52",
          4471 => x"e5",
          4472 => x"cc",
          4473 => x"dc",
          4474 => x"38",
          4475 => x"cf",
          4476 => x"cc",
          4477 => x"88",
          4478 => x"cc",
          4479 => x"38",
          4480 => x"c2",
          4481 => x"cc",
          4482 => x"cc",
          4483 => x"81",
          4484 => x"07",
          4485 => x"55",
          4486 => x"2e",
          4487 => x"80",
          4488 => x"80",
          4489 => x"77",
          4490 => x"3f",
          4491 => x"08",
          4492 => x"38",
          4493 => x"ba",
          4494 => x"dc",
          4495 => x"74",
          4496 => x"0c",
          4497 => x"04",
          4498 => x"82",
          4499 => x"c0",
          4500 => x"3d",
          4501 => x"3f",
          4502 => x"08",
          4503 => x"cc",
          4504 => x"38",
          4505 => x"52",
          4506 => x"52",
          4507 => x"3f",
          4508 => x"08",
          4509 => x"cc",
          4510 => x"88",
          4511 => x"39",
          4512 => x"08",
          4513 => x"81",
          4514 => x"38",
          4515 => x"05",
          4516 => x"2a",
          4517 => x"55",
          4518 => x"81",
          4519 => x"5a",
          4520 => x"3d",
          4521 => x"c1",
          4522 => x"dc",
          4523 => x"55",
          4524 => x"cc",
          4525 => x"87",
          4526 => x"cc",
          4527 => x"09",
          4528 => x"38",
          4529 => x"dc",
          4530 => x"2e",
          4531 => x"86",
          4532 => x"81",
          4533 => x"81",
          4534 => x"dc",
          4535 => x"78",
          4536 => x"3f",
          4537 => x"08",
          4538 => x"cc",
          4539 => x"38",
          4540 => x"52",
          4541 => x"ff",
          4542 => x"78",
          4543 => x"b4",
          4544 => x"54",
          4545 => x"15",
          4546 => x"b2",
          4547 => x"ca",
          4548 => x"b6",
          4549 => x"53",
          4550 => x"53",
          4551 => x"3f",
          4552 => x"b4",
          4553 => x"d4",
          4554 => x"b6",
          4555 => x"54",
          4556 => x"d5",
          4557 => x"53",
          4558 => x"11",
          4559 => x"d7",
          4560 => x"81",
          4561 => x"34",
          4562 => x"a4",
          4563 => x"cc",
          4564 => x"dc",
          4565 => x"38",
          4566 => x"0a",
          4567 => x"05",
          4568 => x"d0",
          4569 => x"64",
          4570 => x"c9",
          4571 => x"54",
          4572 => x"15",
          4573 => x"81",
          4574 => x"34",
          4575 => x"b8",
          4576 => x"dc",
          4577 => x"8b",
          4578 => x"75",
          4579 => x"ff",
          4580 => x"73",
          4581 => x"0c",
          4582 => x"04",
          4583 => x"a9",
          4584 => x"51",
          4585 => x"82",
          4586 => x"ff",
          4587 => x"a9",
          4588 => x"ee",
          4589 => x"cc",
          4590 => x"dc",
          4591 => x"d3",
          4592 => x"a9",
          4593 => x"9d",
          4594 => x"58",
          4595 => x"81",
          4596 => x"55",
          4597 => x"08",
          4598 => x"02",
          4599 => x"33",
          4600 => x"54",
          4601 => x"82",
          4602 => x"53",
          4603 => x"52",
          4604 => x"88",
          4605 => x"b4",
          4606 => x"53",
          4607 => x"3d",
          4608 => x"ff",
          4609 => x"aa",
          4610 => x"73",
          4611 => x"3f",
          4612 => x"08",
          4613 => x"cc",
          4614 => x"63",
          4615 => x"81",
          4616 => x"65",
          4617 => x"2e",
          4618 => x"55",
          4619 => x"81",
          4620 => x"84",
          4621 => x"06",
          4622 => x"73",
          4623 => x"3f",
          4624 => x"08",
          4625 => x"cc",
          4626 => x"38",
          4627 => x"53",
          4628 => x"95",
          4629 => x"16",
          4630 => x"87",
          4631 => x"05",
          4632 => x"34",
          4633 => x"70",
          4634 => x"81",
          4635 => x"55",
          4636 => x"74",
          4637 => x"73",
          4638 => x"78",
          4639 => x"83",
          4640 => x"16",
          4641 => x"2a",
          4642 => x"51",
          4643 => x"80",
          4644 => x"38",
          4645 => x"80",
          4646 => x"52",
          4647 => x"be",
          4648 => x"cc",
          4649 => x"51",
          4650 => x"3f",
          4651 => x"dc",
          4652 => x"2e",
          4653 => x"81",
          4654 => x"52",
          4655 => x"b5",
          4656 => x"dc",
          4657 => x"80",
          4658 => x"58",
          4659 => x"cc",
          4660 => x"38",
          4661 => x"54",
          4662 => x"09",
          4663 => x"38",
          4664 => x"52",
          4665 => x"af",
          4666 => x"81",
          4667 => x"34",
          4668 => x"dc",
          4669 => x"38",
          4670 => x"ca",
          4671 => x"cc",
          4672 => x"dc",
          4673 => x"38",
          4674 => x"b5",
          4675 => x"dc",
          4676 => x"74",
          4677 => x"0c",
          4678 => x"04",
          4679 => x"02",
          4680 => x"33",
          4681 => x"80",
          4682 => x"57",
          4683 => x"95",
          4684 => x"52",
          4685 => x"d2",
          4686 => x"dc",
          4687 => x"81",
          4688 => x"80",
          4689 => x"5a",
          4690 => x"3d",
          4691 => x"c9",
          4692 => x"dc",
          4693 => x"81",
          4694 => x"b8",
          4695 => x"cf",
          4696 => x"a0",
          4697 => x"55",
          4698 => x"75",
          4699 => x"71",
          4700 => x"33",
          4701 => x"74",
          4702 => x"57",
          4703 => x"8b",
          4704 => x"54",
          4705 => x"15",
          4706 => x"ff",
          4707 => x"81",
          4708 => x"55",
          4709 => x"cc",
          4710 => x"0d",
          4711 => x"0d",
          4712 => x"53",
          4713 => x"05",
          4714 => x"51",
          4715 => x"81",
          4716 => x"55",
          4717 => x"08",
          4718 => x"76",
          4719 => x"93",
          4720 => x"51",
          4721 => x"81",
          4722 => x"55",
          4723 => x"08",
          4724 => x"80",
          4725 => x"81",
          4726 => x"86",
          4727 => x"38",
          4728 => x"86",
          4729 => x"90",
          4730 => x"54",
          4731 => x"ff",
          4732 => x"76",
          4733 => x"83",
          4734 => x"51",
          4735 => x"3f",
          4736 => x"08",
          4737 => x"dc",
          4738 => x"3d",
          4739 => x"3d",
          4740 => x"5c",
          4741 => x"98",
          4742 => x"52",
          4743 => x"d1",
          4744 => x"dc",
          4745 => x"dc",
          4746 => x"70",
          4747 => x"08",
          4748 => x"51",
          4749 => x"80",
          4750 => x"38",
          4751 => x"06",
          4752 => x"80",
          4753 => x"38",
          4754 => x"5f",
          4755 => x"3d",
          4756 => x"ff",
          4757 => x"81",
          4758 => x"57",
          4759 => x"08",
          4760 => x"74",
          4761 => x"c3",
          4762 => x"dc",
          4763 => x"81",
          4764 => x"bf",
          4765 => x"cc",
          4766 => x"cc",
          4767 => x"59",
          4768 => x"81",
          4769 => x"56",
          4770 => x"33",
          4771 => x"16",
          4772 => x"27",
          4773 => x"56",
          4774 => x"80",
          4775 => x"80",
          4776 => x"ff",
          4777 => x"70",
          4778 => x"56",
          4779 => x"e8",
          4780 => x"76",
          4781 => x"81",
          4782 => x"80",
          4783 => x"57",
          4784 => x"78",
          4785 => x"51",
          4786 => x"2e",
          4787 => x"73",
          4788 => x"38",
          4789 => x"08",
          4790 => x"b1",
          4791 => x"dc",
          4792 => x"81",
          4793 => x"a7",
          4794 => x"33",
          4795 => x"c3",
          4796 => x"2e",
          4797 => x"e4",
          4798 => x"2e",
          4799 => x"56",
          4800 => x"05",
          4801 => x"e3",
          4802 => x"cc",
          4803 => x"76",
          4804 => x"0c",
          4805 => x"04",
          4806 => x"82",
          4807 => x"ff",
          4808 => x"9d",
          4809 => x"fa",
          4810 => x"cc",
          4811 => x"cc",
          4812 => x"81",
          4813 => x"83",
          4814 => x"53",
          4815 => x"3d",
          4816 => x"ff",
          4817 => x"73",
          4818 => x"70",
          4819 => x"52",
          4820 => x"9f",
          4821 => x"bc",
          4822 => x"74",
          4823 => x"6d",
          4824 => x"70",
          4825 => x"af",
          4826 => x"dc",
          4827 => x"2e",
          4828 => x"70",
          4829 => x"57",
          4830 => x"fd",
          4831 => x"cc",
          4832 => x"8d",
          4833 => x"2b",
          4834 => x"81",
          4835 => x"86",
          4836 => x"cc",
          4837 => x"9f",
          4838 => x"ff",
          4839 => x"54",
          4840 => x"8a",
          4841 => x"70",
          4842 => x"06",
          4843 => x"ff",
          4844 => x"38",
          4845 => x"15",
          4846 => x"80",
          4847 => x"74",
          4848 => x"9c",
          4849 => x"89",
          4850 => x"cc",
          4851 => x"81",
          4852 => x"88",
          4853 => x"26",
          4854 => x"39",
          4855 => x"86",
          4856 => x"81",
          4857 => x"ff",
          4858 => x"38",
          4859 => x"54",
          4860 => x"81",
          4861 => x"81",
          4862 => x"78",
          4863 => x"5a",
          4864 => x"6d",
          4865 => x"81",
          4866 => x"57",
          4867 => x"9f",
          4868 => x"38",
          4869 => x"54",
          4870 => x"81",
          4871 => x"b1",
          4872 => x"2e",
          4873 => x"a7",
          4874 => x"15",
          4875 => x"54",
          4876 => x"09",
          4877 => x"38",
          4878 => x"76",
          4879 => x"41",
          4880 => x"52",
          4881 => x"52",
          4882 => x"b3",
          4883 => x"cc",
          4884 => x"dc",
          4885 => x"f7",
          4886 => x"74",
          4887 => x"e5",
          4888 => x"cc",
          4889 => x"dc",
          4890 => x"38",
          4891 => x"38",
          4892 => x"74",
          4893 => x"39",
          4894 => x"08",
          4895 => x"81",
          4896 => x"38",
          4897 => x"74",
          4898 => x"38",
          4899 => x"51",
          4900 => x"3f",
          4901 => x"08",
          4902 => x"cc",
          4903 => x"a0",
          4904 => x"cc",
          4905 => x"51",
          4906 => x"3f",
          4907 => x"0b",
          4908 => x"8b",
          4909 => x"67",
          4910 => x"a7",
          4911 => x"81",
          4912 => x"34",
          4913 => x"ad",
          4914 => x"dc",
          4915 => x"73",
          4916 => x"dc",
          4917 => x"3d",
          4918 => x"3d",
          4919 => x"02",
          4920 => x"cb",
          4921 => x"3d",
          4922 => x"72",
          4923 => x"5a",
          4924 => x"81",
          4925 => x"58",
          4926 => x"08",
          4927 => x"91",
          4928 => x"77",
          4929 => x"7c",
          4930 => x"38",
          4931 => x"59",
          4932 => x"90",
          4933 => x"81",
          4934 => x"06",
          4935 => x"73",
          4936 => x"54",
          4937 => x"82",
          4938 => x"39",
          4939 => x"8b",
          4940 => x"11",
          4941 => x"2b",
          4942 => x"54",
          4943 => x"fe",
          4944 => x"ff",
          4945 => x"70",
          4946 => x"07",
          4947 => x"dc",
          4948 => x"8c",
          4949 => x"40",
          4950 => x"55",
          4951 => x"88",
          4952 => x"08",
          4953 => x"38",
          4954 => x"77",
          4955 => x"56",
          4956 => x"51",
          4957 => x"3f",
          4958 => x"55",
          4959 => x"08",
          4960 => x"38",
          4961 => x"dc",
          4962 => x"2e",
          4963 => x"81",
          4964 => x"ff",
          4965 => x"38",
          4966 => x"08",
          4967 => x"16",
          4968 => x"2e",
          4969 => x"87",
          4970 => x"74",
          4971 => x"74",
          4972 => x"81",
          4973 => x"38",
          4974 => x"ff",
          4975 => x"2e",
          4976 => x"7b",
          4977 => x"80",
          4978 => x"81",
          4979 => x"81",
          4980 => x"06",
          4981 => x"56",
          4982 => x"52",
          4983 => x"af",
          4984 => x"dc",
          4985 => x"81",
          4986 => x"80",
          4987 => x"81",
          4988 => x"56",
          4989 => x"d3",
          4990 => x"ff",
          4991 => x"7c",
          4992 => x"55",
          4993 => x"b3",
          4994 => x"1b",
          4995 => x"1b",
          4996 => x"33",
          4997 => x"54",
          4998 => x"34",
          4999 => x"fe",
          5000 => x"08",
          5001 => x"74",
          5002 => x"75",
          5003 => x"16",
          5004 => x"33",
          5005 => x"73",
          5006 => x"77",
          5007 => x"dc",
          5008 => x"3d",
          5009 => x"3d",
          5010 => x"02",
          5011 => x"eb",
          5012 => x"3d",
          5013 => x"59",
          5014 => x"8b",
          5015 => x"81",
          5016 => x"24",
          5017 => x"81",
          5018 => x"84",
          5019 => x"e8",
          5020 => x"51",
          5021 => x"2e",
          5022 => x"75",
          5023 => x"cc",
          5024 => x"06",
          5025 => x"7e",
          5026 => x"d0",
          5027 => x"cc",
          5028 => x"06",
          5029 => x"56",
          5030 => x"74",
          5031 => x"76",
          5032 => x"81",
          5033 => x"8a",
          5034 => x"b2",
          5035 => x"fc",
          5036 => x"52",
          5037 => x"a4",
          5038 => x"dc",
          5039 => x"38",
          5040 => x"80",
          5041 => x"74",
          5042 => x"26",
          5043 => x"15",
          5044 => x"74",
          5045 => x"38",
          5046 => x"80",
          5047 => x"84",
          5048 => x"92",
          5049 => x"80",
          5050 => x"38",
          5051 => x"06",
          5052 => x"2e",
          5053 => x"56",
          5054 => x"78",
          5055 => x"89",
          5056 => x"2b",
          5057 => x"43",
          5058 => x"38",
          5059 => x"30",
          5060 => x"77",
          5061 => x"91",
          5062 => x"c2",
          5063 => x"f8",
          5064 => x"52",
          5065 => x"a4",
          5066 => x"56",
          5067 => x"08",
          5068 => x"77",
          5069 => x"77",
          5070 => x"cc",
          5071 => x"45",
          5072 => x"bf",
          5073 => x"8e",
          5074 => x"26",
          5075 => x"74",
          5076 => x"48",
          5077 => x"75",
          5078 => x"38",
          5079 => x"81",
          5080 => x"fa",
          5081 => x"2a",
          5082 => x"56",
          5083 => x"2e",
          5084 => x"87",
          5085 => x"82",
          5086 => x"38",
          5087 => x"55",
          5088 => x"83",
          5089 => x"81",
          5090 => x"56",
          5091 => x"80",
          5092 => x"38",
          5093 => x"83",
          5094 => x"06",
          5095 => x"78",
          5096 => x"91",
          5097 => x"0b",
          5098 => x"22",
          5099 => x"80",
          5100 => x"74",
          5101 => x"38",
          5102 => x"56",
          5103 => x"17",
          5104 => x"57",
          5105 => x"2e",
          5106 => x"75",
          5107 => x"79",
          5108 => x"fe",
          5109 => x"81",
          5110 => x"84",
          5111 => x"05",
          5112 => x"5e",
          5113 => x"80",
          5114 => x"cc",
          5115 => x"8a",
          5116 => x"fd",
          5117 => x"75",
          5118 => x"38",
          5119 => x"78",
          5120 => x"8c",
          5121 => x"0b",
          5122 => x"22",
          5123 => x"80",
          5124 => x"74",
          5125 => x"38",
          5126 => x"56",
          5127 => x"17",
          5128 => x"57",
          5129 => x"2e",
          5130 => x"75",
          5131 => x"79",
          5132 => x"fe",
          5133 => x"81",
          5134 => x"10",
          5135 => x"81",
          5136 => x"9f",
          5137 => x"38",
          5138 => x"dc",
          5139 => x"81",
          5140 => x"05",
          5141 => x"2a",
          5142 => x"56",
          5143 => x"17",
          5144 => x"81",
          5145 => x"60",
          5146 => x"65",
          5147 => x"12",
          5148 => x"30",
          5149 => x"74",
          5150 => x"59",
          5151 => x"7d",
          5152 => x"81",
          5153 => x"76",
          5154 => x"41",
          5155 => x"76",
          5156 => x"90",
          5157 => x"62",
          5158 => x"51",
          5159 => x"26",
          5160 => x"75",
          5161 => x"31",
          5162 => x"65",
          5163 => x"fe",
          5164 => x"81",
          5165 => x"58",
          5166 => x"09",
          5167 => x"38",
          5168 => x"08",
          5169 => x"26",
          5170 => x"78",
          5171 => x"79",
          5172 => x"78",
          5173 => x"86",
          5174 => x"82",
          5175 => x"06",
          5176 => x"83",
          5177 => x"81",
          5178 => x"27",
          5179 => x"8f",
          5180 => x"55",
          5181 => x"26",
          5182 => x"59",
          5183 => x"62",
          5184 => x"74",
          5185 => x"38",
          5186 => x"88",
          5187 => x"cc",
          5188 => x"26",
          5189 => x"86",
          5190 => x"1a",
          5191 => x"79",
          5192 => x"38",
          5193 => x"80",
          5194 => x"2e",
          5195 => x"83",
          5196 => x"9f",
          5197 => x"8b",
          5198 => x"06",
          5199 => x"74",
          5200 => x"84",
          5201 => x"52",
          5202 => x"a2",
          5203 => x"53",
          5204 => x"52",
          5205 => x"a2",
          5206 => x"80",
          5207 => x"51",
          5208 => x"3f",
          5209 => x"34",
          5210 => x"ff",
          5211 => x"1b",
          5212 => x"a2",
          5213 => x"90",
          5214 => x"83",
          5215 => x"70",
          5216 => x"80",
          5217 => x"55",
          5218 => x"ff",
          5219 => x"66",
          5220 => x"ff",
          5221 => x"38",
          5222 => x"ff",
          5223 => x"1b",
          5224 => x"f2",
          5225 => x"74",
          5226 => x"51",
          5227 => x"3f",
          5228 => x"1c",
          5229 => x"98",
          5230 => x"a0",
          5231 => x"ff",
          5232 => x"51",
          5233 => x"3f",
          5234 => x"1b",
          5235 => x"e4",
          5236 => x"2e",
          5237 => x"80",
          5238 => x"88",
          5239 => x"80",
          5240 => x"ff",
          5241 => x"7c",
          5242 => x"51",
          5243 => x"3f",
          5244 => x"1b",
          5245 => x"bc",
          5246 => x"b0",
          5247 => x"a0",
          5248 => x"52",
          5249 => x"ff",
          5250 => x"ff",
          5251 => x"c0",
          5252 => x"0b",
          5253 => x"34",
          5254 => x"cb",
          5255 => x"c7",
          5256 => x"39",
          5257 => x"0a",
          5258 => x"51",
          5259 => x"3f",
          5260 => x"ff",
          5261 => x"1b",
          5262 => x"da",
          5263 => x"0b",
          5264 => x"a9",
          5265 => x"34",
          5266 => x"cb",
          5267 => x"1b",
          5268 => x"8f",
          5269 => x"d5",
          5270 => x"1b",
          5271 => x"ff",
          5272 => x"81",
          5273 => x"7a",
          5274 => x"ff",
          5275 => x"81",
          5276 => x"cc",
          5277 => x"38",
          5278 => x"09",
          5279 => x"ee",
          5280 => x"60",
          5281 => x"7a",
          5282 => x"ff",
          5283 => x"84",
          5284 => x"52",
          5285 => x"9f",
          5286 => x"8b",
          5287 => x"52",
          5288 => x"9f",
          5289 => x"8a",
          5290 => x"52",
          5291 => x"51",
          5292 => x"3f",
          5293 => x"83",
          5294 => x"ff",
          5295 => x"82",
          5296 => x"1b",
          5297 => x"ec",
          5298 => x"d5",
          5299 => x"ff",
          5300 => x"75",
          5301 => x"05",
          5302 => x"7e",
          5303 => x"e5",
          5304 => x"60",
          5305 => x"52",
          5306 => x"9a",
          5307 => x"53",
          5308 => x"51",
          5309 => x"3f",
          5310 => x"58",
          5311 => x"09",
          5312 => x"38",
          5313 => x"51",
          5314 => x"3f",
          5315 => x"1b",
          5316 => x"a0",
          5317 => x"52",
          5318 => x"91",
          5319 => x"ff",
          5320 => x"81",
          5321 => x"f8",
          5322 => x"7a",
          5323 => x"84",
          5324 => x"61",
          5325 => x"26",
          5326 => x"57",
          5327 => x"53",
          5328 => x"51",
          5329 => x"3f",
          5330 => x"08",
          5331 => x"84",
          5332 => x"dc",
          5333 => x"7a",
          5334 => x"aa",
          5335 => x"75",
          5336 => x"56",
          5337 => x"81",
          5338 => x"80",
          5339 => x"38",
          5340 => x"83",
          5341 => x"63",
          5342 => x"74",
          5343 => x"38",
          5344 => x"54",
          5345 => x"52",
          5346 => x"99",
          5347 => x"dc",
          5348 => x"c1",
          5349 => x"75",
          5350 => x"56",
          5351 => x"8c",
          5352 => x"2e",
          5353 => x"56",
          5354 => x"ff",
          5355 => x"84",
          5356 => x"2e",
          5357 => x"56",
          5358 => x"58",
          5359 => x"38",
          5360 => x"77",
          5361 => x"ff",
          5362 => x"82",
          5363 => x"78",
          5364 => x"c2",
          5365 => x"1b",
          5366 => x"34",
          5367 => x"16",
          5368 => x"82",
          5369 => x"83",
          5370 => x"84",
          5371 => x"67",
          5372 => x"fd",
          5373 => x"51",
          5374 => x"3f",
          5375 => x"16",
          5376 => x"cc",
          5377 => x"bf",
          5378 => x"86",
          5379 => x"dc",
          5380 => x"16",
          5381 => x"83",
          5382 => x"ff",
          5383 => x"66",
          5384 => x"1b",
          5385 => x"8c",
          5386 => x"77",
          5387 => x"7e",
          5388 => x"91",
          5389 => x"81",
          5390 => x"a2",
          5391 => x"80",
          5392 => x"ff",
          5393 => x"81",
          5394 => x"cc",
          5395 => x"89",
          5396 => x"8a",
          5397 => x"86",
          5398 => x"cc",
          5399 => x"81",
          5400 => x"99",
          5401 => x"f5",
          5402 => x"60",
          5403 => x"79",
          5404 => x"5a",
          5405 => x"78",
          5406 => x"8d",
          5407 => x"55",
          5408 => x"fc",
          5409 => x"51",
          5410 => x"7a",
          5411 => x"81",
          5412 => x"8c",
          5413 => x"74",
          5414 => x"38",
          5415 => x"81",
          5416 => x"81",
          5417 => x"8a",
          5418 => x"06",
          5419 => x"76",
          5420 => x"76",
          5421 => x"55",
          5422 => x"cc",
          5423 => x"0d",
          5424 => x"0d",
          5425 => x"70",
          5426 => x"74",
          5427 => x"ea",
          5428 => x"74",
          5429 => x"14",
          5430 => x"de",
          5431 => x"55",
          5432 => x"55",
          5433 => x"2e",
          5434 => x"56",
          5435 => x"9f",
          5436 => x"51",
          5437 => x"38",
          5438 => x"09",
          5439 => x"38",
          5440 => x"81",
          5441 => x"72",
          5442 => x"29",
          5443 => x"05",
          5444 => x"70",
          5445 => x"fe",
          5446 => x"81",
          5447 => x"8b",
          5448 => x"33",
          5449 => x"2e",
          5450 => x"81",
          5451 => x"ff",
          5452 => x"96",
          5453 => x"38",
          5454 => x"81",
          5455 => x"88",
          5456 => x"ff",
          5457 => x"52",
          5458 => x"81",
          5459 => x"84",
          5460 => x"fc",
          5461 => x"08",
          5462 => x"e8",
          5463 => x"39",
          5464 => x"51",
          5465 => x"81",
          5466 => x"80",
          5467 => x"cf",
          5468 => x"eb",
          5469 => x"ac",
          5470 => x"39",
          5471 => x"51",
          5472 => x"81",
          5473 => x"80",
          5474 => x"cf",
          5475 => x"cf",
          5476 => x"f8",
          5477 => x"39",
          5478 => x"51",
          5479 => x"81",
          5480 => x"bb",
          5481 => x"c4",
          5482 => x"81",
          5483 => x"af",
          5484 => x"84",
          5485 => x"81",
          5486 => x"a3",
          5487 => x"b8",
          5488 => x"81",
          5489 => x"97",
          5490 => x"e4",
          5491 => x"81",
          5492 => x"8b",
          5493 => x"94",
          5494 => x"81",
          5495 => x"ff",
          5496 => x"83",
          5497 => x"fb",
          5498 => x"79",
          5499 => x"87",
          5500 => x"38",
          5501 => x"87",
          5502 => x"91",
          5503 => x"52",
          5504 => x"ea",
          5505 => x"dc",
          5506 => x"75",
          5507 => x"ea",
          5508 => x"cc",
          5509 => x"53",
          5510 => x"d2",
          5511 => x"8b",
          5512 => x"3d",
          5513 => x"3d",
          5514 => x"84",
          5515 => x"05",
          5516 => x"80",
          5517 => x"70",
          5518 => x"25",
          5519 => x"59",
          5520 => x"87",
          5521 => x"38",
          5522 => x"76",
          5523 => x"ff",
          5524 => x"93",
          5525 => x"ff",
          5526 => x"76",
          5527 => x"70",
          5528 => x"9d",
          5529 => x"cc",
          5530 => x"dc",
          5531 => x"38",
          5532 => x"08",
          5533 => x"88",
          5534 => x"cc",
          5535 => x"3d",
          5536 => x"84",
          5537 => x"52",
          5538 => x"da",
          5539 => x"cc",
          5540 => x"dc",
          5541 => x"38",
          5542 => x"80",
          5543 => x"74",
          5544 => x"59",
          5545 => x"96",
          5546 => x"51",
          5547 => x"76",
          5548 => x"07",
          5549 => x"30",
          5550 => x"72",
          5551 => x"51",
          5552 => x"2e",
          5553 => x"d2",
          5554 => x"c0",
          5555 => x"52",
          5556 => x"93",
          5557 => x"75",
          5558 => x"0c",
          5559 => x"04",
          5560 => x"7b",
          5561 => x"b3",
          5562 => x"58",
          5563 => x"53",
          5564 => x"51",
          5565 => x"81",
          5566 => x"a4",
          5567 => x"2e",
          5568 => x"81",
          5569 => x"98",
          5570 => x"7f",
          5571 => x"cc",
          5572 => x"7d",
          5573 => x"81",
          5574 => x"57",
          5575 => x"04",
          5576 => x"cc",
          5577 => x"0d",
          5578 => x"0d",
          5579 => x"02",
          5580 => x"cf",
          5581 => x"73",
          5582 => x"5f",
          5583 => x"5e",
          5584 => x"81",
          5585 => x"ff",
          5586 => x"81",
          5587 => x"ff",
          5588 => x"80",
          5589 => x"27",
          5590 => x"7b",
          5591 => x"38",
          5592 => x"a7",
          5593 => x"39",
          5594 => x"72",
          5595 => x"38",
          5596 => x"81",
          5597 => x"ff",
          5598 => x"89",
          5599 => x"f4",
          5600 => x"fd",
          5601 => x"55",
          5602 => x"74",
          5603 => x"7a",
          5604 => x"72",
          5605 => x"d2",
          5606 => x"88",
          5607 => x"39",
          5608 => x"51",
          5609 => x"3f",
          5610 => x"a1",
          5611 => x"53",
          5612 => x"8e",
          5613 => x"52",
          5614 => x"51",
          5615 => x"3f",
          5616 => x"d3",
          5617 => x"82",
          5618 => x"15",
          5619 => x"ff",
          5620 => x"ff",
          5621 => x"d3",
          5622 => x"82",
          5623 => x"55",
          5624 => x"bc",
          5625 => x"70",
          5626 => x"80",
          5627 => x"27",
          5628 => x"56",
          5629 => x"74",
          5630 => x"81",
          5631 => x"06",
          5632 => x"06",
          5633 => x"80",
          5634 => x"73",
          5635 => x"85",
          5636 => x"83",
          5637 => x"ff",
          5638 => x"81",
          5639 => x"39",
          5640 => x"51",
          5641 => x"3f",
          5642 => x"1c",
          5643 => x"f6",
          5644 => x"dc",
          5645 => x"2b",
          5646 => x"51",
          5647 => x"2e",
          5648 => x"ab",
          5649 => x"c7",
          5650 => x"cc",
          5651 => x"70",
          5652 => x"a0",
          5653 => x"72",
          5654 => x"30",
          5655 => x"73",
          5656 => x"51",
          5657 => x"57",
          5658 => x"73",
          5659 => x"76",
          5660 => x"81",
          5661 => x"80",
          5662 => x"7c",
          5663 => x"78",
          5664 => x"38",
          5665 => x"81",
          5666 => x"8f",
          5667 => x"fc",
          5668 => x"9b",
          5669 => x"d3",
          5670 => x"d3",
          5671 => x"ff",
          5672 => x"81",
          5673 => x"51",
          5674 => x"3f",
          5675 => x"54",
          5676 => x"53",
          5677 => x"33",
          5678 => x"b4",
          5679 => x"a5",
          5680 => x"2e",
          5681 => x"fa",
          5682 => x"3d",
          5683 => x"3d",
          5684 => x"96",
          5685 => x"fe",
          5686 => x"81",
          5687 => x"c3",
          5688 => x"d0",
          5689 => x"bb",
          5690 => x"fe",
          5691 => x"72",
          5692 => x"81",
          5693 => x"71",
          5694 => x"38",
          5695 => x"f1",
          5696 => x"d3",
          5697 => x"f3",
          5698 => x"51",
          5699 => x"3f",
          5700 => x"70",
          5701 => x"52",
          5702 => x"95",
          5703 => x"fe",
          5704 => x"81",
          5705 => x"fe",
          5706 => x"80",
          5707 => x"f3",
          5708 => x"2a",
          5709 => x"51",
          5710 => x"2e",
          5711 => x"51",
          5712 => x"3f",
          5713 => x"51",
          5714 => x"3f",
          5715 => x"f0",
          5716 => x"84",
          5717 => x"06",
          5718 => x"80",
          5719 => x"81",
          5720 => x"bf",
          5721 => x"a0",
          5722 => x"b7",
          5723 => x"fe",
          5724 => x"72",
          5725 => x"81",
          5726 => x"71",
          5727 => x"38",
          5728 => x"f0",
          5729 => x"d4",
          5730 => x"f2",
          5731 => x"51",
          5732 => x"3f",
          5733 => x"70",
          5734 => x"52",
          5735 => x"95",
          5736 => x"fe",
          5737 => x"81",
          5738 => x"fe",
          5739 => x"80",
          5740 => x"ef",
          5741 => x"2a",
          5742 => x"51",
          5743 => x"2e",
          5744 => x"51",
          5745 => x"3f",
          5746 => x"51",
          5747 => x"3f",
          5748 => x"ef",
          5749 => x"88",
          5750 => x"06",
          5751 => x"80",
          5752 => x"81",
          5753 => x"bb",
          5754 => x"f0",
          5755 => x"b3",
          5756 => x"fe",
          5757 => x"fe",
          5758 => x"84",
          5759 => x"fb",
          5760 => x"79",
          5761 => x"56",
          5762 => x"51",
          5763 => x"3f",
          5764 => x"33",
          5765 => x"38",
          5766 => x"d5",
          5767 => x"f3",
          5768 => x"b9",
          5769 => x"dc",
          5770 => x"70",
          5771 => x"08",
          5772 => x"82",
          5773 => x"51",
          5774 => x"d9",
          5775 => x"d9",
          5776 => x"73",
          5777 => x"81",
          5778 => x"81",
          5779 => x"74",
          5780 => x"f4",
          5781 => x"dc",
          5782 => x"2e",
          5783 => x"dc",
          5784 => x"fe",
          5785 => x"8e",
          5786 => x"d0",
          5787 => x"3f",
          5788 => x"d9",
          5789 => x"d9",
          5790 => x"73",
          5791 => x"81",
          5792 => x"74",
          5793 => x"ff",
          5794 => x"80",
          5795 => x"cc",
          5796 => x"0d",
          5797 => x"0d",
          5798 => x"81",
          5799 => x"5f",
          5800 => x"7c",
          5801 => x"b4",
          5802 => x"cc",
          5803 => x"06",
          5804 => x"2e",
          5805 => x"a2",
          5806 => x"c0",
          5807 => x"70",
          5808 => x"82",
          5809 => x"53",
          5810 => x"dd",
          5811 => x"b7",
          5812 => x"dc",
          5813 => x"2e",
          5814 => x"d5",
          5815 => x"c1",
          5816 => x"5f",
          5817 => x"fc",
          5818 => x"95",
          5819 => x"70",
          5820 => x"f8",
          5821 => x"fe",
          5822 => x"3d",
          5823 => x"51",
          5824 => x"81",
          5825 => x"90",
          5826 => x"2c",
          5827 => x"80",
          5828 => x"b3",
          5829 => x"c2",
          5830 => x"78",
          5831 => x"d5",
          5832 => x"24",
          5833 => x"80",
          5834 => x"38",
          5835 => x"80",
          5836 => x"e9",
          5837 => x"c0",
          5838 => x"38",
          5839 => x"24",
          5840 => x"78",
          5841 => x"92",
          5842 => x"39",
          5843 => x"2e",
          5844 => x"78",
          5845 => x"92",
          5846 => x"c3",
          5847 => x"38",
          5848 => x"2e",
          5849 => x"8a",
          5850 => x"81",
          5851 => x"99",
          5852 => x"83",
          5853 => x"78",
          5854 => x"89",
          5855 => x"9d",
          5856 => x"85",
          5857 => x"38",
          5858 => x"b4",
          5859 => x"11",
          5860 => x"05",
          5861 => x"c2",
          5862 => x"cc",
          5863 => x"fe",
          5864 => x"3d",
          5865 => x"53",
          5866 => x"51",
          5867 => x"3f",
          5868 => x"08",
          5869 => x"ad",
          5870 => x"fe",
          5871 => x"ff",
          5872 => x"ff",
          5873 => x"81",
          5874 => x"86",
          5875 => x"cc",
          5876 => x"d6",
          5877 => x"fa",
          5878 => x"63",
          5879 => x"7b",
          5880 => x"38",
          5881 => x"7a",
          5882 => x"5c",
          5883 => x"26",
          5884 => x"e1",
          5885 => x"ff",
          5886 => x"ff",
          5887 => x"ff",
          5888 => x"81",
          5889 => x"80",
          5890 => x"38",
          5891 => x"fc",
          5892 => x"84",
          5893 => x"81",
          5894 => x"dc",
          5895 => x"2e",
          5896 => x"b4",
          5897 => x"11",
          5898 => x"05",
          5899 => x"aa",
          5900 => x"cc",
          5901 => x"fd",
          5902 => x"d6",
          5903 => x"f9",
          5904 => x"5a",
          5905 => x"81",
          5906 => x"59",
          5907 => x"05",
          5908 => x"34",
          5909 => x"42",
          5910 => x"3d",
          5911 => x"53",
          5912 => x"51",
          5913 => x"3f",
          5914 => x"08",
          5915 => x"f5",
          5916 => x"fe",
          5917 => x"ff",
          5918 => x"ff",
          5919 => x"81",
          5920 => x"80",
          5921 => x"38",
          5922 => x"f8",
          5923 => x"84",
          5924 => x"80",
          5925 => x"dc",
          5926 => x"2e",
          5927 => x"81",
          5928 => x"fe",
          5929 => x"63",
          5930 => x"27",
          5931 => x"70",
          5932 => x"5e",
          5933 => x"7c",
          5934 => x"78",
          5935 => x"79",
          5936 => x"52",
          5937 => x"51",
          5938 => x"3f",
          5939 => x"81",
          5940 => x"d5",
          5941 => x"c4",
          5942 => x"39",
          5943 => x"80",
          5944 => x"84",
          5945 => x"ff",
          5946 => x"dc",
          5947 => x"df",
          5948 => x"c0",
          5949 => x"80",
          5950 => x"81",
          5951 => x"44",
          5952 => x"81",
          5953 => x"59",
          5954 => x"88",
          5955 => x"80",
          5956 => x"39",
          5957 => x"33",
          5958 => x"2e",
          5959 => x"d9",
          5960 => x"ab",
          5961 => x"c3",
          5962 => x"80",
          5963 => x"81",
          5964 => x"44",
          5965 => x"d9",
          5966 => x"78",
          5967 => x"38",
          5968 => x"08",
          5969 => x"81",
          5970 => x"fc",
          5971 => x"b4",
          5972 => x"11",
          5973 => x"05",
          5974 => x"fe",
          5975 => x"cc",
          5976 => x"38",
          5977 => x"33",
          5978 => x"2e",
          5979 => x"d8",
          5980 => x"80",
          5981 => x"d9",
          5982 => x"78",
          5983 => x"38",
          5984 => x"08",
          5985 => x"81",
          5986 => x"59",
          5987 => x"88",
          5988 => x"8c",
          5989 => x"39",
          5990 => x"33",
          5991 => x"2e",
          5992 => x"d9",
          5993 => x"99",
          5994 => x"be",
          5995 => x"80",
          5996 => x"81",
          5997 => x"43",
          5998 => x"d9",
          5999 => x"05",
          6000 => x"fe",
          6001 => x"ff",
          6002 => x"fe",
          6003 => x"81",
          6004 => x"80",
          6005 => x"80",
          6006 => x"7a",
          6007 => x"38",
          6008 => x"90",
          6009 => x"70",
          6010 => x"2a",
          6011 => x"51",
          6012 => x"78",
          6013 => x"38",
          6014 => x"83",
          6015 => x"81",
          6016 => x"fe",
          6017 => x"a0",
          6018 => x"61",
          6019 => x"63",
          6020 => x"3f",
          6021 => x"51",
          6022 => x"3f",
          6023 => x"b4",
          6024 => x"11",
          6025 => x"05",
          6026 => x"ae",
          6027 => x"cc",
          6028 => x"f9",
          6029 => x"3d",
          6030 => x"53",
          6031 => x"51",
          6032 => x"3f",
          6033 => x"08",
          6034 => x"38",
          6035 => x"80",
          6036 => x"79",
          6037 => x"05",
          6038 => x"fe",
          6039 => x"ff",
          6040 => x"fe",
          6041 => x"81",
          6042 => x"e0",
          6043 => x"39",
          6044 => x"54",
          6045 => x"e4",
          6046 => x"e9",
          6047 => x"52",
          6048 => x"fb",
          6049 => x"45",
          6050 => x"78",
          6051 => x"d5",
          6052 => x"27",
          6053 => x"3d",
          6054 => x"53",
          6055 => x"51",
          6056 => x"3f",
          6057 => x"08",
          6058 => x"38",
          6059 => x"80",
          6060 => x"79",
          6061 => x"05",
          6062 => x"39",
          6063 => x"51",
          6064 => x"3f",
          6065 => x"b4",
          6066 => x"11",
          6067 => x"05",
          6068 => x"f8",
          6069 => x"cc",
          6070 => x"f8",
          6071 => x"3d",
          6072 => x"53",
          6073 => x"51",
          6074 => x"3f",
          6075 => x"08",
          6076 => x"38",
          6077 => x"be",
          6078 => x"70",
          6079 => x"23",
          6080 => x"3d",
          6081 => x"53",
          6082 => x"51",
          6083 => x"3f",
          6084 => x"08",
          6085 => x"cd",
          6086 => x"22",
          6087 => x"d6",
          6088 => x"f9",
          6089 => x"f8",
          6090 => x"fe",
          6091 => x"79",
          6092 => x"59",
          6093 => x"f7",
          6094 => x"9f",
          6095 => x"60",
          6096 => x"d5",
          6097 => x"fe",
          6098 => x"ff",
          6099 => x"fe",
          6100 => x"81",
          6101 => x"80",
          6102 => x"60",
          6103 => x"05",
          6104 => x"82",
          6105 => x"78",
          6106 => x"39",
          6107 => x"51",
          6108 => x"3f",
          6109 => x"b4",
          6110 => x"11",
          6111 => x"05",
          6112 => x"c8",
          6113 => x"cc",
          6114 => x"f6",
          6115 => x"3d",
          6116 => x"53",
          6117 => x"51",
          6118 => x"3f",
          6119 => x"08",
          6120 => x"38",
          6121 => x"0c",
          6122 => x"05",
          6123 => x"fe",
          6124 => x"ff",
          6125 => x"fe",
          6126 => x"81",
          6127 => x"e4",
          6128 => x"39",
          6129 => x"54",
          6130 => x"84",
          6131 => x"95",
          6132 => x"52",
          6133 => x"f8",
          6134 => x"45",
          6135 => x"78",
          6136 => x"81",
          6137 => x"27",
          6138 => x"3d",
          6139 => x"53",
          6140 => x"51",
          6141 => x"3f",
          6142 => x"08",
          6143 => x"38",
          6144 => x"0c",
          6145 => x"05",
          6146 => x"39",
          6147 => x"51",
          6148 => x"3f",
          6149 => x"b4",
          6150 => x"11",
          6151 => x"05",
          6152 => x"b6",
          6153 => x"cc",
          6154 => x"f5",
          6155 => x"52",
          6156 => x"51",
          6157 => x"3f",
          6158 => x"04",
          6159 => x"80",
          6160 => x"84",
          6161 => x"f9",
          6162 => x"dc",
          6163 => x"2e",
          6164 => x"63",
          6165 => x"ac",
          6166 => x"89",
          6167 => x"78",
          6168 => x"cc",
          6169 => x"f4",
          6170 => x"dc",
          6171 => x"81",
          6172 => x"fe",
          6173 => x"f4",
          6174 => x"d7",
          6175 => x"f1",
          6176 => x"d5",
          6177 => x"dd",
          6178 => x"80",
          6179 => x"f1",
          6180 => x"ff",
          6181 => x"eb",
          6182 => x"c9",
          6183 => x"33",
          6184 => x"80",
          6185 => x"38",
          6186 => x"59",
          6187 => x"81",
          6188 => x"3d",
          6189 => x"51",
          6190 => x"3f",
          6191 => x"08",
          6192 => x"7a",
          6193 => x"38",
          6194 => x"89",
          6195 => x"2e",
          6196 => x"cd",
          6197 => x"2e",
          6198 => x"c5",
          6199 => x"94",
          6200 => x"81",
          6201 => x"80",
          6202 => x"9c",
          6203 => x"ff",
          6204 => x"fe",
          6205 => x"bb",
          6206 => x"bc",
          6207 => x"ff",
          6208 => x"fe",
          6209 => x"ab",
          6210 => x"81",
          6211 => x"80",
          6212 => x"ac",
          6213 => x"ff",
          6214 => x"fe",
          6215 => x"93",
          6216 => x"80",
          6217 => x"b8",
          6218 => x"ff",
          6219 => x"fe",
          6220 => x"81",
          6221 => x"81",
          6222 => x"80",
          6223 => x"11",
          6224 => x"55",
          6225 => x"80",
          6226 => x"80",
          6227 => x"3d",
          6228 => x"51",
          6229 => x"81",
          6230 => x"81",
          6231 => x"09",
          6232 => x"72",
          6233 => x"51",
          6234 => x"80",
          6235 => x"26",
          6236 => x"5a",
          6237 => x"59",
          6238 => x"8d",
          6239 => x"70",
          6240 => x"5c",
          6241 => x"bb",
          6242 => x"32",
          6243 => x"07",
          6244 => x"38",
          6245 => x"09",
          6246 => x"c9",
          6247 => x"c0",
          6248 => x"c1",
          6249 => x"39",
          6250 => x"80",
          6251 => x"80",
          6252 => x"94",
          6253 => x"54",
          6254 => x"80",
          6255 => x"fe",
          6256 => x"81",
          6257 => x"90",
          6258 => x"55",
          6259 => x"80",
          6260 => x"fe",
          6261 => x"72",
          6262 => x"08",
          6263 => x"87",
          6264 => x"70",
          6265 => x"87",
          6266 => x"72",
          6267 => x"8a",
          6268 => x"cc",
          6269 => x"75",
          6270 => x"87",
          6271 => x"73",
          6272 => x"f6",
          6273 => x"dc",
          6274 => x"75",
          6275 => x"83",
          6276 => x"94",
          6277 => x"80",
          6278 => x"c0",
          6279 => x"a3",
          6280 => x"dc",
          6281 => x"bd",
          6282 => x"e0",
          6283 => x"b7",
          6284 => x"de",
          6285 => x"d0",
          6286 => x"c5",
          6287 => x"dc",
          6288 => x"bd",
          6289 => x"cd",
          6290 => x"c1",
          6291 => x"ec",
          6292 => x"c1",
          6293 => x"00",
          6294 => x"ff",
          6295 => x"ff",
          6296 => x"00",
          6297 => x"ff",
          6298 => x"18",
          6299 => x"18",
          6300 => x"18",
          6301 => x"18",
          6302 => x"18",
          6303 => x"55",
          6304 => x"55",
          6305 => x"55",
          6306 => x"55",
          6307 => x"55",
          6308 => x"55",
          6309 => x"55",
          6310 => x"55",
          6311 => x"55",
          6312 => x"55",
          6313 => x"55",
          6314 => x"55",
          6315 => x"55",
          6316 => x"55",
          6317 => x"55",
          6318 => x"55",
          6319 => x"55",
          6320 => x"55",
          6321 => x"55",
          6322 => x"55",
          6323 => x"2f",
          6324 => x"25",
          6325 => x"64",
          6326 => x"3a",
          6327 => x"25",
          6328 => x"0a",
          6329 => x"43",
          6330 => x"6e",
          6331 => x"75",
          6332 => x"69",
          6333 => x"00",
          6334 => x"66",
          6335 => x"20",
          6336 => x"20",
          6337 => x"66",
          6338 => x"00",
          6339 => x"44",
          6340 => x"63",
          6341 => x"69",
          6342 => x"65",
          6343 => x"74",
          6344 => x"0a",
          6345 => x"20",
          6346 => x"20",
          6347 => x"41",
          6348 => x"28",
          6349 => x"58",
          6350 => x"38",
          6351 => x"0a",
          6352 => x"20",
          6353 => x"52",
          6354 => x"20",
          6355 => x"28",
          6356 => x"58",
          6357 => x"38",
          6358 => x"0a",
          6359 => x"20",
          6360 => x"53",
          6361 => x"52",
          6362 => x"28",
          6363 => x"58",
          6364 => x"38",
          6365 => x"0a",
          6366 => x"20",
          6367 => x"41",
          6368 => x"20",
          6369 => x"28",
          6370 => x"58",
          6371 => x"38",
          6372 => x"0a",
          6373 => x"20",
          6374 => x"4d",
          6375 => x"20",
          6376 => x"28",
          6377 => x"58",
          6378 => x"38",
          6379 => x"0a",
          6380 => x"20",
          6381 => x"20",
          6382 => x"44",
          6383 => x"28",
          6384 => x"69",
          6385 => x"20",
          6386 => x"32",
          6387 => x"0a",
          6388 => x"20",
          6389 => x"4d",
          6390 => x"20",
          6391 => x"28",
          6392 => x"65",
          6393 => x"20",
          6394 => x"32",
          6395 => x"0a",
          6396 => x"20",
          6397 => x"54",
          6398 => x"54",
          6399 => x"28",
          6400 => x"6e",
          6401 => x"73",
          6402 => x"32",
          6403 => x"0a",
          6404 => x"20",
          6405 => x"53",
          6406 => x"4e",
          6407 => x"55",
          6408 => x"00",
          6409 => x"20",
          6410 => x"20",
          6411 => x"0a",
          6412 => x"20",
          6413 => x"43",
          6414 => x"00",
          6415 => x"20",
          6416 => x"32",
          6417 => x"00",
          6418 => x"20",
          6419 => x"49",
          6420 => x"00",
          6421 => x"64",
          6422 => x"73",
          6423 => x"0a",
          6424 => x"20",
          6425 => x"55",
          6426 => x"73",
          6427 => x"56",
          6428 => x"6f",
          6429 => x"64",
          6430 => x"73",
          6431 => x"20",
          6432 => x"58",
          6433 => x"00",
          6434 => x"20",
          6435 => x"55",
          6436 => x"6d",
          6437 => x"20",
          6438 => x"72",
          6439 => x"64",
          6440 => x"73",
          6441 => x"20",
          6442 => x"58",
          6443 => x"00",
          6444 => x"20",
          6445 => x"61",
          6446 => x"53",
          6447 => x"74",
          6448 => x"64",
          6449 => x"73",
          6450 => x"20",
          6451 => x"20",
          6452 => x"58",
          6453 => x"00",
          6454 => x"73",
          6455 => x"00",
          6456 => x"20",
          6457 => x"55",
          6458 => x"20",
          6459 => x"20",
          6460 => x"20",
          6461 => x"20",
          6462 => x"20",
          6463 => x"20",
          6464 => x"58",
          6465 => x"00",
          6466 => x"20",
          6467 => x"73",
          6468 => x"20",
          6469 => x"63",
          6470 => x"72",
          6471 => x"20",
          6472 => x"20",
          6473 => x"20",
          6474 => x"25",
          6475 => x"4d",
          6476 => x"00",
          6477 => x"20",
          6478 => x"52",
          6479 => x"43",
          6480 => x"6b",
          6481 => x"65",
          6482 => x"20",
          6483 => x"20",
          6484 => x"20",
          6485 => x"25",
          6486 => x"4d",
          6487 => x"00",
          6488 => x"20",
          6489 => x"73",
          6490 => x"6e",
          6491 => x"44",
          6492 => x"20",
          6493 => x"63",
          6494 => x"72",
          6495 => x"20",
          6496 => x"25",
          6497 => x"4d",
          6498 => x"00",
          6499 => x"61",
          6500 => x"00",
          6501 => x"64",
          6502 => x"00",
          6503 => x"65",
          6504 => x"00",
          6505 => x"4f",
          6506 => x"4f",
          6507 => x"00",
          6508 => x"6b",
          6509 => x"6e",
          6510 => x"00",
          6511 => x"2b",
          6512 => x"3c",
          6513 => x"5b",
          6514 => x"00",
          6515 => x"54",
          6516 => x"54",
          6517 => x"00",
          6518 => x"90",
          6519 => x"4f",
          6520 => x"30",
          6521 => x"20",
          6522 => x"45",
          6523 => x"20",
          6524 => x"33",
          6525 => x"20",
          6526 => x"20",
          6527 => x"45",
          6528 => x"20",
          6529 => x"20",
          6530 => x"20",
          6531 => x"65",
          6532 => x"00",
          6533 => x"00",
          6534 => x"00",
          6535 => x"45",
          6536 => x"8f",
          6537 => x"45",
          6538 => x"8e",
          6539 => x"92",
          6540 => x"55",
          6541 => x"9a",
          6542 => x"9e",
          6543 => x"4f",
          6544 => x"a6",
          6545 => x"aa",
          6546 => x"ae",
          6547 => x"b2",
          6548 => x"b6",
          6549 => x"ba",
          6550 => x"be",
          6551 => x"c2",
          6552 => x"c6",
          6553 => x"ca",
          6554 => x"ce",
          6555 => x"d2",
          6556 => x"d6",
          6557 => x"da",
          6558 => x"de",
          6559 => x"e2",
          6560 => x"e6",
          6561 => x"ea",
          6562 => x"ee",
          6563 => x"f2",
          6564 => x"f6",
          6565 => x"fa",
          6566 => x"fe",
          6567 => x"2c",
          6568 => x"5d",
          6569 => x"2a",
          6570 => x"3f",
          6571 => x"00",
          6572 => x"00",
          6573 => x"00",
          6574 => x"02",
          6575 => x"00",
          6576 => x"00",
          6577 => x"00",
          6578 => x"00",
          6579 => x"00",
          6580 => x"6e",
          6581 => x"00",
          6582 => x"6f",
          6583 => x"00",
          6584 => x"6e",
          6585 => x"00",
          6586 => x"6f",
          6587 => x"00",
          6588 => x"78",
          6589 => x"00",
          6590 => x"6c",
          6591 => x"00",
          6592 => x"6f",
          6593 => x"00",
          6594 => x"69",
          6595 => x"00",
          6596 => x"75",
          6597 => x"00",
          6598 => x"62",
          6599 => x"68",
          6600 => x"77",
          6601 => x"64",
          6602 => x"65",
          6603 => x"64",
          6604 => x"65",
          6605 => x"6c",
          6606 => x"00",
          6607 => x"70",
          6608 => x"73",
          6609 => x"74",
          6610 => x"73",
          6611 => x"00",
          6612 => x"66",
          6613 => x"00",
          6614 => x"73",
          6615 => x"00",
          6616 => x"61",
          6617 => x"00",
          6618 => x"73",
          6619 => x"72",
          6620 => x"0a",
          6621 => x"74",
          6622 => x"61",
          6623 => x"72",
          6624 => x"2e",
          6625 => x"00",
          6626 => x"73",
          6627 => x"6f",
          6628 => x"65",
          6629 => x"2e",
          6630 => x"00",
          6631 => x"20",
          6632 => x"65",
          6633 => x"75",
          6634 => x"0a",
          6635 => x"20",
          6636 => x"68",
          6637 => x"75",
          6638 => x"0a",
          6639 => x"76",
          6640 => x"64",
          6641 => x"6c",
          6642 => x"6d",
          6643 => x"00",
          6644 => x"63",
          6645 => x"20",
          6646 => x"69",
          6647 => x"0a",
          6648 => x"6c",
          6649 => x"6c",
          6650 => x"64",
          6651 => x"78",
          6652 => x"73",
          6653 => x"00",
          6654 => x"6c",
          6655 => x"61",
          6656 => x"65",
          6657 => x"76",
          6658 => x"64",
          6659 => x"00",
          6660 => x"20",
          6661 => x"77",
          6662 => x"65",
          6663 => x"6f",
          6664 => x"74",
          6665 => x"0a",
          6666 => x"69",
          6667 => x"6e",
          6668 => x"65",
          6669 => x"73",
          6670 => x"76",
          6671 => x"64",
          6672 => x"00",
          6673 => x"73",
          6674 => x"6f",
          6675 => x"6e",
          6676 => x"65",
          6677 => x"00",
          6678 => x"20",
          6679 => x"70",
          6680 => x"62",
          6681 => x"66",
          6682 => x"73",
          6683 => x"65",
          6684 => x"6f",
          6685 => x"20",
          6686 => x"64",
          6687 => x"2e",
          6688 => x"00",
          6689 => x"72",
          6690 => x"20",
          6691 => x"72",
          6692 => x"2e",
          6693 => x"00",
          6694 => x"6d",
          6695 => x"74",
          6696 => x"70",
          6697 => x"74",
          6698 => x"20",
          6699 => x"63",
          6700 => x"65",
          6701 => x"00",
          6702 => x"6c",
          6703 => x"73",
          6704 => x"63",
          6705 => x"2e",
          6706 => x"00",
          6707 => x"73",
          6708 => x"69",
          6709 => x"6e",
          6710 => x"65",
          6711 => x"79",
          6712 => x"00",
          6713 => x"6f",
          6714 => x"6e",
          6715 => x"70",
          6716 => x"66",
          6717 => x"73",
          6718 => x"00",
          6719 => x"72",
          6720 => x"74",
          6721 => x"20",
          6722 => x"6f",
          6723 => x"63",
          6724 => x"00",
          6725 => x"63",
          6726 => x"73",
          6727 => x"00",
          6728 => x"6b",
          6729 => x"6e",
          6730 => x"72",
          6731 => x"0a",
          6732 => x"6c",
          6733 => x"79",
          6734 => x"20",
          6735 => x"61",
          6736 => x"6c",
          6737 => x"79",
          6738 => x"2f",
          6739 => x"2e",
          6740 => x"00",
          6741 => x"61",
          6742 => x"00",
          6743 => x"38",
          6744 => x"00",
          6745 => x"20",
          6746 => x"34",
          6747 => x"00",
          6748 => x"20",
          6749 => x"20",
          6750 => x"00",
          6751 => x"32",
          6752 => x"00",
          6753 => x"00",
          6754 => x"00",
          6755 => x"0a",
          6756 => x"53",
          6757 => x"2a",
          6758 => x"20",
          6759 => x"00",
          6760 => x"2f",
          6761 => x"32",
          6762 => x"00",
          6763 => x"2e",
          6764 => x"00",
          6765 => x"50",
          6766 => x"72",
          6767 => x"25",
          6768 => x"29",
          6769 => x"20",
          6770 => x"2a",
          6771 => x"00",
          6772 => x"55",
          6773 => x"74",
          6774 => x"75",
          6775 => x"48",
          6776 => x"6c",
          6777 => x"00",
          6778 => x"6d",
          6779 => x"69",
          6780 => x"72",
          6781 => x"74",
          6782 => x"00",
          6783 => x"32",
          6784 => x"74",
          6785 => x"75",
          6786 => x"00",
          6787 => x"43",
          6788 => x"52",
          6789 => x"6e",
          6790 => x"72",
          6791 => x"0a",
          6792 => x"43",
          6793 => x"57",
          6794 => x"6e",
          6795 => x"72",
          6796 => x"0a",
          6797 => x"52",
          6798 => x"52",
          6799 => x"6e",
          6800 => x"72",
          6801 => x"0a",
          6802 => x"52",
          6803 => x"54",
          6804 => x"6e",
          6805 => x"72",
          6806 => x"0a",
          6807 => x"52",
          6808 => x"52",
          6809 => x"6e",
          6810 => x"72",
          6811 => x"0a",
          6812 => x"52",
          6813 => x"54",
          6814 => x"6e",
          6815 => x"72",
          6816 => x"0a",
          6817 => x"74",
          6818 => x"67",
          6819 => x"20",
          6820 => x"65",
          6821 => x"2e",
          6822 => x"00",
          6823 => x"61",
          6824 => x"6e",
          6825 => x"69",
          6826 => x"2e",
          6827 => x"00",
          6828 => x"74",
          6829 => x"65",
          6830 => x"61",
          6831 => x"00",
          6832 => x"00",
          6833 => x"69",
          6834 => x"20",
          6835 => x"69",
          6836 => x"69",
          6837 => x"73",
          6838 => x"64",
          6839 => x"72",
          6840 => x"2c",
          6841 => x"65",
          6842 => x"20",
          6843 => x"74",
          6844 => x"6e",
          6845 => x"6c",
          6846 => x"00",
          6847 => x"00",
          6848 => x"65",
          6849 => x"6e",
          6850 => x"2e",
          6851 => x"00",
          6852 => x"70",
          6853 => x"67",
          6854 => x"00",
          6855 => x"6d",
          6856 => x"69",
          6857 => x"2e",
          6858 => x"00",
          6859 => x"38",
          6860 => x"25",
          6861 => x"29",
          6862 => x"30",
          6863 => x"28",
          6864 => x"78",
          6865 => x"00",
          6866 => x"6d",
          6867 => x"65",
          6868 => x"79",
          6869 => x"00",
          6870 => x"6f",
          6871 => x"65",
          6872 => x"0a",
          6873 => x"38",
          6874 => x"30",
          6875 => x"00",
          6876 => x"3f",
          6877 => x"00",
          6878 => x"38",
          6879 => x"30",
          6880 => x"00",
          6881 => x"38",
          6882 => x"30",
          6883 => x"00",
          6884 => x"65",
          6885 => x"69",
          6886 => x"63",
          6887 => x"20",
          6888 => x"30",
          6889 => x"2e",
          6890 => x"00",
          6891 => x"6c",
          6892 => x"67",
          6893 => x"64",
          6894 => x"20",
          6895 => x"78",
          6896 => x"2e",
          6897 => x"00",
          6898 => x"6c",
          6899 => x"65",
          6900 => x"6e",
          6901 => x"63",
          6902 => x"20",
          6903 => x"29",
          6904 => x"00",
          6905 => x"73",
          6906 => x"74",
          6907 => x"20",
          6908 => x"6c",
          6909 => x"74",
          6910 => x"2e",
          6911 => x"00",
          6912 => x"6c",
          6913 => x"65",
          6914 => x"74",
          6915 => x"2e",
          6916 => x"00",
          6917 => x"55",
          6918 => x"6e",
          6919 => x"3a",
          6920 => x"5c",
          6921 => x"25",
          6922 => x"00",
          6923 => x"3a",
          6924 => x"5c",
          6925 => x"00",
          6926 => x"3a",
          6927 => x"00",
          6928 => x"64",
          6929 => x"6d",
          6930 => x"64",
          6931 => x"00",
          6932 => x"6e",
          6933 => x"67",
          6934 => x"0a",
          6935 => x"61",
          6936 => x"6e",
          6937 => x"6e",
          6938 => x"72",
          6939 => x"73",
          6940 => x"0a",
          6941 => x"00",
          6942 => x"00",
          6943 => x"7f",
          6944 => x"00",
          6945 => x"7f",
          6946 => x"00",
          6947 => x"7f",
          6948 => x"00",
          6949 => x"00",
          6950 => x"00",
          6951 => x"ff",
          6952 => x"00",
          6953 => x"00",
          6954 => x"78",
          6955 => x"00",
          6956 => x"e1",
          6957 => x"e1",
          6958 => x"e1",
          6959 => x"00",
          6960 => x"01",
          6961 => x"01",
          6962 => x"10",
          6963 => x"00",
          6964 => x"00",
          6965 => x"00",
          6966 => x"00",
          6967 => x"66",
          6968 => x"01",
          6969 => x"00",
          6970 => x"00",
          6971 => x"66",
          6972 => x"01",
          6973 => x"00",
          6974 => x"00",
          6975 => x"66",
          6976 => x"03",
          6977 => x"00",
          6978 => x"00",
          6979 => x"66",
          6980 => x"03",
          6981 => x"00",
          6982 => x"00",
          6983 => x"66",
          6984 => x"03",
          6985 => x"00",
          6986 => x"00",
          6987 => x"66",
          6988 => x"04",
          6989 => x"00",
          6990 => x"00",
          6991 => x"67",
          6992 => x"04",
          6993 => x"00",
          6994 => x"00",
          6995 => x"67",
          6996 => x"04",
          6997 => x"00",
          6998 => x"00",
          6999 => x"67",
          7000 => x"04",
          7001 => x"00",
          7002 => x"00",
          7003 => x"67",
          7004 => x"04",
          7005 => x"00",
          7006 => x"00",
          7007 => x"67",
          7008 => x"04",
          7009 => x"00",
          7010 => x"00",
          7011 => x"67",
          7012 => x"04",
          7013 => x"00",
          7014 => x"00",
          7015 => x"67",
          7016 => x"05",
          7017 => x"00",
          7018 => x"00",
          7019 => x"67",
          7020 => x"05",
          7021 => x"00",
          7022 => x"00",
          7023 => x"67",
          7024 => x"05",
          7025 => x"00",
          7026 => x"00",
          7027 => x"67",
          7028 => x"05",
          7029 => x"00",
          7030 => x"00",
          7031 => x"67",
          7032 => x"07",
          7033 => x"00",
          7034 => x"00",
          7035 => x"67",
          7036 => x"07",
          7037 => x"00",
          7038 => x"00",
          7039 => x"67",
          7040 => x"08",
          7041 => x"00",
          7042 => x"00",
          7043 => x"67",
          7044 => x"08",
          7045 => x"00",
          7046 => x"00",
          7047 => x"67",
          7048 => x"08",
          7049 => x"00",
          7050 => x"00",
          7051 => x"67",
          7052 => x"08",
          7053 => x"00",
          7054 => x"00",
          7055 => x"67",
          7056 => x"09",
          7057 => x"00",
          7058 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"a6",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"90",
           267 => x"0b",
           268 => x"04",
           269 => x"90",
           270 => x"0b",
           271 => x"04",
           272 => x"90",
           273 => x"0b",
           274 => x"04",
           275 => x"90",
           276 => x"0b",
           277 => x"04",
           278 => x"90",
           279 => x"0b",
           280 => x"04",
           281 => x"91",
           282 => x"0b",
           283 => x"04",
           284 => x"91",
           285 => x"0b",
           286 => x"04",
           287 => x"91",
           288 => x"0b",
           289 => x"04",
           290 => x"91",
           291 => x"0b",
           292 => x"04",
           293 => x"92",
           294 => x"0b",
           295 => x"04",
           296 => x"92",
           297 => x"0b",
           298 => x"04",
           299 => x"92",
           300 => x"0b",
           301 => x"04",
           302 => x"92",
           303 => x"0b",
           304 => x"04",
           305 => x"93",
           306 => x"0b",
           307 => x"04",
           308 => x"93",
           309 => x"0b",
           310 => x"04",
           311 => x"93",
           312 => x"0b",
           313 => x"04",
           314 => x"93",
           315 => x"0b",
           316 => x"04",
           317 => x"94",
           318 => x"0b",
           319 => x"04",
           320 => x"94",
           321 => x"0b",
           322 => x"04",
           323 => x"94",
           324 => x"0b",
           325 => x"04",
           326 => x"94",
           327 => x"0b",
           328 => x"04",
           329 => x"95",
           330 => x"0b",
           331 => x"04",
           332 => x"95",
           333 => x"0b",
           334 => x"04",
           335 => x"95",
           336 => x"0b",
           337 => x"04",
           338 => x"95",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"00",
           386 => x"00",
           387 => x"00",
           388 => x"00",
           389 => x"00",
           390 => x"00",
           391 => x"00",
           392 => x"00",
           393 => x"00",
           394 => x"00",
           395 => x"00",
           396 => x"00",
           397 => x"00",
           398 => x"00",
           399 => x"00",
           400 => x"00",
           401 => x"00",
           402 => x"00",
           403 => x"00",
           404 => x"00",
           405 => x"00",
           406 => x"00",
           407 => x"00",
           408 => x"00",
           409 => x"00",
           410 => x"00",
           411 => x"00",
           412 => x"00",
           413 => x"00",
           414 => x"00",
           415 => x"00",
           416 => x"00",
           417 => x"00",
           418 => x"00",
           419 => x"00",
           420 => x"00",
           421 => x"00",
           422 => x"00",
           423 => x"00",
           424 => x"00",
           425 => x"00",
           426 => x"00",
           427 => x"00",
           428 => x"00",
           429 => x"00",
           430 => x"00",
           431 => x"00",
           432 => x"00",
           433 => x"00",
           434 => x"00",
           435 => x"00",
           436 => x"00",
           437 => x"00",
           438 => x"00",
           439 => x"00",
           440 => x"00",
           441 => x"00",
           442 => x"00",
           443 => x"00",
           444 => x"00",
           445 => x"00",
           446 => x"00",
           447 => x"00",
           448 => x"00",
           449 => x"00",
           450 => x"00",
           451 => x"00",
           452 => x"00",
           453 => x"00",
           454 => x"00",
           455 => x"00",
           456 => x"00",
           457 => x"00",
           458 => x"00",
           459 => x"00",
           460 => x"00",
           461 => x"00",
           462 => x"00",
           463 => x"00",
           464 => x"00",
           465 => x"00",
           466 => x"00",
           467 => x"00",
           468 => x"00",
           469 => x"00",
           470 => x"00",
           471 => x"00",
           472 => x"00",
           473 => x"00",
           474 => x"00",
           475 => x"00",
           476 => x"00",
           477 => x"00",
           478 => x"00",
           479 => x"00",
           480 => x"00",
           481 => x"00",
           482 => x"00",
           483 => x"00",
           484 => x"00",
           485 => x"00",
           486 => x"00",
           487 => x"00",
           488 => x"00",
           489 => x"00",
           490 => x"00",
           491 => x"00",
           492 => x"00",
           493 => x"00",
           494 => x"00",
           495 => x"00",
           496 => x"00",
           497 => x"00",
           498 => x"00",
           499 => x"00",
           500 => x"00",
           501 => x"00",
           502 => x"00",
           503 => x"00",
           504 => x"00",
           505 => x"00",
           506 => x"00",
           507 => x"00",
           508 => x"00",
           509 => x"00",
           510 => x"00",
           511 => x"00",
           512 => x"00",
           513 => x"81",
           514 => x"a4",
           515 => x"dc",
           516 => x"80",
           517 => x"dc",
           518 => x"a3",
           519 => x"d8",
           520 => x"90",
           521 => x"d8",
           522 => x"2d",
           523 => x"08",
           524 => x"04",
           525 => x"0c",
           526 => x"81",
           527 => x"83",
           528 => x"81",
           529 => x"b8",
           530 => x"dc",
           531 => x"80",
           532 => x"dc",
           533 => x"bc",
           534 => x"d8",
           535 => x"90",
           536 => x"d8",
           537 => x"2d",
           538 => x"08",
           539 => x"04",
           540 => x"0c",
           541 => x"81",
           542 => x"83",
           543 => x"81",
           544 => x"bb",
           545 => x"dc",
           546 => x"80",
           547 => x"dc",
           548 => x"e4",
           549 => x"d8",
           550 => x"90",
           551 => x"d8",
           552 => x"2d",
           553 => x"08",
           554 => x"04",
           555 => x"0c",
           556 => x"81",
           557 => x"83",
           558 => x"81",
           559 => x"a6",
           560 => x"dc",
           561 => x"80",
           562 => x"dc",
           563 => x"8e",
           564 => x"d8",
           565 => x"90",
           566 => x"d8",
           567 => x"2d",
           568 => x"08",
           569 => x"04",
           570 => x"0c",
           571 => x"81",
           572 => x"83",
           573 => x"81",
           574 => x"a2",
           575 => x"dc",
           576 => x"80",
           577 => x"dc",
           578 => x"ee",
           579 => x"dc",
           580 => x"80",
           581 => x"dc",
           582 => x"fa",
           583 => x"dc",
           584 => x"80",
           585 => x"dc",
           586 => x"f2",
           587 => x"dc",
           588 => x"80",
           589 => x"dc",
           590 => x"f5",
           591 => x"dc",
           592 => x"80",
           593 => x"dc",
           594 => x"80",
           595 => x"dc",
           596 => x"80",
           597 => x"dc",
           598 => x"88",
           599 => x"dc",
           600 => x"80",
           601 => x"dc",
           602 => x"f9",
           603 => x"dc",
           604 => x"80",
           605 => x"dc",
           606 => x"83",
           607 => x"dc",
           608 => x"80",
           609 => x"dc",
           610 => x"84",
           611 => x"dc",
           612 => x"80",
           613 => x"dc",
           614 => x"84",
           615 => x"dc",
           616 => x"80",
           617 => x"dc",
           618 => x"8c",
           619 => x"dc",
           620 => x"80",
           621 => x"dc",
           622 => x"8a",
           623 => x"dc",
           624 => x"80",
           625 => x"dc",
           626 => x"8f",
           627 => x"dc",
           628 => x"80",
           629 => x"dc",
           630 => x"85",
           631 => x"dc",
           632 => x"80",
           633 => x"dc",
           634 => x"92",
           635 => x"dc",
           636 => x"80",
           637 => x"dc",
           638 => x"93",
           639 => x"dc",
           640 => x"80",
           641 => x"dc",
           642 => x"fb",
           643 => x"dc",
           644 => x"80",
           645 => x"dc",
           646 => x"fb",
           647 => x"dc",
           648 => x"80",
           649 => x"dc",
           650 => x"fc",
           651 => x"dc",
           652 => x"80",
           653 => x"dc",
           654 => x"86",
           655 => x"dc",
           656 => x"80",
           657 => x"dc",
           658 => x"94",
           659 => x"dc",
           660 => x"80",
           661 => x"dc",
           662 => x"96",
           663 => x"dc",
           664 => x"80",
           665 => x"dc",
           666 => x"99",
           667 => x"dc",
           668 => x"80",
           669 => x"dc",
           670 => x"ed",
           671 => x"dc",
           672 => x"80",
           673 => x"dc",
           674 => x"9c",
           675 => x"dc",
           676 => x"80",
           677 => x"dc",
           678 => x"da",
           679 => x"d8",
           680 => x"90",
           681 => x"d8",
           682 => x"c4",
           683 => x"d8",
           684 => x"90",
           685 => x"d8",
           686 => x"a8",
           687 => x"d8",
           688 => x"90",
           689 => x"d8",
           690 => x"2d",
           691 => x"08",
           692 => x"04",
           693 => x"0c",
           694 => x"81",
           695 => x"83",
           696 => x"81",
           697 => x"a3",
           698 => x"dc",
           699 => x"80",
           700 => x"dc",
           701 => x"aa",
           702 => x"dc",
           703 => x"80",
           704 => x"04",
           705 => x"10",
           706 => x"10",
           707 => x"10",
           708 => x"10",
           709 => x"10",
           710 => x"10",
           711 => x"10",
           712 => x"53",
           713 => x"00",
           714 => x"06",
           715 => x"09",
           716 => x"05",
           717 => x"2b",
           718 => x"06",
           719 => x"04",
           720 => x"72",
           721 => x"05",
           722 => x"05",
           723 => x"72",
           724 => x"53",
           725 => x"51",
           726 => x"04",
           727 => x"70",
           728 => x"27",
           729 => x"71",
           730 => x"53",
           731 => x"0b",
           732 => x"90",
           733 => x"c3",
           734 => x"81",
           735 => x"02",
           736 => x"0c",
           737 => x"80",
           738 => x"d8",
           739 => x"08",
           740 => x"d8",
           741 => x"08",
           742 => x"3f",
           743 => x"08",
           744 => x"cc",
           745 => x"3d",
           746 => x"d8",
           747 => x"dc",
           748 => x"81",
           749 => x"fd",
           750 => x"53",
           751 => x"08",
           752 => x"52",
           753 => x"08",
           754 => x"51",
           755 => x"81",
           756 => x"70",
           757 => x"0c",
           758 => x"0d",
           759 => x"0c",
           760 => x"d8",
           761 => x"dc",
           762 => x"3d",
           763 => x"81",
           764 => x"fc",
           765 => x"dc",
           766 => x"05",
           767 => x"b9",
           768 => x"d8",
           769 => x"08",
           770 => x"d8",
           771 => x"0c",
           772 => x"dc",
           773 => x"05",
           774 => x"d8",
           775 => x"08",
           776 => x"0b",
           777 => x"08",
           778 => x"81",
           779 => x"f4",
           780 => x"dc",
           781 => x"05",
           782 => x"d8",
           783 => x"08",
           784 => x"38",
           785 => x"08",
           786 => x"30",
           787 => x"08",
           788 => x"80",
           789 => x"d8",
           790 => x"0c",
           791 => x"08",
           792 => x"8a",
           793 => x"81",
           794 => x"f0",
           795 => x"dc",
           796 => x"05",
           797 => x"d8",
           798 => x"0c",
           799 => x"dc",
           800 => x"05",
           801 => x"dc",
           802 => x"05",
           803 => x"df",
           804 => x"cc",
           805 => x"dc",
           806 => x"05",
           807 => x"dc",
           808 => x"05",
           809 => x"90",
           810 => x"d8",
           811 => x"08",
           812 => x"d8",
           813 => x"0c",
           814 => x"08",
           815 => x"70",
           816 => x"0c",
           817 => x"0d",
           818 => x"0c",
           819 => x"d8",
           820 => x"dc",
           821 => x"3d",
           822 => x"81",
           823 => x"fc",
           824 => x"dc",
           825 => x"05",
           826 => x"99",
           827 => x"d8",
           828 => x"08",
           829 => x"d8",
           830 => x"0c",
           831 => x"dc",
           832 => x"05",
           833 => x"d8",
           834 => x"08",
           835 => x"38",
           836 => x"08",
           837 => x"30",
           838 => x"08",
           839 => x"81",
           840 => x"d8",
           841 => x"08",
           842 => x"d8",
           843 => x"08",
           844 => x"81",
           845 => x"70",
           846 => x"08",
           847 => x"54",
           848 => x"08",
           849 => x"80",
           850 => x"81",
           851 => x"f8",
           852 => x"81",
           853 => x"f8",
           854 => x"dc",
           855 => x"05",
           856 => x"dc",
           857 => x"87",
           858 => x"dc",
           859 => x"81",
           860 => x"02",
           861 => x"0c",
           862 => x"81",
           863 => x"d8",
           864 => x"0c",
           865 => x"dc",
           866 => x"05",
           867 => x"d8",
           868 => x"08",
           869 => x"08",
           870 => x"27",
           871 => x"dc",
           872 => x"05",
           873 => x"ae",
           874 => x"81",
           875 => x"8c",
           876 => x"a2",
           877 => x"d8",
           878 => x"08",
           879 => x"d8",
           880 => x"0c",
           881 => x"08",
           882 => x"10",
           883 => x"08",
           884 => x"ff",
           885 => x"dc",
           886 => x"05",
           887 => x"80",
           888 => x"dc",
           889 => x"05",
           890 => x"d8",
           891 => x"08",
           892 => x"81",
           893 => x"88",
           894 => x"dc",
           895 => x"05",
           896 => x"dc",
           897 => x"05",
           898 => x"d8",
           899 => x"08",
           900 => x"08",
           901 => x"07",
           902 => x"08",
           903 => x"81",
           904 => x"fc",
           905 => x"2a",
           906 => x"08",
           907 => x"81",
           908 => x"8c",
           909 => x"2a",
           910 => x"08",
           911 => x"ff",
           912 => x"dc",
           913 => x"05",
           914 => x"93",
           915 => x"d8",
           916 => x"08",
           917 => x"d8",
           918 => x"0c",
           919 => x"81",
           920 => x"f8",
           921 => x"81",
           922 => x"f4",
           923 => x"81",
           924 => x"f4",
           925 => x"dc",
           926 => x"3d",
           927 => x"d8",
           928 => x"3d",
           929 => x"71",
           930 => x"9f",
           931 => x"55",
           932 => x"72",
           933 => x"74",
           934 => x"70",
           935 => x"38",
           936 => x"71",
           937 => x"38",
           938 => x"81",
           939 => x"ff",
           940 => x"ff",
           941 => x"06",
           942 => x"81",
           943 => x"86",
           944 => x"74",
           945 => x"75",
           946 => x"90",
           947 => x"54",
           948 => x"27",
           949 => x"71",
           950 => x"53",
           951 => x"70",
           952 => x"0c",
           953 => x"84",
           954 => x"72",
           955 => x"05",
           956 => x"12",
           957 => x"26",
           958 => x"72",
           959 => x"72",
           960 => x"05",
           961 => x"12",
           962 => x"26",
           963 => x"53",
           964 => x"fb",
           965 => x"79",
           966 => x"83",
           967 => x"52",
           968 => x"71",
           969 => x"54",
           970 => x"73",
           971 => x"c6",
           972 => x"54",
           973 => x"70",
           974 => x"52",
           975 => x"2e",
           976 => x"33",
           977 => x"2e",
           978 => x"95",
           979 => x"81",
           980 => x"70",
           981 => x"54",
           982 => x"70",
           983 => x"33",
           984 => x"ff",
           985 => x"ff",
           986 => x"31",
           987 => x"0c",
           988 => x"3d",
           989 => x"09",
           990 => x"fd",
           991 => x"70",
           992 => x"81",
           993 => x"51",
           994 => x"38",
           995 => x"16",
           996 => x"56",
           997 => x"08",
           998 => x"73",
           999 => x"ff",
          1000 => x"0b",
          1001 => x"0c",
          1002 => x"04",
          1003 => x"80",
          1004 => x"71",
          1005 => x"87",
          1006 => x"dc",
          1007 => x"ff",
          1008 => x"ff",
          1009 => x"72",
          1010 => x"38",
          1011 => x"cc",
          1012 => x"0d",
          1013 => x"0d",
          1014 => x"70",
          1015 => x"71",
          1016 => x"ca",
          1017 => x"51",
          1018 => x"09",
          1019 => x"38",
          1020 => x"f1",
          1021 => x"84",
          1022 => x"53",
          1023 => x"70",
          1024 => x"53",
          1025 => x"a0",
          1026 => x"81",
          1027 => x"2e",
          1028 => x"e5",
          1029 => x"ff",
          1030 => x"a0",
          1031 => x"06",
          1032 => x"73",
          1033 => x"55",
          1034 => x"0c",
          1035 => x"81",
          1036 => x"87",
          1037 => x"fc",
          1038 => x"53",
          1039 => x"2e",
          1040 => x"3d",
          1041 => x"72",
          1042 => x"3f",
          1043 => x"08",
          1044 => x"53",
          1045 => x"53",
          1046 => x"cc",
          1047 => x"0d",
          1048 => x"0d",
          1049 => x"33",
          1050 => x"53",
          1051 => x"8b",
          1052 => x"38",
          1053 => x"ff",
          1054 => x"52",
          1055 => x"81",
          1056 => x"13",
          1057 => x"52",
          1058 => x"80",
          1059 => x"13",
          1060 => x"52",
          1061 => x"80",
          1062 => x"13",
          1063 => x"52",
          1064 => x"80",
          1065 => x"13",
          1066 => x"52",
          1067 => x"26",
          1068 => x"8a",
          1069 => x"87",
          1070 => x"e7",
          1071 => x"38",
          1072 => x"c0",
          1073 => x"72",
          1074 => x"98",
          1075 => x"13",
          1076 => x"98",
          1077 => x"13",
          1078 => x"98",
          1079 => x"13",
          1080 => x"98",
          1081 => x"13",
          1082 => x"98",
          1083 => x"13",
          1084 => x"98",
          1085 => x"87",
          1086 => x"0c",
          1087 => x"98",
          1088 => x"0b",
          1089 => x"9c",
          1090 => x"71",
          1091 => x"0c",
          1092 => x"04",
          1093 => x"7f",
          1094 => x"98",
          1095 => x"7d",
          1096 => x"98",
          1097 => x"7d",
          1098 => x"c0",
          1099 => x"5a",
          1100 => x"34",
          1101 => x"b4",
          1102 => x"83",
          1103 => x"c0",
          1104 => x"5a",
          1105 => x"34",
          1106 => x"ac",
          1107 => x"85",
          1108 => x"c0",
          1109 => x"5a",
          1110 => x"34",
          1111 => x"a4",
          1112 => x"88",
          1113 => x"c0",
          1114 => x"5a",
          1115 => x"23",
          1116 => x"79",
          1117 => x"06",
          1118 => x"ff",
          1119 => x"86",
          1120 => x"85",
          1121 => x"84",
          1122 => x"83",
          1123 => x"82",
          1124 => x"7d",
          1125 => x"06",
          1126 => x"cc",
          1127 => x"3f",
          1128 => x"04",
          1129 => x"02",
          1130 => x"70",
          1131 => x"2a",
          1132 => x"70",
          1133 => x"d8",
          1134 => x"3d",
          1135 => x"3d",
          1136 => x"0b",
          1137 => x"33",
          1138 => x"06",
          1139 => x"87",
          1140 => x"51",
          1141 => x"86",
          1142 => x"94",
          1143 => x"08",
          1144 => x"70",
          1145 => x"54",
          1146 => x"2e",
          1147 => x"91",
          1148 => x"06",
          1149 => x"d7",
          1150 => x"32",
          1151 => x"51",
          1152 => x"2e",
          1153 => x"93",
          1154 => x"06",
          1155 => x"ff",
          1156 => x"81",
          1157 => x"87",
          1158 => x"52",
          1159 => x"86",
          1160 => x"94",
          1161 => x"72",
          1162 => x"dc",
          1163 => x"3d",
          1164 => x"3d",
          1165 => x"05",
          1166 => x"81",
          1167 => x"70",
          1168 => x"57",
          1169 => x"c0",
          1170 => x"74",
          1171 => x"38",
          1172 => x"94",
          1173 => x"70",
          1174 => x"81",
          1175 => x"52",
          1176 => x"8c",
          1177 => x"2a",
          1178 => x"51",
          1179 => x"38",
          1180 => x"70",
          1181 => x"51",
          1182 => x"8d",
          1183 => x"2a",
          1184 => x"51",
          1185 => x"be",
          1186 => x"ff",
          1187 => x"c0",
          1188 => x"70",
          1189 => x"38",
          1190 => x"90",
          1191 => x"0c",
          1192 => x"04",
          1193 => x"79",
          1194 => x"33",
          1195 => x"06",
          1196 => x"70",
          1197 => x"fe",
          1198 => x"ff",
          1199 => x"0b",
          1200 => x"f4",
          1201 => x"ff",
          1202 => x"55",
          1203 => x"94",
          1204 => x"80",
          1205 => x"87",
          1206 => x"51",
          1207 => x"96",
          1208 => x"06",
          1209 => x"70",
          1210 => x"38",
          1211 => x"70",
          1212 => x"51",
          1213 => x"72",
          1214 => x"81",
          1215 => x"70",
          1216 => x"38",
          1217 => x"70",
          1218 => x"51",
          1219 => x"38",
          1220 => x"06",
          1221 => x"94",
          1222 => x"80",
          1223 => x"87",
          1224 => x"52",
          1225 => x"81",
          1226 => x"70",
          1227 => x"53",
          1228 => x"ff",
          1229 => x"81",
          1230 => x"89",
          1231 => x"fe",
          1232 => x"0b",
          1233 => x"33",
          1234 => x"06",
          1235 => x"c0",
          1236 => x"72",
          1237 => x"38",
          1238 => x"94",
          1239 => x"70",
          1240 => x"81",
          1241 => x"51",
          1242 => x"e2",
          1243 => x"ff",
          1244 => x"c0",
          1245 => x"70",
          1246 => x"38",
          1247 => x"90",
          1248 => x"70",
          1249 => x"81",
          1250 => x"51",
          1251 => x"04",
          1252 => x"0b",
          1253 => x"f4",
          1254 => x"ff",
          1255 => x"87",
          1256 => x"52",
          1257 => x"86",
          1258 => x"94",
          1259 => x"08",
          1260 => x"70",
          1261 => x"51",
          1262 => x"70",
          1263 => x"38",
          1264 => x"06",
          1265 => x"94",
          1266 => x"80",
          1267 => x"87",
          1268 => x"52",
          1269 => x"98",
          1270 => x"2c",
          1271 => x"71",
          1272 => x"0c",
          1273 => x"04",
          1274 => x"87",
          1275 => x"08",
          1276 => x"8a",
          1277 => x"70",
          1278 => x"b4",
          1279 => x"9e",
          1280 => x"d8",
          1281 => x"c0",
          1282 => x"81",
          1283 => x"87",
          1284 => x"08",
          1285 => x"0c",
          1286 => x"98",
          1287 => x"84",
          1288 => x"9e",
          1289 => x"d9",
          1290 => x"c0",
          1291 => x"81",
          1292 => x"87",
          1293 => x"08",
          1294 => x"0c",
          1295 => x"b0",
          1296 => x"94",
          1297 => x"9e",
          1298 => x"d9",
          1299 => x"c0",
          1300 => x"81",
          1301 => x"87",
          1302 => x"08",
          1303 => x"0c",
          1304 => x"c0",
          1305 => x"a4",
          1306 => x"9e",
          1307 => x"d9",
          1308 => x"c0",
          1309 => x"51",
          1310 => x"ac",
          1311 => x"9e",
          1312 => x"d9",
          1313 => x"c0",
          1314 => x"81",
          1315 => x"87",
          1316 => x"08",
          1317 => x"0c",
          1318 => x"d9",
          1319 => x"0b",
          1320 => x"90",
          1321 => x"80",
          1322 => x"52",
          1323 => x"2e",
          1324 => x"52",
          1325 => x"bd",
          1326 => x"87",
          1327 => x"08",
          1328 => x"0a",
          1329 => x"52",
          1330 => x"83",
          1331 => x"71",
          1332 => x"34",
          1333 => x"c0",
          1334 => x"70",
          1335 => x"06",
          1336 => x"70",
          1337 => x"38",
          1338 => x"81",
          1339 => x"80",
          1340 => x"9e",
          1341 => x"88",
          1342 => x"51",
          1343 => x"80",
          1344 => x"81",
          1345 => x"d9",
          1346 => x"0b",
          1347 => x"90",
          1348 => x"80",
          1349 => x"52",
          1350 => x"2e",
          1351 => x"52",
          1352 => x"c1",
          1353 => x"87",
          1354 => x"08",
          1355 => x"80",
          1356 => x"52",
          1357 => x"83",
          1358 => x"71",
          1359 => x"34",
          1360 => x"c0",
          1361 => x"70",
          1362 => x"06",
          1363 => x"70",
          1364 => x"38",
          1365 => x"81",
          1366 => x"80",
          1367 => x"9e",
          1368 => x"82",
          1369 => x"51",
          1370 => x"80",
          1371 => x"81",
          1372 => x"d9",
          1373 => x"0b",
          1374 => x"90",
          1375 => x"80",
          1376 => x"52",
          1377 => x"2e",
          1378 => x"52",
          1379 => x"c5",
          1380 => x"87",
          1381 => x"08",
          1382 => x"80",
          1383 => x"52",
          1384 => x"83",
          1385 => x"71",
          1386 => x"34",
          1387 => x"c0",
          1388 => x"70",
          1389 => x"51",
          1390 => x"80",
          1391 => x"81",
          1392 => x"d9",
          1393 => x"c0",
          1394 => x"70",
          1395 => x"70",
          1396 => x"51",
          1397 => x"d9",
          1398 => x"0b",
          1399 => x"90",
          1400 => x"80",
          1401 => x"52",
          1402 => x"83",
          1403 => x"71",
          1404 => x"34",
          1405 => x"90",
          1406 => x"f0",
          1407 => x"2a",
          1408 => x"70",
          1409 => x"34",
          1410 => x"c0",
          1411 => x"70",
          1412 => x"52",
          1413 => x"2e",
          1414 => x"52",
          1415 => x"cb",
          1416 => x"9e",
          1417 => x"87",
          1418 => x"70",
          1419 => x"34",
          1420 => x"04",
          1421 => x"81",
          1422 => x"85",
          1423 => x"d9",
          1424 => x"73",
          1425 => x"38",
          1426 => x"51",
          1427 => x"81",
          1428 => x"85",
          1429 => x"d9",
          1430 => x"73",
          1431 => x"38",
          1432 => x"08",
          1433 => x"08",
          1434 => x"81",
          1435 => x"8a",
          1436 => x"d9",
          1437 => x"73",
          1438 => x"38",
          1439 => x"08",
          1440 => x"08",
          1441 => x"81",
          1442 => x"8a",
          1443 => x"d9",
          1444 => x"73",
          1445 => x"38",
          1446 => x"08",
          1447 => x"08",
          1448 => x"81",
          1449 => x"8a",
          1450 => x"d9",
          1451 => x"73",
          1452 => x"38",
          1453 => x"08",
          1454 => x"08",
          1455 => x"81",
          1456 => x"8a",
          1457 => x"d9",
          1458 => x"73",
          1459 => x"38",
          1460 => x"08",
          1461 => x"08",
          1462 => x"81",
          1463 => x"8a",
          1464 => x"d9",
          1465 => x"73",
          1466 => x"38",
          1467 => x"33",
          1468 => x"b0",
          1469 => x"3f",
          1470 => x"33",
          1471 => x"2e",
          1472 => x"d9",
          1473 => x"81",
          1474 => x"89",
          1475 => x"d9",
          1476 => x"73",
          1477 => x"38",
          1478 => x"33",
          1479 => x"f0",
          1480 => x"3f",
          1481 => x"33",
          1482 => x"2e",
          1483 => x"c8",
          1484 => x"ce",
          1485 => x"bf",
          1486 => x"80",
          1487 => x"81",
          1488 => x"83",
          1489 => x"d9",
          1490 => x"73",
          1491 => x"38",
          1492 => x"51",
          1493 => x"81",
          1494 => x"54",
          1495 => x"88",
          1496 => x"bc",
          1497 => x"3f",
          1498 => x"33",
          1499 => x"2e",
          1500 => x"c8",
          1501 => x"8a",
          1502 => x"d4",
          1503 => x"3f",
          1504 => x"08",
          1505 => x"e0",
          1506 => x"3f",
          1507 => x"08",
          1508 => x"88",
          1509 => x"3f",
          1510 => x"08",
          1511 => x"b0",
          1512 => x"3f",
          1513 => x"51",
          1514 => x"81",
          1515 => x"52",
          1516 => x"51",
          1517 => x"81",
          1518 => x"56",
          1519 => x"52",
          1520 => x"b7",
          1521 => x"cc",
          1522 => x"c0",
          1523 => x"31",
          1524 => x"dc",
          1525 => x"81",
          1526 => x"88",
          1527 => x"d9",
          1528 => x"73",
          1529 => x"38",
          1530 => x"08",
          1531 => x"c0",
          1532 => x"e7",
          1533 => x"dc",
          1534 => x"84",
          1535 => x"71",
          1536 => x"81",
          1537 => x"52",
          1538 => x"51",
          1539 => x"81",
          1540 => x"54",
          1541 => x"a8",
          1542 => x"b8",
          1543 => x"84",
          1544 => x"51",
          1545 => x"81",
          1546 => x"bd",
          1547 => x"76",
          1548 => x"54",
          1549 => x"08",
          1550 => x"e0",
          1551 => x"3f",
          1552 => x"51",
          1553 => x"87",
          1554 => x"fe",
          1555 => x"92",
          1556 => x"05",
          1557 => x"26",
          1558 => x"84",
          1559 => x"e8",
          1560 => x"08",
          1561 => x"8c",
          1562 => x"81",
          1563 => x"97",
          1564 => x"9c",
          1565 => x"81",
          1566 => x"8b",
          1567 => x"a8",
          1568 => x"81",
          1569 => x"80",
          1570 => x"3d",
          1571 => x"88",
          1572 => x"80",
          1573 => x"96",
          1574 => x"81",
          1575 => x"87",
          1576 => x"0c",
          1577 => x"0d",
          1578 => x"33",
          1579 => x"2e",
          1580 => x"85",
          1581 => x"ed",
          1582 => x"e4",
          1583 => x"80",
          1584 => x"72",
          1585 => x"dc",
          1586 => x"05",
          1587 => x"0c",
          1588 => x"dc",
          1589 => x"71",
          1590 => x"38",
          1591 => x"2d",
          1592 => x"04",
          1593 => x"02",
          1594 => x"81",
          1595 => x"76",
          1596 => x"0c",
          1597 => x"ad",
          1598 => x"dc",
          1599 => x"3d",
          1600 => x"3d",
          1601 => x"73",
          1602 => x"ff",
          1603 => x"71",
          1604 => x"38",
          1605 => x"06",
          1606 => x"54",
          1607 => x"e7",
          1608 => x"0d",
          1609 => x"0d",
          1610 => x"dc",
          1611 => x"dc",
          1612 => x"54",
          1613 => x"81",
          1614 => x"53",
          1615 => x"8e",
          1616 => x"ff",
          1617 => x"14",
          1618 => x"3f",
          1619 => x"81",
          1620 => x"86",
          1621 => x"ec",
          1622 => x"68",
          1623 => x"70",
          1624 => x"33",
          1625 => x"2e",
          1626 => x"75",
          1627 => x"81",
          1628 => x"38",
          1629 => x"70",
          1630 => x"33",
          1631 => x"75",
          1632 => x"81",
          1633 => x"81",
          1634 => x"75",
          1635 => x"81",
          1636 => x"82",
          1637 => x"81",
          1638 => x"56",
          1639 => x"09",
          1640 => x"38",
          1641 => x"71",
          1642 => x"81",
          1643 => x"59",
          1644 => x"9d",
          1645 => x"53",
          1646 => x"95",
          1647 => x"29",
          1648 => x"76",
          1649 => x"79",
          1650 => x"5b",
          1651 => x"e5",
          1652 => x"ec",
          1653 => x"70",
          1654 => x"25",
          1655 => x"32",
          1656 => x"72",
          1657 => x"73",
          1658 => x"58",
          1659 => x"73",
          1660 => x"38",
          1661 => x"79",
          1662 => x"5b",
          1663 => x"75",
          1664 => x"de",
          1665 => x"80",
          1666 => x"89",
          1667 => x"70",
          1668 => x"55",
          1669 => x"cf",
          1670 => x"38",
          1671 => x"24",
          1672 => x"80",
          1673 => x"8e",
          1674 => x"c3",
          1675 => x"73",
          1676 => x"81",
          1677 => x"99",
          1678 => x"c4",
          1679 => x"38",
          1680 => x"73",
          1681 => x"81",
          1682 => x"80",
          1683 => x"38",
          1684 => x"2e",
          1685 => x"f9",
          1686 => x"d8",
          1687 => x"38",
          1688 => x"77",
          1689 => x"08",
          1690 => x"80",
          1691 => x"55",
          1692 => x"8d",
          1693 => x"70",
          1694 => x"51",
          1695 => x"f5",
          1696 => x"2a",
          1697 => x"74",
          1698 => x"53",
          1699 => x"8f",
          1700 => x"fc",
          1701 => x"81",
          1702 => x"80",
          1703 => x"73",
          1704 => x"3f",
          1705 => x"56",
          1706 => x"27",
          1707 => x"a0",
          1708 => x"3f",
          1709 => x"84",
          1710 => x"33",
          1711 => x"93",
          1712 => x"95",
          1713 => x"91",
          1714 => x"8d",
          1715 => x"89",
          1716 => x"fb",
          1717 => x"86",
          1718 => x"2a",
          1719 => x"51",
          1720 => x"2e",
          1721 => x"84",
          1722 => x"86",
          1723 => x"78",
          1724 => x"08",
          1725 => x"32",
          1726 => x"72",
          1727 => x"51",
          1728 => x"74",
          1729 => x"38",
          1730 => x"88",
          1731 => x"7a",
          1732 => x"55",
          1733 => x"3d",
          1734 => x"52",
          1735 => x"8e",
          1736 => x"cc",
          1737 => x"06",
          1738 => x"52",
          1739 => x"3f",
          1740 => x"08",
          1741 => x"27",
          1742 => x"14",
          1743 => x"f8",
          1744 => x"87",
          1745 => x"81",
          1746 => x"b0",
          1747 => x"7d",
          1748 => x"5f",
          1749 => x"75",
          1750 => x"07",
          1751 => x"54",
          1752 => x"26",
          1753 => x"ff",
          1754 => x"84",
          1755 => x"06",
          1756 => x"80",
          1757 => x"96",
          1758 => x"e0",
          1759 => x"73",
          1760 => x"57",
          1761 => x"06",
          1762 => x"54",
          1763 => x"a0",
          1764 => x"2a",
          1765 => x"54",
          1766 => x"38",
          1767 => x"76",
          1768 => x"38",
          1769 => x"fd",
          1770 => x"06",
          1771 => x"38",
          1772 => x"56",
          1773 => x"26",
          1774 => x"3d",
          1775 => x"05",
          1776 => x"ff",
          1777 => x"53",
          1778 => x"d9",
          1779 => x"38",
          1780 => x"56",
          1781 => x"27",
          1782 => x"a0",
          1783 => x"3f",
          1784 => x"3d",
          1785 => x"3d",
          1786 => x"70",
          1787 => x"52",
          1788 => x"73",
          1789 => x"3f",
          1790 => x"04",
          1791 => x"74",
          1792 => x"0c",
          1793 => x"05",
          1794 => x"fa",
          1795 => x"dc",
          1796 => x"80",
          1797 => x"0b",
          1798 => x"0c",
          1799 => x"04",
          1800 => x"81",
          1801 => x"76",
          1802 => x"0c",
          1803 => x"05",
          1804 => x"53",
          1805 => x"72",
          1806 => x"0c",
          1807 => x"04",
          1808 => x"77",
          1809 => x"e0",
          1810 => x"54",
          1811 => x"54",
          1812 => x"80",
          1813 => x"dc",
          1814 => x"71",
          1815 => x"cc",
          1816 => x"06",
          1817 => x"2e",
          1818 => x"72",
          1819 => x"38",
          1820 => x"70",
          1821 => x"25",
          1822 => x"73",
          1823 => x"38",
          1824 => x"86",
          1825 => x"54",
          1826 => x"73",
          1827 => x"ff",
          1828 => x"72",
          1829 => x"74",
          1830 => x"72",
          1831 => x"54",
          1832 => x"81",
          1833 => x"39",
          1834 => x"80",
          1835 => x"51",
          1836 => x"81",
          1837 => x"dc",
          1838 => x"3d",
          1839 => x"3d",
          1840 => x"e0",
          1841 => x"dc",
          1842 => x"53",
          1843 => x"fe",
          1844 => x"81",
          1845 => x"84",
          1846 => x"f8",
          1847 => x"7c",
          1848 => x"70",
          1849 => x"75",
          1850 => x"55",
          1851 => x"2e",
          1852 => x"87",
          1853 => x"76",
          1854 => x"73",
          1855 => x"81",
          1856 => x"81",
          1857 => x"77",
          1858 => x"70",
          1859 => x"58",
          1860 => x"09",
          1861 => x"c2",
          1862 => x"81",
          1863 => x"75",
          1864 => x"55",
          1865 => x"e2",
          1866 => x"90",
          1867 => x"f8",
          1868 => x"8f",
          1869 => x"81",
          1870 => x"75",
          1871 => x"55",
          1872 => x"81",
          1873 => x"27",
          1874 => x"d0",
          1875 => x"55",
          1876 => x"73",
          1877 => x"80",
          1878 => x"14",
          1879 => x"72",
          1880 => x"e0",
          1881 => x"80",
          1882 => x"39",
          1883 => x"55",
          1884 => x"80",
          1885 => x"e0",
          1886 => x"38",
          1887 => x"81",
          1888 => x"53",
          1889 => x"81",
          1890 => x"53",
          1891 => x"8e",
          1892 => x"70",
          1893 => x"55",
          1894 => x"27",
          1895 => x"77",
          1896 => x"74",
          1897 => x"76",
          1898 => x"77",
          1899 => x"70",
          1900 => x"55",
          1901 => x"77",
          1902 => x"38",
          1903 => x"74",
          1904 => x"55",
          1905 => x"cc",
          1906 => x"0d",
          1907 => x"0d",
          1908 => x"56",
          1909 => x"0c",
          1910 => x"70",
          1911 => x"73",
          1912 => x"81",
          1913 => x"81",
          1914 => x"ed",
          1915 => x"2e",
          1916 => x"8e",
          1917 => x"08",
          1918 => x"76",
          1919 => x"56",
          1920 => x"b0",
          1921 => x"06",
          1922 => x"75",
          1923 => x"76",
          1924 => x"70",
          1925 => x"73",
          1926 => x"8b",
          1927 => x"73",
          1928 => x"85",
          1929 => x"82",
          1930 => x"76",
          1931 => x"70",
          1932 => x"ac",
          1933 => x"a0",
          1934 => x"fa",
          1935 => x"53",
          1936 => x"57",
          1937 => x"98",
          1938 => x"39",
          1939 => x"80",
          1940 => x"26",
          1941 => x"86",
          1942 => x"80",
          1943 => x"57",
          1944 => x"74",
          1945 => x"38",
          1946 => x"27",
          1947 => x"14",
          1948 => x"06",
          1949 => x"14",
          1950 => x"06",
          1951 => x"74",
          1952 => x"f9",
          1953 => x"ff",
          1954 => x"89",
          1955 => x"38",
          1956 => x"c5",
          1957 => x"29",
          1958 => x"81",
          1959 => x"76",
          1960 => x"56",
          1961 => x"ba",
          1962 => x"2e",
          1963 => x"30",
          1964 => x"0c",
          1965 => x"81",
          1966 => x"8a",
          1967 => x"ff",
          1968 => x"8f",
          1969 => x"81",
          1970 => x"26",
          1971 => x"d9",
          1972 => x"52",
          1973 => x"cc",
          1974 => x"0d",
          1975 => x"0d",
          1976 => x"33",
          1977 => x"9f",
          1978 => x"53",
          1979 => x"81",
          1980 => x"38",
          1981 => x"87",
          1982 => x"11",
          1983 => x"54",
          1984 => x"84",
          1985 => x"54",
          1986 => x"87",
          1987 => x"11",
          1988 => x"0c",
          1989 => x"c0",
          1990 => x"70",
          1991 => x"70",
          1992 => x"51",
          1993 => x"8a",
          1994 => x"98",
          1995 => x"70",
          1996 => x"08",
          1997 => x"06",
          1998 => x"38",
          1999 => x"8c",
          2000 => x"80",
          2001 => x"71",
          2002 => x"14",
          2003 => x"d4",
          2004 => x"70",
          2005 => x"0c",
          2006 => x"04",
          2007 => x"60",
          2008 => x"8c",
          2009 => x"33",
          2010 => x"5b",
          2011 => x"5a",
          2012 => x"81",
          2013 => x"81",
          2014 => x"52",
          2015 => x"38",
          2016 => x"84",
          2017 => x"92",
          2018 => x"c0",
          2019 => x"87",
          2020 => x"13",
          2021 => x"57",
          2022 => x"0b",
          2023 => x"8c",
          2024 => x"0c",
          2025 => x"75",
          2026 => x"2a",
          2027 => x"51",
          2028 => x"80",
          2029 => x"7b",
          2030 => x"7b",
          2031 => x"5d",
          2032 => x"59",
          2033 => x"06",
          2034 => x"73",
          2035 => x"81",
          2036 => x"ff",
          2037 => x"72",
          2038 => x"38",
          2039 => x"8c",
          2040 => x"c3",
          2041 => x"98",
          2042 => x"71",
          2043 => x"38",
          2044 => x"2e",
          2045 => x"76",
          2046 => x"92",
          2047 => x"72",
          2048 => x"06",
          2049 => x"f7",
          2050 => x"5a",
          2051 => x"80",
          2052 => x"70",
          2053 => x"5a",
          2054 => x"80",
          2055 => x"73",
          2056 => x"06",
          2057 => x"38",
          2058 => x"fe",
          2059 => x"fc",
          2060 => x"52",
          2061 => x"83",
          2062 => x"71",
          2063 => x"dc",
          2064 => x"3d",
          2065 => x"3d",
          2066 => x"64",
          2067 => x"bf",
          2068 => x"40",
          2069 => x"59",
          2070 => x"58",
          2071 => x"81",
          2072 => x"81",
          2073 => x"52",
          2074 => x"09",
          2075 => x"b1",
          2076 => x"84",
          2077 => x"92",
          2078 => x"c0",
          2079 => x"87",
          2080 => x"13",
          2081 => x"56",
          2082 => x"87",
          2083 => x"0c",
          2084 => x"82",
          2085 => x"58",
          2086 => x"84",
          2087 => x"06",
          2088 => x"71",
          2089 => x"38",
          2090 => x"05",
          2091 => x"0c",
          2092 => x"73",
          2093 => x"81",
          2094 => x"71",
          2095 => x"38",
          2096 => x"8c",
          2097 => x"d0",
          2098 => x"98",
          2099 => x"71",
          2100 => x"38",
          2101 => x"2e",
          2102 => x"76",
          2103 => x"92",
          2104 => x"72",
          2105 => x"06",
          2106 => x"f7",
          2107 => x"59",
          2108 => x"1a",
          2109 => x"06",
          2110 => x"59",
          2111 => x"80",
          2112 => x"73",
          2113 => x"06",
          2114 => x"38",
          2115 => x"fe",
          2116 => x"fc",
          2117 => x"52",
          2118 => x"83",
          2119 => x"71",
          2120 => x"dc",
          2121 => x"3d",
          2122 => x"3d",
          2123 => x"84",
          2124 => x"33",
          2125 => x"a7",
          2126 => x"54",
          2127 => x"fa",
          2128 => x"dc",
          2129 => x"06",
          2130 => x"72",
          2131 => x"85",
          2132 => x"98",
          2133 => x"56",
          2134 => x"80",
          2135 => x"76",
          2136 => x"74",
          2137 => x"c0",
          2138 => x"54",
          2139 => x"2e",
          2140 => x"d4",
          2141 => x"2e",
          2142 => x"80",
          2143 => x"08",
          2144 => x"70",
          2145 => x"51",
          2146 => x"2e",
          2147 => x"c0",
          2148 => x"52",
          2149 => x"87",
          2150 => x"08",
          2151 => x"38",
          2152 => x"87",
          2153 => x"14",
          2154 => x"70",
          2155 => x"52",
          2156 => x"96",
          2157 => x"92",
          2158 => x"0a",
          2159 => x"39",
          2160 => x"0c",
          2161 => x"39",
          2162 => x"54",
          2163 => x"cc",
          2164 => x"0d",
          2165 => x"0d",
          2166 => x"33",
          2167 => x"88",
          2168 => x"dc",
          2169 => x"51",
          2170 => x"04",
          2171 => x"75",
          2172 => x"82",
          2173 => x"90",
          2174 => x"2b",
          2175 => x"33",
          2176 => x"88",
          2177 => x"71",
          2178 => x"cc",
          2179 => x"54",
          2180 => x"85",
          2181 => x"ff",
          2182 => x"02",
          2183 => x"05",
          2184 => x"70",
          2185 => x"05",
          2186 => x"88",
          2187 => x"72",
          2188 => x"0d",
          2189 => x"0d",
          2190 => x"52",
          2191 => x"81",
          2192 => x"70",
          2193 => x"70",
          2194 => x"05",
          2195 => x"88",
          2196 => x"72",
          2197 => x"54",
          2198 => x"2a",
          2199 => x"34",
          2200 => x"04",
          2201 => x"76",
          2202 => x"54",
          2203 => x"2e",
          2204 => x"70",
          2205 => x"33",
          2206 => x"05",
          2207 => x"11",
          2208 => x"84",
          2209 => x"fe",
          2210 => x"77",
          2211 => x"53",
          2212 => x"81",
          2213 => x"ff",
          2214 => x"f4",
          2215 => x"0d",
          2216 => x"0d",
          2217 => x"56",
          2218 => x"70",
          2219 => x"33",
          2220 => x"05",
          2221 => x"71",
          2222 => x"56",
          2223 => x"72",
          2224 => x"38",
          2225 => x"e2",
          2226 => x"dc",
          2227 => x"3d",
          2228 => x"3d",
          2229 => x"54",
          2230 => x"71",
          2231 => x"38",
          2232 => x"70",
          2233 => x"f3",
          2234 => x"81",
          2235 => x"84",
          2236 => x"80",
          2237 => x"cc",
          2238 => x"0b",
          2239 => x"0c",
          2240 => x"0d",
          2241 => x"0b",
          2242 => x"56",
          2243 => x"2e",
          2244 => x"81",
          2245 => x"08",
          2246 => x"70",
          2247 => x"33",
          2248 => x"a2",
          2249 => x"cc",
          2250 => x"09",
          2251 => x"38",
          2252 => x"08",
          2253 => x"b0",
          2254 => x"a4",
          2255 => x"9c",
          2256 => x"56",
          2257 => x"27",
          2258 => x"16",
          2259 => x"82",
          2260 => x"06",
          2261 => x"54",
          2262 => x"78",
          2263 => x"33",
          2264 => x"3f",
          2265 => x"5a",
          2266 => x"cc",
          2267 => x"0d",
          2268 => x"0d",
          2269 => x"56",
          2270 => x"b0",
          2271 => x"af",
          2272 => x"fe",
          2273 => x"dc",
          2274 => x"81",
          2275 => x"9f",
          2276 => x"74",
          2277 => x"52",
          2278 => x"51",
          2279 => x"81",
          2280 => x"80",
          2281 => x"ff",
          2282 => x"74",
          2283 => x"76",
          2284 => x"0c",
          2285 => x"04",
          2286 => x"7a",
          2287 => x"fe",
          2288 => x"dc",
          2289 => x"81",
          2290 => x"81",
          2291 => x"33",
          2292 => x"2e",
          2293 => x"80",
          2294 => x"17",
          2295 => x"81",
          2296 => x"06",
          2297 => x"84",
          2298 => x"dc",
          2299 => x"b4",
          2300 => x"56",
          2301 => x"82",
          2302 => x"84",
          2303 => x"fc",
          2304 => x"8b",
          2305 => x"52",
          2306 => x"a9",
          2307 => x"85",
          2308 => x"84",
          2309 => x"fc",
          2310 => x"17",
          2311 => x"9c",
          2312 => x"91",
          2313 => x"08",
          2314 => x"17",
          2315 => x"3f",
          2316 => x"81",
          2317 => x"19",
          2318 => x"53",
          2319 => x"17",
          2320 => x"82",
          2321 => x"18",
          2322 => x"80",
          2323 => x"33",
          2324 => x"3f",
          2325 => x"08",
          2326 => x"38",
          2327 => x"81",
          2328 => x"8a",
          2329 => x"fb",
          2330 => x"fe",
          2331 => x"08",
          2332 => x"56",
          2333 => x"74",
          2334 => x"38",
          2335 => x"75",
          2336 => x"16",
          2337 => x"53",
          2338 => x"cc",
          2339 => x"0d",
          2340 => x"0d",
          2341 => x"08",
          2342 => x"81",
          2343 => x"df",
          2344 => x"15",
          2345 => x"d7",
          2346 => x"33",
          2347 => x"82",
          2348 => x"38",
          2349 => x"89",
          2350 => x"2e",
          2351 => x"bf",
          2352 => x"2e",
          2353 => x"81",
          2354 => x"81",
          2355 => x"89",
          2356 => x"08",
          2357 => x"52",
          2358 => x"3f",
          2359 => x"08",
          2360 => x"74",
          2361 => x"14",
          2362 => x"81",
          2363 => x"2a",
          2364 => x"05",
          2365 => x"57",
          2366 => x"f5",
          2367 => x"cc",
          2368 => x"38",
          2369 => x"06",
          2370 => x"33",
          2371 => x"78",
          2372 => x"06",
          2373 => x"5c",
          2374 => x"53",
          2375 => x"38",
          2376 => x"06",
          2377 => x"39",
          2378 => x"a4",
          2379 => x"52",
          2380 => x"bd",
          2381 => x"cc",
          2382 => x"38",
          2383 => x"fe",
          2384 => x"b4",
          2385 => x"8d",
          2386 => x"cc",
          2387 => x"ff",
          2388 => x"39",
          2389 => x"a4",
          2390 => x"52",
          2391 => x"91",
          2392 => x"cc",
          2393 => x"76",
          2394 => x"fc",
          2395 => x"b4",
          2396 => x"f8",
          2397 => x"cc",
          2398 => x"06",
          2399 => x"81",
          2400 => x"dc",
          2401 => x"3d",
          2402 => x"3d",
          2403 => x"7e",
          2404 => x"82",
          2405 => x"27",
          2406 => x"76",
          2407 => x"27",
          2408 => x"75",
          2409 => x"79",
          2410 => x"38",
          2411 => x"89",
          2412 => x"2e",
          2413 => x"80",
          2414 => x"2e",
          2415 => x"81",
          2416 => x"81",
          2417 => x"89",
          2418 => x"08",
          2419 => x"52",
          2420 => x"3f",
          2421 => x"08",
          2422 => x"cc",
          2423 => x"38",
          2424 => x"06",
          2425 => x"81",
          2426 => x"06",
          2427 => x"77",
          2428 => x"2e",
          2429 => x"84",
          2430 => x"06",
          2431 => x"06",
          2432 => x"53",
          2433 => x"81",
          2434 => x"34",
          2435 => x"a4",
          2436 => x"52",
          2437 => x"d9",
          2438 => x"cc",
          2439 => x"dc",
          2440 => x"94",
          2441 => x"ff",
          2442 => x"05",
          2443 => x"54",
          2444 => x"38",
          2445 => x"74",
          2446 => x"06",
          2447 => x"07",
          2448 => x"74",
          2449 => x"39",
          2450 => x"a4",
          2451 => x"52",
          2452 => x"9d",
          2453 => x"cc",
          2454 => x"dc",
          2455 => x"d8",
          2456 => x"ff",
          2457 => x"76",
          2458 => x"06",
          2459 => x"05",
          2460 => x"3f",
          2461 => x"87",
          2462 => x"08",
          2463 => x"51",
          2464 => x"81",
          2465 => x"59",
          2466 => x"08",
          2467 => x"f0",
          2468 => x"82",
          2469 => x"06",
          2470 => x"05",
          2471 => x"54",
          2472 => x"3f",
          2473 => x"08",
          2474 => x"74",
          2475 => x"51",
          2476 => x"81",
          2477 => x"34",
          2478 => x"cc",
          2479 => x"0d",
          2480 => x"0d",
          2481 => x"72",
          2482 => x"56",
          2483 => x"27",
          2484 => x"98",
          2485 => x"9d",
          2486 => x"2e",
          2487 => x"53",
          2488 => x"51",
          2489 => x"81",
          2490 => x"54",
          2491 => x"08",
          2492 => x"93",
          2493 => x"80",
          2494 => x"54",
          2495 => x"81",
          2496 => x"54",
          2497 => x"74",
          2498 => x"fb",
          2499 => x"dc",
          2500 => x"81",
          2501 => x"80",
          2502 => x"38",
          2503 => x"08",
          2504 => x"38",
          2505 => x"08",
          2506 => x"38",
          2507 => x"52",
          2508 => x"d6",
          2509 => x"cc",
          2510 => x"98",
          2511 => x"11",
          2512 => x"57",
          2513 => x"74",
          2514 => x"81",
          2515 => x"0c",
          2516 => x"81",
          2517 => x"84",
          2518 => x"55",
          2519 => x"ff",
          2520 => x"54",
          2521 => x"cc",
          2522 => x"0d",
          2523 => x"0d",
          2524 => x"08",
          2525 => x"79",
          2526 => x"17",
          2527 => x"80",
          2528 => x"98",
          2529 => x"26",
          2530 => x"58",
          2531 => x"52",
          2532 => x"fd",
          2533 => x"74",
          2534 => x"08",
          2535 => x"38",
          2536 => x"08",
          2537 => x"cc",
          2538 => x"82",
          2539 => x"17",
          2540 => x"cc",
          2541 => x"c7",
          2542 => x"90",
          2543 => x"56",
          2544 => x"2e",
          2545 => x"77",
          2546 => x"81",
          2547 => x"38",
          2548 => x"98",
          2549 => x"26",
          2550 => x"56",
          2551 => x"51",
          2552 => x"80",
          2553 => x"cc",
          2554 => x"09",
          2555 => x"38",
          2556 => x"08",
          2557 => x"cc",
          2558 => x"30",
          2559 => x"80",
          2560 => x"07",
          2561 => x"08",
          2562 => x"55",
          2563 => x"ef",
          2564 => x"cc",
          2565 => x"95",
          2566 => x"08",
          2567 => x"27",
          2568 => x"98",
          2569 => x"89",
          2570 => x"85",
          2571 => x"db",
          2572 => x"81",
          2573 => x"17",
          2574 => x"89",
          2575 => x"75",
          2576 => x"ac",
          2577 => x"7a",
          2578 => x"3f",
          2579 => x"08",
          2580 => x"38",
          2581 => x"dc",
          2582 => x"2e",
          2583 => x"86",
          2584 => x"cc",
          2585 => x"dc",
          2586 => x"70",
          2587 => x"07",
          2588 => x"7c",
          2589 => x"55",
          2590 => x"f8",
          2591 => x"2e",
          2592 => x"ff",
          2593 => x"55",
          2594 => x"ff",
          2595 => x"76",
          2596 => x"3f",
          2597 => x"08",
          2598 => x"08",
          2599 => x"dc",
          2600 => x"80",
          2601 => x"55",
          2602 => x"94",
          2603 => x"2e",
          2604 => x"53",
          2605 => x"51",
          2606 => x"81",
          2607 => x"55",
          2608 => x"75",
          2609 => x"98",
          2610 => x"05",
          2611 => x"56",
          2612 => x"26",
          2613 => x"15",
          2614 => x"84",
          2615 => x"07",
          2616 => x"18",
          2617 => x"ff",
          2618 => x"2e",
          2619 => x"39",
          2620 => x"39",
          2621 => x"08",
          2622 => x"81",
          2623 => x"74",
          2624 => x"0c",
          2625 => x"04",
          2626 => x"7a",
          2627 => x"f3",
          2628 => x"dc",
          2629 => x"81",
          2630 => x"cc",
          2631 => x"38",
          2632 => x"51",
          2633 => x"81",
          2634 => x"81",
          2635 => x"b0",
          2636 => x"84",
          2637 => x"52",
          2638 => x"52",
          2639 => x"3f",
          2640 => x"39",
          2641 => x"8a",
          2642 => x"75",
          2643 => x"38",
          2644 => x"19",
          2645 => x"81",
          2646 => x"ed",
          2647 => x"dc",
          2648 => x"2e",
          2649 => x"15",
          2650 => x"70",
          2651 => x"07",
          2652 => x"53",
          2653 => x"75",
          2654 => x"0c",
          2655 => x"04",
          2656 => x"7a",
          2657 => x"58",
          2658 => x"f0",
          2659 => x"80",
          2660 => x"9f",
          2661 => x"80",
          2662 => x"90",
          2663 => x"17",
          2664 => x"aa",
          2665 => x"53",
          2666 => x"88",
          2667 => x"08",
          2668 => x"38",
          2669 => x"53",
          2670 => x"17",
          2671 => x"72",
          2672 => x"fe",
          2673 => x"08",
          2674 => x"80",
          2675 => x"16",
          2676 => x"2b",
          2677 => x"75",
          2678 => x"73",
          2679 => x"f5",
          2680 => x"dc",
          2681 => x"81",
          2682 => x"ff",
          2683 => x"81",
          2684 => x"cc",
          2685 => x"38",
          2686 => x"81",
          2687 => x"26",
          2688 => x"58",
          2689 => x"73",
          2690 => x"39",
          2691 => x"51",
          2692 => x"81",
          2693 => x"98",
          2694 => x"94",
          2695 => x"17",
          2696 => x"58",
          2697 => x"9a",
          2698 => x"81",
          2699 => x"74",
          2700 => x"98",
          2701 => x"83",
          2702 => x"b4",
          2703 => x"0c",
          2704 => x"81",
          2705 => x"8a",
          2706 => x"f8",
          2707 => x"70",
          2708 => x"08",
          2709 => x"57",
          2710 => x"0a",
          2711 => x"38",
          2712 => x"15",
          2713 => x"08",
          2714 => x"72",
          2715 => x"cb",
          2716 => x"ff",
          2717 => x"81",
          2718 => x"13",
          2719 => x"94",
          2720 => x"74",
          2721 => x"85",
          2722 => x"22",
          2723 => x"73",
          2724 => x"38",
          2725 => x"8a",
          2726 => x"05",
          2727 => x"06",
          2728 => x"8a",
          2729 => x"73",
          2730 => x"3f",
          2731 => x"08",
          2732 => x"81",
          2733 => x"cc",
          2734 => x"ff",
          2735 => x"81",
          2736 => x"ff",
          2737 => x"38",
          2738 => x"81",
          2739 => x"26",
          2740 => x"7b",
          2741 => x"98",
          2742 => x"55",
          2743 => x"94",
          2744 => x"73",
          2745 => x"3f",
          2746 => x"08",
          2747 => x"81",
          2748 => x"80",
          2749 => x"38",
          2750 => x"dc",
          2751 => x"2e",
          2752 => x"55",
          2753 => x"08",
          2754 => x"38",
          2755 => x"08",
          2756 => x"fb",
          2757 => x"dc",
          2758 => x"38",
          2759 => x"0c",
          2760 => x"51",
          2761 => x"81",
          2762 => x"98",
          2763 => x"90",
          2764 => x"16",
          2765 => x"15",
          2766 => x"74",
          2767 => x"0c",
          2768 => x"04",
          2769 => x"7b",
          2770 => x"5b",
          2771 => x"52",
          2772 => x"ac",
          2773 => x"cc",
          2774 => x"dc",
          2775 => x"ec",
          2776 => x"cc",
          2777 => x"17",
          2778 => x"51",
          2779 => x"81",
          2780 => x"54",
          2781 => x"08",
          2782 => x"81",
          2783 => x"9c",
          2784 => x"33",
          2785 => x"72",
          2786 => x"09",
          2787 => x"38",
          2788 => x"dc",
          2789 => x"72",
          2790 => x"55",
          2791 => x"53",
          2792 => x"8e",
          2793 => x"56",
          2794 => x"09",
          2795 => x"38",
          2796 => x"dc",
          2797 => x"81",
          2798 => x"fd",
          2799 => x"dc",
          2800 => x"81",
          2801 => x"80",
          2802 => x"38",
          2803 => x"09",
          2804 => x"38",
          2805 => x"81",
          2806 => x"8b",
          2807 => x"fd",
          2808 => x"9a",
          2809 => x"eb",
          2810 => x"dc",
          2811 => x"ff",
          2812 => x"70",
          2813 => x"53",
          2814 => x"09",
          2815 => x"38",
          2816 => x"eb",
          2817 => x"dc",
          2818 => x"2b",
          2819 => x"72",
          2820 => x"0c",
          2821 => x"04",
          2822 => x"77",
          2823 => x"ff",
          2824 => x"9a",
          2825 => x"55",
          2826 => x"76",
          2827 => x"53",
          2828 => x"09",
          2829 => x"38",
          2830 => x"52",
          2831 => x"eb",
          2832 => x"3d",
          2833 => x"3d",
          2834 => x"5b",
          2835 => x"08",
          2836 => x"15",
          2837 => x"81",
          2838 => x"15",
          2839 => x"51",
          2840 => x"81",
          2841 => x"58",
          2842 => x"08",
          2843 => x"9c",
          2844 => x"33",
          2845 => x"86",
          2846 => x"80",
          2847 => x"13",
          2848 => x"06",
          2849 => x"06",
          2850 => x"72",
          2851 => x"81",
          2852 => x"53",
          2853 => x"2e",
          2854 => x"53",
          2855 => x"a9",
          2856 => x"74",
          2857 => x"72",
          2858 => x"38",
          2859 => x"99",
          2860 => x"cc",
          2861 => x"06",
          2862 => x"88",
          2863 => x"06",
          2864 => x"54",
          2865 => x"a0",
          2866 => x"74",
          2867 => x"3f",
          2868 => x"08",
          2869 => x"cc",
          2870 => x"98",
          2871 => x"fa",
          2872 => x"80",
          2873 => x"0c",
          2874 => x"cc",
          2875 => x"0d",
          2876 => x"0d",
          2877 => x"57",
          2878 => x"73",
          2879 => x"3f",
          2880 => x"08",
          2881 => x"cc",
          2882 => x"98",
          2883 => x"75",
          2884 => x"3f",
          2885 => x"08",
          2886 => x"cc",
          2887 => x"a0",
          2888 => x"cc",
          2889 => x"14",
          2890 => x"db",
          2891 => x"a0",
          2892 => x"14",
          2893 => x"ac",
          2894 => x"83",
          2895 => x"81",
          2896 => x"87",
          2897 => x"fd",
          2898 => x"70",
          2899 => x"08",
          2900 => x"55",
          2901 => x"3f",
          2902 => x"08",
          2903 => x"13",
          2904 => x"73",
          2905 => x"83",
          2906 => x"3d",
          2907 => x"3d",
          2908 => x"57",
          2909 => x"89",
          2910 => x"17",
          2911 => x"81",
          2912 => x"70",
          2913 => x"55",
          2914 => x"08",
          2915 => x"81",
          2916 => x"52",
          2917 => x"a8",
          2918 => x"2e",
          2919 => x"84",
          2920 => x"52",
          2921 => x"09",
          2922 => x"38",
          2923 => x"81",
          2924 => x"81",
          2925 => x"73",
          2926 => x"55",
          2927 => x"55",
          2928 => x"c5",
          2929 => x"88",
          2930 => x"0b",
          2931 => x"9c",
          2932 => x"8b",
          2933 => x"17",
          2934 => x"08",
          2935 => x"52",
          2936 => x"81",
          2937 => x"76",
          2938 => x"51",
          2939 => x"81",
          2940 => x"86",
          2941 => x"12",
          2942 => x"3f",
          2943 => x"08",
          2944 => x"88",
          2945 => x"f3",
          2946 => x"70",
          2947 => x"80",
          2948 => x"51",
          2949 => x"af",
          2950 => x"81",
          2951 => x"dc",
          2952 => x"74",
          2953 => x"38",
          2954 => x"88",
          2955 => x"39",
          2956 => x"80",
          2957 => x"56",
          2958 => x"af",
          2959 => x"06",
          2960 => x"56",
          2961 => x"32",
          2962 => x"80",
          2963 => x"51",
          2964 => x"dc",
          2965 => x"1c",
          2966 => x"33",
          2967 => x"9f",
          2968 => x"ff",
          2969 => x"1c",
          2970 => x"7a",
          2971 => x"3f",
          2972 => x"08",
          2973 => x"39",
          2974 => x"a0",
          2975 => x"5e",
          2976 => x"52",
          2977 => x"ff",
          2978 => x"59",
          2979 => x"33",
          2980 => x"ae",
          2981 => x"06",
          2982 => x"78",
          2983 => x"81",
          2984 => x"32",
          2985 => x"9f",
          2986 => x"26",
          2987 => x"53",
          2988 => x"73",
          2989 => x"17",
          2990 => x"34",
          2991 => x"db",
          2992 => x"32",
          2993 => x"9f",
          2994 => x"54",
          2995 => x"2e",
          2996 => x"80",
          2997 => x"75",
          2998 => x"bd",
          2999 => x"7e",
          3000 => x"a0",
          3001 => x"bd",
          3002 => x"82",
          3003 => x"18",
          3004 => x"1a",
          3005 => x"a0",
          3006 => x"fc",
          3007 => x"32",
          3008 => x"80",
          3009 => x"30",
          3010 => x"71",
          3011 => x"51",
          3012 => x"55",
          3013 => x"ac",
          3014 => x"81",
          3015 => x"78",
          3016 => x"51",
          3017 => x"af",
          3018 => x"06",
          3019 => x"55",
          3020 => x"32",
          3021 => x"80",
          3022 => x"51",
          3023 => x"db",
          3024 => x"39",
          3025 => x"09",
          3026 => x"38",
          3027 => x"7c",
          3028 => x"54",
          3029 => x"a2",
          3030 => x"32",
          3031 => x"ae",
          3032 => x"72",
          3033 => x"9f",
          3034 => x"51",
          3035 => x"74",
          3036 => x"88",
          3037 => x"fe",
          3038 => x"98",
          3039 => x"80",
          3040 => x"75",
          3041 => x"81",
          3042 => x"33",
          3043 => x"51",
          3044 => x"81",
          3045 => x"80",
          3046 => x"78",
          3047 => x"81",
          3048 => x"5a",
          3049 => x"d2",
          3050 => x"cc",
          3051 => x"80",
          3052 => x"1c",
          3053 => x"27",
          3054 => x"79",
          3055 => x"74",
          3056 => x"7a",
          3057 => x"74",
          3058 => x"39",
          3059 => x"cb",
          3060 => x"fe",
          3061 => x"cc",
          3062 => x"ff",
          3063 => x"73",
          3064 => x"38",
          3065 => x"81",
          3066 => x"54",
          3067 => x"75",
          3068 => x"17",
          3069 => x"39",
          3070 => x"0c",
          3071 => x"99",
          3072 => x"54",
          3073 => x"2e",
          3074 => x"84",
          3075 => x"34",
          3076 => x"76",
          3077 => x"8b",
          3078 => x"81",
          3079 => x"56",
          3080 => x"80",
          3081 => x"1b",
          3082 => x"08",
          3083 => x"51",
          3084 => x"81",
          3085 => x"56",
          3086 => x"08",
          3087 => x"98",
          3088 => x"76",
          3089 => x"3f",
          3090 => x"08",
          3091 => x"cc",
          3092 => x"38",
          3093 => x"70",
          3094 => x"73",
          3095 => x"be",
          3096 => x"33",
          3097 => x"73",
          3098 => x"8b",
          3099 => x"83",
          3100 => x"06",
          3101 => x"73",
          3102 => x"53",
          3103 => x"51",
          3104 => x"81",
          3105 => x"80",
          3106 => x"75",
          3107 => x"f3",
          3108 => x"9f",
          3109 => x"1c",
          3110 => x"74",
          3111 => x"38",
          3112 => x"09",
          3113 => x"e7",
          3114 => x"2a",
          3115 => x"77",
          3116 => x"51",
          3117 => x"2e",
          3118 => x"81",
          3119 => x"80",
          3120 => x"38",
          3121 => x"ab",
          3122 => x"55",
          3123 => x"75",
          3124 => x"73",
          3125 => x"55",
          3126 => x"82",
          3127 => x"06",
          3128 => x"ab",
          3129 => x"33",
          3130 => x"70",
          3131 => x"55",
          3132 => x"2e",
          3133 => x"1b",
          3134 => x"06",
          3135 => x"52",
          3136 => x"db",
          3137 => x"cc",
          3138 => x"0c",
          3139 => x"74",
          3140 => x"0c",
          3141 => x"04",
          3142 => x"7c",
          3143 => x"08",
          3144 => x"55",
          3145 => x"59",
          3146 => x"81",
          3147 => x"70",
          3148 => x"33",
          3149 => x"52",
          3150 => x"2e",
          3151 => x"ee",
          3152 => x"2e",
          3153 => x"81",
          3154 => x"33",
          3155 => x"81",
          3156 => x"52",
          3157 => x"26",
          3158 => x"14",
          3159 => x"06",
          3160 => x"52",
          3161 => x"80",
          3162 => x"0b",
          3163 => x"59",
          3164 => x"7a",
          3165 => x"70",
          3166 => x"33",
          3167 => x"05",
          3168 => x"9f",
          3169 => x"53",
          3170 => x"89",
          3171 => x"70",
          3172 => x"54",
          3173 => x"12",
          3174 => x"26",
          3175 => x"12",
          3176 => x"06",
          3177 => x"30",
          3178 => x"51",
          3179 => x"2e",
          3180 => x"85",
          3181 => x"be",
          3182 => x"74",
          3183 => x"30",
          3184 => x"9f",
          3185 => x"2a",
          3186 => x"54",
          3187 => x"2e",
          3188 => x"15",
          3189 => x"55",
          3190 => x"ff",
          3191 => x"39",
          3192 => x"86",
          3193 => x"7c",
          3194 => x"51",
          3195 => x"dc",
          3196 => x"70",
          3197 => x"0c",
          3198 => x"04",
          3199 => x"78",
          3200 => x"83",
          3201 => x"0b",
          3202 => x"79",
          3203 => x"e2",
          3204 => x"55",
          3205 => x"08",
          3206 => x"84",
          3207 => x"df",
          3208 => x"dc",
          3209 => x"ff",
          3210 => x"83",
          3211 => x"d4",
          3212 => x"81",
          3213 => x"38",
          3214 => x"17",
          3215 => x"74",
          3216 => x"09",
          3217 => x"38",
          3218 => x"81",
          3219 => x"30",
          3220 => x"79",
          3221 => x"54",
          3222 => x"74",
          3223 => x"09",
          3224 => x"38",
          3225 => x"cb",
          3226 => x"ea",
          3227 => x"b1",
          3228 => x"cc",
          3229 => x"dc",
          3230 => x"2e",
          3231 => x"53",
          3232 => x"52",
          3233 => x"51",
          3234 => x"81",
          3235 => x"55",
          3236 => x"08",
          3237 => x"38",
          3238 => x"81",
          3239 => x"88",
          3240 => x"f2",
          3241 => x"02",
          3242 => x"cb",
          3243 => x"55",
          3244 => x"60",
          3245 => x"3f",
          3246 => x"08",
          3247 => x"80",
          3248 => x"cc",
          3249 => x"fc",
          3250 => x"cc",
          3251 => x"81",
          3252 => x"70",
          3253 => x"8c",
          3254 => x"2e",
          3255 => x"73",
          3256 => x"81",
          3257 => x"33",
          3258 => x"80",
          3259 => x"81",
          3260 => x"d7",
          3261 => x"dc",
          3262 => x"ff",
          3263 => x"06",
          3264 => x"98",
          3265 => x"2e",
          3266 => x"74",
          3267 => x"81",
          3268 => x"8a",
          3269 => x"ac",
          3270 => x"39",
          3271 => x"77",
          3272 => x"81",
          3273 => x"33",
          3274 => x"3f",
          3275 => x"08",
          3276 => x"70",
          3277 => x"55",
          3278 => x"86",
          3279 => x"80",
          3280 => x"74",
          3281 => x"81",
          3282 => x"8a",
          3283 => x"f4",
          3284 => x"53",
          3285 => x"fd",
          3286 => x"dc",
          3287 => x"ff",
          3288 => x"82",
          3289 => x"06",
          3290 => x"8c",
          3291 => x"58",
          3292 => x"f6",
          3293 => x"58",
          3294 => x"2e",
          3295 => x"fa",
          3296 => x"e8",
          3297 => x"cc",
          3298 => x"78",
          3299 => x"5a",
          3300 => x"90",
          3301 => x"75",
          3302 => x"38",
          3303 => x"3d",
          3304 => x"70",
          3305 => x"08",
          3306 => x"7a",
          3307 => x"38",
          3308 => x"51",
          3309 => x"81",
          3310 => x"81",
          3311 => x"81",
          3312 => x"38",
          3313 => x"83",
          3314 => x"38",
          3315 => x"84",
          3316 => x"38",
          3317 => x"81",
          3318 => x"38",
          3319 => x"db",
          3320 => x"dc",
          3321 => x"ff",
          3322 => x"72",
          3323 => x"09",
          3324 => x"d0",
          3325 => x"14",
          3326 => x"3f",
          3327 => x"08",
          3328 => x"06",
          3329 => x"38",
          3330 => x"51",
          3331 => x"81",
          3332 => x"58",
          3333 => x"0c",
          3334 => x"33",
          3335 => x"80",
          3336 => x"ff",
          3337 => x"ff",
          3338 => x"55",
          3339 => x"81",
          3340 => x"38",
          3341 => x"06",
          3342 => x"80",
          3343 => x"52",
          3344 => x"8a",
          3345 => x"80",
          3346 => x"ff",
          3347 => x"53",
          3348 => x"86",
          3349 => x"83",
          3350 => x"c5",
          3351 => x"f5",
          3352 => x"cc",
          3353 => x"dc",
          3354 => x"15",
          3355 => x"06",
          3356 => x"76",
          3357 => x"80",
          3358 => x"da",
          3359 => x"dc",
          3360 => x"ff",
          3361 => x"74",
          3362 => x"d4",
          3363 => x"dc",
          3364 => x"cc",
          3365 => x"c2",
          3366 => x"b9",
          3367 => x"cc",
          3368 => x"ff",
          3369 => x"56",
          3370 => x"83",
          3371 => x"14",
          3372 => x"71",
          3373 => x"5a",
          3374 => x"26",
          3375 => x"8a",
          3376 => x"74",
          3377 => x"ff",
          3378 => x"81",
          3379 => x"55",
          3380 => x"08",
          3381 => x"ec",
          3382 => x"cc",
          3383 => x"ff",
          3384 => x"83",
          3385 => x"74",
          3386 => x"26",
          3387 => x"57",
          3388 => x"26",
          3389 => x"57",
          3390 => x"56",
          3391 => x"82",
          3392 => x"15",
          3393 => x"0c",
          3394 => x"0c",
          3395 => x"a4",
          3396 => x"1d",
          3397 => x"54",
          3398 => x"2e",
          3399 => x"af",
          3400 => x"14",
          3401 => x"3f",
          3402 => x"08",
          3403 => x"06",
          3404 => x"72",
          3405 => x"79",
          3406 => x"80",
          3407 => x"d9",
          3408 => x"dc",
          3409 => x"15",
          3410 => x"2b",
          3411 => x"8d",
          3412 => x"2e",
          3413 => x"77",
          3414 => x"0c",
          3415 => x"76",
          3416 => x"38",
          3417 => x"70",
          3418 => x"81",
          3419 => x"53",
          3420 => x"89",
          3421 => x"56",
          3422 => x"08",
          3423 => x"38",
          3424 => x"15",
          3425 => x"8c",
          3426 => x"80",
          3427 => x"34",
          3428 => x"09",
          3429 => x"92",
          3430 => x"14",
          3431 => x"3f",
          3432 => x"08",
          3433 => x"06",
          3434 => x"2e",
          3435 => x"80",
          3436 => x"1b",
          3437 => x"db",
          3438 => x"dc",
          3439 => x"ea",
          3440 => x"cc",
          3441 => x"34",
          3442 => x"51",
          3443 => x"81",
          3444 => x"83",
          3445 => x"53",
          3446 => x"d5",
          3447 => x"06",
          3448 => x"b4",
          3449 => x"84",
          3450 => x"cc",
          3451 => x"85",
          3452 => x"09",
          3453 => x"38",
          3454 => x"51",
          3455 => x"81",
          3456 => x"86",
          3457 => x"f2",
          3458 => x"06",
          3459 => x"9c",
          3460 => x"d8",
          3461 => x"cc",
          3462 => x"0c",
          3463 => x"51",
          3464 => x"81",
          3465 => x"8c",
          3466 => x"74",
          3467 => x"f8",
          3468 => x"53",
          3469 => x"f8",
          3470 => x"15",
          3471 => x"94",
          3472 => x"56",
          3473 => x"cc",
          3474 => x"0d",
          3475 => x"0d",
          3476 => x"55",
          3477 => x"b9",
          3478 => x"53",
          3479 => x"b1",
          3480 => x"52",
          3481 => x"a9",
          3482 => x"22",
          3483 => x"57",
          3484 => x"2e",
          3485 => x"99",
          3486 => x"33",
          3487 => x"3f",
          3488 => x"08",
          3489 => x"71",
          3490 => x"74",
          3491 => x"83",
          3492 => x"78",
          3493 => x"52",
          3494 => x"cc",
          3495 => x"0d",
          3496 => x"0d",
          3497 => x"33",
          3498 => x"3d",
          3499 => x"56",
          3500 => x"8b",
          3501 => x"81",
          3502 => x"24",
          3503 => x"dc",
          3504 => x"29",
          3505 => x"05",
          3506 => x"55",
          3507 => x"84",
          3508 => x"34",
          3509 => x"80",
          3510 => x"80",
          3511 => x"75",
          3512 => x"75",
          3513 => x"38",
          3514 => x"3d",
          3515 => x"05",
          3516 => x"3f",
          3517 => x"08",
          3518 => x"dc",
          3519 => x"3d",
          3520 => x"3d",
          3521 => x"84",
          3522 => x"05",
          3523 => x"89",
          3524 => x"2e",
          3525 => x"77",
          3526 => x"54",
          3527 => x"05",
          3528 => x"84",
          3529 => x"f6",
          3530 => x"dc",
          3531 => x"81",
          3532 => x"84",
          3533 => x"5c",
          3534 => x"3d",
          3535 => x"ed",
          3536 => x"dc",
          3537 => x"81",
          3538 => x"92",
          3539 => x"d7",
          3540 => x"98",
          3541 => x"73",
          3542 => x"38",
          3543 => x"9c",
          3544 => x"80",
          3545 => x"38",
          3546 => x"95",
          3547 => x"2e",
          3548 => x"aa",
          3549 => x"ea",
          3550 => x"dc",
          3551 => x"9e",
          3552 => x"05",
          3553 => x"54",
          3554 => x"38",
          3555 => x"70",
          3556 => x"54",
          3557 => x"8e",
          3558 => x"83",
          3559 => x"88",
          3560 => x"83",
          3561 => x"83",
          3562 => x"06",
          3563 => x"80",
          3564 => x"38",
          3565 => x"51",
          3566 => x"81",
          3567 => x"56",
          3568 => x"0a",
          3569 => x"05",
          3570 => x"3f",
          3571 => x"0b",
          3572 => x"80",
          3573 => x"7a",
          3574 => x"3f",
          3575 => x"9c",
          3576 => x"d1",
          3577 => x"81",
          3578 => x"34",
          3579 => x"80",
          3580 => x"b0",
          3581 => x"54",
          3582 => x"52",
          3583 => x"05",
          3584 => x"3f",
          3585 => x"08",
          3586 => x"cc",
          3587 => x"38",
          3588 => x"82",
          3589 => x"b2",
          3590 => x"84",
          3591 => x"06",
          3592 => x"73",
          3593 => x"38",
          3594 => x"ad",
          3595 => x"2a",
          3596 => x"51",
          3597 => x"2e",
          3598 => x"81",
          3599 => x"80",
          3600 => x"87",
          3601 => x"39",
          3602 => x"51",
          3603 => x"81",
          3604 => x"7b",
          3605 => x"12",
          3606 => x"81",
          3607 => x"81",
          3608 => x"83",
          3609 => x"06",
          3610 => x"80",
          3611 => x"77",
          3612 => x"58",
          3613 => x"08",
          3614 => x"63",
          3615 => x"63",
          3616 => x"57",
          3617 => x"81",
          3618 => x"81",
          3619 => x"88",
          3620 => x"9c",
          3621 => x"d2",
          3622 => x"dc",
          3623 => x"dc",
          3624 => x"1b",
          3625 => x"0c",
          3626 => x"22",
          3627 => x"77",
          3628 => x"80",
          3629 => x"34",
          3630 => x"1a",
          3631 => x"94",
          3632 => x"85",
          3633 => x"06",
          3634 => x"80",
          3635 => x"38",
          3636 => x"08",
          3637 => x"84",
          3638 => x"cc",
          3639 => x"0c",
          3640 => x"70",
          3641 => x"52",
          3642 => x"39",
          3643 => x"51",
          3644 => x"81",
          3645 => x"57",
          3646 => x"08",
          3647 => x"38",
          3648 => x"dc",
          3649 => x"2e",
          3650 => x"83",
          3651 => x"75",
          3652 => x"74",
          3653 => x"07",
          3654 => x"54",
          3655 => x"8a",
          3656 => x"75",
          3657 => x"73",
          3658 => x"98",
          3659 => x"a9",
          3660 => x"ff",
          3661 => x"80",
          3662 => x"76",
          3663 => x"d6",
          3664 => x"dc",
          3665 => x"38",
          3666 => x"39",
          3667 => x"81",
          3668 => x"05",
          3669 => x"84",
          3670 => x"0c",
          3671 => x"81",
          3672 => x"97",
          3673 => x"f2",
          3674 => x"63",
          3675 => x"40",
          3676 => x"7e",
          3677 => x"fc",
          3678 => x"51",
          3679 => x"81",
          3680 => x"55",
          3681 => x"08",
          3682 => x"19",
          3683 => x"80",
          3684 => x"74",
          3685 => x"39",
          3686 => x"81",
          3687 => x"56",
          3688 => x"82",
          3689 => x"39",
          3690 => x"1a",
          3691 => x"82",
          3692 => x"0b",
          3693 => x"81",
          3694 => x"39",
          3695 => x"94",
          3696 => x"55",
          3697 => x"83",
          3698 => x"7b",
          3699 => x"89",
          3700 => x"08",
          3701 => x"06",
          3702 => x"81",
          3703 => x"8a",
          3704 => x"05",
          3705 => x"06",
          3706 => x"a8",
          3707 => x"38",
          3708 => x"55",
          3709 => x"19",
          3710 => x"51",
          3711 => x"81",
          3712 => x"55",
          3713 => x"ff",
          3714 => x"ff",
          3715 => x"38",
          3716 => x"0c",
          3717 => x"52",
          3718 => x"cb",
          3719 => x"cc",
          3720 => x"ff",
          3721 => x"dc",
          3722 => x"7c",
          3723 => x"57",
          3724 => x"80",
          3725 => x"1a",
          3726 => x"22",
          3727 => x"75",
          3728 => x"38",
          3729 => x"58",
          3730 => x"53",
          3731 => x"1b",
          3732 => x"88",
          3733 => x"cc",
          3734 => x"38",
          3735 => x"33",
          3736 => x"80",
          3737 => x"b0",
          3738 => x"31",
          3739 => x"27",
          3740 => x"80",
          3741 => x"52",
          3742 => x"77",
          3743 => x"7d",
          3744 => x"e0",
          3745 => x"2b",
          3746 => x"76",
          3747 => x"94",
          3748 => x"ff",
          3749 => x"71",
          3750 => x"7b",
          3751 => x"38",
          3752 => x"19",
          3753 => x"51",
          3754 => x"81",
          3755 => x"fe",
          3756 => x"53",
          3757 => x"83",
          3758 => x"b4",
          3759 => x"51",
          3760 => x"7b",
          3761 => x"08",
          3762 => x"76",
          3763 => x"08",
          3764 => x"0c",
          3765 => x"f3",
          3766 => x"75",
          3767 => x"0c",
          3768 => x"04",
          3769 => x"60",
          3770 => x"40",
          3771 => x"80",
          3772 => x"3d",
          3773 => x"77",
          3774 => x"3f",
          3775 => x"08",
          3776 => x"cc",
          3777 => x"91",
          3778 => x"74",
          3779 => x"38",
          3780 => x"b8",
          3781 => x"33",
          3782 => x"70",
          3783 => x"56",
          3784 => x"74",
          3785 => x"a4",
          3786 => x"82",
          3787 => x"34",
          3788 => x"98",
          3789 => x"91",
          3790 => x"56",
          3791 => x"94",
          3792 => x"11",
          3793 => x"76",
          3794 => x"75",
          3795 => x"80",
          3796 => x"38",
          3797 => x"70",
          3798 => x"56",
          3799 => x"fd",
          3800 => x"11",
          3801 => x"77",
          3802 => x"5c",
          3803 => x"38",
          3804 => x"88",
          3805 => x"74",
          3806 => x"52",
          3807 => x"18",
          3808 => x"51",
          3809 => x"81",
          3810 => x"55",
          3811 => x"08",
          3812 => x"ab",
          3813 => x"2e",
          3814 => x"74",
          3815 => x"95",
          3816 => x"19",
          3817 => x"08",
          3818 => x"88",
          3819 => x"55",
          3820 => x"9c",
          3821 => x"09",
          3822 => x"38",
          3823 => x"c1",
          3824 => x"cc",
          3825 => x"38",
          3826 => x"52",
          3827 => x"97",
          3828 => x"cc",
          3829 => x"fe",
          3830 => x"dc",
          3831 => x"7c",
          3832 => x"57",
          3833 => x"80",
          3834 => x"1b",
          3835 => x"22",
          3836 => x"75",
          3837 => x"38",
          3838 => x"59",
          3839 => x"53",
          3840 => x"1a",
          3841 => x"be",
          3842 => x"cc",
          3843 => x"38",
          3844 => x"08",
          3845 => x"56",
          3846 => x"9b",
          3847 => x"53",
          3848 => x"77",
          3849 => x"7d",
          3850 => x"16",
          3851 => x"3f",
          3852 => x"0b",
          3853 => x"78",
          3854 => x"80",
          3855 => x"18",
          3856 => x"08",
          3857 => x"7e",
          3858 => x"3f",
          3859 => x"08",
          3860 => x"7e",
          3861 => x"0c",
          3862 => x"19",
          3863 => x"08",
          3864 => x"84",
          3865 => x"57",
          3866 => x"27",
          3867 => x"56",
          3868 => x"52",
          3869 => x"f9",
          3870 => x"cc",
          3871 => x"38",
          3872 => x"52",
          3873 => x"83",
          3874 => x"b4",
          3875 => x"d4",
          3876 => x"81",
          3877 => x"34",
          3878 => x"7e",
          3879 => x"0c",
          3880 => x"1a",
          3881 => x"94",
          3882 => x"1b",
          3883 => x"5e",
          3884 => x"27",
          3885 => x"55",
          3886 => x"0c",
          3887 => x"90",
          3888 => x"c0",
          3889 => x"90",
          3890 => x"56",
          3891 => x"cc",
          3892 => x"0d",
          3893 => x"0d",
          3894 => x"fc",
          3895 => x"52",
          3896 => x"3f",
          3897 => x"08",
          3898 => x"cc",
          3899 => x"38",
          3900 => x"70",
          3901 => x"81",
          3902 => x"55",
          3903 => x"80",
          3904 => x"16",
          3905 => x"51",
          3906 => x"81",
          3907 => x"57",
          3908 => x"08",
          3909 => x"a4",
          3910 => x"11",
          3911 => x"55",
          3912 => x"16",
          3913 => x"08",
          3914 => x"75",
          3915 => x"e8",
          3916 => x"08",
          3917 => x"51",
          3918 => x"82",
          3919 => x"52",
          3920 => x"c9",
          3921 => x"52",
          3922 => x"c9",
          3923 => x"54",
          3924 => x"15",
          3925 => x"cc",
          3926 => x"dc",
          3927 => x"17",
          3928 => x"06",
          3929 => x"90",
          3930 => x"81",
          3931 => x"8a",
          3932 => x"fc",
          3933 => x"70",
          3934 => x"d9",
          3935 => x"cc",
          3936 => x"dc",
          3937 => x"38",
          3938 => x"05",
          3939 => x"f1",
          3940 => x"dc",
          3941 => x"81",
          3942 => x"87",
          3943 => x"cc",
          3944 => x"72",
          3945 => x"0c",
          3946 => x"04",
          3947 => x"84",
          3948 => x"e4",
          3949 => x"80",
          3950 => x"cc",
          3951 => x"38",
          3952 => x"08",
          3953 => x"34",
          3954 => x"81",
          3955 => x"83",
          3956 => x"ef",
          3957 => x"53",
          3958 => x"05",
          3959 => x"51",
          3960 => x"81",
          3961 => x"55",
          3962 => x"08",
          3963 => x"76",
          3964 => x"93",
          3965 => x"51",
          3966 => x"81",
          3967 => x"55",
          3968 => x"08",
          3969 => x"80",
          3970 => x"70",
          3971 => x"56",
          3972 => x"89",
          3973 => x"94",
          3974 => x"b2",
          3975 => x"05",
          3976 => x"2a",
          3977 => x"51",
          3978 => x"80",
          3979 => x"76",
          3980 => x"52",
          3981 => x"3f",
          3982 => x"08",
          3983 => x"8e",
          3984 => x"cc",
          3985 => x"09",
          3986 => x"38",
          3987 => x"81",
          3988 => x"93",
          3989 => x"e4",
          3990 => x"6f",
          3991 => x"7a",
          3992 => x"9e",
          3993 => x"05",
          3994 => x"51",
          3995 => x"81",
          3996 => x"57",
          3997 => x"08",
          3998 => x"7b",
          3999 => x"94",
          4000 => x"55",
          4001 => x"73",
          4002 => x"ed",
          4003 => x"93",
          4004 => x"55",
          4005 => x"81",
          4006 => x"57",
          4007 => x"08",
          4008 => x"68",
          4009 => x"c9",
          4010 => x"dc",
          4011 => x"81",
          4012 => x"82",
          4013 => x"52",
          4014 => x"a3",
          4015 => x"cc",
          4016 => x"52",
          4017 => x"b8",
          4018 => x"cc",
          4019 => x"dc",
          4020 => x"a2",
          4021 => x"74",
          4022 => x"3f",
          4023 => x"08",
          4024 => x"cc",
          4025 => x"69",
          4026 => x"d9",
          4027 => x"81",
          4028 => x"2e",
          4029 => x"52",
          4030 => x"cf",
          4031 => x"cc",
          4032 => x"dc",
          4033 => x"2e",
          4034 => x"84",
          4035 => x"06",
          4036 => x"57",
          4037 => x"76",
          4038 => x"9e",
          4039 => x"05",
          4040 => x"dc",
          4041 => x"90",
          4042 => x"81",
          4043 => x"56",
          4044 => x"80",
          4045 => x"02",
          4046 => x"81",
          4047 => x"70",
          4048 => x"56",
          4049 => x"81",
          4050 => x"78",
          4051 => x"38",
          4052 => x"99",
          4053 => x"81",
          4054 => x"18",
          4055 => x"18",
          4056 => x"58",
          4057 => x"33",
          4058 => x"ee",
          4059 => x"6f",
          4060 => x"af",
          4061 => x"8d",
          4062 => x"2e",
          4063 => x"8a",
          4064 => x"6f",
          4065 => x"af",
          4066 => x"0b",
          4067 => x"33",
          4068 => x"81",
          4069 => x"70",
          4070 => x"52",
          4071 => x"56",
          4072 => x"8d",
          4073 => x"70",
          4074 => x"51",
          4075 => x"f5",
          4076 => x"54",
          4077 => x"a7",
          4078 => x"74",
          4079 => x"38",
          4080 => x"73",
          4081 => x"81",
          4082 => x"81",
          4083 => x"39",
          4084 => x"81",
          4085 => x"74",
          4086 => x"81",
          4087 => x"91",
          4088 => x"6e",
          4089 => x"59",
          4090 => x"7a",
          4091 => x"5c",
          4092 => x"26",
          4093 => x"7a",
          4094 => x"dc",
          4095 => x"3d",
          4096 => x"3d",
          4097 => x"8d",
          4098 => x"54",
          4099 => x"55",
          4100 => x"81",
          4101 => x"53",
          4102 => x"08",
          4103 => x"91",
          4104 => x"72",
          4105 => x"8c",
          4106 => x"73",
          4107 => x"38",
          4108 => x"70",
          4109 => x"81",
          4110 => x"57",
          4111 => x"73",
          4112 => x"08",
          4113 => x"94",
          4114 => x"75",
          4115 => x"97",
          4116 => x"11",
          4117 => x"2b",
          4118 => x"73",
          4119 => x"38",
          4120 => x"16",
          4121 => x"93",
          4122 => x"cc",
          4123 => x"78",
          4124 => x"55",
          4125 => x"83",
          4126 => x"cc",
          4127 => x"96",
          4128 => x"70",
          4129 => x"94",
          4130 => x"71",
          4131 => x"08",
          4132 => x"53",
          4133 => x"15",
          4134 => x"a6",
          4135 => x"74",
          4136 => x"3f",
          4137 => x"08",
          4138 => x"cc",
          4139 => x"81",
          4140 => x"dc",
          4141 => x"2e",
          4142 => x"81",
          4143 => x"88",
          4144 => x"98",
          4145 => x"80",
          4146 => x"38",
          4147 => x"80",
          4148 => x"77",
          4149 => x"08",
          4150 => x"0c",
          4151 => x"70",
          4152 => x"81",
          4153 => x"5a",
          4154 => x"2e",
          4155 => x"52",
          4156 => x"f9",
          4157 => x"cc",
          4158 => x"dc",
          4159 => x"38",
          4160 => x"08",
          4161 => x"73",
          4162 => x"c7",
          4163 => x"dc",
          4164 => x"73",
          4165 => x"38",
          4166 => x"af",
          4167 => x"73",
          4168 => x"27",
          4169 => x"98",
          4170 => x"a0",
          4171 => x"08",
          4172 => x"0c",
          4173 => x"06",
          4174 => x"2e",
          4175 => x"52",
          4176 => x"a3",
          4177 => x"cc",
          4178 => x"82",
          4179 => x"34",
          4180 => x"c4",
          4181 => x"91",
          4182 => x"53",
          4183 => x"89",
          4184 => x"cc",
          4185 => x"94",
          4186 => x"8c",
          4187 => x"27",
          4188 => x"8c",
          4189 => x"15",
          4190 => x"07",
          4191 => x"16",
          4192 => x"ff",
          4193 => x"80",
          4194 => x"77",
          4195 => x"2e",
          4196 => x"9c",
          4197 => x"53",
          4198 => x"cc",
          4199 => x"0d",
          4200 => x"0d",
          4201 => x"54",
          4202 => x"81",
          4203 => x"53",
          4204 => x"05",
          4205 => x"84",
          4206 => x"e7",
          4207 => x"cc",
          4208 => x"dc",
          4209 => x"ea",
          4210 => x"0c",
          4211 => x"51",
          4212 => x"81",
          4213 => x"55",
          4214 => x"08",
          4215 => x"ab",
          4216 => x"98",
          4217 => x"80",
          4218 => x"38",
          4219 => x"70",
          4220 => x"81",
          4221 => x"57",
          4222 => x"ad",
          4223 => x"08",
          4224 => x"d3",
          4225 => x"dc",
          4226 => x"17",
          4227 => x"86",
          4228 => x"17",
          4229 => x"75",
          4230 => x"3f",
          4231 => x"08",
          4232 => x"2e",
          4233 => x"85",
          4234 => x"86",
          4235 => x"2e",
          4236 => x"76",
          4237 => x"73",
          4238 => x"0c",
          4239 => x"04",
          4240 => x"76",
          4241 => x"05",
          4242 => x"53",
          4243 => x"81",
          4244 => x"87",
          4245 => x"cc",
          4246 => x"86",
          4247 => x"fb",
          4248 => x"79",
          4249 => x"05",
          4250 => x"56",
          4251 => x"3f",
          4252 => x"08",
          4253 => x"cc",
          4254 => x"38",
          4255 => x"81",
          4256 => x"52",
          4257 => x"f8",
          4258 => x"cc",
          4259 => x"ca",
          4260 => x"cc",
          4261 => x"51",
          4262 => x"81",
          4263 => x"53",
          4264 => x"08",
          4265 => x"81",
          4266 => x"80",
          4267 => x"81",
          4268 => x"a6",
          4269 => x"73",
          4270 => x"3f",
          4271 => x"51",
          4272 => x"81",
          4273 => x"84",
          4274 => x"70",
          4275 => x"2c",
          4276 => x"cc",
          4277 => x"51",
          4278 => x"81",
          4279 => x"87",
          4280 => x"ee",
          4281 => x"57",
          4282 => x"3d",
          4283 => x"3d",
          4284 => x"af",
          4285 => x"cc",
          4286 => x"dc",
          4287 => x"38",
          4288 => x"51",
          4289 => x"81",
          4290 => x"55",
          4291 => x"08",
          4292 => x"80",
          4293 => x"70",
          4294 => x"58",
          4295 => x"85",
          4296 => x"8d",
          4297 => x"2e",
          4298 => x"52",
          4299 => x"be",
          4300 => x"dc",
          4301 => x"3d",
          4302 => x"3d",
          4303 => x"55",
          4304 => x"92",
          4305 => x"52",
          4306 => x"de",
          4307 => x"dc",
          4308 => x"81",
          4309 => x"82",
          4310 => x"74",
          4311 => x"98",
          4312 => x"11",
          4313 => x"59",
          4314 => x"75",
          4315 => x"38",
          4316 => x"81",
          4317 => x"5b",
          4318 => x"82",
          4319 => x"39",
          4320 => x"08",
          4321 => x"59",
          4322 => x"09",
          4323 => x"38",
          4324 => x"57",
          4325 => x"3d",
          4326 => x"c1",
          4327 => x"dc",
          4328 => x"2e",
          4329 => x"dc",
          4330 => x"2e",
          4331 => x"dc",
          4332 => x"70",
          4333 => x"08",
          4334 => x"7a",
          4335 => x"7f",
          4336 => x"54",
          4337 => x"77",
          4338 => x"80",
          4339 => x"15",
          4340 => x"cc",
          4341 => x"75",
          4342 => x"52",
          4343 => x"52",
          4344 => x"8d",
          4345 => x"cc",
          4346 => x"dc",
          4347 => x"d6",
          4348 => x"33",
          4349 => x"1a",
          4350 => x"54",
          4351 => x"09",
          4352 => x"38",
          4353 => x"ff",
          4354 => x"81",
          4355 => x"83",
          4356 => x"70",
          4357 => x"25",
          4358 => x"59",
          4359 => x"9b",
          4360 => x"51",
          4361 => x"3f",
          4362 => x"08",
          4363 => x"70",
          4364 => x"25",
          4365 => x"59",
          4366 => x"75",
          4367 => x"7a",
          4368 => x"ff",
          4369 => x"7c",
          4370 => x"90",
          4371 => x"11",
          4372 => x"56",
          4373 => x"15",
          4374 => x"dc",
          4375 => x"3d",
          4376 => x"3d",
          4377 => x"3d",
          4378 => x"70",
          4379 => x"dd",
          4380 => x"cc",
          4381 => x"dc",
          4382 => x"a8",
          4383 => x"33",
          4384 => x"a0",
          4385 => x"33",
          4386 => x"70",
          4387 => x"55",
          4388 => x"73",
          4389 => x"8e",
          4390 => x"08",
          4391 => x"18",
          4392 => x"80",
          4393 => x"38",
          4394 => x"08",
          4395 => x"08",
          4396 => x"c4",
          4397 => x"dc",
          4398 => x"88",
          4399 => x"80",
          4400 => x"17",
          4401 => x"51",
          4402 => x"3f",
          4403 => x"08",
          4404 => x"81",
          4405 => x"81",
          4406 => x"cc",
          4407 => x"09",
          4408 => x"38",
          4409 => x"39",
          4410 => x"77",
          4411 => x"cc",
          4412 => x"08",
          4413 => x"98",
          4414 => x"81",
          4415 => x"52",
          4416 => x"bd",
          4417 => x"cc",
          4418 => x"17",
          4419 => x"0c",
          4420 => x"80",
          4421 => x"73",
          4422 => x"75",
          4423 => x"38",
          4424 => x"34",
          4425 => x"81",
          4426 => x"89",
          4427 => x"e2",
          4428 => x"53",
          4429 => x"a4",
          4430 => x"3d",
          4431 => x"3f",
          4432 => x"08",
          4433 => x"cc",
          4434 => x"38",
          4435 => x"3d",
          4436 => x"3d",
          4437 => x"d1",
          4438 => x"dc",
          4439 => x"81",
          4440 => x"81",
          4441 => x"80",
          4442 => x"70",
          4443 => x"81",
          4444 => x"56",
          4445 => x"81",
          4446 => x"98",
          4447 => x"74",
          4448 => x"38",
          4449 => x"05",
          4450 => x"06",
          4451 => x"55",
          4452 => x"38",
          4453 => x"51",
          4454 => x"81",
          4455 => x"74",
          4456 => x"81",
          4457 => x"56",
          4458 => x"80",
          4459 => x"54",
          4460 => x"08",
          4461 => x"2e",
          4462 => x"73",
          4463 => x"cc",
          4464 => x"52",
          4465 => x"52",
          4466 => x"3f",
          4467 => x"08",
          4468 => x"cc",
          4469 => x"38",
          4470 => x"08",
          4471 => x"cc",
          4472 => x"dc",
          4473 => x"81",
          4474 => x"86",
          4475 => x"80",
          4476 => x"dc",
          4477 => x"2e",
          4478 => x"dc",
          4479 => x"c0",
          4480 => x"ce",
          4481 => x"dc",
          4482 => x"dc",
          4483 => x"70",
          4484 => x"08",
          4485 => x"51",
          4486 => x"80",
          4487 => x"73",
          4488 => x"38",
          4489 => x"52",
          4490 => x"95",
          4491 => x"cc",
          4492 => x"8c",
          4493 => x"ff",
          4494 => x"81",
          4495 => x"55",
          4496 => x"cc",
          4497 => x"0d",
          4498 => x"0d",
          4499 => x"3d",
          4500 => x"9a",
          4501 => x"cb",
          4502 => x"cc",
          4503 => x"dc",
          4504 => x"b0",
          4505 => x"69",
          4506 => x"70",
          4507 => x"97",
          4508 => x"cc",
          4509 => x"dc",
          4510 => x"38",
          4511 => x"94",
          4512 => x"cc",
          4513 => x"09",
          4514 => x"88",
          4515 => x"df",
          4516 => x"85",
          4517 => x"51",
          4518 => x"74",
          4519 => x"78",
          4520 => x"8a",
          4521 => x"57",
          4522 => x"81",
          4523 => x"75",
          4524 => x"dc",
          4525 => x"38",
          4526 => x"dc",
          4527 => x"2e",
          4528 => x"83",
          4529 => x"81",
          4530 => x"ff",
          4531 => x"06",
          4532 => x"54",
          4533 => x"73",
          4534 => x"81",
          4535 => x"52",
          4536 => x"a4",
          4537 => x"cc",
          4538 => x"dc",
          4539 => x"9a",
          4540 => x"a0",
          4541 => x"51",
          4542 => x"3f",
          4543 => x"0b",
          4544 => x"78",
          4545 => x"bf",
          4546 => x"88",
          4547 => x"80",
          4548 => x"ff",
          4549 => x"75",
          4550 => x"11",
          4551 => x"f8",
          4552 => x"78",
          4553 => x"80",
          4554 => x"ff",
          4555 => x"78",
          4556 => x"80",
          4557 => x"7f",
          4558 => x"d4",
          4559 => x"c9",
          4560 => x"54",
          4561 => x"15",
          4562 => x"cb",
          4563 => x"dc",
          4564 => x"81",
          4565 => x"b2",
          4566 => x"b2",
          4567 => x"96",
          4568 => x"b5",
          4569 => x"53",
          4570 => x"51",
          4571 => x"64",
          4572 => x"8b",
          4573 => x"54",
          4574 => x"15",
          4575 => x"ff",
          4576 => x"81",
          4577 => x"54",
          4578 => x"53",
          4579 => x"51",
          4580 => x"3f",
          4581 => x"cc",
          4582 => x"0d",
          4583 => x"0d",
          4584 => x"05",
          4585 => x"3f",
          4586 => x"3d",
          4587 => x"52",
          4588 => x"d5",
          4589 => x"dc",
          4590 => x"81",
          4591 => x"82",
          4592 => x"4d",
          4593 => x"52",
          4594 => x"52",
          4595 => x"3f",
          4596 => x"08",
          4597 => x"cc",
          4598 => x"38",
          4599 => x"05",
          4600 => x"06",
          4601 => x"73",
          4602 => x"a0",
          4603 => x"08",
          4604 => x"ff",
          4605 => x"ff",
          4606 => x"ac",
          4607 => x"92",
          4608 => x"54",
          4609 => x"3f",
          4610 => x"52",
          4611 => x"f7",
          4612 => x"cc",
          4613 => x"dc",
          4614 => x"38",
          4615 => x"09",
          4616 => x"38",
          4617 => x"08",
          4618 => x"88",
          4619 => x"39",
          4620 => x"08",
          4621 => x"81",
          4622 => x"38",
          4623 => x"b1",
          4624 => x"cc",
          4625 => x"dc",
          4626 => x"c8",
          4627 => x"93",
          4628 => x"ff",
          4629 => x"8d",
          4630 => x"b4",
          4631 => x"af",
          4632 => x"17",
          4633 => x"33",
          4634 => x"70",
          4635 => x"55",
          4636 => x"38",
          4637 => x"54",
          4638 => x"34",
          4639 => x"0b",
          4640 => x"8b",
          4641 => x"84",
          4642 => x"06",
          4643 => x"73",
          4644 => x"e5",
          4645 => x"2e",
          4646 => x"75",
          4647 => x"c6",
          4648 => x"dc",
          4649 => x"78",
          4650 => x"bb",
          4651 => x"81",
          4652 => x"80",
          4653 => x"38",
          4654 => x"08",
          4655 => x"ff",
          4656 => x"81",
          4657 => x"79",
          4658 => x"58",
          4659 => x"dc",
          4660 => x"c0",
          4661 => x"33",
          4662 => x"2e",
          4663 => x"99",
          4664 => x"75",
          4665 => x"c6",
          4666 => x"54",
          4667 => x"15",
          4668 => x"81",
          4669 => x"9c",
          4670 => x"c8",
          4671 => x"dc",
          4672 => x"81",
          4673 => x"8c",
          4674 => x"ff",
          4675 => x"81",
          4676 => x"55",
          4677 => x"cc",
          4678 => x"0d",
          4679 => x"0d",
          4680 => x"05",
          4681 => x"05",
          4682 => x"33",
          4683 => x"53",
          4684 => x"05",
          4685 => x"51",
          4686 => x"81",
          4687 => x"55",
          4688 => x"08",
          4689 => x"78",
          4690 => x"95",
          4691 => x"51",
          4692 => x"81",
          4693 => x"55",
          4694 => x"08",
          4695 => x"80",
          4696 => x"81",
          4697 => x"86",
          4698 => x"38",
          4699 => x"61",
          4700 => x"12",
          4701 => x"7a",
          4702 => x"51",
          4703 => x"74",
          4704 => x"78",
          4705 => x"83",
          4706 => x"51",
          4707 => x"3f",
          4708 => x"08",
          4709 => x"dc",
          4710 => x"3d",
          4711 => x"3d",
          4712 => x"82",
          4713 => x"d0",
          4714 => x"3d",
          4715 => x"3f",
          4716 => x"08",
          4717 => x"cc",
          4718 => x"38",
          4719 => x"52",
          4720 => x"05",
          4721 => x"3f",
          4722 => x"08",
          4723 => x"cc",
          4724 => x"02",
          4725 => x"33",
          4726 => x"54",
          4727 => x"a6",
          4728 => x"22",
          4729 => x"71",
          4730 => x"53",
          4731 => x"51",
          4732 => x"3f",
          4733 => x"0b",
          4734 => x"76",
          4735 => x"b8",
          4736 => x"cc",
          4737 => x"81",
          4738 => x"93",
          4739 => x"ea",
          4740 => x"6b",
          4741 => x"53",
          4742 => x"05",
          4743 => x"51",
          4744 => x"81",
          4745 => x"81",
          4746 => x"30",
          4747 => x"cc",
          4748 => x"25",
          4749 => x"79",
          4750 => x"85",
          4751 => x"75",
          4752 => x"73",
          4753 => x"f9",
          4754 => x"80",
          4755 => x"8d",
          4756 => x"54",
          4757 => x"3f",
          4758 => x"08",
          4759 => x"cc",
          4760 => x"38",
          4761 => x"51",
          4762 => x"81",
          4763 => x"57",
          4764 => x"08",
          4765 => x"dc",
          4766 => x"dc",
          4767 => x"5b",
          4768 => x"18",
          4769 => x"18",
          4770 => x"74",
          4771 => x"81",
          4772 => x"78",
          4773 => x"8b",
          4774 => x"54",
          4775 => x"75",
          4776 => x"38",
          4777 => x"1b",
          4778 => x"55",
          4779 => x"2e",
          4780 => x"39",
          4781 => x"09",
          4782 => x"38",
          4783 => x"80",
          4784 => x"70",
          4785 => x"25",
          4786 => x"80",
          4787 => x"38",
          4788 => x"bc",
          4789 => x"11",
          4790 => x"ff",
          4791 => x"81",
          4792 => x"57",
          4793 => x"08",
          4794 => x"70",
          4795 => x"80",
          4796 => x"83",
          4797 => x"80",
          4798 => x"84",
          4799 => x"a7",
          4800 => x"b4",
          4801 => x"ad",
          4802 => x"dc",
          4803 => x"0c",
          4804 => x"cc",
          4805 => x"0d",
          4806 => x"0d",
          4807 => x"3d",
          4808 => x"52",
          4809 => x"ce",
          4810 => x"dc",
          4811 => x"dc",
          4812 => x"54",
          4813 => x"08",
          4814 => x"8b",
          4815 => x"8b",
          4816 => x"59",
          4817 => x"3f",
          4818 => x"33",
          4819 => x"06",
          4820 => x"57",
          4821 => x"81",
          4822 => x"58",
          4823 => x"06",
          4824 => x"4e",
          4825 => x"ff",
          4826 => x"81",
          4827 => x"80",
          4828 => x"6c",
          4829 => x"53",
          4830 => x"ae",
          4831 => x"dc",
          4832 => x"2e",
          4833 => x"88",
          4834 => x"6d",
          4835 => x"55",
          4836 => x"dc",
          4837 => x"ff",
          4838 => x"83",
          4839 => x"51",
          4840 => x"26",
          4841 => x"15",
          4842 => x"ff",
          4843 => x"80",
          4844 => x"87",
          4845 => x"9c",
          4846 => x"74",
          4847 => x"38",
          4848 => x"cd",
          4849 => x"ae",
          4850 => x"dc",
          4851 => x"38",
          4852 => x"27",
          4853 => x"89",
          4854 => x"8b",
          4855 => x"27",
          4856 => x"55",
          4857 => x"81",
          4858 => x"8f",
          4859 => x"2a",
          4860 => x"70",
          4861 => x"34",
          4862 => x"74",
          4863 => x"05",
          4864 => x"17",
          4865 => x"70",
          4866 => x"52",
          4867 => x"73",
          4868 => x"c8",
          4869 => x"33",
          4870 => x"73",
          4871 => x"81",
          4872 => x"80",
          4873 => x"02",
          4874 => x"76",
          4875 => x"51",
          4876 => x"2e",
          4877 => x"87",
          4878 => x"57",
          4879 => x"79",
          4880 => x"80",
          4881 => x"70",
          4882 => x"ba",
          4883 => x"dc",
          4884 => x"81",
          4885 => x"80",
          4886 => x"52",
          4887 => x"bf",
          4888 => x"dc",
          4889 => x"81",
          4890 => x"8d",
          4891 => x"c4",
          4892 => x"e5",
          4893 => x"c6",
          4894 => x"cc",
          4895 => x"09",
          4896 => x"cc",
          4897 => x"76",
          4898 => x"c4",
          4899 => x"74",
          4900 => x"b0",
          4901 => x"cc",
          4902 => x"dc",
          4903 => x"38",
          4904 => x"dc",
          4905 => x"67",
          4906 => x"db",
          4907 => x"88",
          4908 => x"34",
          4909 => x"52",
          4910 => x"ab",
          4911 => x"54",
          4912 => x"15",
          4913 => x"ff",
          4914 => x"81",
          4915 => x"54",
          4916 => x"81",
          4917 => x"9c",
          4918 => x"f2",
          4919 => x"62",
          4920 => x"80",
          4921 => x"93",
          4922 => x"55",
          4923 => x"5e",
          4924 => x"3f",
          4925 => x"08",
          4926 => x"cc",
          4927 => x"38",
          4928 => x"58",
          4929 => x"38",
          4930 => x"97",
          4931 => x"08",
          4932 => x"38",
          4933 => x"70",
          4934 => x"81",
          4935 => x"55",
          4936 => x"87",
          4937 => x"39",
          4938 => x"90",
          4939 => x"82",
          4940 => x"8a",
          4941 => x"89",
          4942 => x"7f",
          4943 => x"56",
          4944 => x"3f",
          4945 => x"06",
          4946 => x"72",
          4947 => x"81",
          4948 => x"05",
          4949 => x"7c",
          4950 => x"55",
          4951 => x"27",
          4952 => x"16",
          4953 => x"83",
          4954 => x"76",
          4955 => x"80",
          4956 => x"79",
          4957 => x"99",
          4958 => x"7f",
          4959 => x"14",
          4960 => x"83",
          4961 => x"81",
          4962 => x"81",
          4963 => x"38",
          4964 => x"08",
          4965 => x"95",
          4966 => x"cc",
          4967 => x"81",
          4968 => x"7b",
          4969 => x"06",
          4970 => x"39",
          4971 => x"56",
          4972 => x"09",
          4973 => x"b9",
          4974 => x"80",
          4975 => x"80",
          4976 => x"78",
          4977 => x"7a",
          4978 => x"38",
          4979 => x"73",
          4980 => x"81",
          4981 => x"ff",
          4982 => x"74",
          4983 => x"ff",
          4984 => x"81",
          4985 => x"58",
          4986 => x"08",
          4987 => x"74",
          4988 => x"16",
          4989 => x"73",
          4990 => x"39",
          4991 => x"7e",
          4992 => x"0c",
          4993 => x"2e",
          4994 => x"88",
          4995 => x"8c",
          4996 => x"1a",
          4997 => x"07",
          4998 => x"1b",
          4999 => x"08",
          5000 => x"16",
          5001 => x"75",
          5002 => x"38",
          5003 => x"90",
          5004 => x"15",
          5005 => x"54",
          5006 => x"34",
          5007 => x"81",
          5008 => x"90",
          5009 => x"e9",
          5010 => x"6d",
          5011 => x"80",
          5012 => x"9d",
          5013 => x"5c",
          5014 => x"3f",
          5015 => x"0b",
          5016 => x"08",
          5017 => x"38",
          5018 => x"08",
          5019 => x"dc",
          5020 => x"08",
          5021 => x"80",
          5022 => x"80",
          5023 => x"dc",
          5024 => x"ff",
          5025 => x"52",
          5026 => x"a0",
          5027 => x"dc",
          5028 => x"ff",
          5029 => x"06",
          5030 => x"56",
          5031 => x"38",
          5032 => x"70",
          5033 => x"55",
          5034 => x"8b",
          5035 => x"3d",
          5036 => x"83",
          5037 => x"ff",
          5038 => x"81",
          5039 => x"99",
          5040 => x"74",
          5041 => x"38",
          5042 => x"80",
          5043 => x"ff",
          5044 => x"55",
          5045 => x"83",
          5046 => x"78",
          5047 => x"38",
          5048 => x"26",
          5049 => x"81",
          5050 => x"8b",
          5051 => x"79",
          5052 => x"80",
          5053 => x"93",
          5054 => x"39",
          5055 => x"6e",
          5056 => x"89",
          5057 => x"48",
          5058 => x"83",
          5059 => x"61",
          5060 => x"25",
          5061 => x"55",
          5062 => x"8a",
          5063 => x"3d",
          5064 => x"81",
          5065 => x"ff",
          5066 => x"81",
          5067 => x"cc",
          5068 => x"38",
          5069 => x"70",
          5070 => x"dc",
          5071 => x"56",
          5072 => x"38",
          5073 => x"55",
          5074 => x"75",
          5075 => x"38",
          5076 => x"70",
          5077 => x"ff",
          5078 => x"83",
          5079 => x"78",
          5080 => x"89",
          5081 => x"81",
          5082 => x"06",
          5083 => x"80",
          5084 => x"77",
          5085 => x"74",
          5086 => x"8d",
          5087 => x"06",
          5088 => x"2e",
          5089 => x"77",
          5090 => x"93",
          5091 => x"74",
          5092 => x"cb",
          5093 => x"7d",
          5094 => x"81",
          5095 => x"38",
          5096 => x"66",
          5097 => x"81",
          5098 => x"c0",
          5099 => x"74",
          5100 => x"38",
          5101 => x"98",
          5102 => x"c0",
          5103 => x"82",
          5104 => x"57",
          5105 => x"80",
          5106 => x"76",
          5107 => x"38",
          5108 => x"51",
          5109 => x"3f",
          5110 => x"08",
          5111 => x"87",
          5112 => x"2a",
          5113 => x"5c",
          5114 => x"dc",
          5115 => x"80",
          5116 => x"44",
          5117 => x"0a",
          5118 => x"ec",
          5119 => x"39",
          5120 => x"66",
          5121 => x"81",
          5122 => x"b0",
          5123 => x"74",
          5124 => x"38",
          5125 => x"98",
          5126 => x"b0",
          5127 => x"82",
          5128 => x"57",
          5129 => x"80",
          5130 => x"76",
          5131 => x"38",
          5132 => x"51",
          5133 => x"3f",
          5134 => x"08",
          5135 => x"57",
          5136 => x"08",
          5137 => x"96",
          5138 => x"81",
          5139 => x"10",
          5140 => x"08",
          5141 => x"72",
          5142 => x"59",
          5143 => x"ff",
          5144 => x"5d",
          5145 => x"44",
          5146 => x"11",
          5147 => x"70",
          5148 => x"71",
          5149 => x"06",
          5150 => x"52",
          5151 => x"40",
          5152 => x"09",
          5153 => x"38",
          5154 => x"18",
          5155 => x"39",
          5156 => x"79",
          5157 => x"70",
          5158 => x"58",
          5159 => x"76",
          5160 => x"38",
          5161 => x"7d",
          5162 => x"70",
          5163 => x"55",
          5164 => x"3f",
          5165 => x"08",
          5166 => x"2e",
          5167 => x"9b",
          5168 => x"cc",
          5169 => x"f5",
          5170 => x"38",
          5171 => x"38",
          5172 => x"59",
          5173 => x"38",
          5174 => x"7d",
          5175 => x"81",
          5176 => x"38",
          5177 => x"0b",
          5178 => x"08",
          5179 => x"78",
          5180 => x"1a",
          5181 => x"c0",
          5182 => x"74",
          5183 => x"39",
          5184 => x"55",
          5185 => x"8f",
          5186 => x"fd",
          5187 => x"dc",
          5188 => x"f5",
          5189 => x"78",
          5190 => x"79",
          5191 => x"80",
          5192 => x"f1",
          5193 => x"39",
          5194 => x"81",
          5195 => x"06",
          5196 => x"55",
          5197 => x"27",
          5198 => x"81",
          5199 => x"56",
          5200 => x"38",
          5201 => x"80",
          5202 => x"ff",
          5203 => x"8b",
          5204 => x"d8",
          5205 => x"ff",
          5206 => x"84",
          5207 => x"1b",
          5208 => x"b3",
          5209 => x"1c",
          5210 => x"ff",
          5211 => x"8e",
          5212 => x"a1",
          5213 => x"0b",
          5214 => x"7d",
          5215 => x"30",
          5216 => x"84",
          5217 => x"51",
          5218 => x"51",
          5219 => x"3f",
          5220 => x"83",
          5221 => x"90",
          5222 => x"ff",
          5223 => x"93",
          5224 => x"a0",
          5225 => x"39",
          5226 => x"1b",
          5227 => x"85",
          5228 => x"95",
          5229 => x"52",
          5230 => x"ff",
          5231 => x"81",
          5232 => x"1b",
          5233 => x"cf",
          5234 => x"9c",
          5235 => x"a0",
          5236 => x"83",
          5237 => x"06",
          5238 => x"82",
          5239 => x"52",
          5240 => x"51",
          5241 => x"3f",
          5242 => x"1b",
          5243 => x"c5",
          5244 => x"ac",
          5245 => x"a0",
          5246 => x"52",
          5247 => x"ff",
          5248 => x"86",
          5249 => x"51",
          5250 => x"3f",
          5251 => x"80",
          5252 => x"a9",
          5253 => x"1c",
          5254 => x"81",
          5255 => x"80",
          5256 => x"ae",
          5257 => x"b2",
          5258 => x"1b",
          5259 => x"85",
          5260 => x"ff",
          5261 => x"96",
          5262 => x"9f",
          5263 => x"80",
          5264 => x"34",
          5265 => x"1c",
          5266 => x"81",
          5267 => x"ab",
          5268 => x"a0",
          5269 => x"d4",
          5270 => x"fe",
          5271 => x"59",
          5272 => x"3f",
          5273 => x"53",
          5274 => x"51",
          5275 => x"3f",
          5276 => x"dc",
          5277 => x"e7",
          5278 => x"2e",
          5279 => x"80",
          5280 => x"54",
          5281 => x"53",
          5282 => x"51",
          5283 => x"3f",
          5284 => x"80",
          5285 => x"ff",
          5286 => x"84",
          5287 => x"d2",
          5288 => x"ff",
          5289 => x"86",
          5290 => x"f2",
          5291 => x"1b",
          5292 => x"81",
          5293 => x"52",
          5294 => x"51",
          5295 => x"3f",
          5296 => x"ec",
          5297 => x"9e",
          5298 => x"d4",
          5299 => x"51",
          5300 => x"3f",
          5301 => x"87",
          5302 => x"52",
          5303 => x"9a",
          5304 => x"54",
          5305 => x"7a",
          5306 => x"ff",
          5307 => x"65",
          5308 => x"7a",
          5309 => x"8f",
          5310 => x"80",
          5311 => x"2e",
          5312 => x"9a",
          5313 => x"7a",
          5314 => x"a9",
          5315 => x"84",
          5316 => x"9e",
          5317 => x"0a",
          5318 => x"51",
          5319 => x"ff",
          5320 => x"7d",
          5321 => x"38",
          5322 => x"52",
          5323 => x"9e",
          5324 => x"55",
          5325 => x"62",
          5326 => x"74",
          5327 => x"75",
          5328 => x"7e",
          5329 => x"fe",
          5330 => x"cc",
          5331 => x"38",
          5332 => x"81",
          5333 => x"52",
          5334 => x"9e",
          5335 => x"16",
          5336 => x"56",
          5337 => x"38",
          5338 => x"77",
          5339 => x"8d",
          5340 => x"7d",
          5341 => x"38",
          5342 => x"57",
          5343 => x"83",
          5344 => x"76",
          5345 => x"7a",
          5346 => x"ff",
          5347 => x"81",
          5348 => x"81",
          5349 => x"16",
          5350 => x"56",
          5351 => x"38",
          5352 => x"83",
          5353 => x"86",
          5354 => x"ff",
          5355 => x"38",
          5356 => x"82",
          5357 => x"81",
          5358 => x"06",
          5359 => x"fe",
          5360 => x"53",
          5361 => x"51",
          5362 => x"3f",
          5363 => x"52",
          5364 => x"9c",
          5365 => x"be",
          5366 => x"75",
          5367 => x"81",
          5368 => x"0b",
          5369 => x"77",
          5370 => x"75",
          5371 => x"60",
          5372 => x"80",
          5373 => x"75",
          5374 => x"ff",
          5375 => x"85",
          5376 => x"dc",
          5377 => x"2a",
          5378 => x"75",
          5379 => x"81",
          5380 => x"87",
          5381 => x"52",
          5382 => x"51",
          5383 => x"3f",
          5384 => x"ca",
          5385 => x"9c",
          5386 => x"54",
          5387 => x"52",
          5388 => x"98",
          5389 => x"56",
          5390 => x"08",
          5391 => x"53",
          5392 => x"51",
          5393 => x"3f",
          5394 => x"dc",
          5395 => x"38",
          5396 => x"56",
          5397 => x"56",
          5398 => x"dc",
          5399 => x"75",
          5400 => x"0c",
          5401 => x"04",
          5402 => x"7d",
          5403 => x"80",
          5404 => x"05",
          5405 => x"76",
          5406 => x"38",
          5407 => x"11",
          5408 => x"53",
          5409 => x"79",
          5410 => x"3f",
          5411 => x"09",
          5412 => x"38",
          5413 => x"55",
          5414 => x"db",
          5415 => x"70",
          5416 => x"34",
          5417 => x"74",
          5418 => x"81",
          5419 => x"80",
          5420 => x"55",
          5421 => x"76",
          5422 => x"dc",
          5423 => x"3d",
          5424 => x"3d",
          5425 => x"08",
          5426 => x"57",
          5427 => x"80",
          5428 => x"39",
          5429 => x"85",
          5430 => x"80",
          5431 => x"15",
          5432 => x"33",
          5433 => x"a0",
          5434 => x"81",
          5435 => x"70",
          5436 => x"06",
          5437 => x"e6",
          5438 => x"2e",
          5439 => x"88",
          5440 => x"70",
          5441 => x"34",
          5442 => x"90",
          5443 => x"dc",
          5444 => x"53",
          5445 => x"54",
          5446 => x"3f",
          5447 => x"08",
          5448 => x"14",
          5449 => x"81",
          5450 => x"38",
          5451 => x"81",
          5452 => x"53",
          5453 => x"d2",
          5454 => x"72",
          5455 => x"0c",
          5456 => x"04",
          5457 => x"73",
          5458 => x"26",
          5459 => x"71",
          5460 => x"c4",
          5461 => x"71",
          5462 => x"ce",
          5463 => x"80",
          5464 => x"f4",
          5465 => x"39",
          5466 => x"51",
          5467 => x"81",
          5468 => x"80",
          5469 => x"cf",
          5470 => x"e4",
          5471 => x"bc",
          5472 => x"39",
          5473 => x"51",
          5474 => x"81",
          5475 => x"80",
          5476 => x"cf",
          5477 => x"c8",
          5478 => x"90",
          5479 => x"39",
          5480 => x"51",
          5481 => x"d0",
          5482 => x"39",
          5483 => x"51",
          5484 => x"d1",
          5485 => x"39",
          5486 => x"51",
          5487 => x"d1",
          5488 => x"39",
          5489 => x"51",
          5490 => x"d1",
          5491 => x"39",
          5492 => x"51",
          5493 => x"d2",
          5494 => x"39",
          5495 => x"51",
          5496 => x"3f",
          5497 => x"04",
          5498 => x"77",
          5499 => x"74",
          5500 => x"8a",
          5501 => x"75",
          5502 => x"51",
          5503 => x"e8",
          5504 => x"fe",
          5505 => x"81",
          5506 => x"52",
          5507 => x"ea",
          5508 => x"dc",
          5509 => x"79",
          5510 => x"81",
          5511 => x"ff",
          5512 => x"87",
          5513 => x"ec",
          5514 => x"02",
          5515 => x"e3",
          5516 => x"57",
          5517 => x"30",
          5518 => x"73",
          5519 => x"59",
          5520 => x"77",
          5521 => x"83",
          5522 => x"74",
          5523 => x"81",
          5524 => x"55",
          5525 => x"80",
          5526 => x"53",
          5527 => x"3d",
          5528 => x"c1",
          5529 => x"dc",
          5530 => x"81",
          5531 => x"b8",
          5532 => x"cc",
          5533 => x"98",
          5534 => x"dc",
          5535 => x"96",
          5536 => x"54",
          5537 => x"77",
          5538 => x"c5",
          5539 => x"dc",
          5540 => x"81",
          5541 => x"90",
          5542 => x"74",
          5543 => x"38",
          5544 => x"19",
          5545 => x"39",
          5546 => x"05",
          5547 => x"3f",
          5548 => x"78",
          5549 => x"7b",
          5550 => x"2a",
          5551 => x"57",
          5552 => x"80",
          5553 => x"81",
          5554 => x"87",
          5555 => x"08",
          5556 => x"fe",
          5557 => x"56",
          5558 => x"cc",
          5559 => x"0d",
          5560 => x"0d",
          5561 => x"05",
          5562 => x"57",
          5563 => x"80",
          5564 => x"79",
          5565 => x"3f",
          5566 => x"08",
          5567 => x"80",
          5568 => x"75",
          5569 => x"38",
          5570 => x"55",
          5571 => x"dc",
          5572 => x"52",
          5573 => x"2d",
          5574 => x"08",
          5575 => x"77",
          5576 => x"dc",
          5577 => x"3d",
          5578 => x"3d",
          5579 => x"63",
          5580 => x"80",
          5581 => x"73",
          5582 => x"41",
          5583 => x"5e",
          5584 => x"52",
          5585 => x"51",
          5586 => x"3f",
          5587 => x"51",
          5588 => x"3f",
          5589 => x"79",
          5590 => x"38",
          5591 => x"89",
          5592 => x"2e",
          5593 => x"c6",
          5594 => x"53",
          5595 => x"8e",
          5596 => x"52",
          5597 => x"51",
          5598 => x"3f",
          5599 => x"d2",
          5600 => x"82",
          5601 => x"15",
          5602 => x"39",
          5603 => x"72",
          5604 => x"38",
          5605 => x"81",
          5606 => x"ff",
          5607 => x"89",
          5608 => x"f0",
          5609 => x"da",
          5610 => x"55",
          5611 => x"18",
          5612 => x"27",
          5613 => x"33",
          5614 => x"fc",
          5615 => x"a6",
          5616 => x"81",
          5617 => x"ff",
          5618 => x"81",
          5619 => x"51",
          5620 => x"3f",
          5621 => x"81",
          5622 => x"ff",
          5623 => x"80",
          5624 => x"27",
          5625 => x"18",
          5626 => x"53",
          5627 => x"7a",
          5628 => x"81",
          5629 => x"9f",
          5630 => x"38",
          5631 => x"73",
          5632 => x"ff",
          5633 => x"72",
          5634 => x"38",
          5635 => x"26",
          5636 => x"51",
          5637 => x"51",
          5638 => x"3f",
          5639 => x"c1",
          5640 => x"8c",
          5641 => x"da",
          5642 => x"79",
          5643 => x"fe",
          5644 => x"81",
          5645 => x"98",
          5646 => x"2c",
          5647 => x"a0",
          5648 => x"06",
          5649 => x"f6",
          5650 => x"dc",
          5651 => x"2b",
          5652 => x"70",
          5653 => x"30",
          5654 => x"70",
          5655 => x"07",
          5656 => x"06",
          5657 => x"59",
          5658 => x"80",
          5659 => x"38",
          5660 => x"09",
          5661 => x"38",
          5662 => x"39",
          5663 => x"72",
          5664 => x"be",
          5665 => x"72",
          5666 => x"0c",
          5667 => x"04",
          5668 => x"02",
          5669 => x"81",
          5670 => x"81",
          5671 => x"55",
          5672 => x"3f",
          5673 => x"22",
          5674 => x"9f",
          5675 => x"a0",
          5676 => x"ac",
          5677 => x"ad",
          5678 => x"d3",
          5679 => x"86",
          5680 => x"80",
          5681 => x"fe",
          5682 => x"86",
          5683 => x"fe",
          5684 => x"c0",
          5685 => x"53",
          5686 => x"3f",
          5687 => x"f1",
          5688 => x"d3",
          5689 => x"f3",
          5690 => x"51",
          5691 => x"3f",
          5692 => x"70",
          5693 => x"52",
          5694 => x"95",
          5695 => x"fe",
          5696 => x"81",
          5697 => x"fe",
          5698 => x"80",
          5699 => x"94",
          5700 => x"2a",
          5701 => x"51",
          5702 => x"2e",
          5703 => x"51",
          5704 => x"3f",
          5705 => x"51",
          5706 => x"3f",
          5707 => x"f0",
          5708 => x"83",
          5709 => x"06",
          5710 => x"80",
          5711 => x"81",
          5712 => x"e0",
          5713 => x"8c",
          5714 => x"d8",
          5715 => x"fe",
          5716 => x"72",
          5717 => x"81",
          5718 => x"71",
          5719 => x"38",
          5720 => x"f0",
          5721 => x"d4",
          5722 => x"f2",
          5723 => x"51",
          5724 => x"3f",
          5725 => x"70",
          5726 => x"52",
          5727 => x"95",
          5728 => x"fe",
          5729 => x"81",
          5730 => x"fe",
          5731 => x"80",
          5732 => x"90",
          5733 => x"2a",
          5734 => x"51",
          5735 => x"2e",
          5736 => x"51",
          5737 => x"3f",
          5738 => x"51",
          5739 => x"3f",
          5740 => x"ef",
          5741 => x"87",
          5742 => x"06",
          5743 => x"80",
          5744 => x"81",
          5745 => x"dc",
          5746 => x"dc",
          5747 => x"d4",
          5748 => x"fe",
          5749 => x"72",
          5750 => x"81",
          5751 => x"71",
          5752 => x"38",
          5753 => x"ef",
          5754 => x"d4",
          5755 => x"f1",
          5756 => x"51",
          5757 => x"3f",
          5758 => x"3f",
          5759 => x"04",
          5760 => x"77",
          5761 => x"56",
          5762 => x"75",
          5763 => x"f2",
          5764 => x"d8",
          5765 => x"a7",
          5766 => x"81",
          5767 => x"81",
          5768 => x"ff",
          5769 => x"81",
          5770 => x"30",
          5771 => x"cc",
          5772 => x"25",
          5773 => x"51",
          5774 => x"81",
          5775 => x"81",
          5776 => x"54",
          5777 => x"09",
          5778 => x"38",
          5779 => x"53",
          5780 => x"51",
          5781 => x"81",
          5782 => x"80",
          5783 => x"81",
          5784 => x"51",
          5785 => x"3f",
          5786 => x"f3",
          5787 => x"83",
          5788 => x"81",
          5789 => x"81",
          5790 => x"54",
          5791 => x"09",
          5792 => x"38",
          5793 => x"51",
          5794 => x"3f",
          5795 => x"dc",
          5796 => x"3d",
          5797 => x"3d",
          5798 => x"71",
          5799 => x"0c",
          5800 => x"52",
          5801 => x"88",
          5802 => x"dc",
          5803 => x"ff",
          5804 => x"7d",
          5805 => x"06",
          5806 => x"d5",
          5807 => x"3d",
          5808 => x"ff",
          5809 => x"7c",
          5810 => x"81",
          5811 => x"ff",
          5812 => x"81",
          5813 => x"7d",
          5814 => x"81",
          5815 => x"8d",
          5816 => x"70",
          5817 => x"d5",
          5818 => x"fc",
          5819 => x"3d",
          5820 => x"80",
          5821 => x"51",
          5822 => x"b4",
          5823 => x"05",
          5824 => x"3f",
          5825 => x"08",
          5826 => x"90",
          5827 => x"78",
          5828 => x"87",
          5829 => x"80",
          5830 => x"38",
          5831 => x"81",
          5832 => x"bd",
          5833 => x"78",
          5834 => x"ba",
          5835 => x"2e",
          5836 => x"8a",
          5837 => x"80",
          5838 => x"a1",
          5839 => x"c0",
          5840 => x"38",
          5841 => x"82",
          5842 => x"d2",
          5843 => x"f9",
          5844 => x"38",
          5845 => x"24",
          5846 => x"80",
          5847 => x"98",
          5848 => x"f8",
          5849 => x"38",
          5850 => x"78",
          5851 => x"8a",
          5852 => x"81",
          5853 => x"38",
          5854 => x"2e",
          5855 => x"8a",
          5856 => x"81",
          5857 => x"8f",
          5858 => x"39",
          5859 => x"80",
          5860 => x"84",
          5861 => x"82",
          5862 => x"dc",
          5863 => x"2e",
          5864 => x"b4",
          5865 => x"11",
          5866 => x"05",
          5867 => x"ab",
          5868 => x"cc",
          5869 => x"fe",
          5870 => x"3d",
          5871 => x"53",
          5872 => x"51",
          5873 => x"3f",
          5874 => x"08",
          5875 => x"dc",
          5876 => x"81",
          5877 => x"fe",
          5878 => x"63",
          5879 => x"79",
          5880 => x"f2",
          5881 => x"78",
          5882 => x"05",
          5883 => x"7a",
          5884 => x"81",
          5885 => x"3d",
          5886 => x"53",
          5887 => x"51",
          5888 => x"3f",
          5889 => x"08",
          5890 => x"da",
          5891 => x"fe",
          5892 => x"ff",
          5893 => x"ff",
          5894 => x"81",
          5895 => x"80",
          5896 => x"38",
          5897 => x"f8",
          5898 => x"84",
          5899 => x"81",
          5900 => x"dc",
          5901 => x"2e",
          5902 => x"81",
          5903 => x"fe",
          5904 => x"63",
          5905 => x"27",
          5906 => x"61",
          5907 => x"81",
          5908 => x"79",
          5909 => x"05",
          5910 => x"b4",
          5911 => x"11",
          5912 => x"05",
          5913 => x"f3",
          5914 => x"cc",
          5915 => x"fc",
          5916 => x"3d",
          5917 => x"53",
          5918 => x"51",
          5919 => x"3f",
          5920 => x"08",
          5921 => x"de",
          5922 => x"fe",
          5923 => x"ff",
          5924 => x"ff",
          5925 => x"81",
          5926 => x"80",
          5927 => x"38",
          5928 => x"51",
          5929 => x"3f",
          5930 => x"63",
          5931 => x"61",
          5932 => x"33",
          5933 => x"78",
          5934 => x"38",
          5935 => x"54",
          5936 => x"79",
          5937 => x"ac",
          5938 => x"9a",
          5939 => x"62",
          5940 => x"5a",
          5941 => x"d6",
          5942 => x"bd",
          5943 => x"ff",
          5944 => x"ff",
          5945 => x"fe",
          5946 => x"81",
          5947 => x"80",
          5948 => x"d9",
          5949 => x"78",
          5950 => x"38",
          5951 => x"08",
          5952 => x"39",
          5953 => x"33",
          5954 => x"2e",
          5955 => x"d9",
          5956 => x"bc",
          5957 => x"c2",
          5958 => x"80",
          5959 => x"81",
          5960 => x"44",
          5961 => x"d9",
          5962 => x"78",
          5963 => x"38",
          5964 => x"08",
          5965 => x"81",
          5966 => x"59",
          5967 => x"88",
          5968 => x"98",
          5969 => x"39",
          5970 => x"08",
          5971 => x"44",
          5972 => x"fc",
          5973 => x"84",
          5974 => x"fe",
          5975 => x"dc",
          5976 => x"de",
          5977 => x"c0",
          5978 => x"80",
          5979 => x"81",
          5980 => x"43",
          5981 => x"81",
          5982 => x"59",
          5983 => x"88",
          5984 => x"84",
          5985 => x"39",
          5986 => x"33",
          5987 => x"2e",
          5988 => x"d9",
          5989 => x"aa",
          5990 => x"c3",
          5991 => x"80",
          5992 => x"81",
          5993 => x"43",
          5994 => x"d9",
          5995 => x"78",
          5996 => x"38",
          5997 => x"08",
          5998 => x"81",
          5999 => x"88",
          6000 => x"3d",
          6001 => x"53",
          6002 => x"51",
          6003 => x"3f",
          6004 => x"08",
          6005 => x"38",
          6006 => x"5c",
          6007 => x"83",
          6008 => x"7a",
          6009 => x"30",
          6010 => x"9f",
          6011 => x"06",
          6012 => x"5a",
          6013 => x"88",
          6014 => x"2e",
          6015 => x"42",
          6016 => x"51",
          6017 => x"3f",
          6018 => x"54",
          6019 => x"52",
          6020 => x"96",
          6021 => x"d8",
          6022 => x"e6",
          6023 => x"39",
          6024 => x"80",
          6025 => x"84",
          6026 => x"fd",
          6027 => x"dc",
          6028 => x"2e",
          6029 => x"b4",
          6030 => x"11",
          6031 => x"05",
          6032 => x"97",
          6033 => x"cc",
          6034 => x"a5",
          6035 => x"02",
          6036 => x"33",
          6037 => x"81",
          6038 => x"3d",
          6039 => x"53",
          6040 => x"51",
          6041 => x"3f",
          6042 => x"08",
          6043 => x"f6",
          6044 => x"33",
          6045 => x"d6",
          6046 => x"fa",
          6047 => x"f8",
          6048 => x"fe",
          6049 => x"79",
          6050 => x"59",
          6051 => x"f8",
          6052 => x"79",
          6053 => x"b4",
          6054 => x"11",
          6055 => x"05",
          6056 => x"b7",
          6057 => x"cc",
          6058 => x"91",
          6059 => x"02",
          6060 => x"33",
          6061 => x"81",
          6062 => x"b5",
          6063 => x"f0",
          6064 => x"be",
          6065 => x"39",
          6066 => x"f4",
          6067 => x"84",
          6068 => x"fd",
          6069 => x"dc",
          6070 => x"2e",
          6071 => x"b4",
          6072 => x"11",
          6073 => x"05",
          6074 => x"e1",
          6075 => x"cc",
          6076 => x"a6",
          6077 => x"02",
          6078 => x"79",
          6079 => x"5b",
          6080 => x"b4",
          6081 => x"11",
          6082 => x"05",
          6083 => x"bd",
          6084 => x"cc",
          6085 => x"f7",
          6086 => x"70",
          6087 => x"81",
          6088 => x"fe",
          6089 => x"80",
          6090 => x"51",
          6091 => x"3f",
          6092 => x"33",
          6093 => x"2e",
          6094 => x"78",
          6095 => x"38",
          6096 => x"41",
          6097 => x"3d",
          6098 => x"53",
          6099 => x"51",
          6100 => x"3f",
          6101 => x"08",
          6102 => x"38",
          6103 => x"be",
          6104 => x"70",
          6105 => x"23",
          6106 => x"ae",
          6107 => x"f0",
          6108 => x"8e",
          6109 => x"39",
          6110 => x"f4",
          6111 => x"84",
          6112 => x"fc",
          6113 => x"dc",
          6114 => x"2e",
          6115 => x"b4",
          6116 => x"11",
          6117 => x"05",
          6118 => x"b1",
          6119 => x"cc",
          6120 => x"a1",
          6121 => x"71",
          6122 => x"84",
          6123 => x"3d",
          6124 => x"53",
          6125 => x"51",
          6126 => x"3f",
          6127 => x"08",
          6128 => x"a2",
          6129 => x"08",
          6130 => x"d7",
          6131 => x"f8",
          6132 => x"f8",
          6133 => x"fe",
          6134 => x"79",
          6135 => x"59",
          6136 => x"f6",
          6137 => x"79",
          6138 => x"b4",
          6139 => x"11",
          6140 => x"05",
          6141 => x"d5",
          6142 => x"cc",
          6143 => x"8d",
          6144 => x"71",
          6145 => x"84",
          6146 => x"b9",
          6147 => x"f0",
          6148 => x"ee",
          6149 => x"39",
          6150 => x"80",
          6151 => x"84",
          6152 => x"f9",
          6153 => x"dc",
          6154 => x"2e",
          6155 => x"63",
          6156 => x"90",
          6157 => x"ae",
          6158 => x"78",
          6159 => x"ff",
          6160 => x"ff",
          6161 => x"fe",
          6162 => x"81",
          6163 => x"80",
          6164 => x"38",
          6165 => x"d7",
          6166 => x"f7",
          6167 => x"59",
          6168 => x"dc",
          6169 => x"2e",
          6170 => x"81",
          6171 => x"52",
          6172 => x"51",
          6173 => x"3f",
          6174 => x"81",
          6175 => x"fe",
          6176 => x"fe",
          6177 => x"f4",
          6178 => x"d8",
          6179 => x"f0",
          6180 => x"59",
          6181 => x"fe",
          6182 => x"f4",
          6183 => x"70",
          6184 => x"78",
          6185 => x"be",
          6186 => x"06",
          6187 => x"2e",
          6188 => x"b4",
          6189 => x"05",
          6190 => x"99",
          6191 => x"cc",
          6192 => x"5b",
          6193 => x"b2",
          6194 => x"24",
          6195 => x"81",
          6196 => x"80",
          6197 => x"83",
          6198 => x"80",
          6199 => x"d8",
          6200 => x"55",
          6201 => x"54",
          6202 => x"d8",
          6203 => x"3d",
          6204 => x"51",
          6205 => x"3f",
          6206 => x"d8",
          6207 => x"3d",
          6208 => x"51",
          6209 => x"3f",
          6210 => x"55",
          6211 => x"54",
          6212 => x"d8",
          6213 => x"3d",
          6214 => x"51",
          6215 => x"3f",
          6216 => x"54",
          6217 => x"d8",
          6218 => x"3d",
          6219 => x"51",
          6220 => x"3f",
          6221 => x"58",
          6222 => x"57",
          6223 => x"81",
          6224 => x"05",
          6225 => x"83",
          6226 => x"83",
          6227 => x"b4",
          6228 => x"05",
          6229 => x"3f",
          6230 => x"08",
          6231 => x"08",
          6232 => x"70",
          6233 => x"25",
          6234 => x"5f",
          6235 => x"83",
          6236 => x"81",
          6237 => x"06",
          6238 => x"2e",
          6239 => x"1b",
          6240 => x"06",
          6241 => x"fe",
          6242 => x"81",
          6243 => x"32",
          6244 => x"8a",
          6245 => x"2e",
          6246 => x"f2",
          6247 => x"d8",
          6248 => x"f4",
          6249 => x"be",
          6250 => x"0d",
          6251 => x"dd",
          6252 => x"c0",
          6253 => x"08",
          6254 => x"84",
          6255 => x"51",
          6256 => x"3f",
          6257 => x"08",
          6258 => x"08",
          6259 => x"84",
          6260 => x"51",
          6261 => x"3f",
          6262 => x"cc",
          6263 => x"0c",
          6264 => x"9c",
          6265 => x"55",
          6266 => x"52",
          6267 => x"d3",
          6268 => x"dc",
          6269 => x"2b",
          6270 => x"53",
          6271 => x"52",
          6272 => x"d2",
          6273 => x"81",
          6274 => x"07",
          6275 => x"80",
          6276 => x"c0",
          6277 => x"8c",
          6278 => x"87",
          6279 => x"0c",
          6280 => x"81",
          6281 => x"a6",
          6282 => x"dc",
          6283 => x"e3",
          6284 => x"ec",
          6285 => x"d8",
          6286 => x"ed",
          6287 => x"d8",
          6288 => x"ed",
          6289 => x"b1",
          6290 => x"ec",
          6291 => x"51",
          6292 => x"f0",
          6293 => x"04",
          6294 => x"ff",
          6295 => x"00",
          6296 => x"ff",
          6297 => x"ff",
          6298 => x"00",
          6299 => x"00",
          6300 => x"00",
          6301 => x"00",
          6302 => x"00",
          6303 => x"00",
          6304 => x"00",
          6305 => x"00",
          6306 => x"00",
          6307 => x"00",
          6308 => x"00",
          6309 => x"00",
          6310 => x"00",
          6311 => x"00",
          6312 => x"00",
          6313 => x"00",
          6314 => x"00",
          6315 => x"00",
          6316 => x"00",
          6317 => x"00",
          6318 => x"00",
          6319 => x"00",
          6320 => x"00",
          6321 => x"00",
          6322 => x"00",
          6323 => x"64",
          6324 => x"2f",
          6325 => x"25",
          6326 => x"64",
          6327 => x"2e",
          6328 => x"64",
          6329 => x"6f",
          6330 => x"6f",
          6331 => x"67",
          6332 => x"74",
          6333 => x"00",
          6334 => x"28",
          6335 => x"6d",
          6336 => x"43",
          6337 => x"6e",
          6338 => x"29",
          6339 => x"0a",
          6340 => x"69",
          6341 => x"20",
          6342 => x"6c",
          6343 => x"6e",
          6344 => x"3a",
          6345 => x"20",
          6346 => x"42",
          6347 => x"52",
          6348 => x"20",
          6349 => x"38",
          6350 => x"30",
          6351 => x"2e",
          6352 => x"20",
          6353 => x"44",
          6354 => x"20",
          6355 => x"20",
          6356 => x"38",
          6357 => x"30",
          6358 => x"2e",
          6359 => x"20",
          6360 => x"4e",
          6361 => x"42",
          6362 => x"20",
          6363 => x"38",
          6364 => x"30",
          6365 => x"2e",
          6366 => x"20",
          6367 => x"52",
          6368 => x"20",
          6369 => x"20",
          6370 => x"38",
          6371 => x"30",
          6372 => x"2e",
          6373 => x"20",
          6374 => x"41",
          6375 => x"20",
          6376 => x"20",
          6377 => x"38",
          6378 => x"30",
          6379 => x"2e",
          6380 => x"20",
          6381 => x"44",
          6382 => x"52",
          6383 => x"20",
          6384 => x"76",
          6385 => x"73",
          6386 => x"30",
          6387 => x"2e",
          6388 => x"20",
          6389 => x"49",
          6390 => x"31",
          6391 => x"20",
          6392 => x"6d",
          6393 => x"20",
          6394 => x"30",
          6395 => x"2e",
          6396 => x"20",
          6397 => x"4e",
          6398 => x"43",
          6399 => x"20",
          6400 => x"61",
          6401 => x"6c",
          6402 => x"30",
          6403 => x"2e",
          6404 => x"20",
          6405 => x"49",
          6406 => x"4f",
          6407 => x"42",
          6408 => x"00",
          6409 => x"20",
          6410 => x"42",
          6411 => x"43",
          6412 => x"20",
          6413 => x"4f",
          6414 => x"0a",
          6415 => x"20",
          6416 => x"53",
          6417 => x"00",
          6418 => x"20",
          6419 => x"50",
          6420 => x"00",
          6421 => x"64",
          6422 => x"73",
          6423 => x"3a",
          6424 => x"20",
          6425 => x"50",
          6426 => x"65",
          6427 => x"20",
          6428 => x"74",
          6429 => x"41",
          6430 => x"65",
          6431 => x"3d",
          6432 => x"38",
          6433 => x"00",
          6434 => x"20",
          6435 => x"50",
          6436 => x"65",
          6437 => x"79",
          6438 => x"61",
          6439 => x"41",
          6440 => x"65",
          6441 => x"3d",
          6442 => x"38",
          6443 => x"00",
          6444 => x"20",
          6445 => x"74",
          6446 => x"20",
          6447 => x"72",
          6448 => x"64",
          6449 => x"73",
          6450 => x"20",
          6451 => x"3d",
          6452 => x"38",
          6453 => x"00",
          6454 => x"69",
          6455 => x"0a",
          6456 => x"20",
          6457 => x"50",
          6458 => x"64",
          6459 => x"20",
          6460 => x"20",
          6461 => x"20",
          6462 => x"20",
          6463 => x"3d",
          6464 => x"34",
          6465 => x"00",
          6466 => x"20",
          6467 => x"79",
          6468 => x"6d",
          6469 => x"6f",
          6470 => x"46",
          6471 => x"20",
          6472 => x"20",
          6473 => x"3d",
          6474 => x"2e",
          6475 => x"64",
          6476 => x"0a",
          6477 => x"20",
          6478 => x"44",
          6479 => x"20",
          6480 => x"63",
          6481 => x"72",
          6482 => x"20",
          6483 => x"20",
          6484 => x"3d",
          6485 => x"2e",
          6486 => x"64",
          6487 => x"0a",
          6488 => x"20",
          6489 => x"69",
          6490 => x"6f",
          6491 => x"53",
          6492 => x"4d",
          6493 => x"6f",
          6494 => x"46",
          6495 => x"3d",
          6496 => x"2e",
          6497 => x"64",
          6498 => x"0a",
          6499 => x"6d",
          6500 => x"00",
          6501 => x"65",
          6502 => x"6d",
          6503 => x"6c",
          6504 => x"00",
          6505 => x"56",
          6506 => x"56",
          6507 => x"6e",
          6508 => x"6e",
          6509 => x"77",
          6510 => x"44",
          6511 => x"2a",
          6512 => x"3b",
          6513 => x"3f",
          6514 => x"7f",
          6515 => x"41",
          6516 => x"41",
          6517 => x"00",
          6518 => x"fe",
          6519 => x"44",
          6520 => x"2e",
          6521 => x"4f",
          6522 => x"4d",
          6523 => x"20",
          6524 => x"54",
          6525 => x"20",
          6526 => x"4f",
          6527 => x"4d",
          6528 => x"20",
          6529 => x"54",
          6530 => x"20",
          6531 => x"00",
          6532 => x"00",
          6533 => x"00",
          6534 => x"00",
          6535 => x"9a",
          6536 => x"41",
          6537 => x"45",
          6538 => x"49",
          6539 => x"92",
          6540 => x"4f",
          6541 => x"99",
          6542 => x"9d",
          6543 => x"49",
          6544 => x"a5",
          6545 => x"a9",
          6546 => x"ad",
          6547 => x"b1",
          6548 => x"b5",
          6549 => x"b9",
          6550 => x"bd",
          6551 => x"c1",
          6552 => x"c5",
          6553 => x"c9",
          6554 => x"cd",
          6555 => x"d1",
          6556 => x"d5",
          6557 => x"d9",
          6558 => x"dd",
          6559 => x"e1",
          6560 => x"e5",
          6561 => x"e9",
          6562 => x"ed",
          6563 => x"f1",
          6564 => x"f5",
          6565 => x"f9",
          6566 => x"fd",
          6567 => x"2e",
          6568 => x"5b",
          6569 => x"22",
          6570 => x"3e",
          6571 => x"00",
          6572 => x"01",
          6573 => x"10",
          6574 => x"00",
          6575 => x"00",
          6576 => x"01",
          6577 => x"04",
          6578 => x"10",
          6579 => x"00",
          6580 => x"69",
          6581 => x"00",
          6582 => x"69",
          6583 => x"6c",
          6584 => x"69",
          6585 => x"00",
          6586 => x"6c",
          6587 => x"00",
          6588 => x"65",
          6589 => x"00",
          6590 => x"63",
          6591 => x"72",
          6592 => x"63",
          6593 => x"00",
          6594 => x"64",
          6595 => x"00",
          6596 => x"64",
          6597 => x"00",
          6598 => x"65",
          6599 => x"65",
          6600 => x"65",
          6601 => x"69",
          6602 => x"69",
          6603 => x"66",
          6604 => x"66",
          6605 => x"61",
          6606 => x"00",
          6607 => x"6d",
          6608 => x"65",
          6609 => x"72",
          6610 => x"65",
          6611 => x"00",
          6612 => x"6e",
          6613 => x"00",
          6614 => x"65",
          6615 => x"00",
          6616 => x"62",
          6617 => x"63",
          6618 => x"69",
          6619 => x"45",
          6620 => x"72",
          6621 => x"6e",
          6622 => x"6e",
          6623 => x"65",
          6624 => x"72",
          6625 => x"00",
          6626 => x"69",
          6627 => x"6e",
          6628 => x"72",
          6629 => x"79",
          6630 => x"00",
          6631 => x"6f",
          6632 => x"6c",
          6633 => x"6f",
          6634 => x"2e",
          6635 => x"6f",
          6636 => x"74",
          6637 => x"6f",
          6638 => x"2e",
          6639 => x"6e",
          6640 => x"69",
          6641 => x"69",
          6642 => x"61",
          6643 => x"0a",
          6644 => x"63",
          6645 => x"73",
          6646 => x"6e",
          6647 => x"2e",
          6648 => x"69",
          6649 => x"61",
          6650 => x"61",
          6651 => x"65",
          6652 => x"74",
          6653 => x"00",
          6654 => x"69",
          6655 => x"68",
          6656 => x"6c",
          6657 => x"6e",
          6658 => x"69",
          6659 => x"00",
          6660 => x"44",
          6661 => x"20",
          6662 => x"74",
          6663 => x"72",
          6664 => x"63",
          6665 => x"2e",
          6666 => x"72",
          6667 => x"20",
          6668 => x"62",
          6669 => x"69",
          6670 => x"6e",
          6671 => x"69",
          6672 => x"00",
          6673 => x"69",
          6674 => x"6e",
          6675 => x"65",
          6676 => x"6c",
          6677 => x"0a",
          6678 => x"6f",
          6679 => x"6d",
          6680 => x"69",
          6681 => x"20",
          6682 => x"65",
          6683 => x"74",
          6684 => x"66",
          6685 => x"64",
          6686 => x"20",
          6687 => x"6b",
          6688 => x"00",
          6689 => x"6f",
          6690 => x"74",
          6691 => x"6f",
          6692 => x"64",
          6693 => x"00",
          6694 => x"69",
          6695 => x"75",
          6696 => x"6f",
          6697 => x"61",
          6698 => x"6e",
          6699 => x"6e",
          6700 => x"6c",
          6701 => x"0a",
          6702 => x"69",
          6703 => x"69",
          6704 => x"6f",
          6705 => x"64",
          6706 => x"00",
          6707 => x"6e",
          6708 => x"66",
          6709 => x"65",
          6710 => x"6d",
          6711 => x"72",
          6712 => x"00",
          6713 => x"6f",
          6714 => x"61",
          6715 => x"6f",
          6716 => x"20",
          6717 => x"65",
          6718 => x"00",
          6719 => x"61",
          6720 => x"65",
          6721 => x"73",
          6722 => x"63",
          6723 => x"65",
          6724 => x"0a",
          6725 => x"75",
          6726 => x"73",
          6727 => x"00",
          6728 => x"6e",
          6729 => x"77",
          6730 => x"72",
          6731 => x"2e",
          6732 => x"25",
          6733 => x"62",
          6734 => x"73",
          6735 => x"20",
          6736 => x"25",
          6737 => x"62",
          6738 => x"73",
          6739 => x"63",
          6740 => x"00",
          6741 => x"65",
          6742 => x"00",
          6743 => x"30",
          6744 => x"00",
          6745 => x"20",
          6746 => x"30",
          6747 => x"00",
          6748 => x"20",
          6749 => x"20",
          6750 => x"00",
          6751 => x"30",
          6752 => x"00",
          6753 => x"20",
          6754 => x"7c",
          6755 => x"0d",
          6756 => x"4f",
          6757 => x"2a",
          6758 => x"73",
          6759 => x"00",
          6760 => x"30",
          6761 => x"2f",
          6762 => x"30",
          6763 => x"31",
          6764 => x"00",
          6765 => x"5a",
          6766 => x"20",
          6767 => x"20",
          6768 => x"78",
          6769 => x"73",
          6770 => x"20",
          6771 => x"0a",
          6772 => x"50",
          6773 => x"6e",
          6774 => x"72",
          6775 => x"20",
          6776 => x"64",
          6777 => x"0a",
          6778 => x"69",
          6779 => x"20",
          6780 => x"65",
          6781 => x"70",
          6782 => x"00",
          6783 => x"53",
          6784 => x"6e",
          6785 => x"72",
          6786 => x"0a",
          6787 => x"4f",
          6788 => x"20",
          6789 => x"69",
          6790 => x"72",
          6791 => x"74",
          6792 => x"4f",
          6793 => x"20",
          6794 => x"69",
          6795 => x"72",
          6796 => x"74",
          6797 => x"41",
          6798 => x"20",
          6799 => x"69",
          6800 => x"72",
          6801 => x"74",
          6802 => x"41",
          6803 => x"20",
          6804 => x"69",
          6805 => x"72",
          6806 => x"74",
          6807 => x"41",
          6808 => x"20",
          6809 => x"69",
          6810 => x"72",
          6811 => x"74",
          6812 => x"41",
          6813 => x"20",
          6814 => x"69",
          6815 => x"72",
          6816 => x"74",
          6817 => x"65",
          6818 => x"6e",
          6819 => x"70",
          6820 => x"6d",
          6821 => x"2e",
          6822 => x"00",
          6823 => x"6e",
          6824 => x"69",
          6825 => x"74",
          6826 => x"72",
          6827 => x"0a",
          6828 => x"75",
          6829 => x"78",
          6830 => x"62",
          6831 => x"00",
          6832 => x"3a",
          6833 => x"61",
          6834 => x"64",
          6835 => x"20",
          6836 => x"74",
          6837 => x"69",
          6838 => x"73",
          6839 => x"61",
          6840 => x"30",
          6841 => x"6c",
          6842 => x"65",
          6843 => x"69",
          6844 => x"61",
          6845 => x"6c",
          6846 => x"0a",
          6847 => x"20",
          6848 => x"6c",
          6849 => x"69",
          6850 => x"2e",
          6851 => x"00",
          6852 => x"6f",
          6853 => x"6e",
          6854 => x"2e",
          6855 => x"6f",
          6856 => x"72",
          6857 => x"2e",
          6858 => x"00",
          6859 => x"30",
          6860 => x"28",
          6861 => x"78",
          6862 => x"25",
          6863 => x"78",
          6864 => x"38",
          6865 => x"00",
          6866 => x"75",
          6867 => x"4d",
          6868 => x"72",
          6869 => x"00",
          6870 => x"43",
          6871 => x"6c",
          6872 => x"2e",
          6873 => x"30",
          6874 => x"25",
          6875 => x"2d",
          6876 => x"3f",
          6877 => x"00",
          6878 => x"30",
          6879 => x"25",
          6880 => x"2d",
          6881 => x"30",
          6882 => x"25",
          6883 => x"2d",
          6884 => x"78",
          6885 => x"74",
          6886 => x"20",
          6887 => x"65",
          6888 => x"25",
          6889 => x"20",
          6890 => x"0a",
          6891 => x"61",
          6892 => x"6e",
          6893 => x"6f",
          6894 => x"40",
          6895 => x"38",
          6896 => x"2e",
          6897 => x"00",
          6898 => x"61",
          6899 => x"72",
          6900 => x"72",
          6901 => x"20",
          6902 => x"65",
          6903 => x"64",
          6904 => x"00",
          6905 => x"65",
          6906 => x"72",
          6907 => x"67",
          6908 => x"70",
          6909 => x"61",
          6910 => x"6e",
          6911 => x"0a",
          6912 => x"6f",
          6913 => x"72",
          6914 => x"6f",
          6915 => x"67",
          6916 => x"0a",
          6917 => x"50",
          6918 => x"69",
          6919 => x"64",
          6920 => x"73",
          6921 => x"2e",
          6922 => x"00",
          6923 => x"64",
          6924 => x"73",
          6925 => x"00",
          6926 => x"64",
          6927 => x"73",
          6928 => x"61",
          6929 => x"6f",
          6930 => x"6e",
          6931 => x"00",
          6932 => x"75",
          6933 => x"6e",
          6934 => x"2e",
          6935 => x"6e",
          6936 => x"69",
          6937 => x"69",
          6938 => x"72",
          6939 => x"74",
          6940 => x"2e",
          6941 => x"00",
          6942 => x"00",
          6943 => x"00",
          6944 => x"00",
          6945 => x"00",
          6946 => x"01",
          6947 => x"00",
          6948 => x"01",
          6949 => x"81",
          6950 => x"00",
          6951 => x"7f",
          6952 => x"00",
          6953 => x"00",
          6954 => x"00",
          6955 => x"00",
          6956 => x"f5",
          6957 => x"f5",
          6958 => x"f5",
          6959 => x"00",
          6960 => x"01",
          6961 => x"01",
          6962 => x"01",
          6963 => x"00",
          6964 => x"00",
          6965 => x"00",
          6966 => x"00",
          6967 => x"00",
          6968 => x"02",
          6969 => x"00",
          6970 => x"00",
          6971 => x"00",
          6972 => x"04",
          6973 => x"00",
          6974 => x"00",
          6975 => x"00",
          6976 => x"14",
          6977 => x"00",
          6978 => x"00",
          6979 => x"00",
          6980 => x"2b",
          6981 => x"00",
          6982 => x"00",
          6983 => x"00",
          6984 => x"30",
          6985 => x"00",
          6986 => x"00",
          6987 => x"00",
          6988 => x"3c",
          6989 => x"00",
          6990 => x"00",
          6991 => x"00",
          6992 => x"3d",
          6993 => x"00",
          6994 => x"00",
          6995 => x"00",
          6996 => x"3f",
          6997 => x"00",
          6998 => x"00",
          6999 => x"00",
          7000 => x"40",
          7001 => x"00",
          7002 => x"00",
          7003 => x"00",
          7004 => x"41",
          7005 => x"00",
          7006 => x"00",
          7007 => x"00",
          7008 => x"42",
          7009 => x"00",
          7010 => x"00",
          7011 => x"00",
          7012 => x"43",
          7013 => x"00",
          7014 => x"00",
          7015 => x"00",
          7016 => x"50",
          7017 => x"00",
          7018 => x"00",
          7019 => x"00",
          7020 => x"51",
          7021 => x"00",
          7022 => x"00",
          7023 => x"00",
          7024 => x"54",
          7025 => x"00",
          7026 => x"00",
          7027 => x"00",
          7028 => x"55",
          7029 => x"00",
          7030 => x"00",
          7031 => x"00",
          7032 => x"79",
          7033 => x"00",
          7034 => x"00",
          7035 => x"00",
          7036 => x"78",
          7037 => x"00",
          7038 => x"00",
          7039 => x"00",
          7040 => x"82",
          7041 => x"00",
          7042 => x"00",
          7043 => x"00",
          7044 => x"83",
          7045 => x"00",
          7046 => x"00",
          7047 => x"00",
          7048 => x"85",
          7049 => x"00",
          7050 => x"00",
          7051 => x"00",
          7052 => x"87",
          7053 => x"00",
          7054 => x"00",
          7055 => x"00",
          7056 => x"8c",
          7057 => x"00",
          7058 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"da",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"be",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"d8",
           163 => x"10",
           164 => x"06",
           165 => x"96",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"df",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"cb",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"94",
           269 => x"0b",
           270 => x"0b",
           271 => x"b2",
           272 => x"0b",
           273 => x"0b",
           274 => x"d0",
           275 => x"0b",
           276 => x"0b",
           277 => x"ee",
           278 => x"0b",
           279 => x"0b",
           280 => x"8c",
           281 => x"0b",
           282 => x"0b",
           283 => x"aa",
           284 => x"0b",
           285 => x"0b",
           286 => x"c8",
           287 => x"0b",
           288 => x"0b",
           289 => x"e6",
           290 => x"0b",
           291 => x"0b",
           292 => x"84",
           293 => x"0b",
           294 => x"0b",
           295 => x"a4",
           296 => x"0b",
           297 => x"0b",
           298 => x"c4",
           299 => x"0b",
           300 => x"0b",
           301 => x"e4",
           302 => x"0b",
           303 => x"0b",
           304 => x"84",
           305 => x"0b",
           306 => x"0b",
           307 => x"a4",
           308 => x"0b",
           309 => x"0b",
           310 => x"c4",
           311 => x"0b",
           312 => x"0b",
           313 => x"e4",
           314 => x"0b",
           315 => x"0b",
           316 => x"84",
           317 => x"0b",
           318 => x"0b",
           319 => x"a4",
           320 => x"0b",
           321 => x"0b",
           322 => x"c4",
           323 => x"0b",
           324 => x"0b",
           325 => x"e4",
           326 => x"0b",
           327 => x"0b",
           328 => x"84",
           329 => x"0b",
           330 => x"0b",
           331 => x"a3",
           332 => x"0b",
           333 => x"0b",
           334 => x"c3",
           335 => x"0b",
           336 => x"0b",
           337 => x"e1",
           338 => x"0b",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"00",
           386 => x"00",
           387 => x"00",
           388 => x"00",
           389 => x"00",
           390 => x"00",
           391 => x"00",
           392 => x"00",
           393 => x"00",
           394 => x"00",
           395 => x"00",
           396 => x"00",
           397 => x"00",
           398 => x"00",
           399 => x"00",
           400 => x"00",
           401 => x"00",
           402 => x"00",
           403 => x"00",
           404 => x"00",
           405 => x"00",
           406 => x"00",
           407 => x"00",
           408 => x"00",
           409 => x"00",
           410 => x"00",
           411 => x"00",
           412 => x"00",
           413 => x"00",
           414 => x"00",
           415 => x"00",
           416 => x"00",
           417 => x"00",
           418 => x"00",
           419 => x"00",
           420 => x"00",
           421 => x"00",
           422 => x"00",
           423 => x"00",
           424 => x"00",
           425 => x"00",
           426 => x"00",
           427 => x"00",
           428 => x"00",
           429 => x"00",
           430 => x"00",
           431 => x"00",
           432 => x"00",
           433 => x"00",
           434 => x"00",
           435 => x"00",
           436 => x"00",
           437 => x"00",
           438 => x"00",
           439 => x"00",
           440 => x"00",
           441 => x"00",
           442 => x"00",
           443 => x"00",
           444 => x"00",
           445 => x"00",
           446 => x"00",
           447 => x"00",
           448 => x"00",
           449 => x"00",
           450 => x"00",
           451 => x"00",
           452 => x"00",
           453 => x"00",
           454 => x"00",
           455 => x"00",
           456 => x"00",
           457 => x"00",
           458 => x"00",
           459 => x"00",
           460 => x"00",
           461 => x"00",
           462 => x"00",
           463 => x"00",
           464 => x"00",
           465 => x"00",
           466 => x"00",
           467 => x"00",
           468 => x"00",
           469 => x"00",
           470 => x"00",
           471 => x"00",
           472 => x"00",
           473 => x"00",
           474 => x"00",
           475 => x"00",
           476 => x"00",
           477 => x"00",
           478 => x"00",
           479 => x"00",
           480 => x"00",
           481 => x"00",
           482 => x"00",
           483 => x"00",
           484 => x"00",
           485 => x"00",
           486 => x"00",
           487 => x"00",
           488 => x"00",
           489 => x"00",
           490 => x"00",
           491 => x"00",
           492 => x"00",
           493 => x"00",
           494 => x"00",
           495 => x"00",
           496 => x"00",
           497 => x"00",
           498 => x"00",
           499 => x"00",
           500 => x"00",
           501 => x"00",
           502 => x"00",
           503 => x"00",
           504 => x"00",
           505 => x"00",
           506 => x"00",
           507 => x"00",
           508 => x"00",
           509 => x"00",
           510 => x"00",
           511 => x"00",
           512 => x"04",
           513 => x"04",
           514 => x"0c",
           515 => x"81",
           516 => x"83",
           517 => x"81",
           518 => x"b1",
           519 => x"dc",
           520 => x"80",
           521 => x"dc",
           522 => x"e2",
           523 => x"d8",
           524 => x"90",
           525 => x"d8",
           526 => x"2d",
           527 => x"08",
           528 => x"04",
           529 => x"0c",
           530 => x"81",
           531 => x"83",
           532 => x"81",
           533 => x"b9",
           534 => x"dc",
           535 => x"80",
           536 => x"dc",
           537 => x"a3",
           538 => x"d8",
           539 => x"90",
           540 => x"d8",
           541 => x"2d",
           542 => x"08",
           543 => x"04",
           544 => x"0c",
           545 => x"81",
           546 => x"83",
           547 => x"81",
           548 => x"b7",
           549 => x"dc",
           550 => x"80",
           551 => x"dc",
           552 => x"fa",
           553 => x"d8",
           554 => x"90",
           555 => x"d8",
           556 => x"2d",
           557 => x"08",
           558 => x"04",
           559 => x"0c",
           560 => x"81",
           561 => x"83",
           562 => x"81",
           563 => x"a7",
           564 => x"dc",
           565 => x"80",
           566 => x"dc",
           567 => x"aa",
           568 => x"d8",
           569 => x"90",
           570 => x"d8",
           571 => x"2d",
           572 => x"08",
           573 => x"04",
           574 => x"0c",
           575 => x"81",
           576 => x"83",
           577 => x"81",
           578 => x"80",
           579 => x"81",
           580 => x"83",
           581 => x"81",
           582 => x"80",
           583 => x"81",
           584 => x"83",
           585 => x"81",
           586 => x"80",
           587 => x"81",
           588 => x"83",
           589 => x"81",
           590 => x"80",
           591 => x"81",
           592 => x"83",
           593 => x"81",
           594 => x"81",
           595 => x"81",
           596 => x"83",
           597 => x"81",
           598 => x"81",
           599 => x"81",
           600 => x"83",
           601 => x"81",
           602 => x"80",
           603 => x"81",
           604 => x"83",
           605 => x"81",
           606 => x"81",
           607 => x"81",
           608 => x"83",
           609 => x"81",
           610 => x"81",
           611 => x"81",
           612 => x"83",
           613 => x"81",
           614 => x"81",
           615 => x"81",
           616 => x"83",
           617 => x"81",
           618 => x"81",
           619 => x"81",
           620 => x"83",
           621 => x"81",
           622 => x"81",
           623 => x"81",
           624 => x"83",
           625 => x"81",
           626 => x"81",
           627 => x"81",
           628 => x"83",
           629 => x"81",
           630 => x"81",
           631 => x"81",
           632 => x"83",
           633 => x"81",
           634 => x"81",
           635 => x"81",
           636 => x"83",
           637 => x"81",
           638 => x"81",
           639 => x"81",
           640 => x"83",
           641 => x"81",
           642 => x"80",
           643 => x"81",
           644 => x"83",
           645 => x"81",
           646 => x"80",
           647 => x"81",
           648 => x"83",
           649 => x"81",
           650 => x"80",
           651 => x"81",
           652 => x"83",
           653 => x"81",
           654 => x"81",
           655 => x"81",
           656 => x"83",
           657 => x"81",
           658 => x"81",
           659 => x"81",
           660 => x"83",
           661 => x"81",
           662 => x"81",
           663 => x"81",
           664 => x"83",
           665 => x"81",
           666 => x"81",
           667 => x"81",
           668 => x"83",
           669 => x"81",
           670 => x"80",
           671 => x"81",
           672 => x"83",
           673 => x"81",
           674 => x"81",
           675 => x"81",
           676 => x"83",
           677 => x"81",
           678 => x"be",
           679 => x"dc",
           680 => x"80",
           681 => x"dc",
           682 => x"c0",
           683 => x"dc",
           684 => x"80",
           685 => x"dc",
           686 => x"c2",
           687 => x"dc",
           688 => x"80",
           689 => x"dc",
           690 => x"d3",
           691 => x"d8",
           692 => x"90",
           693 => x"d8",
           694 => x"2d",
           695 => x"08",
           696 => x"04",
           697 => x"0c",
           698 => x"81",
           699 => x"83",
           700 => x"81",
           701 => x"81",
           702 => x"81",
           703 => x"83",
           704 => x"3c",
           705 => x"10",
           706 => x"10",
           707 => x"10",
           708 => x"10",
           709 => x"10",
           710 => x"10",
           711 => x"10",
           712 => x"10",
           713 => x"00",
           714 => x"ff",
           715 => x"06",
           716 => x"83",
           717 => x"10",
           718 => x"fc",
           719 => x"51",
           720 => x"80",
           721 => x"ff",
           722 => x"06",
           723 => x"52",
           724 => x"0a",
           725 => x"38",
           726 => x"51",
           727 => x"cc",
           728 => x"f8",
           729 => x"80",
           730 => x"05",
           731 => x"0b",
           732 => x"04",
           733 => x"81",
           734 => x"00",
           735 => x"08",
           736 => x"d8",
           737 => x"0d",
           738 => x"dc",
           739 => x"05",
           740 => x"dc",
           741 => x"05",
           742 => x"d4",
           743 => x"cc",
           744 => x"dc",
           745 => x"85",
           746 => x"dc",
           747 => x"81",
           748 => x"02",
           749 => x"0c",
           750 => x"81",
           751 => x"d8",
           752 => x"08",
           753 => x"d8",
           754 => x"08",
           755 => x"3f",
           756 => x"08",
           757 => x"cc",
           758 => x"3d",
           759 => x"d8",
           760 => x"dc",
           761 => x"81",
           762 => x"f9",
           763 => x"0b",
           764 => x"08",
           765 => x"81",
           766 => x"88",
           767 => x"25",
           768 => x"dc",
           769 => x"05",
           770 => x"dc",
           771 => x"05",
           772 => x"81",
           773 => x"f4",
           774 => x"dc",
           775 => x"05",
           776 => x"81",
           777 => x"d8",
           778 => x"0c",
           779 => x"08",
           780 => x"81",
           781 => x"fc",
           782 => x"dc",
           783 => x"05",
           784 => x"b9",
           785 => x"d8",
           786 => x"08",
           787 => x"d8",
           788 => x"0c",
           789 => x"dc",
           790 => x"05",
           791 => x"d8",
           792 => x"08",
           793 => x"0b",
           794 => x"08",
           795 => x"81",
           796 => x"f0",
           797 => x"dc",
           798 => x"05",
           799 => x"81",
           800 => x"8c",
           801 => x"81",
           802 => x"88",
           803 => x"81",
           804 => x"dc",
           805 => x"81",
           806 => x"f8",
           807 => x"81",
           808 => x"fc",
           809 => x"2e",
           810 => x"dc",
           811 => x"05",
           812 => x"dc",
           813 => x"05",
           814 => x"d8",
           815 => x"08",
           816 => x"cc",
           817 => x"3d",
           818 => x"d8",
           819 => x"dc",
           820 => x"81",
           821 => x"fb",
           822 => x"0b",
           823 => x"08",
           824 => x"81",
           825 => x"88",
           826 => x"25",
           827 => x"dc",
           828 => x"05",
           829 => x"dc",
           830 => x"05",
           831 => x"81",
           832 => x"fc",
           833 => x"dc",
           834 => x"05",
           835 => x"90",
           836 => x"d8",
           837 => x"08",
           838 => x"d8",
           839 => x"0c",
           840 => x"dc",
           841 => x"05",
           842 => x"dc",
           843 => x"05",
           844 => x"3f",
           845 => x"08",
           846 => x"d8",
           847 => x"0c",
           848 => x"d8",
           849 => x"08",
           850 => x"38",
           851 => x"08",
           852 => x"30",
           853 => x"08",
           854 => x"81",
           855 => x"f8",
           856 => x"81",
           857 => x"54",
           858 => x"81",
           859 => x"04",
           860 => x"08",
           861 => x"d8",
           862 => x"0d",
           863 => x"dc",
           864 => x"05",
           865 => x"81",
           866 => x"f8",
           867 => x"dc",
           868 => x"05",
           869 => x"d8",
           870 => x"08",
           871 => x"81",
           872 => x"fc",
           873 => x"2e",
           874 => x"0b",
           875 => x"08",
           876 => x"24",
           877 => x"dc",
           878 => x"05",
           879 => x"dc",
           880 => x"05",
           881 => x"d8",
           882 => x"08",
           883 => x"d8",
           884 => x"0c",
           885 => x"81",
           886 => x"fc",
           887 => x"2e",
           888 => x"81",
           889 => x"8c",
           890 => x"dc",
           891 => x"05",
           892 => x"38",
           893 => x"08",
           894 => x"81",
           895 => x"8c",
           896 => x"81",
           897 => x"88",
           898 => x"dc",
           899 => x"05",
           900 => x"d8",
           901 => x"08",
           902 => x"d8",
           903 => x"0c",
           904 => x"08",
           905 => x"81",
           906 => x"d8",
           907 => x"0c",
           908 => x"08",
           909 => x"81",
           910 => x"d8",
           911 => x"0c",
           912 => x"81",
           913 => x"90",
           914 => x"2e",
           915 => x"dc",
           916 => x"05",
           917 => x"dc",
           918 => x"05",
           919 => x"39",
           920 => x"08",
           921 => x"70",
           922 => x"08",
           923 => x"51",
           924 => x"08",
           925 => x"81",
           926 => x"85",
           927 => x"dc",
           928 => x"fc",
           929 => x"79",
           930 => x"05",
           931 => x"57",
           932 => x"83",
           933 => x"38",
           934 => x"51",
           935 => x"a4",
           936 => x"52",
           937 => x"93",
           938 => x"70",
           939 => x"34",
           940 => x"71",
           941 => x"81",
           942 => x"74",
           943 => x"0c",
           944 => x"04",
           945 => x"2b",
           946 => x"71",
           947 => x"51",
           948 => x"72",
           949 => x"72",
           950 => x"05",
           951 => x"71",
           952 => x"53",
           953 => x"70",
           954 => x"0c",
           955 => x"84",
           956 => x"f0",
           957 => x"8f",
           958 => x"83",
           959 => x"38",
           960 => x"84",
           961 => x"fc",
           962 => x"83",
           963 => x"70",
           964 => x"39",
           965 => x"77",
           966 => x"07",
           967 => x"54",
           968 => x"38",
           969 => x"08",
           970 => x"71",
           971 => x"80",
           972 => x"75",
           973 => x"33",
           974 => x"06",
           975 => x"80",
           976 => x"72",
           977 => x"75",
           978 => x"06",
           979 => x"12",
           980 => x"33",
           981 => x"06",
           982 => x"52",
           983 => x"72",
           984 => x"81",
           985 => x"81",
           986 => x"71",
           987 => x"cc",
           988 => x"87",
           989 => x"71",
           990 => x"fb",
           991 => x"06",
           992 => x"82",
           993 => x"51",
           994 => x"97",
           995 => x"84",
           996 => x"54",
           997 => x"75",
           998 => x"38",
           999 => x"52",
          1000 => x"80",
          1001 => x"cc",
          1002 => x"0d",
          1003 => x"0d",
          1004 => x"53",
          1005 => x"52",
          1006 => x"81",
          1007 => x"81",
          1008 => x"07",
          1009 => x"52",
          1010 => x"e8",
          1011 => x"dc",
          1012 => x"3d",
          1013 => x"3d",
          1014 => x"08",
          1015 => x"56",
          1016 => x"80",
          1017 => x"33",
          1018 => x"2e",
          1019 => x"86",
          1020 => x"52",
          1021 => x"53",
          1022 => x"13",
          1023 => x"33",
          1024 => x"06",
          1025 => x"70",
          1026 => x"38",
          1027 => x"80",
          1028 => x"74",
          1029 => x"81",
          1030 => x"70",
          1031 => x"81",
          1032 => x"80",
          1033 => x"05",
          1034 => x"76",
          1035 => x"70",
          1036 => x"0c",
          1037 => x"04",
          1038 => x"76",
          1039 => x"80",
          1040 => x"86",
          1041 => x"52",
          1042 => x"82",
          1043 => x"cc",
          1044 => x"80",
          1045 => x"74",
          1046 => x"dc",
          1047 => x"3d",
          1048 => x"3d",
          1049 => x"11",
          1050 => x"52",
          1051 => x"70",
          1052 => x"98",
          1053 => x"33",
          1054 => x"82",
          1055 => x"26",
          1056 => x"84",
          1057 => x"83",
          1058 => x"26",
          1059 => x"85",
          1060 => x"84",
          1061 => x"26",
          1062 => x"86",
          1063 => x"85",
          1064 => x"26",
          1065 => x"88",
          1066 => x"86",
          1067 => x"e7",
          1068 => x"38",
          1069 => x"54",
          1070 => x"87",
          1071 => x"cc",
          1072 => x"87",
          1073 => x"0c",
          1074 => x"c0",
          1075 => x"82",
          1076 => x"c0",
          1077 => x"83",
          1078 => x"c0",
          1079 => x"84",
          1080 => x"c0",
          1081 => x"85",
          1082 => x"c0",
          1083 => x"86",
          1084 => x"c0",
          1085 => x"74",
          1086 => x"a4",
          1087 => x"c0",
          1088 => x"80",
          1089 => x"98",
          1090 => x"52",
          1091 => x"cc",
          1092 => x"0d",
          1093 => x"0d",
          1094 => x"c0",
          1095 => x"81",
          1096 => x"c0",
          1097 => x"5e",
          1098 => x"87",
          1099 => x"08",
          1100 => x"1c",
          1101 => x"98",
          1102 => x"79",
          1103 => x"87",
          1104 => x"08",
          1105 => x"1c",
          1106 => x"98",
          1107 => x"79",
          1108 => x"87",
          1109 => x"08",
          1110 => x"1c",
          1111 => x"98",
          1112 => x"7b",
          1113 => x"87",
          1114 => x"08",
          1115 => x"1c",
          1116 => x"0c",
          1117 => x"ff",
          1118 => x"83",
          1119 => x"58",
          1120 => x"57",
          1121 => x"56",
          1122 => x"55",
          1123 => x"54",
          1124 => x"53",
          1125 => x"ff",
          1126 => x"c5",
          1127 => x"c7",
          1128 => x"0d",
          1129 => x"0d",
          1130 => x"33",
          1131 => x"9f",
          1132 => x"52",
          1133 => x"81",
          1134 => x"83",
          1135 => x"fb",
          1136 => x"0b",
          1137 => x"f4",
          1138 => x"ff",
          1139 => x"56",
          1140 => x"84",
          1141 => x"2e",
          1142 => x"c0",
          1143 => x"70",
          1144 => x"2a",
          1145 => x"53",
          1146 => x"80",
          1147 => x"71",
          1148 => x"81",
          1149 => x"70",
          1150 => x"81",
          1151 => x"06",
          1152 => x"80",
          1153 => x"71",
          1154 => x"81",
          1155 => x"70",
          1156 => x"73",
          1157 => x"51",
          1158 => x"80",
          1159 => x"2e",
          1160 => x"c0",
          1161 => x"75",
          1162 => x"81",
          1163 => x"87",
          1164 => x"fb",
          1165 => x"9f",
          1166 => x"0b",
          1167 => x"33",
          1168 => x"06",
          1169 => x"87",
          1170 => x"51",
          1171 => x"86",
          1172 => x"94",
          1173 => x"08",
          1174 => x"70",
          1175 => x"54",
          1176 => x"2e",
          1177 => x"91",
          1178 => x"06",
          1179 => x"d7",
          1180 => x"32",
          1181 => x"51",
          1182 => x"2e",
          1183 => x"93",
          1184 => x"06",
          1185 => x"ff",
          1186 => x"81",
          1187 => x"87",
          1188 => x"52",
          1189 => x"86",
          1190 => x"94",
          1191 => x"72",
          1192 => x"0d",
          1193 => x"0d",
          1194 => x"74",
          1195 => x"ff",
          1196 => x"57",
          1197 => x"80",
          1198 => x"81",
          1199 => x"15",
          1200 => x"d8",
          1201 => x"81",
          1202 => x"57",
          1203 => x"c0",
          1204 => x"75",
          1205 => x"38",
          1206 => x"94",
          1207 => x"70",
          1208 => x"81",
          1209 => x"52",
          1210 => x"8c",
          1211 => x"2a",
          1212 => x"51",
          1213 => x"38",
          1214 => x"70",
          1215 => x"51",
          1216 => x"8d",
          1217 => x"2a",
          1218 => x"51",
          1219 => x"be",
          1220 => x"ff",
          1221 => x"c0",
          1222 => x"70",
          1223 => x"38",
          1224 => x"90",
          1225 => x"0c",
          1226 => x"33",
          1227 => x"06",
          1228 => x"70",
          1229 => x"76",
          1230 => x"0c",
          1231 => x"04",
          1232 => x"0b",
          1233 => x"f4",
          1234 => x"ff",
          1235 => x"87",
          1236 => x"51",
          1237 => x"86",
          1238 => x"94",
          1239 => x"08",
          1240 => x"70",
          1241 => x"51",
          1242 => x"2e",
          1243 => x"81",
          1244 => x"87",
          1245 => x"52",
          1246 => x"86",
          1247 => x"94",
          1248 => x"08",
          1249 => x"06",
          1250 => x"0c",
          1251 => x"0d",
          1252 => x"0d",
          1253 => x"d8",
          1254 => x"81",
          1255 => x"53",
          1256 => x"84",
          1257 => x"2e",
          1258 => x"c0",
          1259 => x"71",
          1260 => x"2a",
          1261 => x"51",
          1262 => x"52",
          1263 => x"a0",
          1264 => x"ff",
          1265 => x"c0",
          1266 => x"70",
          1267 => x"38",
          1268 => x"90",
          1269 => x"70",
          1270 => x"98",
          1271 => x"51",
          1272 => x"cc",
          1273 => x"0d",
          1274 => x"0d",
          1275 => x"80",
          1276 => x"2a",
          1277 => x"51",
          1278 => x"84",
          1279 => x"c0",
          1280 => x"81",
          1281 => x"87",
          1282 => x"08",
          1283 => x"0c",
          1284 => x"94",
          1285 => x"80",
          1286 => x"9e",
          1287 => x"d9",
          1288 => x"c0",
          1289 => x"81",
          1290 => x"87",
          1291 => x"08",
          1292 => x"0c",
          1293 => x"ac",
          1294 => x"90",
          1295 => x"9e",
          1296 => x"d9",
          1297 => x"c0",
          1298 => x"81",
          1299 => x"87",
          1300 => x"08",
          1301 => x"0c",
          1302 => x"bc",
          1303 => x"a0",
          1304 => x"9e",
          1305 => x"d9",
          1306 => x"c0",
          1307 => x"81",
          1308 => x"87",
          1309 => x"08",
          1310 => x"d9",
          1311 => x"c0",
          1312 => x"81",
          1313 => x"87",
          1314 => x"08",
          1315 => x"0c",
          1316 => x"8c",
          1317 => x"b8",
          1318 => x"81",
          1319 => x"80",
          1320 => x"9e",
          1321 => x"84",
          1322 => x"51",
          1323 => x"80",
          1324 => x"81",
          1325 => x"d9",
          1326 => x"0b",
          1327 => x"90",
          1328 => x"80",
          1329 => x"52",
          1330 => x"2e",
          1331 => x"52",
          1332 => x"be",
          1333 => x"87",
          1334 => x"08",
          1335 => x"0a",
          1336 => x"52",
          1337 => x"83",
          1338 => x"71",
          1339 => x"34",
          1340 => x"c0",
          1341 => x"70",
          1342 => x"06",
          1343 => x"70",
          1344 => x"38",
          1345 => x"81",
          1346 => x"80",
          1347 => x"9e",
          1348 => x"a0",
          1349 => x"51",
          1350 => x"80",
          1351 => x"81",
          1352 => x"d9",
          1353 => x"0b",
          1354 => x"90",
          1355 => x"80",
          1356 => x"52",
          1357 => x"2e",
          1358 => x"52",
          1359 => x"c2",
          1360 => x"87",
          1361 => x"08",
          1362 => x"80",
          1363 => x"52",
          1364 => x"83",
          1365 => x"71",
          1366 => x"34",
          1367 => x"c0",
          1368 => x"70",
          1369 => x"06",
          1370 => x"70",
          1371 => x"38",
          1372 => x"81",
          1373 => x"80",
          1374 => x"9e",
          1375 => x"81",
          1376 => x"51",
          1377 => x"80",
          1378 => x"81",
          1379 => x"d9",
          1380 => x"0b",
          1381 => x"90",
          1382 => x"c0",
          1383 => x"52",
          1384 => x"2e",
          1385 => x"52",
          1386 => x"c6",
          1387 => x"87",
          1388 => x"08",
          1389 => x"06",
          1390 => x"70",
          1391 => x"38",
          1392 => x"81",
          1393 => x"87",
          1394 => x"08",
          1395 => x"06",
          1396 => x"51",
          1397 => x"81",
          1398 => x"80",
          1399 => x"9e",
          1400 => x"84",
          1401 => x"52",
          1402 => x"2e",
          1403 => x"52",
          1404 => x"c9",
          1405 => x"9e",
          1406 => x"83",
          1407 => x"84",
          1408 => x"51",
          1409 => x"ca",
          1410 => x"87",
          1411 => x"08",
          1412 => x"51",
          1413 => x"80",
          1414 => x"81",
          1415 => x"d9",
          1416 => x"c0",
          1417 => x"70",
          1418 => x"51",
          1419 => x"cc",
          1420 => x"0d",
          1421 => x"0d",
          1422 => x"51",
          1423 => x"81",
          1424 => x"54",
          1425 => x"88",
          1426 => x"f8",
          1427 => x"3f",
          1428 => x"51",
          1429 => x"81",
          1430 => x"54",
          1431 => x"93",
          1432 => x"98",
          1433 => x"9c",
          1434 => x"52",
          1435 => x"51",
          1436 => x"81",
          1437 => x"54",
          1438 => x"93",
          1439 => x"90",
          1440 => x"94",
          1441 => x"52",
          1442 => x"51",
          1443 => x"81",
          1444 => x"54",
          1445 => x"93",
          1446 => x"f8",
          1447 => x"fc",
          1448 => x"52",
          1449 => x"51",
          1450 => x"81",
          1451 => x"54",
          1452 => x"93",
          1453 => x"80",
          1454 => x"84",
          1455 => x"52",
          1456 => x"51",
          1457 => x"81",
          1458 => x"54",
          1459 => x"93",
          1460 => x"88",
          1461 => x"8c",
          1462 => x"52",
          1463 => x"51",
          1464 => x"81",
          1465 => x"54",
          1466 => x"8d",
          1467 => x"c8",
          1468 => x"c7",
          1469 => x"ef",
          1470 => x"cb",
          1471 => x"80",
          1472 => x"81",
          1473 => x"52",
          1474 => x"51",
          1475 => x"81",
          1476 => x"54",
          1477 => x"8d",
          1478 => x"ca",
          1479 => x"c7",
          1480 => x"c3",
          1481 => x"bd",
          1482 => x"80",
          1483 => x"81",
          1484 => x"83",
          1485 => x"d9",
          1486 => x"73",
          1487 => x"38",
          1488 => x"51",
          1489 => x"81",
          1490 => x"54",
          1491 => x"88",
          1492 => x"b0",
          1493 => x"3f",
          1494 => x"33",
          1495 => x"2e",
          1496 => x"c8",
          1497 => x"9b",
          1498 => x"c6",
          1499 => x"80",
          1500 => x"81",
          1501 => x"83",
          1502 => x"c8",
          1503 => x"83",
          1504 => x"a0",
          1505 => x"c8",
          1506 => x"db",
          1507 => x"a4",
          1508 => x"c9",
          1509 => x"cf",
          1510 => x"a8",
          1511 => x"c9",
          1512 => x"c3",
          1513 => x"d8",
          1514 => x"3f",
          1515 => x"22",
          1516 => x"e0",
          1517 => x"3f",
          1518 => x"08",
          1519 => x"c0",
          1520 => x"e7",
          1521 => x"dc",
          1522 => x"84",
          1523 => x"71",
          1524 => x"81",
          1525 => x"52",
          1526 => x"51",
          1527 => x"81",
          1528 => x"54",
          1529 => x"a8",
          1530 => x"b4",
          1531 => x"84",
          1532 => x"51",
          1533 => x"81",
          1534 => x"bd",
          1535 => x"76",
          1536 => x"54",
          1537 => x"08",
          1538 => x"b4",
          1539 => x"3f",
          1540 => x"33",
          1541 => x"2e",
          1542 => x"d9",
          1543 => x"bd",
          1544 => x"75",
          1545 => x"3f",
          1546 => x"08",
          1547 => x"29",
          1548 => x"54",
          1549 => x"cc",
          1550 => x"ca",
          1551 => x"a7",
          1552 => x"c4",
          1553 => x"3f",
          1554 => x"04",
          1555 => x"02",
          1556 => x"ff",
          1557 => x"84",
          1558 => x"71",
          1559 => x"c4",
          1560 => x"71",
          1561 => x"cb",
          1562 => x"39",
          1563 => x"51",
          1564 => x"cb",
          1565 => x"39",
          1566 => x"51",
          1567 => x"cb",
          1568 => x"39",
          1569 => x"51",
          1570 => x"84",
          1571 => x"71",
          1572 => x"04",
          1573 => x"c0",
          1574 => x"04",
          1575 => x"08",
          1576 => x"84",
          1577 => x"3d",
          1578 => x"05",
          1579 => x"8a",
          1580 => x"06",
          1581 => x"51",
          1582 => x"dc",
          1583 => x"71",
          1584 => x"38",
          1585 => x"81",
          1586 => x"81",
          1587 => x"e4",
          1588 => x"81",
          1589 => x"52",
          1590 => x"85",
          1591 => x"71",
          1592 => x"0d",
          1593 => x"0d",
          1594 => x"33",
          1595 => x"08",
          1596 => x"dc",
          1597 => x"ff",
          1598 => x"81",
          1599 => x"84",
          1600 => x"fd",
          1601 => x"54",
          1602 => x"81",
          1603 => x"53",
          1604 => x"8e",
          1605 => x"ff",
          1606 => x"14",
          1607 => x"3f",
          1608 => x"3d",
          1609 => x"3d",
          1610 => x"dc",
          1611 => x"81",
          1612 => x"56",
          1613 => x"70",
          1614 => x"53",
          1615 => x"2e",
          1616 => x"81",
          1617 => x"81",
          1618 => x"da",
          1619 => x"74",
          1620 => x"0c",
          1621 => x"04",
          1622 => x"66",
          1623 => x"78",
          1624 => x"5a",
          1625 => x"80",
          1626 => x"38",
          1627 => x"09",
          1628 => x"de",
          1629 => x"7a",
          1630 => x"5c",
          1631 => x"5b",
          1632 => x"09",
          1633 => x"38",
          1634 => x"39",
          1635 => x"09",
          1636 => x"38",
          1637 => x"70",
          1638 => x"33",
          1639 => x"2e",
          1640 => x"92",
          1641 => x"19",
          1642 => x"70",
          1643 => x"33",
          1644 => x"53",
          1645 => x"16",
          1646 => x"26",
          1647 => x"88",
          1648 => x"05",
          1649 => x"05",
          1650 => x"05",
          1651 => x"5b",
          1652 => x"80",
          1653 => x"30",
          1654 => x"80",
          1655 => x"cc",
          1656 => x"70",
          1657 => x"25",
          1658 => x"54",
          1659 => x"53",
          1660 => x"8c",
          1661 => x"07",
          1662 => x"05",
          1663 => x"5a",
          1664 => x"83",
          1665 => x"54",
          1666 => x"27",
          1667 => x"16",
          1668 => x"06",
          1669 => x"80",
          1670 => x"aa",
          1671 => x"cf",
          1672 => x"73",
          1673 => x"81",
          1674 => x"80",
          1675 => x"38",
          1676 => x"2e",
          1677 => x"81",
          1678 => x"80",
          1679 => x"8a",
          1680 => x"39",
          1681 => x"2e",
          1682 => x"73",
          1683 => x"8a",
          1684 => x"d3",
          1685 => x"80",
          1686 => x"80",
          1687 => x"ee",
          1688 => x"39",
          1689 => x"71",
          1690 => x"53",
          1691 => x"54",
          1692 => x"2e",
          1693 => x"15",
          1694 => x"33",
          1695 => x"72",
          1696 => x"81",
          1697 => x"39",
          1698 => x"56",
          1699 => x"27",
          1700 => x"51",
          1701 => x"75",
          1702 => x"72",
          1703 => x"38",
          1704 => x"df",
          1705 => x"16",
          1706 => x"7b",
          1707 => x"38",
          1708 => x"f2",
          1709 => x"77",
          1710 => x"12",
          1711 => x"53",
          1712 => x"5c",
          1713 => x"5c",
          1714 => x"5c",
          1715 => x"5c",
          1716 => x"51",
          1717 => x"fd",
          1718 => x"82",
          1719 => x"06",
          1720 => x"80",
          1721 => x"77",
          1722 => x"53",
          1723 => x"18",
          1724 => x"72",
          1725 => x"c4",
          1726 => x"70",
          1727 => x"25",
          1728 => x"55",
          1729 => x"8d",
          1730 => x"2e",
          1731 => x"30",
          1732 => x"5b",
          1733 => x"8f",
          1734 => x"7b",
          1735 => x"e1",
          1736 => x"dc",
          1737 => x"ff",
          1738 => x"75",
          1739 => x"cc",
          1740 => x"cc",
          1741 => x"74",
          1742 => x"a7",
          1743 => x"80",
          1744 => x"38",
          1745 => x"72",
          1746 => x"54",
          1747 => x"72",
          1748 => x"05",
          1749 => x"17",
          1750 => x"77",
          1751 => x"51",
          1752 => x"9f",
          1753 => x"72",
          1754 => x"79",
          1755 => x"81",
          1756 => x"72",
          1757 => x"38",
          1758 => x"05",
          1759 => x"ad",
          1760 => x"17",
          1761 => x"81",
          1762 => x"b0",
          1763 => x"38",
          1764 => x"81",
          1765 => x"06",
          1766 => x"9f",
          1767 => x"55",
          1768 => x"97",
          1769 => x"f9",
          1770 => x"81",
          1771 => x"8b",
          1772 => x"16",
          1773 => x"73",
          1774 => x"96",
          1775 => x"e0",
          1776 => x"17",
          1777 => x"33",
          1778 => x"f9",
          1779 => x"f2",
          1780 => x"16",
          1781 => x"7b",
          1782 => x"38",
          1783 => x"c6",
          1784 => x"96",
          1785 => x"fd",
          1786 => x"3d",
          1787 => x"05",
          1788 => x"52",
          1789 => x"e0",
          1790 => x"0d",
          1791 => x"0d",
          1792 => x"e4",
          1793 => x"88",
          1794 => x"51",
          1795 => x"81",
          1796 => x"53",
          1797 => x"80",
          1798 => x"e4",
          1799 => x"0d",
          1800 => x"0d",
          1801 => x"08",
          1802 => x"dc",
          1803 => x"88",
          1804 => x"52",
          1805 => x"3f",
          1806 => x"dc",
          1807 => x"0d",
          1808 => x"0d",
          1809 => x"dc",
          1810 => x"56",
          1811 => x"80",
          1812 => x"2e",
          1813 => x"81",
          1814 => x"52",
          1815 => x"dc",
          1816 => x"ff",
          1817 => x"80",
          1818 => x"38",
          1819 => x"b9",
          1820 => x"32",
          1821 => x"80",
          1822 => x"52",
          1823 => x"8b",
          1824 => x"2e",
          1825 => x"14",
          1826 => x"9f",
          1827 => x"38",
          1828 => x"73",
          1829 => x"38",
          1830 => x"72",
          1831 => x"14",
          1832 => x"f8",
          1833 => x"af",
          1834 => x"52",
          1835 => x"8a",
          1836 => x"3f",
          1837 => x"81",
          1838 => x"87",
          1839 => x"fe",
          1840 => x"dc",
          1841 => x"81",
          1842 => x"77",
          1843 => x"53",
          1844 => x"72",
          1845 => x"0c",
          1846 => x"04",
          1847 => x"7a",
          1848 => x"80",
          1849 => x"58",
          1850 => x"33",
          1851 => x"a0",
          1852 => x"06",
          1853 => x"13",
          1854 => x"39",
          1855 => x"09",
          1856 => x"38",
          1857 => x"11",
          1858 => x"08",
          1859 => x"54",
          1860 => x"2e",
          1861 => x"80",
          1862 => x"08",
          1863 => x"0c",
          1864 => x"33",
          1865 => x"80",
          1866 => x"38",
          1867 => x"80",
          1868 => x"38",
          1869 => x"57",
          1870 => x"0c",
          1871 => x"33",
          1872 => x"39",
          1873 => x"74",
          1874 => x"38",
          1875 => x"80",
          1876 => x"89",
          1877 => x"38",
          1878 => x"d0",
          1879 => x"55",
          1880 => x"80",
          1881 => x"39",
          1882 => x"d9",
          1883 => x"80",
          1884 => x"27",
          1885 => x"80",
          1886 => x"89",
          1887 => x"70",
          1888 => x"55",
          1889 => x"70",
          1890 => x"55",
          1891 => x"27",
          1892 => x"14",
          1893 => x"06",
          1894 => x"74",
          1895 => x"73",
          1896 => x"38",
          1897 => x"14",
          1898 => x"05",
          1899 => x"08",
          1900 => x"54",
          1901 => x"39",
          1902 => x"84",
          1903 => x"55",
          1904 => x"81",
          1905 => x"dc",
          1906 => x"3d",
          1907 => x"3d",
          1908 => x"5a",
          1909 => x"7a",
          1910 => x"08",
          1911 => x"53",
          1912 => x"09",
          1913 => x"38",
          1914 => x"0c",
          1915 => x"ad",
          1916 => x"06",
          1917 => x"76",
          1918 => x"0c",
          1919 => x"33",
          1920 => x"73",
          1921 => x"81",
          1922 => x"38",
          1923 => x"05",
          1924 => x"08",
          1925 => x"53",
          1926 => x"2e",
          1927 => x"57",
          1928 => x"2e",
          1929 => x"39",
          1930 => x"13",
          1931 => x"08",
          1932 => x"53",
          1933 => x"55",
          1934 => x"80",
          1935 => x"14",
          1936 => x"88",
          1937 => x"27",
          1938 => x"eb",
          1939 => x"53",
          1940 => x"89",
          1941 => x"38",
          1942 => x"55",
          1943 => x"8a",
          1944 => x"a0",
          1945 => x"c2",
          1946 => x"74",
          1947 => x"e0",
          1948 => x"ff",
          1949 => x"d0",
          1950 => x"ff",
          1951 => x"90",
          1952 => x"38",
          1953 => x"81",
          1954 => x"53",
          1955 => x"ca",
          1956 => x"27",
          1957 => x"77",
          1958 => x"08",
          1959 => x"0c",
          1960 => x"33",
          1961 => x"ff",
          1962 => x"80",
          1963 => x"74",
          1964 => x"79",
          1965 => x"74",
          1966 => x"0c",
          1967 => x"04",
          1968 => x"02",
          1969 => x"51",
          1970 => x"72",
          1971 => x"81",
          1972 => x"33",
          1973 => x"dc",
          1974 => x"3d",
          1975 => x"3d",
          1976 => x"05",
          1977 => x"05",
          1978 => x"56",
          1979 => x"72",
          1980 => x"e0",
          1981 => x"2b",
          1982 => x"8c",
          1983 => x"88",
          1984 => x"2e",
          1985 => x"88",
          1986 => x"0c",
          1987 => x"8c",
          1988 => x"71",
          1989 => x"87",
          1990 => x"0c",
          1991 => x"08",
          1992 => x"51",
          1993 => x"2e",
          1994 => x"c0",
          1995 => x"51",
          1996 => x"71",
          1997 => x"80",
          1998 => x"92",
          1999 => x"98",
          2000 => x"70",
          2001 => x"38",
          2002 => x"d4",
          2003 => x"d9",
          2004 => x"51",
          2005 => x"cc",
          2006 => x"0d",
          2007 => x"0d",
          2008 => x"02",
          2009 => x"05",
          2010 => x"58",
          2011 => x"52",
          2012 => x"3f",
          2013 => x"08",
          2014 => x"54",
          2015 => x"be",
          2016 => x"75",
          2017 => x"c0",
          2018 => x"87",
          2019 => x"12",
          2020 => x"84",
          2021 => x"40",
          2022 => x"85",
          2023 => x"98",
          2024 => x"7d",
          2025 => x"0c",
          2026 => x"85",
          2027 => x"06",
          2028 => x"71",
          2029 => x"38",
          2030 => x"71",
          2031 => x"05",
          2032 => x"19",
          2033 => x"a2",
          2034 => x"71",
          2035 => x"38",
          2036 => x"83",
          2037 => x"38",
          2038 => x"8a",
          2039 => x"98",
          2040 => x"71",
          2041 => x"c0",
          2042 => x"52",
          2043 => x"87",
          2044 => x"80",
          2045 => x"81",
          2046 => x"c0",
          2047 => x"53",
          2048 => x"82",
          2049 => x"71",
          2050 => x"1a",
          2051 => x"84",
          2052 => x"19",
          2053 => x"06",
          2054 => x"79",
          2055 => x"38",
          2056 => x"80",
          2057 => x"87",
          2058 => x"26",
          2059 => x"73",
          2060 => x"06",
          2061 => x"2e",
          2062 => x"52",
          2063 => x"81",
          2064 => x"8f",
          2065 => x"f3",
          2066 => x"62",
          2067 => x"05",
          2068 => x"57",
          2069 => x"83",
          2070 => x"52",
          2071 => x"3f",
          2072 => x"08",
          2073 => x"54",
          2074 => x"2e",
          2075 => x"81",
          2076 => x"74",
          2077 => x"c0",
          2078 => x"87",
          2079 => x"12",
          2080 => x"84",
          2081 => x"5f",
          2082 => x"0b",
          2083 => x"8c",
          2084 => x"0c",
          2085 => x"80",
          2086 => x"70",
          2087 => x"81",
          2088 => x"54",
          2089 => x"8c",
          2090 => x"81",
          2091 => x"7c",
          2092 => x"58",
          2093 => x"70",
          2094 => x"52",
          2095 => x"8a",
          2096 => x"98",
          2097 => x"71",
          2098 => x"c0",
          2099 => x"52",
          2100 => x"87",
          2101 => x"80",
          2102 => x"81",
          2103 => x"c0",
          2104 => x"53",
          2105 => x"82",
          2106 => x"71",
          2107 => x"19",
          2108 => x"81",
          2109 => x"ff",
          2110 => x"19",
          2111 => x"78",
          2112 => x"38",
          2113 => x"80",
          2114 => x"87",
          2115 => x"26",
          2116 => x"73",
          2117 => x"06",
          2118 => x"2e",
          2119 => x"52",
          2120 => x"81",
          2121 => x"8f",
          2122 => x"fa",
          2123 => x"02",
          2124 => x"05",
          2125 => x"05",
          2126 => x"71",
          2127 => x"57",
          2128 => x"81",
          2129 => x"81",
          2130 => x"54",
          2131 => x"38",
          2132 => x"c0",
          2133 => x"81",
          2134 => x"2e",
          2135 => x"71",
          2136 => x"38",
          2137 => x"87",
          2138 => x"11",
          2139 => x"80",
          2140 => x"80",
          2141 => x"83",
          2142 => x"38",
          2143 => x"72",
          2144 => x"2a",
          2145 => x"51",
          2146 => x"80",
          2147 => x"87",
          2148 => x"08",
          2149 => x"38",
          2150 => x"8c",
          2151 => x"96",
          2152 => x"0c",
          2153 => x"8c",
          2154 => x"08",
          2155 => x"51",
          2156 => x"38",
          2157 => x"56",
          2158 => x"80",
          2159 => x"85",
          2160 => x"77",
          2161 => x"83",
          2162 => x"75",
          2163 => x"dc",
          2164 => x"3d",
          2165 => x"3d",
          2166 => x"11",
          2167 => x"71",
          2168 => x"81",
          2169 => x"53",
          2170 => x"0d",
          2171 => x"0d",
          2172 => x"33",
          2173 => x"71",
          2174 => x"88",
          2175 => x"14",
          2176 => x"07",
          2177 => x"33",
          2178 => x"dc",
          2179 => x"53",
          2180 => x"52",
          2181 => x"04",
          2182 => x"73",
          2183 => x"92",
          2184 => x"52",
          2185 => x"81",
          2186 => x"70",
          2187 => x"70",
          2188 => x"3d",
          2189 => x"3d",
          2190 => x"52",
          2191 => x"70",
          2192 => x"34",
          2193 => x"51",
          2194 => x"81",
          2195 => x"70",
          2196 => x"70",
          2197 => x"05",
          2198 => x"88",
          2199 => x"72",
          2200 => x"0d",
          2201 => x"0d",
          2202 => x"54",
          2203 => x"80",
          2204 => x"71",
          2205 => x"53",
          2206 => x"81",
          2207 => x"ff",
          2208 => x"39",
          2209 => x"04",
          2210 => x"75",
          2211 => x"52",
          2212 => x"70",
          2213 => x"34",
          2214 => x"70",
          2215 => x"3d",
          2216 => x"3d",
          2217 => x"79",
          2218 => x"74",
          2219 => x"56",
          2220 => x"81",
          2221 => x"71",
          2222 => x"16",
          2223 => x"52",
          2224 => x"86",
          2225 => x"2e",
          2226 => x"81",
          2227 => x"86",
          2228 => x"fe",
          2229 => x"76",
          2230 => x"39",
          2231 => x"8a",
          2232 => x"51",
          2233 => x"71",
          2234 => x"33",
          2235 => x"0c",
          2236 => x"04",
          2237 => x"dc",
          2238 => x"80",
          2239 => x"cc",
          2240 => x"3d",
          2241 => x"80",
          2242 => x"33",
          2243 => x"7a",
          2244 => x"38",
          2245 => x"16",
          2246 => x"16",
          2247 => x"17",
          2248 => x"fa",
          2249 => x"dc",
          2250 => x"2e",
          2251 => x"b7",
          2252 => x"cc",
          2253 => x"34",
          2254 => x"70",
          2255 => x"31",
          2256 => x"59",
          2257 => x"77",
          2258 => x"82",
          2259 => x"74",
          2260 => x"81",
          2261 => x"81",
          2262 => x"53",
          2263 => x"16",
          2264 => x"e3",
          2265 => x"81",
          2266 => x"dc",
          2267 => x"3d",
          2268 => x"3d",
          2269 => x"56",
          2270 => x"74",
          2271 => x"2e",
          2272 => x"51",
          2273 => x"81",
          2274 => x"57",
          2275 => x"08",
          2276 => x"54",
          2277 => x"16",
          2278 => x"33",
          2279 => x"3f",
          2280 => x"08",
          2281 => x"38",
          2282 => x"57",
          2283 => x"0c",
          2284 => x"cc",
          2285 => x"0d",
          2286 => x"0d",
          2287 => x"57",
          2288 => x"81",
          2289 => x"58",
          2290 => x"08",
          2291 => x"76",
          2292 => x"83",
          2293 => x"06",
          2294 => x"84",
          2295 => x"78",
          2296 => x"81",
          2297 => x"38",
          2298 => x"81",
          2299 => x"52",
          2300 => x"52",
          2301 => x"3f",
          2302 => x"52",
          2303 => x"51",
          2304 => x"84",
          2305 => x"d2",
          2306 => x"fc",
          2307 => x"8a",
          2308 => x"52",
          2309 => x"51",
          2310 => x"90",
          2311 => x"84",
          2312 => x"fc",
          2313 => x"17",
          2314 => x"a0",
          2315 => x"86",
          2316 => x"08",
          2317 => x"b0",
          2318 => x"55",
          2319 => x"81",
          2320 => x"f8",
          2321 => x"84",
          2322 => x"53",
          2323 => x"17",
          2324 => x"d7",
          2325 => x"cc",
          2326 => x"83",
          2327 => x"77",
          2328 => x"0c",
          2329 => x"04",
          2330 => x"77",
          2331 => x"12",
          2332 => x"55",
          2333 => x"56",
          2334 => x"8d",
          2335 => x"22",
          2336 => x"ac",
          2337 => x"57",
          2338 => x"dc",
          2339 => x"3d",
          2340 => x"3d",
          2341 => x"70",
          2342 => x"57",
          2343 => x"81",
          2344 => x"98",
          2345 => x"81",
          2346 => x"74",
          2347 => x"72",
          2348 => x"f5",
          2349 => x"24",
          2350 => x"81",
          2351 => x"81",
          2352 => x"83",
          2353 => x"38",
          2354 => x"76",
          2355 => x"70",
          2356 => x"16",
          2357 => x"74",
          2358 => x"96",
          2359 => x"cc",
          2360 => x"38",
          2361 => x"06",
          2362 => x"33",
          2363 => x"89",
          2364 => x"08",
          2365 => x"54",
          2366 => x"fc",
          2367 => x"dc",
          2368 => x"fe",
          2369 => x"ff",
          2370 => x"11",
          2371 => x"2b",
          2372 => x"81",
          2373 => x"2a",
          2374 => x"51",
          2375 => x"e2",
          2376 => x"ff",
          2377 => x"da",
          2378 => x"2a",
          2379 => x"05",
          2380 => x"fc",
          2381 => x"dc",
          2382 => x"c6",
          2383 => x"83",
          2384 => x"05",
          2385 => x"f9",
          2386 => x"dc",
          2387 => x"ff",
          2388 => x"ae",
          2389 => x"2a",
          2390 => x"05",
          2391 => x"fc",
          2392 => x"dc",
          2393 => x"38",
          2394 => x"83",
          2395 => x"05",
          2396 => x"f8",
          2397 => x"dc",
          2398 => x"0a",
          2399 => x"39",
          2400 => x"81",
          2401 => x"89",
          2402 => x"f8",
          2403 => x"7c",
          2404 => x"56",
          2405 => x"77",
          2406 => x"38",
          2407 => x"08",
          2408 => x"38",
          2409 => x"72",
          2410 => x"9d",
          2411 => x"24",
          2412 => x"81",
          2413 => x"82",
          2414 => x"83",
          2415 => x"38",
          2416 => x"76",
          2417 => x"70",
          2418 => x"18",
          2419 => x"76",
          2420 => x"9e",
          2421 => x"cc",
          2422 => x"dc",
          2423 => x"d9",
          2424 => x"ff",
          2425 => x"05",
          2426 => x"81",
          2427 => x"54",
          2428 => x"80",
          2429 => x"77",
          2430 => x"f0",
          2431 => x"8f",
          2432 => x"51",
          2433 => x"34",
          2434 => x"17",
          2435 => x"2a",
          2436 => x"05",
          2437 => x"fa",
          2438 => x"dc",
          2439 => x"81",
          2440 => x"81",
          2441 => x"83",
          2442 => x"b4",
          2443 => x"2a",
          2444 => x"8f",
          2445 => x"2a",
          2446 => x"f0",
          2447 => x"06",
          2448 => x"72",
          2449 => x"ec",
          2450 => x"2a",
          2451 => x"05",
          2452 => x"fa",
          2453 => x"dc",
          2454 => x"81",
          2455 => x"80",
          2456 => x"83",
          2457 => x"52",
          2458 => x"fe",
          2459 => x"b4",
          2460 => x"a4",
          2461 => x"76",
          2462 => x"17",
          2463 => x"75",
          2464 => x"3f",
          2465 => x"08",
          2466 => x"cc",
          2467 => x"77",
          2468 => x"77",
          2469 => x"fc",
          2470 => x"b4",
          2471 => x"51",
          2472 => x"c9",
          2473 => x"cc",
          2474 => x"06",
          2475 => x"72",
          2476 => x"3f",
          2477 => x"17",
          2478 => x"dc",
          2479 => x"3d",
          2480 => x"3d",
          2481 => x"7e",
          2482 => x"56",
          2483 => x"75",
          2484 => x"74",
          2485 => x"27",
          2486 => x"80",
          2487 => x"ff",
          2488 => x"75",
          2489 => x"3f",
          2490 => x"08",
          2491 => x"cc",
          2492 => x"38",
          2493 => x"54",
          2494 => x"81",
          2495 => x"39",
          2496 => x"08",
          2497 => x"39",
          2498 => x"51",
          2499 => x"81",
          2500 => x"58",
          2501 => x"08",
          2502 => x"c7",
          2503 => x"cc",
          2504 => x"d2",
          2505 => x"cc",
          2506 => x"cf",
          2507 => x"74",
          2508 => x"fc",
          2509 => x"dc",
          2510 => x"38",
          2511 => x"fe",
          2512 => x"08",
          2513 => x"74",
          2514 => x"38",
          2515 => x"17",
          2516 => x"33",
          2517 => x"73",
          2518 => x"77",
          2519 => x"26",
          2520 => x"80",
          2521 => x"dc",
          2522 => x"3d",
          2523 => x"3d",
          2524 => x"71",
          2525 => x"5b",
          2526 => x"8c",
          2527 => x"77",
          2528 => x"38",
          2529 => x"78",
          2530 => x"81",
          2531 => x"79",
          2532 => x"f9",
          2533 => x"55",
          2534 => x"cc",
          2535 => x"e0",
          2536 => x"cc",
          2537 => x"dc",
          2538 => x"2e",
          2539 => x"98",
          2540 => x"dc",
          2541 => x"82",
          2542 => x"58",
          2543 => x"70",
          2544 => x"80",
          2545 => x"38",
          2546 => x"09",
          2547 => x"e2",
          2548 => x"56",
          2549 => x"76",
          2550 => x"82",
          2551 => x"7a",
          2552 => x"3f",
          2553 => x"dc",
          2554 => x"2e",
          2555 => x"86",
          2556 => x"cc",
          2557 => x"dc",
          2558 => x"70",
          2559 => x"07",
          2560 => x"7c",
          2561 => x"cc",
          2562 => x"51",
          2563 => x"81",
          2564 => x"dc",
          2565 => x"2e",
          2566 => x"17",
          2567 => x"74",
          2568 => x"73",
          2569 => x"27",
          2570 => x"58",
          2571 => x"80",
          2572 => x"56",
          2573 => x"98",
          2574 => x"26",
          2575 => x"56",
          2576 => x"81",
          2577 => x"52",
          2578 => x"c6",
          2579 => x"cc",
          2580 => x"b8",
          2581 => x"81",
          2582 => x"81",
          2583 => x"06",
          2584 => x"dc",
          2585 => x"81",
          2586 => x"09",
          2587 => x"72",
          2588 => x"70",
          2589 => x"51",
          2590 => x"80",
          2591 => x"78",
          2592 => x"06",
          2593 => x"73",
          2594 => x"39",
          2595 => x"52",
          2596 => x"f7",
          2597 => x"cc",
          2598 => x"cc",
          2599 => x"81",
          2600 => x"07",
          2601 => x"55",
          2602 => x"2e",
          2603 => x"80",
          2604 => x"75",
          2605 => x"76",
          2606 => x"3f",
          2607 => x"08",
          2608 => x"38",
          2609 => x"0c",
          2610 => x"fe",
          2611 => x"08",
          2612 => x"74",
          2613 => x"ff",
          2614 => x"0c",
          2615 => x"81",
          2616 => x"84",
          2617 => x"39",
          2618 => x"81",
          2619 => x"8c",
          2620 => x"8c",
          2621 => x"cc",
          2622 => x"39",
          2623 => x"55",
          2624 => x"cc",
          2625 => x"0d",
          2626 => x"0d",
          2627 => x"55",
          2628 => x"81",
          2629 => x"58",
          2630 => x"dc",
          2631 => x"d8",
          2632 => x"74",
          2633 => x"3f",
          2634 => x"08",
          2635 => x"08",
          2636 => x"59",
          2637 => x"77",
          2638 => x"70",
          2639 => x"c8",
          2640 => x"84",
          2641 => x"56",
          2642 => x"58",
          2643 => x"97",
          2644 => x"75",
          2645 => x"52",
          2646 => x"51",
          2647 => x"81",
          2648 => x"80",
          2649 => x"8a",
          2650 => x"32",
          2651 => x"72",
          2652 => x"2a",
          2653 => x"56",
          2654 => x"cc",
          2655 => x"0d",
          2656 => x"0d",
          2657 => x"08",
          2658 => x"74",
          2659 => x"26",
          2660 => x"74",
          2661 => x"72",
          2662 => x"74",
          2663 => x"88",
          2664 => x"73",
          2665 => x"33",
          2666 => x"27",
          2667 => x"16",
          2668 => x"9b",
          2669 => x"2a",
          2670 => x"88",
          2671 => x"58",
          2672 => x"80",
          2673 => x"16",
          2674 => x"0c",
          2675 => x"8a",
          2676 => x"89",
          2677 => x"72",
          2678 => x"38",
          2679 => x"51",
          2680 => x"81",
          2681 => x"54",
          2682 => x"08",
          2683 => x"38",
          2684 => x"dc",
          2685 => x"8b",
          2686 => x"08",
          2687 => x"08",
          2688 => x"82",
          2689 => x"74",
          2690 => x"cb",
          2691 => x"75",
          2692 => x"3f",
          2693 => x"08",
          2694 => x"73",
          2695 => x"98",
          2696 => x"82",
          2697 => x"2e",
          2698 => x"39",
          2699 => x"39",
          2700 => x"13",
          2701 => x"74",
          2702 => x"16",
          2703 => x"18",
          2704 => x"77",
          2705 => x"0c",
          2706 => x"04",
          2707 => x"7a",
          2708 => x"12",
          2709 => x"59",
          2710 => x"80",
          2711 => x"86",
          2712 => x"98",
          2713 => x"14",
          2714 => x"55",
          2715 => x"81",
          2716 => x"83",
          2717 => x"77",
          2718 => x"81",
          2719 => x"0c",
          2720 => x"55",
          2721 => x"76",
          2722 => x"17",
          2723 => x"74",
          2724 => x"9b",
          2725 => x"39",
          2726 => x"ff",
          2727 => x"2a",
          2728 => x"81",
          2729 => x"52",
          2730 => x"e6",
          2731 => x"cc",
          2732 => x"55",
          2733 => x"dc",
          2734 => x"80",
          2735 => x"55",
          2736 => x"08",
          2737 => x"f4",
          2738 => x"08",
          2739 => x"08",
          2740 => x"38",
          2741 => x"77",
          2742 => x"84",
          2743 => x"39",
          2744 => x"52",
          2745 => x"86",
          2746 => x"cc",
          2747 => x"55",
          2748 => x"08",
          2749 => x"c4",
          2750 => x"81",
          2751 => x"81",
          2752 => x"81",
          2753 => x"cc",
          2754 => x"b0",
          2755 => x"cc",
          2756 => x"51",
          2757 => x"81",
          2758 => x"a0",
          2759 => x"15",
          2760 => x"75",
          2761 => x"3f",
          2762 => x"08",
          2763 => x"76",
          2764 => x"77",
          2765 => x"9c",
          2766 => x"55",
          2767 => x"cc",
          2768 => x"0d",
          2769 => x"0d",
          2770 => x"08",
          2771 => x"80",
          2772 => x"fc",
          2773 => x"dc",
          2774 => x"81",
          2775 => x"80",
          2776 => x"dc",
          2777 => x"98",
          2778 => x"78",
          2779 => x"3f",
          2780 => x"08",
          2781 => x"cc",
          2782 => x"38",
          2783 => x"08",
          2784 => x"70",
          2785 => x"58",
          2786 => x"2e",
          2787 => x"83",
          2788 => x"81",
          2789 => x"55",
          2790 => x"81",
          2791 => x"07",
          2792 => x"2e",
          2793 => x"16",
          2794 => x"2e",
          2795 => x"88",
          2796 => x"81",
          2797 => x"56",
          2798 => x"51",
          2799 => x"81",
          2800 => x"54",
          2801 => x"08",
          2802 => x"9b",
          2803 => x"2e",
          2804 => x"83",
          2805 => x"73",
          2806 => x"0c",
          2807 => x"04",
          2808 => x"76",
          2809 => x"54",
          2810 => x"81",
          2811 => x"83",
          2812 => x"76",
          2813 => x"53",
          2814 => x"2e",
          2815 => x"90",
          2816 => x"51",
          2817 => x"81",
          2818 => x"90",
          2819 => x"53",
          2820 => x"cc",
          2821 => x"0d",
          2822 => x"0d",
          2823 => x"83",
          2824 => x"54",
          2825 => x"55",
          2826 => x"3f",
          2827 => x"51",
          2828 => x"2e",
          2829 => x"8b",
          2830 => x"2a",
          2831 => x"51",
          2832 => x"86",
          2833 => x"f7",
          2834 => x"7d",
          2835 => x"75",
          2836 => x"98",
          2837 => x"2e",
          2838 => x"98",
          2839 => x"78",
          2840 => x"3f",
          2841 => x"08",
          2842 => x"cc",
          2843 => x"38",
          2844 => x"70",
          2845 => x"73",
          2846 => x"58",
          2847 => x"8b",
          2848 => x"bf",
          2849 => x"ff",
          2850 => x"53",
          2851 => x"34",
          2852 => x"08",
          2853 => x"e5",
          2854 => x"81",
          2855 => x"2e",
          2856 => x"70",
          2857 => x"57",
          2858 => x"9e",
          2859 => x"2e",
          2860 => x"dc",
          2861 => x"df",
          2862 => x"72",
          2863 => x"81",
          2864 => x"76",
          2865 => x"2e",
          2866 => x"52",
          2867 => x"fc",
          2868 => x"cc",
          2869 => x"dc",
          2870 => x"38",
          2871 => x"fe",
          2872 => x"39",
          2873 => x"16",
          2874 => x"dc",
          2875 => x"3d",
          2876 => x"3d",
          2877 => x"08",
          2878 => x"52",
          2879 => x"c5",
          2880 => x"cc",
          2881 => x"dc",
          2882 => x"38",
          2883 => x"52",
          2884 => x"de",
          2885 => x"cc",
          2886 => x"dc",
          2887 => x"38",
          2888 => x"dc",
          2889 => x"9c",
          2890 => x"ea",
          2891 => x"53",
          2892 => x"9c",
          2893 => x"ea",
          2894 => x"0b",
          2895 => x"74",
          2896 => x"0c",
          2897 => x"04",
          2898 => x"75",
          2899 => x"12",
          2900 => x"53",
          2901 => x"9a",
          2902 => x"cc",
          2903 => x"9c",
          2904 => x"e5",
          2905 => x"0b",
          2906 => x"85",
          2907 => x"fa",
          2908 => x"7a",
          2909 => x"0b",
          2910 => x"98",
          2911 => x"2e",
          2912 => x"80",
          2913 => x"55",
          2914 => x"17",
          2915 => x"33",
          2916 => x"51",
          2917 => x"2e",
          2918 => x"85",
          2919 => x"06",
          2920 => x"e5",
          2921 => x"2e",
          2922 => x"8b",
          2923 => x"70",
          2924 => x"34",
          2925 => x"71",
          2926 => x"05",
          2927 => x"15",
          2928 => x"27",
          2929 => x"15",
          2930 => x"80",
          2931 => x"34",
          2932 => x"52",
          2933 => x"88",
          2934 => x"17",
          2935 => x"52",
          2936 => x"3f",
          2937 => x"08",
          2938 => x"12",
          2939 => x"3f",
          2940 => x"08",
          2941 => x"98",
          2942 => x"da",
          2943 => x"cc",
          2944 => x"23",
          2945 => x"04",
          2946 => x"7f",
          2947 => x"5b",
          2948 => x"33",
          2949 => x"73",
          2950 => x"38",
          2951 => x"80",
          2952 => x"38",
          2953 => x"8c",
          2954 => x"08",
          2955 => x"aa",
          2956 => x"41",
          2957 => x"33",
          2958 => x"73",
          2959 => x"81",
          2960 => x"81",
          2961 => x"dc",
          2962 => x"70",
          2963 => x"07",
          2964 => x"73",
          2965 => x"88",
          2966 => x"70",
          2967 => x"73",
          2968 => x"38",
          2969 => x"ab",
          2970 => x"52",
          2971 => x"91",
          2972 => x"cc",
          2973 => x"98",
          2974 => x"61",
          2975 => x"5a",
          2976 => x"a0",
          2977 => x"e7",
          2978 => x"70",
          2979 => x"79",
          2980 => x"73",
          2981 => x"81",
          2982 => x"38",
          2983 => x"33",
          2984 => x"ae",
          2985 => x"70",
          2986 => x"82",
          2987 => x"51",
          2988 => x"54",
          2989 => x"79",
          2990 => x"74",
          2991 => x"57",
          2992 => x"af",
          2993 => x"70",
          2994 => x"51",
          2995 => x"dc",
          2996 => x"73",
          2997 => x"38",
          2998 => x"82",
          2999 => x"19",
          3000 => x"54",
          3001 => x"82",
          3002 => x"54",
          3003 => x"78",
          3004 => x"81",
          3005 => x"54",
          3006 => x"81",
          3007 => x"af",
          3008 => x"77",
          3009 => x"70",
          3010 => x"25",
          3011 => x"07",
          3012 => x"51",
          3013 => x"2e",
          3014 => x"39",
          3015 => x"80",
          3016 => x"33",
          3017 => x"73",
          3018 => x"81",
          3019 => x"81",
          3020 => x"dc",
          3021 => x"70",
          3022 => x"07",
          3023 => x"73",
          3024 => x"b5",
          3025 => x"2e",
          3026 => x"83",
          3027 => x"76",
          3028 => x"07",
          3029 => x"2e",
          3030 => x"8b",
          3031 => x"77",
          3032 => x"30",
          3033 => x"71",
          3034 => x"53",
          3035 => x"55",
          3036 => x"38",
          3037 => x"5c",
          3038 => x"75",
          3039 => x"73",
          3040 => x"38",
          3041 => x"06",
          3042 => x"11",
          3043 => x"75",
          3044 => x"3f",
          3045 => x"08",
          3046 => x"38",
          3047 => x"33",
          3048 => x"54",
          3049 => x"e6",
          3050 => x"dc",
          3051 => x"2e",
          3052 => x"ff",
          3053 => x"74",
          3054 => x"38",
          3055 => x"75",
          3056 => x"17",
          3057 => x"57",
          3058 => x"a7",
          3059 => x"81",
          3060 => x"e5",
          3061 => x"dc",
          3062 => x"38",
          3063 => x"54",
          3064 => x"89",
          3065 => x"70",
          3066 => x"57",
          3067 => x"54",
          3068 => x"81",
          3069 => x"f7",
          3070 => x"7e",
          3071 => x"2e",
          3072 => x"33",
          3073 => x"e5",
          3074 => x"06",
          3075 => x"7a",
          3076 => x"a0",
          3077 => x"38",
          3078 => x"55",
          3079 => x"84",
          3080 => x"39",
          3081 => x"8b",
          3082 => x"7b",
          3083 => x"7a",
          3084 => x"3f",
          3085 => x"08",
          3086 => x"cc",
          3087 => x"38",
          3088 => x"52",
          3089 => x"aa",
          3090 => x"cc",
          3091 => x"dc",
          3092 => x"c2",
          3093 => x"08",
          3094 => x"55",
          3095 => x"ff",
          3096 => x"15",
          3097 => x"54",
          3098 => x"34",
          3099 => x"70",
          3100 => x"81",
          3101 => x"58",
          3102 => x"8b",
          3103 => x"74",
          3104 => x"3f",
          3105 => x"08",
          3106 => x"38",
          3107 => x"51",
          3108 => x"ff",
          3109 => x"ab",
          3110 => x"55",
          3111 => x"bb",
          3112 => x"2e",
          3113 => x"80",
          3114 => x"85",
          3115 => x"06",
          3116 => x"58",
          3117 => x"80",
          3118 => x"75",
          3119 => x"73",
          3120 => x"b5",
          3121 => x"0b",
          3122 => x"80",
          3123 => x"39",
          3124 => x"54",
          3125 => x"85",
          3126 => x"75",
          3127 => x"81",
          3128 => x"73",
          3129 => x"1b",
          3130 => x"2a",
          3131 => x"51",
          3132 => x"80",
          3133 => x"90",
          3134 => x"ff",
          3135 => x"05",
          3136 => x"f5",
          3137 => x"dc",
          3138 => x"1c",
          3139 => x"39",
          3140 => x"cc",
          3141 => x"0d",
          3142 => x"0d",
          3143 => x"7b",
          3144 => x"73",
          3145 => x"55",
          3146 => x"2e",
          3147 => x"75",
          3148 => x"57",
          3149 => x"26",
          3150 => x"ba",
          3151 => x"70",
          3152 => x"ba",
          3153 => x"06",
          3154 => x"73",
          3155 => x"70",
          3156 => x"51",
          3157 => x"89",
          3158 => x"82",
          3159 => x"ff",
          3160 => x"56",
          3161 => x"2e",
          3162 => x"80",
          3163 => x"8c",
          3164 => x"08",
          3165 => x"76",
          3166 => x"58",
          3167 => x"81",
          3168 => x"ff",
          3169 => x"53",
          3170 => x"26",
          3171 => x"13",
          3172 => x"06",
          3173 => x"9f",
          3174 => x"99",
          3175 => x"e0",
          3176 => x"ff",
          3177 => x"72",
          3178 => x"2a",
          3179 => x"72",
          3180 => x"06",
          3181 => x"ff",
          3182 => x"30",
          3183 => x"70",
          3184 => x"07",
          3185 => x"9f",
          3186 => x"54",
          3187 => x"80",
          3188 => x"81",
          3189 => x"59",
          3190 => x"25",
          3191 => x"8b",
          3192 => x"24",
          3193 => x"76",
          3194 => x"78",
          3195 => x"81",
          3196 => x"51",
          3197 => x"cc",
          3198 => x"0d",
          3199 => x"0d",
          3200 => x"0b",
          3201 => x"ff",
          3202 => x"0c",
          3203 => x"51",
          3204 => x"84",
          3205 => x"cc",
          3206 => x"38",
          3207 => x"51",
          3208 => x"81",
          3209 => x"83",
          3210 => x"54",
          3211 => x"82",
          3212 => x"09",
          3213 => x"e3",
          3214 => x"b4",
          3215 => x"57",
          3216 => x"2e",
          3217 => x"83",
          3218 => x"74",
          3219 => x"70",
          3220 => x"25",
          3221 => x"51",
          3222 => x"38",
          3223 => x"2e",
          3224 => x"b5",
          3225 => x"81",
          3226 => x"80",
          3227 => x"e0",
          3228 => x"dc",
          3229 => x"81",
          3230 => x"80",
          3231 => x"85",
          3232 => x"d0",
          3233 => x"16",
          3234 => x"3f",
          3235 => x"08",
          3236 => x"cc",
          3237 => x"83",
          3238 => x"74",
          3239 => x"0c",
          3240 => x"04",
          3241 => x"61",
          3242 => x"80",
          3243 => x"58",
          3244 => x"0c",
          3245 => x"e1",
          3246 => x"cc",
          3247 => x"56",
          3248 => x"dc",
          3249 => x"86",
          3250 => x"dc",
          3251 => x"29",
          3252 => x"05",
          3253 => x"53",
          3254 => x"80",
          3255 => x"38",
          3256 => x"76",
          3257 => x"74",
          3258 => x"72",
          3259 => x"38",
          3260 => x"51",
          3261 => x"81",
          3262 => x"81",
          3263 => x"81",
          3264 => x"72",
          3265 => x"80",
          3266 => x"38",
          3267 => x"70",
          3268 => x"53",
          3269 => x"86",
          3270 => x"a7",
          3271 => x"34",
          3272 => x"34",
          3273 => x"14",
          3274 => x"b2",
          3275 => x"cc",
          3276 => x"06",
          3277 => x"54",
          3278 => x"72",
          3279 => x"76",
          3280 => x"38",
          3281 => x"70",
          3282 => x"53",
          3283 => x"85",
          3284 => x"70",
          3285 => x"5b",
          3286 => x"81",
          3287 => x"81",
          3288 => x"76",
          3289 => x"81",
          3290 => x"38",
          3291 => x"56",
          3292 => x"83",
          3293 => x"70",
          3294 => x"80",
          3295 => x"83",
          3296 => x"dc",
          3297 => x"dc",
          3298 => x"76",
          3299 => x"05",
          3300 => x"16",
          3301 => x"56",
          3302 => x"d7",
          3303 => x"8d",
          3304 => x"72",
          3305 => x"54",
          3306 => x"57",
          3307 => x"95",
          3308 => x"73",
          3309 => x"3f",
          3310 => x"08",
          3311 => x"57",
          3312 => x"89",
          3313 => x"56",
          3314 => x"d7",
          3315 => x"76",
          3316 => x"f1",
          3317 => x"76",
          3318 => x"e9",
          3319 => x"51",
          3320 => x"81",
          3321 => x"83",
          3322 => x"53",
          3323 => x"2e",
          3324 => x"84",
          3325 => x"ca",
          3326 => x"da",
          3327 => x"cc",
          3328 => x"ff",
          3329 => x"8d",
          3330 => x"14",
          3331 => x"3f",
          3332 => x"08",
          3333 => x"15",
          3334 => x"14",
          3335 => x"34",
          3336 => x"33",
          3337 => x"81",
          3338 => x"54",
          3339 => x"72",
          3340 => x"91",
          3341 => x"ff",
          3342 => x"29",
          3343 => x"33",
          3344 => x"72",
          3345 => x"72",
          3346 => x"38",
          3347 => x"06",
          3348 => x"2e",
          3349 => x"56",
          3350 => x"80",
          3351 => x"da",
          3352 => x"dc",
          3353 => x"81",
          3354 => x"88",
          3355 => x"8f",
          3356 => x"56",
          3357 => x"38",
          3358 => x"51",
          3359 => x"81",
          3360 => x"83",
          3361 => x"55",
          3362 => x"80",
          3363 => x"da",
          3364 => x"dc",
          3365 => x"80",
          3366 => x"da",
          3367 => x"dc",
          3368 => x"ff",
          3369 => x"8d",
          3370 => x"2e",
          3371 => x"88",
          3372 => x"14",
          3373 => x"05",
          3374 => x"75",
          3375 => x"38",
          3376 => x"52",
          3377 => x"51",
          3378 => x"3f",
          3379 => x"08",
          3380 => x"cc",
          3381 => x"82",
          3382 => x"dc",
          3383 => x"ff",
          3384 => x"26",
          3385 => x"57",
          3386 => x"f5",
          3387 => x"82",
          3388 => x"f5",
          3389 => x"81",
          3390 => x"8d",
          3391 => x"2e",
          3392 => x"82",
          3393 => x"16",
          3394 => x"16",
          3395 => x"70",
          3396 => x"7a",
          3397 => x"0c",
          3398 => x"83",
          3399 => x"06",
          3400 => x"de",
          3401 => x"ae",
          3402 => x"cc",
          3403 => x"ff",
          3404 => x"56",
          3405 => x"38",
          3406 => x"38",
          3407 => x"51",
          3408 => x"81",
          3409 => x"a8",
          3410 => x"82",
          3411 => x"39",
          3412 => x"80",
          3413 => x"38",
          3414 => x"15",
          3415 => x"53",
          3416 => x"8d",
          3417 => x"15",
          3418 => x"76",
          3419 => x"51",
          3420 => x"13",
          3421 => x"8d",
          3422 => x"15",
          3423 => x"c5",
          3424 => x"90",
          3425 => x"0b",
          3426 => x"ff",
          3427 => x"15",
          3428 => x"2e",
          3429 => x"81",
          3430 => x"e4",
          3431 => x"b6",
          3432 => x"cc",
          3433 => x"ff",
          3434 => x"81",
          3435 => x"06",
          3436 => x"81",
          3437 => x"51",
          3438 => x"81",
          3439 => x"80",
          3440 => x"dc",
          3441 => x"15",
          3442 => x"14",
          3443 => x"3f",
          3444 => x"08",
          3445 => x"06",
          3446 => x"d4",
          3447 => x"81",
          3448 => x"38",
          3449 => x"d8",
          3450 => x"dc",
          3451 => x"8b",
          3452 => x"2e",
          3453 => x"b3",
          3454 => x"14",
          3455 => x"3f",
          3456 => x"08",
          3457 => x"e4",
          3458 => x"81",
          3459 => x"84",
          3460 => x"d7",
          3461 => x"dc",
          3462 => x"15",
          3463 => x"14",
          3464 => x"3f",
          3465 => x"08",
          3466 => x"76",
          3467 => x"dc",
          3468 => x"05",
          3469 => x"dc",
          3470 => x"86",
          3471 => x"0b",
          3472 => x"80",
          3473 => x"dc",
          3474 => x"3d",
          3475 => x"3d",
          3476 => x"89",
          3477 => x"2e",
          3478 => x"08",
          3479 => x"2e",
          3480 => x"33",
          3481 => x"2e",
          3482 => x"13",
          3483 => x"22",
          3484 => x"76",
          3485 => x"06",
          3486 => x"13",
          3487 => x"c0",
          3488 => x"cc",
          3489 => x"52",
          3490 => x"71",
          3491 => x"55",
          3492 => x"53",
          3493 => x"0c",
          3494 => x"dc",
          3495 => x"3d",
          3496 => x"3d",
          3497 => x"05",
          3498 => x"89",
          3499 => x"52",
          3500 => x"3f",
          3501 => x"0b",
          3502 => x"08",
          3503 => x"81",
          3504 => x"84",
          3505 => x"e8",
          3506 => x"55",
          3507 => x"2e",
          3508 => x"74",
          3509 => x"73",
          3510 => x"38",
          3511 => x"78",
          3512 => x"54",
          3513 => x"92",
          3514 => x"89",
          3515 => x"84",
          3516 => x"b0",
          3517 => x"cc",
          3518 => x"81",
          3519 => x"88",
          3520 => x"eb",
          3521 => x"02",
          3522 => x"e7",
          3523 => x"59",
          3524 => x"80",
          3525 => x"38",
          3526 => x"70",
          3527 => x"d0",
          3528 => x"3d",
          3529 => x"58",
          3530 => x"81",
          3531 => x"55",
          3532 => x"08",
          3533 => x"7a",
          3534 => x"8c",
          3535 => x"56",
          3536 => x"81",
          3537 => x"55",
          3538 => x"08",
          3539 => x"80",
          3540 => x"70",
          3541 => x"57",
          3542 => x"83",
          3543 => x"77",
          3544 => x"73",
          3545 => x"ab",
          3546 => x"2e",
          3547 => x"84",
          3548 => x"06",
          3549 => x"51",
          3550 => x"81",
          3551 => x"55",
          3552 => x"b2",
          3553 => x"06",
          3554 => x"b8",
          3555 => x"2a",
          3556 => x"51",
          3557 => x"2e",
          3558 => x"55",
          3559 => x"77",
          3560 => x"74",
          3561 => x"77",
          3562 => x"81",
          3563 => x"73",
          3564 => x"af",
          3565 => x"7a",
          3566 => x"3f",
          3567 => x"08",
          3568 => x"b2",
          3569 => x"8e",
          3570 => x"ea",
          3571 => x"a0",
          3572 => x"34",
          3573 => x"52",
          3574 => x"bd",
          3575 => x"62",
          3576 => x"d4",
          3577 => x"54",
          3578 => x"15",
          3579 => x"2e",
          3580 => x"7a",
          3581 => x"51",
          3582 => x"75",
          3583 => x"d4",
          3584 => x"be",
          3585 => x"cc",
          3586 => x"dc",
          3587 => x"ca",
          3588 => x"74",
          3589 => x"02",
          3590 => x"70",
          3591 => x"81",
          3592 => x"56",
          3593 => x"86",
          3594 => x"82",
          3595 => x"81",
          3596 => x"06",
          3597 => x"80",
          3598 => x"75",
          3599 => x"73",
          3600 => x"38",
          3601 => x"92",
          3602 => x"7a",
          3603 => x"3f",
          3604 => x"08",
          3605 => x"8c",
          3606 => x"55",
          3607 => x"08",
          3608 => x"77",
          3609 => x"81",
          3610 => x"73",
          3611 => x"38",
          3612 => x"07",
          3613 => x"11",
          3614 => x"0c",
          3615 => x"0c",
          3616 => x"52",
          3617 => x"3f",
          3618 => x"08",
          3619 => x"08",
          3620 => x"63",
          3621 => x"5a",
          3622 => x"81",
          3623 => x"81",
          3624 => x"8c",
          3625 => x"7a",
          3626 => x"17",
          3627 => x"23",
          3628 => x"34",
          3629 => x"1a",
          3630 => x"9c",
          3631 => x"0b",
          3632 => x"77",
          3633 => x"81",
          3634 => x"73",
          3635 => x"8d",
          3636 => x"cc",
          3637 => x"81",
          3638 => x"dc",
          3639 => x"1a",
          3640 => x"22",
          3641 => x"7b",
          3642 => x"a8",
          3643 => x"78",
          3644 => x"3f",
          3645 => x"08",
          3646 => x"cc",
          3647 => x"83",
          3648 => x"81",
          3649 => x"ff",
          3650 => x"06",
          3651 => x"55",
          3652 => x"56",
          3653 => x"76",
          3654 => x"51",
          3655 => x"27",
          3656 => x"70",
          3657 => x"5a",
          3658 => x"76",
          3659 => x"74",
          3660 => x"83",
          3661 => x"73",
          3662 => x"38",
          3663 => x"51",
          3664 => x"81",
          3665 => x"85",
          3666 => x"8e",
          3667 => x"2a",
          3668 => x"08",
          3669 => x"0c",
          3670 => x"79",
          3671 => x"73",
          3672 => x"0c",
          3673 => x"04",
          3674 => x"60",
          3675 => x"40",
          3676 => x"80",
          3677 => x"3d",
          3678 => x"78",
          3679 => x"3f",
          3680 => x"08",
          3681 => x"cc",
          3682 => x"91",
          3683 => x"74",
          3684 => x"38",
          3685 => x"c4",
          3686 => x"33",
          3687 => x"87",
          3688 => x"2e",
          3689 => x"95",
          3690 => x"91",
          3691 => x"56",
          3692 => x"81",
          3693 => x"34",
          3694 => x"a0",
          3695 => x"08",
          3696 => x"31",
          3697 => x"27",
          3698 => x"5c",
          3699 => x"82",
          3700 => x"19",
          3701 => x"ff",
          3702 => x"74",
          3703 => x"7e",
          3704 => x"ff",
          3705 => x"2a",
          3706 => x"79",
          3707 => x"87",
          3708 => x"08",
          3709 => x"98",
          3710 => x"78",
          3711 => x"3f",
          3712 => x"08",
          3713 => x"27",
          3714 => x"74",
          3715 => x"a3",
          3716 => x"1a",
          3717 => x"08",
          3718 => x"d4",
          3719 => x"dc",
          3720 => x"2e",
          3721 => x"81",
          3722 => x"1a",
          3723 => x"59",
          3724 => x"2e",
          3725 => x"77",
          3726 => x"11",
          3727 => x"55",
          3728 => x"85",
          3729 => x"31",
          3730 => x"76",
          3731 => x"81",
          3732 => x"ca",
          3733 => x"dc",
          3734 => x"d7",
          3735 => x"11",
          3736 => x"74",
          3737 => x"38",
          3738 => x"77",
          3739 => x"78",
          3740 => x"84",
          3741 => x"16",
          3742 => x"08",
          3743 => x"2b",
          3744 => x"cf",
          3745 => x"89",
          3746 => x"39",
          3747 => x"0c",
          3748 => x"83",
          3749 => x"80",
          3750 => x"55",
          3751 => x"83",
          3752 => x"9c",
          3753 => x"7e",
          3754 => x"3f",
          3755 => x"08",
          3756 => x"75",
          3757 => x"08",
          3758 => x"1f",
          3759 => x"7c",
          3760 => x"3f",
          3761 => x"7e",
          3762 => x"0c",
          3763 => x"1b",
          3764 => x"1c",
          3765 => x"fd",
          3766 => x"56",
          3767 => x"cc",
          3768 => x"0d",
          3769 => x"0d",
          3770 => x"64",
          3771 => x"58",
          3772 => x"90",
          3773 => x"52",
          3774 => x"d2",
          3775 => x"cc",
          3776 => x"dc",
          3777 => x"38",
          3778 => x"55",
          3779 => x"86",
          3780 => x"83",
          3781 => x"18",
          3782 => x"2a",
          3783 => x"51",
          3784 => x"56",
          3785 => x"83",
          3786 => x"39",
          3787 => x"19",
          3788 => x"83",
          3789 => x"0b",
          3790 => x"81",
          3791 => x"39",
          3792 => x"7c",
          3793 => x"74",
          3794 => x"38",
          3795 => x"7b",
          3796 => x"ec",
          3797 => x"08",
          3798 => x"06",
          3799 => x"81",
          3800 => x"8a",
          3801 => x"05",
          3802 => x"06",
          3803 => x"bf",
          3804 => x"38",
          3805 => x"55",
          3806 => x"7a",
          3807 => x"98",
          3808 => x"77",
          3809 => x"3f",
          3810 => x"08",
          3811 => x"cc",
          3812 => x"82",
          3813 => x"81",
          3814 => x"38",
          3815 => x"ff",
          3816 => x"98",
          3817 => x"18",
          3818 => x"74",
          3819 => x"7e",
          3820 => x"08",
          3821 => x"2e",
          3822 => x"8d",
          3823 => x"ce",
          3824 => x"dc",
          3825 => x"ee",
          3826 => x"08",
          3827 => x"d1",
          3828 => x"dc",
          3829 => x"2e",
          3830 => x"81",
          3831 => x"1b",
          3832 => x"5a",
          3833 => x"2e",
          3834 => x"78",
          3835 => x"11",
          3836 => x"55",
          3837 => x"85",
          3838 => x"31",
          3839 => x"76",
          3840 => x"81",
          3841 => x"c8",
          3842 => x"dc",
          3843 => x"a6",
          3844 => x"11",
          3845 => x"56",
          3846 => x"27",
          3847 => x"80",
          3848 => x"08",
          3849 => x"2b",
          3850 => x"b4",
          3851 => x"b5",
          3852 => x"80",
          3853 => x"34",
          3854 => x"56",
          3855 => x"8c",
          3856 => x"19",
          3857 => x"38",
          3858 => x"b6",
          3859 => x"cc",
          3860 => x"38",
          3861 => x"12",
          3862 => x"9c",
          3863 => x"18",
          3864 => x"06",
          3865 => x"31",
          3866 => x"76",
          3867 => x"7b",
          3868 => x"08",
          3869 => x"cd",
          3870 => x"dc",
          3871 => x"b6",
          3872 => x"7c",
          3873 => x"08",
          3874 => x"1f",
          3875 => x"cb",
          3876 => x"55",
          3877 => x"16",
          3878 => x"31",
          3879 => x"7f",
          3880 => x"94",
          3881 => x"70",
          3882 => x"8c",
          3883 => x"58",
          3884 => x"76",
          3885 => x"75",
          3886 => x"19",
          3887 => x"39",
          3888 => x"80",
          3889 => x"74",
          3890 => x"80",
          3891 => x"dc",
          3892 => x"3d",
          3893 => x"3d",
          3894 => x"3d",
          3895 => x"70",
          3896 => x"ea",
          3897 => x"cc",
          3898 => x"dc",
          3899 => x"fb",
          3900 => x"33",
          3901 => x"70",
          3902 => x"55",
          3903 => x"2e",
          3904 => x"a0",
          3905 => x"78",
          3906 => x"3f",
          3907 => x"08",
          3908 => x"cc",
          3909 => x"38",
          3910 => x"8b",
          3911 => x"07",
          3912 => x"8b",
          3913 => x"16",
          3914 => x"52",
          3915 => x"dd",
          3916 => x"16",
          3917 => x"15",
          3918 => x"3f",
          3919 => x"0a",
          3920 => x"51",
          3921 => x"76",
          3922 => x"51",
          3923 => x"78",
          3924 => x"83",
          3925 => x"51",
          3926 => x"81",
          3927 => x"90",
          3928 => x"bf",
          3929 => x"73",
          3930 => x"76",
          3931 => x"0c",
          3932 => x"04",
          3933 => x"76",
          3934 => x"fe",
          3935 => x"dc",
          3936 => x"81",
          3937 => x"9c",
          3938 => x"fc",
          3939 => x"51",
          3940 => x"81",
          3941 => x"53",
          3942 => x"08",
          3943 => x"dc",
          3944 => x"0c",
          3945 => x"cc",
          3946 => x"0d",
          3947 => x"0d",
          3948 => x"e6",
          3949 => x"52",
          3950 => x"dc",
          3951 => x"8b",
          3952 => x"cc",
          3953 => x"fc",
          3954 => x"71",
          3955 => x"0c",
          3956 => x"04",
          3957 => x"80",
          3958 => x"d0",
          3959 => x"3d",
          3960 => x"3f",
          3961 => x"08",
          3962 => x"cc",
          3963 => x"38",
          3964 => x"52",
          3965 => x"05",
          3966 => x"3f",
          3967 => x"08",
          3968 => x"cc",
          3969 => x"02",
          3970 => x"33",
          3971 => x"55",
          3972 => x"25",
          3973 => x"7a",
          3974 => x"54",
          3975 => x"a2",
          3976 => x"84",
          3977 => x"06",
          3978 => x"73",
          3979 => x"38",
          3980 => x"70",
          3981 => x"a8",
          3982 => x"cc",
          3983 => x"0c",
          3984 => x"dc",
          3985 => x"2e",
          3986 => x"83",
          3987 => x"74",
          3988 => x"0c",
          3989 => x"04",
          3990 => x"6f",
          3991 => x"80",
          3992 => x"53",
          3993 => x"b8",
          3994 => x"3d",
          3995 => x"3f",
          3996 => x"08",
          3997 => x"cc",
          3998 => x"38",
          3999 => x"7c",
          4000 => x"47",
          4001 => x"54",
          4002 => x"81",
          4003 => x"52",
          4004 => x"52",
          4005 => x"3f",
          4006 => x"08",
          4007 => x"cc",
          4008 => x"38",
          4009 => x"51",
          4010 => x"81",
          4011 => x"57",
          4012 => x"08",
          4013 => x"69",
          4014 => x"da",
          4015 => x"dc",
          4016 => x"76",
          4017 => x"d5",
          4018 => x"dc",
          4019 => x"81",
          4020 => x"82",
          4021 => x"52",
          4022 => x"eb",
          4023 => x"cc",
          4024 => x"dc",
          4025 => x"38",
          4026 => x"51",
          4027 => x"73",
          4028 => x"08",
          4029 => x"76",
          4030 => x"d6",
          4031 => x"dc",
          4032 => x"81",
          4033 => x"80",
          4034 => x"76",
          4035 => x"81",
          4036 => x"82",
          4037 => x"39",
          4038 => x"38",
          4039 => x"bc",
          4040 => x"51",
          4041 => x"76",
          4042 => x"11",
          4043 => x"51",
          4044 => x"73",
          4045 => x"38",
          4046 => x"55",
          4047 => x"16",
          4048 => x"56",
          4049 => x"38",
          4050 => x"73",
          4051 => x"90",
          4052 => x"2e",
          4053 => x"16",
          4054 => x"ff",
          4055 => x"ff",
          4056 => x"58",
          4057 => x"74",
          4058 => x"75",
          4059 => x"18",
          4060 => x"58",
          4061 => x"fe",
          4062 => x"7b",
          4063 => x"06",
          4064 => x"18",
          4065 => x"58",
          4066 => x"80",
          4067 => x"fc",
          4068 => x"29",
          4069 => x"05",
          4070 => x"33",
          4071 => x"56",
          4072 => x"2e",
          4073 => x"16",
          4074 => x"33",
          4075 => x"73",
          4076 => x"16",
          4077 => x"26",
          4078 => x"55",
          4079 => x"91",
          4080 => x"54",
          4081 => x"70",
          4082 => x"34",
          4083 => x"ec",
          4084 => x"70",
          4085 => x"34",
          4086 => x"09",
          4087 => x"38",
          4088 => x"39",
          4089 => x"19",
          4090 => x"33",
          4091 => x"05",
          4092 => x"78",
          4093 => x"80",
          4094 => x"81",
          4095 => x"9e",
          4096 => x"f7",
          4097 => x"7d",
          4098 => x"05",
          4099 => x"57",
          4100 => x"3f",
          4101 => x"08",
          4102 => x"cc",
          4103 => x"38",
          4104 => x"53",
          4105 => x"38",
          4106 => x"54",
          4107 => x"92",
          4108 => x"33",
          4109 => x"70",
          4110 => x"54",
          4111 => x"38",
          4112 => x"15",
          4113 => x"70",
          4114 => x"58",
          4115 => x"82",
          4116 => x"8a",
          4117 => x"89",
          4118 => x"53",
          4119 => x"b7",
          4120 => x"ff",
          4121 => x"96",
          4122 => x"dc",
          4123 => x"15",
          4124 => x"53",
          4125 => x"96",
          4126 => x"dc",
          4127 => x"26",
          4128 => x"30",
          4129 => x"70",
          4130 => x"77",
          4131 => x"18",
          4132 => x"51",
          4133 => x"88",
          4134 => x"73",
          4135 => x"52",
          4136 => x"ca",
          4137 => x"cc",
          4138 => x"dc",
          4139 => x"2e",
          4140 => x"81",
          4141 => x"ff",
          4142 => x"38",
          4143 => x"08",
          4144 => x"73",
          4145 => x"73",
          4146 => x"9c",
          4147 => x"27",
          4148 => x"75",
          4149 => x"16",
          4150 => x"17",
          4151 => x"33",
          4152 => x"70",
          4153 => x"55",
          4154 => x"80",
          4155 => x"73",
          4156 => x"cc",
          4157 => x"dc",
          4158 => x"81",
          4159 => x"94",
          4160 => x"cc",
          4161 => x"39",
          4162 => x"51",
          4163 => x"81",
          4164 => x"54",
          4165 => x"be",
          4166 => x"27",
          4167 => x"53",
          4168 => x"08",
          4169 => x"73",
          4170 => x"ff",
          4171 => x"15",
          4172 => x"16",
          4173 => x"ff",
          4174 => x"80",
          4175 => x"73",
          4176 => x"c6",
          4177 => x"dc",
          4178 => x"38",
          4179 => x"16",
          4180 => x"80",
          4181 => x"0b",
          4182 => x"81",
          4183 => x"75",
          4184 => x"dc",
          4185 => x"58",
          4186 => x"54",
          4187 => x"74",
          4188 => x"73",
          4189 => x"90",
          4190 => x"c0",
          4191 => x"90",
          4192 => x"83",
          4193 => x"72",
          4194 => x"38",
          4195 => x"08",
          4196 => x"77",
          4197 => x"80",
          4198 => x"dc",
          4199 => x"3d",
          4200 => x"3d",
          4201 => x"89",
          4202 => x"2e",
          4203 => x"80",
          4204 => x"fc",
          4205 => x"3d",
          4206 => x"e1",
          4207 => x"dc",
          4208 => x"81",
          4209 => x"80",
          4210 => x"76",
          4211 => x"75",
          4212 => x"3f",
          4213 => x"08",
          4214 => x"cc",
          4215 => x"38",
          4216 => x"70",
          4217 => x"57",
          4218 => x"a2",
          4219 => x"33",
          4220 => x"70",
          4221 => x"55",
          4222 => x"2e",
          4223 => x"16",
          4224 => x"51",
          4225 => x"81",
          4226 => x"88",
          4227 => x"54",
          4228 => x"84",
          4229 => x"52",
          4230 => x"e5",
          4231 => x"cc",
          4232 => x"84",
          4233 => x"06",
          4234 => x"55",
          4235 => x"80",
          4236 => x"80",
          4237 => x"54",
          4238 => x"cc",
          4239 => x"0d",
          4240 => x"0d",
          4241 => x"fc",
          4242 => x"52",
          4243 => x"3f",
          4244 => x"08",
          4245 => x"dc",
          4246 => x"0c",
          4247 => x"04",
          4248 => x"77",
          4249 => x"fc",
          4250 => x"53",
          4251 => x"de",
          4252 => x"cc",
          4253 => x"dc",
          4254 => x"df",
          4255 => x"38",
          4256 => x"08",
          4257 => x"cd",
          4258 => x"dc",
          4259 => x"80",
          4260 => x"dc",
          4261 => x"73",
          4262 => x"3f",
          4263 => x"08",
          4264 => x"cc",
          4265 => x"09",
          4266 => x"38",
          4267 => x"39",
          4268 => x"08",
          4269 => x"52",
          4270 => x"b3",
          4271 => x"73",
          4272 => x"3f",
          4273 => x"08",
          4274 => x"30",
          4275 => x"9f",
          4276 => x"dc",
          4277 => x"51",
          4278 => x"72",
          4279 => x"0c",
          4280 => x"04",
          4281 => x"65",
          4282 => x"89",
          4283 => x"96",
          4284 => x"df",
          4285 => x"dc",
          4286 => x"81",
          4287 => x"b2",
          4288 => x"75",
          4289 => x"3f",
          4290 => x"08",
          4291 => x"cc",
          4292 => x"02",
          4293 => x"33",
          4294 => x"55",
          4295 => x"25",
          4296 => x"55",
          4297 => x"80",
          4298 => x"76",
          4299 => x"d4",
          4300 => x"81",
          4301 => x"94",
          4302 => x"f0",
          4303 => x"65",
          4304 => x"53",
          4305 => x"05",
          4306 => x"51",
          4307 => x"81",
          4308 => x"5b",
          4309 => x"08",
          4310 => x"7c",
          4311 => x"08",
          4312 => x"fe",
          4313 => x"08",
          4314 => x"55",
          4315 => x"91",
          4316 => x"0c",
          4317 => x"81",
          4318 => x"39",
          4319 => x"c7",
          4320 => x"cc",
          4321 => x"55",
          4322 => x"2e",
          4323 => x"bf",
          4324 => x"5f",
          4325 => x"92",
          4326 => x"51",
          4327 => x"81",
          4328 => x"ff",
          4329 => x"81",
          4330 => x"81",
          4331 => x"81",
          4332 => x"30",
          4333 => x"cc",
          4334 => x"25",
          4335 => x"19",
          4336 => x"5a",
          4337 => x"08",
          4338 => x"38",
          4339 => x"a4",
          4340 => x"dc",
          4341 => x"58",
          4342 => x"77",
          4343 => x"7d",
          4344 => x"bf",
          4345 => x"dc",
          4346 => x"81",
          4347 => x"80",
          4348 => x"70",
          4349 => x"ff",
          4350 => x"56",
          4351 => x"2e",
          4352 => x"9e",
          4353 => x"51",
          4354 => x"3f",
          4355 => x"08",
          4356 => x"06",
          4357 => x"80",
          4358 => x"19",
          4359 => x"54",
          4360 => x"14",
          4361 => x"c5",
          4362 => x"cc",
          4363 => x"06",
          4364 => x"80",
          4365 => x"19",
          4366 => x"54",
          4367 => x"06",
          4368 => x"79",
          4369 => x"78",
          4370 => x"79",
          4371 => x"84",
          4372 => x"07",
          4373 => x"84",
          4374 => x"81",
          4375 => x"92",
          4376 => x"f9",
          4377 => x"8a",
          4378 => x"53",
          4379 => x"e3",
          4380 => x"dc",
          4381 => x"81",
          4382 => x"81",
          4383 => x"17",
          4384 => x"81",
          4385 => x"17",
          4386 => x"2a",
          4387 => x"51",
          4388 => x"55",
          4389 => x"81",
          4390 => x"17",
          4391 => x"8c",
          4392 => x"81",
          4393 => x"9b",
          4394 => x"cc",
          4395 => x"17",
          4396 => x"51",
          4397 => x"81",
          4398 => x"74",
          4399 => x"56",
          4400 => x"98",
          4401 => x"76",
          4402 => x"c6",
          4403 => x"cc",
          4404 => x"09",
          4405 => x"38",
          4406 => x"dc",
          4407 => x"2e",
          4408 => x"85",
          4409 => x"a3",
          4410 => x"38",
          4411 => x"dc",
          4412 => x"15",
          4413 => x"38",
          4414 => x"53",
          4415 => x"08",
          4416 => x"c3",
          4417 => x"dc",
          4418 => x"94",
          4419 => x"18",
          4420 => x"33",
          4421 => x"54",
          4422 => x"34",
          4423 => x"85",
          4424 => x"18",
          4425 => x"74",
          4426 => x"0c",
          4427 => x"04",
          4428 => x"82",
          4429 => x"ff",
          4430 => x"a1",
          4431 => x"e4",
          4432 => x"cc",
          4433 => x"dc",
          4434 => x"f5",
          4435 => x"a1",
          4436 => x"95",
          4437 => x"58",
          4438 => x"81",
          4439 => x"55",
          4440 => x"08",
          4441 => x"02",
          4442 => x"33",
          4443 => x"70",
          4444 => x"55",
          4445 => x"73",
          4446 => x"75",
          4447 => x"80",
          4448 => x"bd",
          4449 => x"d6",
          4450 => x"81",
          4451 => x"87",
          4452 => x"ad",
          4453 => x"78",
          4454 => x"3f",
          4455 => x"08",
          4456 => x"70",
          4457 => x"55",
          4458 => x"2e",
          4459 => x"78",
          4460 => x"cc",
          4461 => x"08",
          4462 => x"38",
          4463 => x"dc",
          4464 => x"76",
          4465 => x"70",
          4466 => x"b5",
          4467 => x"cc",
          4468 => x"dc",
          4469 => x"e9",
          4470 => x"cc",
          4471 => x"51",
          4472 => x"81",
          4473 => x"55",
          4474 => x"08",
          4475 => x"55",
          4476 => x"81",
          4477 => x"84",
          4478 => x"81",
          4479 => x"80",
          4480 => x"51",
          4481 => x"81",
          4482 => x"81",
          4483 => x"30",
          4484 => x"cc",
          4485 => x"25",
          4486 => x"75",
          4487 => x"38",
          4488 => x"8f",
          4489 => x"75",
          4490 => x"c1",
          4491 => x"dc",
          4492 => x"74",
          4493 => x"51",
          4494 => x"3f",
          4495 => x"08",
          4496 => x"dc",
          4497 => x"3d",
          4498 => x"3d",
          4499 => x"99",
          4500 => x"52",
          4501 => x"d8",
          4502 => x"dc",
          4503 => x"81",
          4504 => x"82",
          4505 => x"5e",
          4506 => x"3d",
          4507 => x"cf",
          4508 => x"dc",
          4509 => x"81",
          4510 => x"86",
          4511 => x"82",
          4512 => x"dc",
          4513 => x"2e",
          4514 => x"82",
          4515 => x"80",
          4516 => x"70",
          4517 => x"06",
          4518 => x"54",
          4519 => x"38",
          4520 => x"52",
          4521 => x"52",
          4522 => x"3f",
          4523 => x"08",
          4524 => x"81",
          4525 => x"83",
          4526 => x"81",
          4527 => x"81",
          4528 => x"06",
          4529 => x"54",
          4530 => x"08",
          4531 => x"81",
          4532 => x"81",
          4533 => x"39",
          4534 => x"38",
          4535 => x"08",
          4536 => x"c4",
          4537 => x"dc",
          4538 => x"81",
          4539 => x"81",
          4540 => x"53",
          4541 => x"19",
          4542 => x"8c",
          4543 => x"ae",
          4544 => x"34",
          4545 => x"0b",
          4546 => x"82",
          4547 => x"52",
          4548 => x"51",
          4549 => x"3f",
          4550 => x"b4",
          4551 => x"c9",
          4552 => x"53",
          4553 => x"53",
          4554 => x"51",
          4555 => x"3f",
          4556 => x"0b",
          4557 => x"34",
          4558 => x"80",
          4559 => x"51",
          4560 => x"78",
          4561 => x"83",
          4562 => x"51",
          4563 => x"81",
          4564 => x"54",
          4565 => x"08",
          4566 => x"88",
          4567 => x"64",
          4568 => x"ff",
          4569 => x"75",
          4570 => x"78",
          4571 => x"3f",
          4572 => x"0b",
          4573 => x"78",
          4574 => x"83",
          4575 => x"51",
          4576 => x"3f",
          4577 => x"08",
          4578 => x"80",
          4579 => x"76",
          4580 => x"ae",
          4581 => x"dc",
          4582 => x"3d",
          4583 => x"3d",
          4584 => x"84",
          4585 => x"f1",
          4586 => x"a8",
          4587 => x"05",
          4588 => x"51",
          4589 => x"81",
          4590 => x"55",
          4591 => x"08",
          4592 => x"78",
          4593 => x"08",
          4594 => x"70",
          4595 => x"b8",
          4596 => x"cc",
          4597 => x"dc",
          4598 => x"b9",
          4599 => x"9b",
          4600 => x"a0",
          4601 => x"55",
          4602 => x"38",
          4603 => x"3d",
          4604 => x"3d",
          4605 => x"51",
          4606 => x"3f",
          4607 => x"52",
          4608 => x"52",
          4609 => x"dd",
          4610 => x"08",
          4611 => x"cb",
          4612 => x"dc",
          4613 => x"81",
          4614 => x"95",
          4615 => x"2e",
          4616 => x"88",
          4617 => x"3d",
          4618 => x"38",
          4619 => x"e5",
          4620 => x"cc",
          4621 => x"09",
          4622 => x"b8",
          4623 => x"c9",
          4624 => x"dc",
          4625 => x"81",
          4626 => x"81",
          4627 => x"56",
          4628 => x"3d",
          4629 => x"52",
          4630 => x"ff",
          4631 => x"02",
          4632 => x"8b",
          4633 => x"16",
          4634 => x"2a",
          4635 => x"51",
          4636 => x"89",
          4637 => x"07",
          4638 => x"17",
          4639 => x"81",
          4640 => x"34",
          4641 => x"70",
          4642 => x"81",
          4643 => x"55",
          4644 => x"80",
          4645 => x"64",
          4646 => x"38",
          4647 => x"51",
          4648 => x"81",
          4649 => x"52",
          4650 => x"b7",
          4651 => x"55",
          4652 => x"08",
          4653 => x"dd",
          4654 => x"cc",
          4655 => x"51",
          4656 => x"3f",
          4657 => x"08",
          4658 => x"11",
          4659 => x"81",
          4660 => x"80",
          4661 => x"16",
          4662 => x"ae",
          4663 => x"06",
          4664 => x"53",
          4665 => x"51",
          4666 => x"78",
          4667 => x"83",
          4668 => x"39",
          4669 => x"08",
          4670 => x"51",
          4671 => x"81",
          4672 => x"55",
          4673 => x"08",
          4674 => x"51",
          4675 => x"3f",
          4676 => x"08",
          4677 => x"dc",
          4678 => x"3d",
          4679 => x"3d",
          4680 => x"db",
          4681 => x"84",
          4682 => x"05",
          4683 => x"82",
          4684 => x"d0",
          4685 => x"3d",
          4686 => x"3f",
          4687 => x"08",
          4688 => x"cc",
          4689 => x"38",
          4690 => x"52",
          4691 => x"05",
          4692 => x"3f",
          4693 => x"08",
          4694 => x"cc",
          4695 => x"02",
          4696 => x"33",
          4697 => x"54",
          4698 => x"aa",
          4699 => x"06",
          4700 => x"8b",
          4701 => x"06",
          4702 => x"07",
          4703 => x"56",
          4704 => x"34",
          4705 => x"0b",
          4706 => x"78",
          4707 => x"a9",
          4708 => x"cc",
          4709 => x"81",
          4710 => x"95",
          4711 => x"ef",
          4712 => x"56",
          4713 => x"3d",
          4714 => x"94",
          4715 => x"f4",
          4716 => x"cc",
          4717 => x"dc",
          4718 => x"cb",
          4719 => x"63",
          4720 => x"d4",
          4721 => x"c0",
          4722 => x"cc",
          4723 => x"dc",
          4724 => x"38",
          4725 => x"05",
          4726 => x"06",
          4727 => x"73",
          4728 => x"16",
          4729 => x"22",
          4730 => x"07",
          4731 => x"1f",
          4732 => x"c2",
          4733 => x"81",
          4734 => x"34",
          4735 => x"b3",
          4736 => x"dc",
          4737 => x"74",
          4738 => x"0c",
          4739 => x"04",
          4740 => x"69",
          4741 => x"80",
          4742 => x"d0",
          4743 => x"3d",
          4744 => x"3f",
          4745 => x"08",
          4746 => x"08",
          4747 => x"dc",
          4748 => x"80",
          4749 => x"57",
          4750 => x"81",
          4751 => x"70",
          4752 => x"55",
          4753 => x"80",
          4754 => x"5d",
          4755 => x"52",
          4756 => x"52",
          4757 => x"a9",
          4758 => x"cc",
          4759 => x"dc",
          4760 => x"d1",
          4761 => x"73",
          4762 => x"3f",
          4763 => x"08",
          4764 => x"cc",
          4765 => x"81",
          4766 => x"81",
          4767 => x"65",
          4768 => x"78",
          4769 => x"7b",
          4770 => x"55",
          4771 => x"34",
          4772 => x"8a",
          4773 => x"38",
          4774 => x"1a",
          4775 => x"34",
          4776 => x"9e",
          4777 => x"70",
          4778 => x"51",
          4779 => x"a0",
          4780 => x"8e",
          4781 => x"2e",
          4782 => x"86",
          4783 => x"34",
          4784 => x"30",
          4785 => x"80",
          4786 => x"7a",
          4787 => x"c1",
          4788 => x"2e",
          4789 => x"a0",
          4790 => x"51",
          4791 => x"3f",
          4792 => x"08",
          4793 => x"cc",
          4794 => x"7b",
          4795 => x"55",
          4796 => x"73",
          4797 => x"38",
          4798 => x"73",
          4799 => x"38",
          4800 => x"15",
          4801 => x"ff",
          4802 => x"81",
          4803 => x"7b",
          4804 => x"dc",
          4805 => x"3d",
          4806 => x"3d",
          4807 => x"9c",
          4808 => x"05",
          4809 => x"51",
          4810 => x"81",
          4811 => x"81",
          4812 => x"56",
          4813 => x"cc",
          4814 => x"38",
          4815 => x"52",
          4816 => x"52",
          4817 => x"c0",
          4818 => x"70",
          4819 => x"ff",
          4820 => x"55",
          4821 => x"27",
          4822 => x"78",
          4823 => x"ff",
          4824 => x"05",
          4825 => x"55",
          4826 => x"3f",
          4827 => x"08",
          4828 => x"38",
          4829 => x"70",
          4830 => x"ff",
          4831 => x"81",
          4832 => x"80",
          4833 => x"74",
          4834 => x"07",
          4835 => x"4e",
          4836 => x"81",
          4837 => x"55",
          4838 => x"70",
          4839 => x"06",
          4840 => x"99",
          4841 => x"e0",
          4842 => x"ff",
          4843 => x"54",
          4844 => x"27",
          4845 => x"cb",
          4846 => x"55",
          4847 => x"a3",
          4848 => x"81",
          4849 => x"ff",
          4850 => x"81",
          4851 => x"93",
          4852 => x"75",
          4853 => x"76",
          4854 => x"38",
          4855 => x"77",
          4856 => x"86",
          4857 => x"39",
          4858 => x"27",
          4859 => x"88",
          4860 => x"78",
          4861 => x"5a",
          4862 => x"57",
          4863 => x"81",
          4864 => x"81",
          4865 => x"33",
          4866 => x"06",
          4867 => x"57",
          4868 => x"fe",
          4869 => x"3d",
          4870 => x"55",
          4871 => x"2e",
          4872 => x"76",
          4873 => x"38",
          4874 => x"55",
          4875 => x"33",
          4876 => x"a0",
          4877 => x"06",
          4878 => x"17",
          4879 => x"38",
          4880 => x"43",
          4881 => x"3d",
          4882 => x"ff",
          4883 => x"81",
          4884 => x"54",
          4885 => x"08",
          4886 => x"81",
          4887 => x"ff",
          4888 => x"81",
          4889 => x"54",
          4890 => x"08",
          4891 => x"80",
          4892 => x"54",
          4893 => x"80",
          4894 => x"dc",
          4895 => x"2e",
          4896 => x"80",
          4897 => x"54",
          4898 => x"80",
          4899 => x"52",
          4900 => x"bd",
          4901 => x"dc",
          4902 => x"81",
          4903 => x"b1",
          4904 => x"81",
          4905 => x"52",
          4906 => x"ab",
          4907 => x"54",
          4908 => x"15",
          4909 => x"78",
          4910 => x"ff",
          4911 => x"79",
          4912 => x"83",
          4913 => x"51",
          4914 => x"3f",
          4915 => x"08",
          4916 => x"74",
          4917 => x"0c",
          4918 => x"04",
          4919 => x"60",
          4920 => x"05",
          4921 => x"33",
          4922 => x"05",
          4923 => x"40",
          4924 => x"da",
          4925 => x"cc",
          4926 => x"dc",
          4927 => x"bd",
          4928 => x"33",
          4929 => x"b5",
          4930 => x"2e",
          4931 => x"1a",
          4932 => x"90",
          4933 => x"33",
          4934 => x"70",
          4935 => x"55",
          4936 => x"38",
          4937 => x"97",
          4938 => x"82",
          4939 => x"58",
          4940 => x"7e",
          4941 => x"70",
          4942 => x"55",
          4943 => x"56",
          4944 => x"b8",
          4945 => x"7d",
          4946 => x"70",
          4947 => x"2a",
          4948 => x"08",
          4949 => x"08",
          4950 => x"5d",
          4951 => x"77",
          4952 => x"98",
          4953 => x"26",
          4954 => x"57",
          4955 => x"59",
          4956 => x"52",
          4957 => x"ae",
          4958 => x"15",
          4959 => x"98",
          4960 => x"26",
          4961 => x"55",
          4962 => x"08",
          4963 => x"99",
          4964 => x"cc",
          4965 => x"ff",
          4966 => x"dc",
          4967 => x"38",
          4968 => x"75",
          4969 => x"81",
          4970 => x"93",
          4971 => x"80",
          4972 => x"2e",
          4973 => x"ff",
          4974 => x"58",
          4975 => x"7d",
          4976 => x"38",
          4977 => x"55",
          4978 => x"b4",
          4979 => x"56",
          4980 => x"09",
          4981 => x"38",
          4982 => x"53",
          4983 => x"51",
          4984 => x"3f",
          4985 => x"08",
          4986 => x"cc",
          4987 => x"38",
          4988 => x"ff",
          4989 => x"5c",
          4990 => x"84",
          4991 => x"5c",
          4992 => x"12",
          4993 => x"80",
          4994 => x"78",
          4995 => x"7c",
          4996 => x"90",
          4997 => x"c0",
          4998 => x"90",
          4999 => x"15",
          5000 => x"90",
          5001 => x"54",
          5002 => x"91",
          5003 => x"31",
          5004 => x"84",
          5005 => x"07",
          5006 => x"16",
          5007 => x"73",
          5008 => x"0c",
          5009 => x"04",
          5010 => x"6b",
          5011 => x"05",
          5012 => x"33",
          5013 => x"5a",
          5014 => x"bd",
          5015 => x"80",
          5016 => x"cc",
          5017 => x"f8",
          5018 => x"cc",
          5019 => x"81",
          5020 => x"70",
          5021 => x"74",
          5022 => x"38",
          5023 => x"81",
          5024 => x"81",
          5025 => x"81",
          5026 => x"ff",
          5027 => x"81",
          5028 => x"81",
          5029 => x"81",
          5030 => x"83",
          5031 => x"c0",
          5032 => x"2a",
          5033 => x"51",
          5034 => x"74",
          5035 => x"99",
          5036 => x"53",
          5037 => x"51",
          5038 => x"3f",
          5039 => x"08",
          5040 => x"55",
          5041 => x"92",
          5042 => x"80",
          5043 => x"38",
          5044 => x"06",
          5045 => x"2e",
          5046 => x"48",
          5047 => x"87",
          5048 => x"79",
          5049 => x"78",
          5050 => x"26",
          5051 => x"19",
          5052 => x"74",
          5053 => x"38",
          5054 => x"e4",
          5055 => x"2a",
          5056 => x"70",
          5057 => x"59",
          5058 => x"7a",
          5059 => x"56",
          5060 => x"80",
          5061 => x"51",
          5062 => x"74",
          5063 => x"99",
          5064 => x"53",
          5065 => x"51",
          5066 => x"3f",
          5067 => x"dc",
          5068 => x"ac",
          5069 => x"2a",
          5070 => x"81",
          5071 => x"43",
          5072 => x"83",
          5073 => x"66",
          5074 => x"60",
          5075 => x"90",
          5076 => x"31",
          5077 => x"80",
          5078 => x"8a",
          5079 => x"56",
          5080 => x"26",
          5081 => x"77",
          5082 => x"81",
          5083 => x"74",
          5084 => x"38",
          5085 => x"55",
          5086 => x"83",
          5087 => x"81",
          5088 => x"80",
          5089 => x"38",
          5090 => x"55",
          5091 => x"5e",
          5092 => x"89",
          5093 => x"5a",
          5094 => x"09",
          5095 => x"e1",
          5096 => x"38",
          5097 => x"57",
          5098 => x"cd",
          5099 => x"5a",
          5100 => x"9d",
          5101 => x"26",
          5102 => x"cd",
          5103 => x"10",
          5104 => x"22",
          5105 => x"74",
          5106 => x"38",
          5107 => x"ee",
          5108 => x"66",
          5109 => x"a4",
          5110 => x"cc",
          5111 => x"84",
          5112 => x"89",
          5113 => x"a0",
          5114 => x"81",
          5115 => x"fc",
          5116 => x"56",
          5117 => x"f0",
          5118 => x"80",
          5119 => x"d3",
          5120 => x"38",
          5121 => x"57",
          5122 => x"cd",
          5123 => x"5a",
          5124 => x"9d",
          5125 => x"26",
          5126 => x"cd",
          5127 => x"10",
          5128 => x"22",
          5129 => x"74",
          5130 => x"38",
          5131 => x"ee",
          5132 => x"66",
          5133 => x"c4",
          5134 => x"cc",
          5135 => x"05",
          5136 => x"cc",
          5137 => x"26",
          5138 => x"0b",
          5139 => x"08",
          5140 => x"cc",
          5141 => x"11",
          5142 => x"05",
          5143 => x"83",
          5144 => x"2a",
          5145 => x"a0",
          5146 => x"7d",
          5147 => x"69",
          5148 => x"05",
          5149 => x"72",
          5150 => x"5c",
          5151 => x"59",
          5152 => x"2e",
          5153 => x"89",
          5154 => x"60",
          5155 => x"84",
          5156 => x"5d",
          5157 => x"18",
          5158 => x"68",
          5159 => x"74",
          5160 => x"af",
          5161 => x"31",
          5162 => x"53",
          5163 => x"52",
          5164 => x"c8",
          5165 => x"cc",
          5166 => x"83",
          5167 => x"06",
          5168 => x"dc",
          5169 => x"ff",
          5170 => x"dd",
          5171 => x"83",
          5172 => x"2a",
          5173 => x"be",
          5174 => x"39",
          5175 => x"09",
          5176 => x"c5",
          5177 => x"f5",
          5178 => x"cc",
          5179 => x"38",
          5180 => x"79",
          5181 => x"80",
          5182 => x"38",
          5183 => x"96",
          5184 => x"06",
          5185 => x"2e",
          5186 => x"5e",
          5187 => x"81",
          5188 => x"9f",
          5189 => x"38",
          5190 => x"38",
          5191 => x"81",
          5192 => x"fc",
          5193 => x"ab",
          5194 => x"7d",
          5195 => x"81",
          5196 => x"7d",
          5197 => x"78",
          5198 => x"74",
          5199 => x"8e",
          5200 => x"9c",
          5201 => x"53",
          5202 => x"51",
          5203 => x"3f",
          5204 => x"cb",
          5205 => x"51",
          5206 => x"3f",
          5207 => x"8b",
          5208 => x"a1",
          5209 => x"8d",
          5210 => x"83",
          5211 => x"52",
          5212 => x"ff",
          5213 => x"81",
          5214 => x"34",
          5215 => x"70",
          5216 => x"2a",
          5217 => x"54",
          5218 => x"1b",
          5219 => x"88",
          5220 => x"74",
          5221 => x"26",
          5222 => x"83",
          5223 => x"52",
          5224 => x"ff",
          5225 => x"8a",
          5226 => x"a0",
          5227 => x"a1",
          5228 => x"0b",
          5229 => x"bf",
          5230 => x"51",
          5231 => x"3f",
          5232 => x"9a",
          5233 => x"a0",
          5234 => x"52",
          5235 => x"ff",
          5236 => x"7d",
          5237 => x"81",
          5238 => x"38",
          5239 => x"0a",
          5240 => x"1b",
          5241 => x"ce",
          5242 => x"a4",
          5243 => x"a0",
          5244 => x"52",
          5245 => x"ff",
          5246 => x"81",
          5247 => x"51",
          5248 => x"3f",
          5249 => x"1b",
          5250 => x"8c",
          5251 => x"0b",
          5252 => x"34",
          5253 => x"c2",
          5254 => x"53",
          5255 => x"52",
          5256 => x"51",
          5257 => x"88",
          5258 => x"a7",
          5259 => x"a0",
          5260 => x"83",
          5261 => x"52",
          5262 => x"ff",
          5263 => x"ff",
          5264 => x"1c",
          5265 => x"a6",
          5266 => x"53",
          5267 => x"52",
          5268 => x"ff",
          5269 => x"82",
          5270 => x"83",
          5271 => x"52",
          5272 => x"b4",
          5273 => x"60",
          5274 => x"7e",
          5275 => x"d7",
          5276 => x"81",
          5277 => x"83",
          5278 => x"83",
          5279 => x"06",
          5280 => x"75",
          5281 => x"05",
          5282 => x"7e",
          5283 => x"b7",
          5284 => x"53",
          5285 => x"51",
          5286 => x"3f",
          5287 => x"a4",
          5288 => x"51",
          5289 => x"3f",
          5290 => x"e4",
          5291 => x"e4",
          5292 => x"9f",
          5293 => x"18",
          5294 => x"1b",
          5295 => x"f6",
          5296 => x"83",
          5297 => x"ff",
          5298 => x"82",
          5299 => x"78",
          5300 => x"c4",
          5301 => x"60",
          5302 => x"7a",
          5303 => x"ff",
          5304 => x"75",
          5305 => x"53",
          5306 => x"51",
          5307 => x"3f",
          5308 => x"52",
          5309 => x"9f",
          5310 => x"56",
          5311 => x"83",
          5312 => x"06",
          5313 => x"52",
          5314 => x"9e",
          5315 => x"52",
          5316 => x"ff",
          5317 => x"f0",
          5318 => x"1b",
          5319 => x"87",
          5320 => x"55",
          5321 => x"83",
          5322 => x"74",
          5323 => x"ff",
          5324 => x"7c",
          5325 => x"74",
          5326 => x"38",
          5327 => x"54",
          5328 => x"52",
          5329 => x"99",
          5330 => x"dc",
          5331 => x"87",
          5332 => x"53",
          5333 => x"08",
          5334 => x"ff",
          5335 => x"76",
          5336 => x"31",
          5337 => x"cd",
          5338 => x"58",
          5339 => x"ff",
          5340 => x"55",
          5341 => x"83",
          5342 => x"61",
          5343 => x"26",
          5344 => x"57",
          5345 => x"53",
          5346 => x"51",
          5347 => x"3f",
          5348 => x"08",
          5349 => x"76",
          5350 => x"31",
          5351 => x"db",
          5352 => x"7d",
          5353 => x"38",
          5354 => x"83",
          5355 => x"8a",
          5356 => x"7d",
          5357 => x"38",
          5358 => x"81",
          5359 => x"80",
          5360 => x"80",
          5361 => x"7a",
          5362 => x"bc",
          5363 => x"d5",
          5364 => x"ff",
          5365 => x"83",
          5366 => x"77",
          5367 => x"0b",
          5368 => x"81",
          5369 => x"34",
          5370 => x"34",
          5371 => x"34",
          5372 => x"56",
          5373 => x"52",
          5374 => x"ee",
          5375 => x"0b",
          5376 => x"81",
          5377 => x"82",
          5378 => x"56",
          5379 => x"34",
          5380 => x"08",
          5381 => x"60",
          5382 => x"1b",
          5383 => x"96",
          5384 => x"83",
          5385 => x"ff",
          5386 => x"81",
          5387 => x"7a",
          5388 => x"ff",
          5389 => x"81",
          5390 => x"cc",
          5391 => x"80",
          5392 => x"7e",
          5393 => x"e3",
          5394 => x"81",
          5395 => x"90",
          5396 => x"8e",
          5397 => x"81",
          5398 => x"81",
          5399 => x"56",
          5400 => x"cc",
          5401 => x"0d",
          5402 => x"0d",
          5403 => x"59",
          5404 => x"ff",
          5405 => x"57",
          5406 => x"b4",
          5407 => x"f8",
          5408 => x"81",
          5409 => x"52",
          5410 => x"dc",
          5411 => x"2e",
          5412 => x"9c",
          5413 => x"33",
          5414 => x"2e",
          5415 => x"76",
          5416 => x"58",
          5417 => x"57",
          5418 => x"09",
          5419 => x"38",
          5420 => x"78",
          5421 => x"38",
          5422 => x"81",
          5423 => x"8d",
          5424 => x"fa",
          5425 => x"70",
          5426 => x"56",
          5427 => x"2e",
          5428 => x"8e",
          5429 => x"0c",
          5430 => x"53",
          5431 => x"81",
          5432 => x"75",
          5433 => x"73",
          5434 => x"38",
          5435 => x"30",
          5436 => x"77",
          5437 => x"72",
          5438 => x"a0",
          5439 => x"06",
          5440 => x"75",
          5441 => x"57",
          5442 => x"75",
          5443 => x"d9",
          5444 => x"08",
          5445 => x"52",
          5446 => x"f8",
          5447 => x"cc",
          5448 => x"84",
          5449 => x"72",
          5450 => x"a9",
          5451 => x"70",
          5452 => x"57",
          5453 => x"27",
          5454 => x"53",
          5455 => x"cc",
          5456 => x"0d",
          5457 => x"0d",
          5458 => x"93",
          5459 => x"38",
          5460 => x"81",
          5461 => x"52",
          5462 => x"81",
          5463 => x"81",
          5464 => x"ce",
          5465 => x"f9",
          5466 => x"88",
          5467 => x"39",
          5468 => x"51",
          5469 => x"81",
          5470 => x"80",
          5471 => x"cf",
          5472 => x"dd",
          5473 => x"d0",
          5474 => x"39",
          5475 => x"51",
          5476 => x"81",
          5477 => x"80",
          5478 => x"d0",
          5479 => x"c1",
          5480 => x"a8",
          5481 => x"81",
          5482 => x"b5",
          5483 => x"d8",
          5484 => x"81",
          5485 => x"a9",
          5486 => x"98",
          5487 => x"81",
          5488 => x"9d",
          5489 => x"cc",
          5490 => x"81",
          5491 => x"91",
          5492 => x"fc",
          5493 => x"81",
          5494 => x"85",
          5495 => x"a0",
          5496 => x"9f",
          5497 => x"0d",
          5498 => x"0d",
          5499 => x"56",
          5500 => x"26",
          5501 => x"52",
          5502 => x"29",
          5503 => x"87",
          5504 => x"51",
          5505 => x"3f",
          5506 => x"08",
          5507 => x"fe",
          5508 => x"81",
          5509 => x"54",
          5510 => x"52",
          5511 => x"51",
          5512 => x"3f",
          5513 => x"04",
          5514 => x"66",
          5515 => x"80",
          5516 => x"5b",
          5517 => x"78",
          5518 => x"07",
          5519 => x"57",
          5520 => x"56",
          5521 => x"26",
          5522 => x"56",
          5523 => x"70",
          5524 => x"51",
          5525 => x"74",
          5526 => x"81",
          5527 => x"8c",
          5528 => x"56",
          5529 => x"81",
          5530 => x"57",
          5531 => x"08",
          5532 => x"dc",
          5533 => x"c0",
          5534 => x"81",
          5535 => x"59",
          5536 => x"05",
          5537 => x"53",
          5538 => x"51",
          5539 => x"81",
          5540 => x"57",
          5541 => x"08",
          5542 => x"55",
          5543 => x"89",
          5544 => x"75",
          5545 => x"d8",
          5546 => x"d8",
          5547 => x"c4",
          5548 => x"70",
          5549 => x"25",
          5550 => x"9f",
          5551 => x"51",
          5552 => x"74",
          5553 => x"38",
          5554 => x"53",
          5555 => x"88",
          5556 => x"51",
          5557 => x"76",
          5558 => x"dc",
          5559 => x"3d",
          5560 => x"3d",
          5561 => x"84",
          5562 => x"33",
          5563 => x"57",
          5564 => x"52",
          5565 => x"b0",
          5566 => x"cc",
          5567 => x"75",
          5568 => x"38",
          5569 => x"98",
          5570 => x"60",
          5571 => x"81",
          5572 => x"7e",
          5573 => x"77",
          5574 => x"cc",
          5575 => x"39",
          5576 => x"81",
          5577 => x"89",
          5578 => x"f3",
          5579 => x"61",
          5580 => x"05",
          5581 => x"33",
          5582 => x"68",
          5583 => x"5c",
          5584 => x"7a",
          5585 => x"dc",
          5586 => x"9b",
          5587 => x"e4",
          5588 => x"af",
          5589 => x"74",
          5590 => x"fc",
          5591 => x"2e",
          5592 => x"a0",
          5593 => x"80",
          5594 => x"18",
          5595 => x"27",
          5596 => x"22",
          5597 => x"e8",
          5598 => x"eb",
          5599 => x"81",
          5600 => x"ff",
          5601 => x"82",
          5602 => x"c3",
          5603 => x"53",
          5604 => x"8e",
          5605 => x"52",
          5606 => x"51",
          5607 => x"3f",
          5608 => x"d2",
          5609 => x"82",
          5610 => x"15",
          5611 => x"74",
          5612 => x"7a",
          5613 => x"72",
          5614 => x"d2",
          5615 => x"88",
          5616 => x"39",
          5617 => x"51",
          5618 => x"3f",
          5619 => x"a0",
          5620 => x"d2",
          5621 => x"39",
          5622 => x"51",
          5623 => x"3f",
          5624 => x"79",
          5625 => x"74",
          5626 => x"55",
          5627 => x"72",
          5628 => x"38",
          5629 => x"53",
          5630 => x"83",
          5631 => x"75",
          5632 => x"81",
          5633 => x"53",
          5634 => x"8b",
          5635 => x"fe",
          5636 => x"73",
          5637 => x"a0",
          5638 => x"8a",
          5639 => x"55",
          5640 => x"d3",
          5641 => x"81",
          5642 => x"18",
          5643 => x"58",
          5644 => x"3f",
          5645 => x"08",
          5646 => x"98",
          5647 => x"76",
          5648 => x"81",
          5649 => x"fe",
          5650 => x"81",
          5651 => x"98",
          5652 => x"2c",
          5653 => x"70",
          5654 => x"32",
          5655 => x"72",
          5656 => x"07",
          5657 => x"58",
          5658 => x"57",
          5659 => x"d7",
          5660 => x"2e",
          5661 => x"85",
          5662 => x"8c",
          5663 => x"53",
          5664 => x"fd",
          5665 => x"53",
          5666 => x"cc",
          5667 => x"0d",
          5668 => x"0d",
          5669 => x"33",
          5670 => x"53",
          5671 => x"52",
          5672 => x"c3",
          5673 => x"ac",
          5674 => x"ff",
          5675 => x"d3",
          5676 => x"d3",
          5677 => x"d9",
          5678 => x"81",
          5679 => x"ff",
          5680 => x"74",
          5681 => x"38",
          5682 => x"3f",
          5683 => x"04",
          5684 => x"87",
          5685 => x"08",
          5686 => x"b8",
          5687 => x"fe",
          5688 => x"81",
          5689 => x"fe",
          5690 => x"80",
          5691 => x"b5",
          5692 => x"2a",
          5693 => x"51",
          5694 => x"2e",
          5695 => x"51",
          5696 => x"3f",
          5697 => x"51",
          5698 => x"3f",
          5699 => x"f1",
          5700 => x"82",
          5701 => x"06",
          5702 => x"80",
          5703 => x"81",
          5704 => x"81",
          5705 => x"fc",
          5706 => x"f9",
          5707 => x"fe",
          5708 => x"72",
          5709 => x"81",
          5710 => x"71",
          5711 => x"38",
          5712 => x"f0",
          5713 => x"d4",
          5714 => x"f2",
          5715 => x"51",
          5716 => x"3f",
          5717 => x"70",
          5718 => x"52",
          5719 => x"95",
          5720 => x"fe",
          5721 => x"81",
          5722 => x"fe",
          5723 => x"80",
          5724 => x"b1",
          5725 => x"2a",
          5726 => x"51",
          5727 => x"2e",
          5728 => x"51",
          5729 => x"3f",
          5730 => x"51",
          5731 => x"3f",
          5732 => x"f0",
          5733 => x"86",
          5734 => x"06",
          5735 => x"80",
          5736 => x"81",
          5737 => x"fd",
          5738 => x"c8",
          5739 => x"f5",
          5740 => x"fe",
          5741 => x"72",
          5742 => x"81",
          5743 => x"71",
          5744 => x"38",
          5745 => x"ef",
          5746 => x"d4",
          5747 => x"f1",
          5748 => x"51",
          5749 => x"3f",
          5750 => x"70",
          5751 => x"52",
          5752 => x"95",
          5753 => x"fe",
          5754 => x"81",
          5755 => x"fe",
          5756 => x"80",
          5757 => x"ad",
          5758 => x"a0",
          5759 => x"0d",
          5760 => x"0d",
          5761 => x"55",
          5762 => x"52",
          5763 => x"e8",
          5764 => x"d9",
          5765 => x"73",
          5766 => x"53",
          5767 => x"52",
          5768 => x"51",
          5769 => x"3f",
          5770 => x"08",
          5771 => x"dc",
          5772 => x"80",
          5773 => x"31",
          5774 => x"73",
          5775 => x"34",
          5776 => x"33",
          5777 => x"2e",
          5778 => x"ac",
          5779 => x"d0",
          5780 => x"75",
          5781 => x"3f",
          5782 => x"08",
          5783 => x"38",
          5784 => x"08",
          5785 => x"9b",
          5786 => x"81",
          5787 => x"c6",
          5788 => x"0b",
          5789 => x"34",
          5790 => x"33",
          5791 => x"2e",
          5792 => x"89",
          5793 => x"75",
          5794 => x"b5",
          5795 => x"81",
          5796 => x"87",
          5797 => x"ce",
          5798 => x"70",
          5799 => x"cc",
          5800 => x"81",
          5801 => x"ff",
          5802 => x"81",
          5803 => x"81",
          5804 => x"78",
          5805 => x"81",
          5806 => x"81",
          5807 => x"96",
          5808 => x"59",
          5809 => x"3f",
          5810 => x"52",
          5811 => x"51",
          5812 => x"3f",
          5813 => x"08",
          5814 => x"38",
          5815 => x"51",
          5816 => x"81",
          5817 => x"81",
          5818 => x"fe",
          5819 => x"96",
          5820 => x"5a",
          5821 => x"79",
          5822 => x"3f",
          5823 => x"84",
          5824 => x"bf",
          5825 => x"cc",
          5826 => x"70",
          5827 => x"59",
          5828 => x"2e",
          5829 => x"78",
          5830 => x"b2",
          5831 => x"2e",
          5832 => x"78",
          5833 => x"38",
          5834 => x"ff",
          5835 => x"bc",
          5836 => x"38",
          5837 => x"78",
          5838 => x"83",
          5839 => x"80",
          5840 => x"dd",
          5841 => x"2e",
          5842 => x"8a",
          5843 => x"80",
          5844 => x"ea",
          5845 => x"f9",
          5846 => x"78",
          5847 => x"88",
          5848 => x"80",
          5849 => x"b1",
          5850 => x"39",
          5851 => x"2e",
          5852 => x"78",
          5853 => x"8b",
          5854 => x"82",
          5855 => x"38",
          5856 => x"78",
          5857 => x"8a",
          5858 => x"93",
          5859 => x"ff",
          5860 => x"ff",
          5861 => x"ff",
          5862 => x"81",
          5863 => x"80",
          5864 => x"38",
          5865 => x"fc",
          5866 => x"84",
          5867 => x"82",
          5868 => x"dc",
          5869 => x"2e",
          5870 => x"b4",
          5871 => x"11",
          5872 => x"05",
          5873 => x"94",
          5874 => x"cc",
          5875 => x"81",
          5876 => x"42",
          5877 => x"51",
          5878 => x"3f",
          5879 => x"5a",
          5880 => x"81",
          5881 => x"59",
          5882 => x"84",
          5883 => x"7a",
          5884 => x"38",
          5885 => x"b4",
          5886 => x"11",
          5887 => x"05",
          5888 => x"d8",
          5889 => x"cc",
          5890 => x"fd",
          5891 => x"3d",
          5892 => x"53",
          5893 => x"51",
          5894 => x"3f",
          5895 => x"08",
          5896 => x"c3",
          5897 => x"fe",
          5898 => x"ff",
          5899 => x"ff",
          5900 => x"81",
          5901 => x"80",
          5902 => x"38",
          5903 => x"51",
          5904 => x"3f",
          5905 => x"63",
          5906 => x"38",
          5907 => x"70",
          5908 => x"33",
          5909 => x"81",
          5910 => x"39",
          5911 => x"80",
          5912 => x"84",
          5913 => x"80",
          5914 => x"dc",
          5915 => x"2e",
          5916 => x"b4",
          5917 => x"11",
          5918 => x"05",
          5919 => x"dc",
          5920 => x"cc",
          5921 => x"fc",
          5922 => x"3d",
          5923 => x"53",
          5924 => x"51",
          5925 => x"3f",
          5926 => x"08",
          5927 => x"c7",
          5928 => x"9c",
          5929 => x"db",
          5930 => x"79",
          5931 => x"38",
          5932 => x"7b",
          5933 => x"5b",
          5934 => x"92",
          5935 => x"7a",
          5936 => x"53",
          5937 => x"d6",
          5938 => x"fe",
          5939 => x"1a",
          5940 => x"43",
          5941 => x"81",
          5942 => x"82",
          5943 => x"3d",
          5944 => x"53",
          5945 => x"51",
          5946 => x"3f",
          5947 => x"08",
          5948 => x"81",
          5949 => x"59",
          5950 => x"89",
          5951 => x"f8",
          5952 => x"cd",
          5953 => x"c1",
          5954 => x"80",
          5955 => x"81",
          5956 => x"44",
          5957 => x"d9",
          5958 => x"78",
          5959 => x"38",
          5960 => x"08",
          5961 => x"81",
          5962 => x"59",
          5963 => x"88",
          5964 => x"90",
          5965 => x"39",
          5966 => x"33",
          5967 => x"2e",
          5968 => x"d9",
          5969 => x"89",
          5970 => x"a8",
          5971 => x"05",
          5972 => x"fe",
          5973 => x"ff",
          5974 => x"fe",
          5975 => x"81",
          5976 => x"80",
          5977 => x"d9",
          5978 => x"78",
          5979 => x"38",
          5980 => x"08",
          5981 => x"39",
          5982 => x"33",
          5983 => x"2e",
          5984 => x"d9",
          5985 => x"bb",
          5986 => x"c2",
          5987 => x"80",
          5988 => x"81",
          5989 => x"43",
          5990 => x"d9",
          5991 => x"78",
          5992 => x"38",
          5993 => x"08",
          5994 => x"81",
          5995 => x"59",
          5996 => x"88",
          5997 => x"9c",
          5998 => x"39",
          5999 => x"08",
          6000 => x"b4",
          6001 => x"11",
          6002 => x"05",
          6003 => x"8c",
          6004 => x"cc",
          6005 => x"a7",
          6006 => x"5c",
          6007 => x"2e",
          6008 => x"5c",
          6009 => x"70",
          6010 => x"07",
          6011 => x"7f",
          6012 => x"5a",
          6013 => x"2e",
          6014 => x"a0",
          6015 => x"88",
          6016 => x"c8",
          6017 => x"fb",
          6018 => x"63",
          6019 => x"62",
          6020 => x"f2",
          6021 => x"d6",
          6022 => x"f5",
          6023 => x"c7",
          6024 => x"ff",
          6025 => x"ff",
          6026 => x"fe",
          6027 => x"81",
          6028 => x"80",
          6029 => x"38",
          6030 => x"fc",
          6031 => x"84",
          6032 => x"fd",
          6033 => x"dc",
          6034 => x"2e",
          6035 => x"59",
          6036 => x"05",
          6037 => x"63",
          6038 => x"b4",
          6039 => x"11",
          6040 => x"05",
          6041 => x"f4",
          6042 => x"cc",
          6043 => x"f8",
          6044 => x"70",
          6045 => x"81",
          6046 => x"fe",
          6047 => x"80",
          6048 => x"51",
          6049 => x"3f",
          6050 => x"33",
          6051 => x"2e",
          6052 => x"9f",
          6053 => x"38",
          6054 => x"fc",
          6055 => x"84",
          6056 => x"fc",
          6057 => x"dc",
          6058 => x"2e",
          6059 => x"59",
          6060 => x"05",
          6061 => x"63",
          6062 => x"ff",
          6063 => x"d6",
          6064 => x"f4",
          6065 => x"aa",
          6066 => x"fe",
          6067 => x"ff",
          6068 => x"fe",
          6069 => x"81",
          6070 => x"80",
          6071 => x"38",
          6072 => x"f0",
          6073 => x"84",
          6074 => x"fd",
          6075 => x"dc",
          6076 => x"2e",
          6077 => x"59",
          6078 => x"22",
          6079 => x"05",
          6080 => x"41",
          6081 => x"f0",
          6082 => x"84",
          6083 => x"fd",
          6084 => x"dc",
          6085 => x"38",
          6086 => x"60",
          6087 => x"52",
          6088 => x"51",
          6089 => x"3f",
          6090 => x"79",
          6091 => x"91",
          6092 => x"79",
          6093 => x"ae",
          6094 => x"38",
          6095 => x"87",
          6096 => x"05",
          6097 => x"b4",
          6098 => x"11",
          6099 => x"05",
          6100 => x"fa",
          6101 => x"cc",
          6102 => x"92",
          6103 => x"02",
          6104 => x"79",
          6105 => x"5b",
          6106 => x"ff",
          6107 => x"d6",
          6108 => x"f3",
          6109 => x"a3",
          6110 => x"fe",
          6111 => x"ff",
          6112 => x"fe",
          6113 => x"81",
          6114 => x"80",
          6115 => x"38",
          6116 => x"f0",
          6117 => x"84",
          6118 => x"fc",
          6119 => x"dc",
          6120 => x"2e",
          6121 => x"60",
          6122 => x"60",
          6123 => x"b4",
          6124 => x"11",
          6125 => x"05",
          6126 => x"92",
          6127 => x"cc",
          6128 => x"f6",
          6129 => x"70",
          6130 => x"81",
          6131 => x"fe",
          6132 => x"80",
          6133 => x"51",
          6134 => x"3f",
          6135 => x"33",
          6136 => x"2e",
          6137 => x"9f",
          6138 => x"38",
          6139 => x"f0",
          6140 => x"84",
          6141 => x"fb",
          6142 => x"dc",
          6143 => x"2e",
          6144 => x"60",
          6145 => x"60",
          6146 => x"ff",
          6147 => x"d6",
          6148 => x"f1",
          6149 => x"ae",
          6150 => x"ff",
          6151 => x"ff",
          6152 => x"fe",
          6153 => x"81",
          6154 => x"80",
          6155 => x"38",
          6156 => x"d7",
          6157 => x"f7",
          6158 => x"59",
          6159 => x"3d",
          6160 => x"53",
          6161 => x"51",
          6162 => x"3f",
          6163 => x"08",
          6164 => x"93",
          6165 => x"81",
          6166 => x"fe",
          6167 => x"63",
          6168 => x"81",
          6169 => x"80",
          6170 => x"38",
          6171 => x"08",
          6172 => x"c8",
          6173 => x"ef",
          6174 => x"39",
          6175 => x"51",
          6176 => x"3f",
          6177 => x"3f",
          6178 => x"81",
          6179 => x"fe",
          6180 => x"80",
          6181 => x"39",
          6182 => x"3f",
          6183 => x"64",
          6184 => x"59",
          6185 => x"f4",
          6186 => x"7d",
          6187 => x"80",
          6188 => x"38",
          6189 => x"84",
          6190 => x"de",
          6191 => x"dc",
          6192 => x"81",
          6193 => x"2e",
          6194 => x"82",
          6195 => x"7a",
          6196 => x"38",
          6197 => x"7a",
          6198 => x"38",
          6199 => x"81",
          6200 => x"7b",
          6201 => x"98",
          6202 => x"81",
          6203 => x"b4",
          6204 => x"05",
          6205 => x"85",
          6206 => x"81",
          6207 => x"b4",
          6208 => x"05",
          6209 => x"f5",
          6210 => x"7b",
          6211 => x"98",
          6212 => x"81",
          6213 => x"b4",
          6214 => x"05",
          6215 => x"dd",
          6216 => x"7b",
          6217 => x"81",
          6218 => x"b4",
          6219 => x"05",
          6220 => x"c9",
          6221 => x"f8",
          6222 => x"80",
          6223 => x"64",
          6224 => x"81",
          6225 => x"54",
          6226 => x"53",
          6227 => x"52",
          6228 => x"b0",
          6229 => x"8a",
          6230 => x"cc",
          6231 => x"cc",
          6232 => x"30",
          6233 => x"80",
          6234 => x"5b",
          6235 => x"7a",
          6236 => x"38",
          6237 => x"7a",
          6238 => x"80",
          6239 => x"81",
          6240 => x"ff",
          6241 => x"7a",
          6242 => x"7d",
          6243 => x"81",
          6244 => x"78",
          6245 => x"ff",
          6246 => x"06",
          6247 => x"81",
          6248 => x"fe",
          6249 => x"f2",
          6250 => x"3d",
          6251 => x"81",
          6252 => x"87",
          6253 => x"70",
          6254 => x"87",
          6255 => x"72",
          6256 => x"b8",
          6257 => x"cc",
          6258 => x"75",
          6259 => x"87",
          6260 => x"73",
          6261 => x"a4",
          6262 => x"dc",
          6263 => x"75",
          6264 => x"94",
          6265 => x"54",
          6266 => x"80",
          6267 => x"fe",
          6268 => x"81",
          6269 => x"90",
          6270 => x"55",
          6271 => x"80",
          6272 => x"fe",
          6273 => x"72",
          6274 => x"08",
          6275 => x"8c",
          6276 => x"87",
          6277 => x"0c",
          6278 => x"0b",
          6279 => x"94",
          6280 => x"0b",
          6281 => x"0c",
          6282 => x"81",
          6283 => x"fe",
          6284 => x"fe",
          6285 => x"81",
          6286 => x"fe",
          6287 => x"81",
          6288 => x"fe",
          6289 => x"81",
          6290 => x"fe",
          6291 => x"81",
          6292 => x"3f",
          6293 => x"80",
          6294 => x"00",
          6295 => x"ff",
          6296 => x"ff",
          6297 => x"ff",
          6298 => x"00",
          6299 => x"00",
          6300 => x"00",
          6301 => x"00",
          6302 => x"00",
          6303 => x"00",
          6304 => x"00",
          6305 => x"00",
          6306 => x"00",
          6307 => x"00",
          6308 => x"00",
          6309 => x"00",
          6310 => x"00",
          6311 => x"00",
          6312 => x"00",
          6313 => x"00",
          6314 => x"00",
          6315 => x"00",
          6316 => x"00",
          6317 => x"00",
          6318 => x"00",
          6319 => x"00",
          6320 => x"00",
          6321 => x"00",
          6322 => x"00",
          6323 => x"25",
          6324 => x"64",
          6325 => x"20",
          6326 => x"25",
          6327 => x"64",
          6328 => x"25",
          6329 => x"53",
          6330 => x"43",
          6331 => x"69",
          6332 => x"61",
          6333 => x"6e",
          6334 => x"20",
          6335 => x"6f",
          6336 => x"6f",
          6337 => x"6f",
          6338 => x"67",
          6339 => x"3a",
          6340 => x"76",
          6341 => x"73",
          6342 => x"70",
          6343 => x"65",
          6344 => x"64",
          6345 => x"20",
          6346 => x"57",
          6347 => x"44",
          6348 => x"20",
          6349 => x"30",
          6350 => x"25",
          6351 => x"29",
          6352 => x"20",
          6353 => x"53",
          6354 => x"4d",
          6355 => x"20",
          6356 => x"30",
          6357 => x"25",
          6358 => x"29",
          6359 => x"20",
          6360 => x"49",
          6361 => x"20",
          6362 => x"4d",
          6363 => x"30",
          6364 => x"25",
          6365 => x"29",
          6366 => x"20",
          6367 => x"42",
          6368 => x"20",
          6369 => x"20",
          6370 => x"30",
          6371 => x"25",
          6372 => x"29",
          6373 => x"20",
          6374 => x"52",
          6375 => x"20",
          6376 => x"20",
          6377 => x"30",
          6378 => x"25",
          6379 => x"29",
          6380 => x"20",
          6381 => x"53",
          6382 => x"41",
          6383 => x"20",
          6384 => x"65",
          6385 => x"65",
          6386 => x"25",
          6387 => x"29",
          6388 => x"20",
          6389 => x"54",
          6390 => x"52",
          6391 => x"20",
          6392 => x"69",
          6393 => x"73",
          6394 => x"25",
          6395 => x"29",
          6396 => x"20",
          6397 => x"49",
          6398 => x"20",
          6399 => x"4c",
          6400 => x"68",
          6401 => x"65",
          6402 => x"25",
          6403 => x"29",
          6404 => x"20",
          6405 => x"57",
          6406 => x"42",
          6407 => x"20",
          6408 => x"0a",
          6409 => x"20",
          6410 => x"57",
          6411 => x"32",
          6412 => x"20",
          6413 => x"49",
          6414 => x"4c",
          6415 => x"20",
          6416 => x"50",
          6417 => x"00",
          6418 => x"20",
          6419 => x"53",
          6420 => x"00",
          6421 => x"41",
          6422 => x"65",
          6423 => x"73",
          6424 => x"20",
          6425 => x"43",
          6426 => x"52",
          6427 => x"74",
          6428 => x"63",
          6429 => x"20",
          6430 => x"72",
          6431 => x"20",
          6432 => x"30",
          6433 => x"00",
          6434 => x"20",
          6435 => x"43",
          6436 => x"4d",
          6437 => x"72",
          6438 => x"74",
          6439 => x"20",
          6440 => x"72",
          6441 => x"20",
          6442 => x"30",
          6443 => x"00",
          6444 => x"20",
          6445 => x"53",
          6446 => x"6b",
          6447 => x"61",
          6448 => x"41",
          6449 => x"65",
          6450 => x"20",
          6451 => x"20",
          6452 => x"30",
          6453 => x"00",
          6454 => x"4d",
          6455 => x"3a",
          6456 => x"20",
          6457 => x"5a",
          6458 => x"49",
          6459 => x"20",
          6460 => x"20",
          6461 => x"20",
          6462 => x"20",
          6463 => x"20",
          6464 => x"30",
          6465 => x"00",
          6466 => x"20",
          6467 => x"53",
          6468 => x"65",
          6469 => x"6c",
          6470 => x"20",
          6471 => x"71",
          6472 => x"20",
          6473 => x"20",
          6474 => x"64",
          6475 => x"34",
          6476 => x"7a",
          6477 => x"20",
          6478 => x"53",
          6479 => x"4d",
          6480 => x"6f",
          6481 => x"46",
          6482 => x"20",
          6483 => x"20",
          6484 => x"20",
          6485 => x"64",
          6486 => x"34",
          6487 => x"7a",
          6488 => x"20",
          6489 => x"57",
          6490 => x"62",
          6491 => x"20",
          6492 => x"41",
          6493 => x"6c",
          6494 => x"20",
          6495 => x"71",
          6496 => x"64",
          6497 => x"34",
          6498 => x"7a",
          6499 => x"53",
          6500 => x"6c",
          6501 => x"4d",
          6502 => x"75",
          6503 => x"46",
          6504 => x"00",
          6505 => x"45",
          6506 => x"45",
          6507 => x"69",
          6508 => x"55",
          6509 => x"6f",
          6510 => x"53",
          6511 => x"22",
          6512 => x"3a",
          6513 => x"3e",
          6514 => x"7c",
          6515 => x"46",
          6516 => x"46",
          6517 => x"32",
          6518 => x"eb",
          6519 => x"53",
          6520 => x"35",
          6521 => x"4e",
          6522 => x"41",
          6523 => x"20",
          6524 => x"41",
          6525 => x"20",
          6526 => x"4e",
          6527 => x"41",
          6528 => x"20",
          6529 => x"41",
          6530 => x"20",
          6531 => x"00",
          6532 => x"00",
          6533 => x"00",
          6534 => x"00",
          6535 => x"80",
          6536 => x"8e",
          6537 => x"45",
          6538 => x"49",
          6539 => x"90",
          6540 => x"99",
          6541 => x"59",
          6542 => x"9c",
          6543 => x"41",
          6544 => x"a5",
          6545 => x"a8",
          6546 => x"ac",
          6547 => x"b0",
          6548 => x"b4",
          6549 => x"b8",
          6550 => x"bc",
          6551 => x"c0",
          6552 => x"c4",
          6553 => x"c8",
          6554 => x"cc",
          6555 => x"d0",
          6556 => x"d4",
          6557 => x"d8",
          6558 => x"dc",
          6559 => x"e0",
          6560 => x"e4",
          6561 => x"e8",
          6562 => x"ec",
          6563 => x"f0",
          6564 => x"f4",
          6565 => x"f8",
          6566 => x"fc",
          6567 => x"2b",
          6568 => x"3d",
          6569 => x"5c",
          6570 => x"3c",
          6571 => x"7f",
          6572 => x"00",
          6573 => x"00",
          6574 => x"01",
          6575 => x"00",
          6576 => x"00",
          6577 => x"00",
          6578 => x"00",
          6579 => x"00",
          6580 => x"64",
          6581 => x"74",
          6582 => x"64",
          6583 => x"74",
          6584 => x"66",
          6585 => x"74",
          6586 => x"66",
          6587 => x"64",
          6588 => x"66",
          6589 => x"63",
          6590 => x"6d",
          6591 => x"61",
          6592 => x"6d",
          6593 => x"79",
          6594 => x"6d",
          6595 => x"66",
          6596 => x"6d",
          6597 => x"70",
          6598 => x"6d",
          6599 => x"6d",
          6600 => x"6d",
          6601 => x"68",
          6602 => x"68",
          6603 => x"68",
          6604 => x"68",
          6605 => x"63",
          6606 => x"00",
          6607 => x"6a",
          6608 => x"72",
          6609 => x"61",
          6610 => x"72",
          6611 => x"74",
          6612 => x"69",
          6613 => x"00",
          6614 => x"74",
          6615 => x"00",
          6616 => x"74",
          6617 => x"69",
          6618 => x"44",
          6619 => x"20",
          6620 => x"6f",
          6621 => x"49",
          6622 => x"72",
          6623 => x"20",
          6624 => x"6f",
          6625 => x"00",
          6626 => x"44",
          6627 => x"20",
          6628 => x"20",
          6629 => x"64",
          6630 => x"00",
          6631 => x"4e",
          6632 => x"69",
          6633 => x"66",
          6634 => x"64",
          6635 => x"4e",
          6636 => x"61",
          6637 => x"66",
          6638 => x"64",
          6639 => x"49",
          6640 => x"6c",
          6641 => x"66",
          6642 => x"6e",
          6643 => x"2e",
          6644 => x"41",
          6645 => x"73",
          6646 => x"65",
          6647 => x"64",
          6648 => x"46",
          6649 => x"20",
          6650 => x"65",
          6651 => x"20",
          6652 => x"73",
          6653 => x"0a",
          6654 => x"46",
          6655 => x"20",
          6656 => x"64",
          6657 => x"69",
          6658 => x"6c",
          6659 => x"0a",
          6660 => x"53",
          6661 => x"73",
          6662 => x"69",
          6663 => x"70",
          6664 => x"65",
          6665 => x"64",
          6666 => x"44",
          6667 => x"65",
          6668 => x"6d",
          6669 => x"20",
          6670 => x"69",
          6671 => x"6c",
          6672 => x"0a",
          6673 => x"44",
          6674 => x"20",
          6675 => x"20",
          6676 => x"62",
          6677 => x"2e",
          6678 => x"4e",
          6679 => x"6f",
          6680 => x"74",
          6681 => x"65",
          6682 => x"6c",
          6683 => x"73",
          6684 => x"20",
          6685 => x"6e",
          6686 => x"6e",
          6687 => x"73",
          6688 => x"00",
          6689 => x"46",
          6690 => x"61",
          6691 => x"62",
          6692 => x"65",
          6693 => x"00",
          6694 => x"54",
          6695 => x"6f",
          6696 => x"20",
          6697 => x"72",
          6698 => x"6f",
          6699 => x"61",
          6700 => x"6c",
          6701 => x"2e",
          6702 => x"46",
          6703 => x"20",
          6704 => x"6c",
          6705 => x"65",
          6706 => x"00",
          6707 => x"49",
          6708 => x"66",
          6709 => x"69",
          6710 => x"20",
          6711 => x"6f",
          6712 => x"0a",
          6713 => x"54",
          6714 => x"6d",
          6715 => x"20",
          6716 => x"6e",
          6717 => x"6c",
          6718 => x"0a",
          6719 => x"50",
          6720 => x"6d",
          6721 => x"72",
          6722 => x"6e",
          6723 => x"72",
          6724 => x"2e",
          6725 => x"53",
          6726 => x"65",
          6727 => x"0a",
          6728 => x"55",
          6729 => x"6f",
          6730 => x"65",
          6731 => x"72",
          6732 => x"0a",
          6733 => x"20",
          6734 => x"65",
          6735 => x"73",
          6736 => x"20",
          6737 => x"20",
          6738 => x"65",
          6739 => x"65",
          6740 => x"00",
          6741 => x"72",
          6742 => x"00",
          6743 => x"25",
          6744 => x"00",
          6745 => x"3a",
          6746 => x"25",
          6747 => x"00",
          6748 => x"20",
          6749 => x"20",
          6750 => x"00",
          6751 => x"25",
          6752 => x"00",
          6753 => x"20",
          6754 => x"20",
          6755 => x"7c",
          6756 => x"7a",
          6757 => x"0a",
          6758 => x"25",
          6759 => x"00",
          6760 => x"31",
          6761 => x"34",
          6762 => x"32",
          6763 => x"76",
          6764 => x"00",
          6765 => x"20",
          6766 => x"2c",
          6767 => x"76",
          6768 => x"32",
          6769 => x"25",
          6770 => x"73",
          6771 => x"0a",
          6772 => x"5a",
          6773 => x"49",
          6774 => x"72",
          6775 => x"74",
          6776 => x"6e",
          6777 => x"72",
          6778 => x"54",
          6779 => x"72",
          6780 => x"74",
          6781 => x"75",
          6782 => x"00",
          6783 => x"50",
          6784 => x"69",
          6785 => x"72",
          6786 => x"74",
          6787 => x"49",
          6788 => x"4c",
          6789 => x"20",
          6790 => x"65",
          6791 => x"70",
          6792 => x"49",
          6793 => x"4c",
          6794 => x"20",
          6795 => x"65",
          6796 => x"70",
          6797 => x"55",
          6798 => x"30",
          6799 => x"20",
          6800 => x"65",
          6801 => x"70",
          6802 => x"55",
          6803 => x"30",
          6804 => x"20",
          6805 => x"65",
          6806 => x"70",
          6807 => x"55",
          6808 => x"31",
          6809 => x"20",
          6810 => x"65",
          6811 => x"70",
          6812 => x"55",
          6813 => x"31",
          6814 => x"20",
          6815 => x"65",
          6816 => x"70",
          6817 => x"53",
          6818 => x"69",
          6819 => x"75",
          6820 => x"69",
          6821 => x"2e",
          6822 => x"00",
          6823 => x"45",
          6824 => x"6c",
          6825 => x"20",
          6826 => x"65",
          6827 => x"2e",
          6828 => x"61",
          6829 => x"65",
          6830 => x"2e",
          6831 => x"00",
          6832 => x"30",
          6833 => x"46",
          6834 => x"65",
          6835 => x"6f",
          6836 => x"69",
          6837 => x"6c",
          6838 => x"20",
          6839 => x"63",
          6840 => x"20",
          6841 => x"70",
          6842 => x"73",
          6843 => x"6e",
          6844 => x"6d",
          6845 => x"61",
          6846 => x"2e",
          6847 => x"2a",
          6848 => x"43",
          6849 => x"72",
          6850 => x"2e",
          6851 => x"00",
          6852 => x"43",
          6853 => x"69",
          6854 => x"2e",
          6855 => x"43",
          6856 => x"61",
          6857 => x"67",
          6858 => x"00",
          6859 => x"25",
          6860 => x"78",
          6861 => x"38",
          6862 => x"3e",
          6863 => x"6c",
          6864 => x"30",
          6865 => x"0a",
          6866 => x"44",
          6867 => x"20",
          6868 => x"6f",
          6869 => x"00",
          6870 => x"0a",
          6871 => x"70",
          6872 => x"65",
          6873 => x"25",
          6874 => x"20",
          6875 => x"58",
          6876 => x"3f",
          6877 => x"00",
          6878 => x"25",
          6879 => x"20",
          6880 => x"58",
          6881 => x"25",
          6882 => x"20",
          6883 => x"58",
          6884 => x"45",
          6885 => x"75",
          6886 => x"67",
          6887 => x"64",
          6888 => x"20",
          6889 => x"78",
          6890 => x"2e",
          6891 => x"43",
          6892 => x"69",
          6893 => x"63",
          6894 => x"20",
          6895 => x"30",
          6896 => x"2e",
          6897 => x"00",
          6898 => x"43",
          6899 => x"20",
          6900 => x"75",
          6901 => x"64",
          6902 => x"64",
          6903 => x"25",
          6904 => x"0a",
          6905 => x"52",
          6906 => x"61",
          6907 => x"6e",
          6908 => x"70",
          6909 => x"63",
          6910 => x"6f",
          6911 => x"2e",
          6912 => x"43",
          6913 => x"20",
          6914 => x"6f",
          6915 => x"6e",
          6916 => x"2e",
          6917 => x"5a",
          6918 => x"62",
          6919 => x"25",
          6920 => x"25",
          6921 => x"73",
          6922 => x"00",
          6923 => x"25",
          6924 => x"25",
          6925 => x"73",
          6926 => x"25",
          6927 => x"25",
          6928 => x"42",
          6929 => x"63",
          6930 => x"61",
          6931 => x"0a",
          6932 => x"52",
          6933 => x"69",
          6934 => x"2e",
          6935 => x"45",
          6936 => x"6c",
          6937 => x"20",
          6938 => x"65",
          6939 => x"70",
          6940 => x"2e",
          6941 => x"00",
          6942 => x"00",
          6943 => x"00",
          6944 => x"00",
          6945 => x"00",
          6946 => x"00",
          6947 => x"00",
          6948 => x"00",
          6949 => x"00",
          6950 => x"01",
          6951 => x"01",
          6952 => x"00",
          6953 => x"00",
          6954 => x"00",
          6955 => x"00",
          6956 => x"05",
          6957 => x"05",
          6958 => x"05",
          6959 => x"00",
          6960 => x"01",
          6961 => x"01",
          6962 => x"01",
          6963 => x"01",
          6964 => x"00",
          6965 => x"01",
          6966 => x"00",
          6967 => x"00",
          6968 => x"01",
          6969 => x"00",
          6970 => x"00",
          6971 => x"00",
          6972 => x"01",
          6973 => x"00",
          6974 => x"00",
          6975 => x"00",
          6976 => x"01",
          6977 => x"00",
          6978 => x"00",
          6979 => x"00",
          6980 => x"01",
          6981 => x"00",
          6982 => x"00",
          6983 => x"00",
          6984 => x"01",
          6985 => x"00",
          6986 => x"00",
          6987 => x"00",
          6988 => x"01",
          6989 => x"00",
          6990 => x"00",
          6991 => x"00",
          6992 => x"01",
          6993 => x"00",
          6994 => x"00",
          6995 => x"00",
          6996 => x"01",
          6997 => x"00",
          6998 => x"00",
          6999 => x"00",
          7000 => x"01",
          7001 => x"00",
          7002 => x"00",
          7003 => x"00",
          7004 => x"01",
          7005 => x"00",
          7006 => x"00",
          7007 => x"00",
          7008 => x"01",
          7009 => x"00",
          7010 => x"00",
          7011 => x"00",
          7012 => x"01",
          7013 => x"00",
          7014 => x"00",
          7015 => x"00",
          7016 => x"01",
          7017 => x"00",
          7018 => x"00",
          7019 => x"00",
          7020 => x"01",
          7021 => x"00",
          7022 => x"00",
          7023 => x"00",
          7024 => x"01",
          7025 => x"00",
          7026 => x"00",
          7027 => x"00",
          7028 => x"01",
          7029 => x"00",
          7030 => x"00",
          7031 => x"00",
          7032 => x"01",
          7033 => x"00",
          7034 => x"00",
          7035 => x"00",
          7036 => x"01",
          7037 => x"00",
          7038 => x"00",
          7039 => x"00",
          7040 => x"01",
          7041 => x"00",
          7042 => x"00",
          7043 => x"00",
          7044 => x"01",
          7045 => x"00",
          7046 => x"00",
          7047 => x"00",
          7048 => x"01",
          7049 => x"00",
          7050 => x"00",
          7051 => x"00",
          7052 => x"01",
          7053 => x"00",
          7054 => x"00",
          7055 => x"00",
          7056 => x"01",
          7057 => x"00",
          7058 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
