-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"88",
             1 => x"0b",
             2 => x"04",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"88",
             9 => x"0b",
            10 => x"04",
            11 => x"88",
            12 => x"0b",
            13 => x"04",
            14 => x"88",
            15 => x"0b",
            16 => x"04",
            17 => x"88",
            18 => x"0b",
            19 => x"04",
            20 => x"88",
            21 => x"0b",
            22 => x"04",
            23 => x"89",
            24 => x"0b",
            25 => x"04",
            26 => x"89",
            27 => x"0b",
            28 => x"04",
            29 => x"89",
            30 => x"0b",
            31 => x"04",
            32 => x"89",
            33 => x"0b",
            34 => x"04",
            35 => x"8a",
            36 => x"0b",
            37 => x"04",
            38 => x"8a",
            39 => x"0b",
            40 => x"04",
            41 => x"8a",
            42 => x"0b",
            43 => x"04",
            44 => x"8a",
            45 => x"0b",
            46 => x"04",
            47 => x"8b",
            48 => x"0b",
            49 => x"04",
            50 => x"8b",
            51 => x"0b",
            52 => x"04",
            53 => x"8b",
            54 => x"0b",
            55 => x"04",
            56 => x"8b",
            57 => x"0b",
            58 => x"04",
            59 => x"8c",
            60 => x"0b",
            61 => x"04",
            62 => x"8c",
            63 => x"0b",
            64 => x"04",
            65 => x"8c",
            66 => x"0b",
            67 => x"04",
            68 => x"8c",
            69 => x"0b",
            70 => x"04",
            71 => x"8d",
            72 => x"0b",
            73 => x"04",
            74 => x"8d",
            75 => x"0b",
            76 => x"04",
            77 => x"8d",
            78 => x"0b",
            79 => x"04",
            80 => x"8d",
            81 => x"0b",
            82 => x"04",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"00",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"00",
           137 => x"00",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"00",
           145 => x"00",
           146 => x"00",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"00",
           153 => x"00",
           154 => x"00",
           155 => x"00",
           156 => x"00",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"00",
           161 => x"00",
           162 => x"00",
           163 => x"00",
           164 => x"00",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"00",
           169 => x"00",
           170 => x"00",
           171 => x"00",
           172 => x"00",
           173 => x"00",
           174 => x"00",
           175 => x"00",
           176 => x"00",
           177 => x"00",
           178 => x"00",
           179 => x"00",
           180 => x"00",
           181 => x"00",
           182 => x"00",
           183 => x"00",
           184 => x"00",
           185 => x"00",
           186 => x"00",
           187 => x"00",
           188 => x"00",
           189 => x"00",
           190 => x"00",
           191 => x"00",
           192 => x"00",
           193 => x"00",
           194 => x"00",
           195 => x"00",
           196 => x"00",
           197 => x"00",
           198 => x"00",
           199 => x"00",
           200 => x"00",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"00",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"00",
           233 => x"00",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"00",
           249 => x"00",
           250 => x"00",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"0c",
           258 => x"81",
           259 => x"81",
           260 => x"81",
           261 => x"a2",
           262 => x"cb",
           263 => x"e4",
           264 => x"cb",
           265 => x"b4",
           266 => x"b0",
           267 => x"90",
           268 => x"b0",
           269 => x"2d",
           270 => x"08",
           271 => x"04",
           272 => x"0c",
           273 => x"81",
           274 => x"81",
           275 => x"81",
           276 => x"ab",
           277 => x"cb",
           278 => x"e4",
           279 => x"cb",
           280 => x"f5",
           281 => x"b0",
           282 => x"90",
           283 => x"b0",
           284 => x"2d",
           285 => x"08",
           286 => x"04",
           287 => x"0c",
           288 => x"81",
           289 => x"81",
           290 => x"81",
           291 => x"a9",
           292 => x"cb",
           293 => x"e4",
           294 => x"cb",
           295 => x"cc",
           296 => x"b0",
           297 => x"90",
           298 => x"b0",
           299 => x"2d",
           300 => x"08",
           301 => x"04",
           302 => x"0c",
           303 => x"81",
           304 => x"81",
           305 => x"81",
           306 => x"9b",
           307 => x"cb",
           308 => x"e4",
           309 => x"cb",
           310 => x"bf",
           311 => x"b0",
           312 => x"90",
           313 => x"b0",
           314 => x"2d",
           315 => x"08",
           316 => x"04",
           317 => x"0c",
           318 => x"81",
           319 => x"81",
           320 => x"81",
           321 => x"80",
           322 => x"81",
           323 => x"81",
           324 => x"81",
           325 => x"80",
           326 => x"81",
           327 => x"81",
           328 => x"81",
           329 => x"80",
           330 => x"81",
           331 => x"81",
           332 => x"81",
           333 => x"80",
           334 => x"81",
           335 => x"81",
           336 => x"81",
           337 => x"80",
           338 => x"81",
           339 => x"81",
           340 => x"81",
           341 => x"80",
           342 => x"81",
           343 => x"81",
           344 => x"81",
           345 => x"80",
           346 => x"81",
           347 => x"81",
           348 => x"81",
           349 => x"80",
           350 => x"81",
           351 => x"81",
           352 => x"81",
           353 => x"80",
           354 => x"81",
           355 => x"81",
           356 => x"81",
           357 => x"80",
           358 => x"81",
           359 => x"81",
           360 => x"81",
           361 => x"80",
           362 => x"81",
           363 => x"81",
           364 => x"81",
           365 => x"80",
           366 => x"81",
           367 => x"81",
           368 => x"81",
           369 => x"81",
           370 => x"81",
           371 => x"81",
           372 => x"81",
           373 => x"80",
           374 => x"81",
           375 => x"81",
           376 => x"81",
           377 => x"81",
           378 => x"81",
           379 => x"81",
           380 => x"81",
           381 => x"81",
           382 => x"81",
           383 => x"81",
           384 => x"81",
           385 => x"80",
           386 => x"81",
           387 => x"81",
           388 => x"81",
           389 => x"80",
           390 => x"81",
           391 => x"81",
           392 => x"81",
           393 => x"80",
           394 => x"81",
           395 => x"81",
           396 => x"81",
           397 => x"80",
           398 => x"81",
           399 => x"81",
           400 => x"81",
           401 => x"81",
           402 => x"81",
           403 => x"81",
           404 => x"81",
           405 => x"81",
           406 => x"81",
           407 => x"81",
           408 => x"81",
           409 => x"81",
           410 => x"81",
           411 => x"81",
           412 => x"81",
           413 => x"80",
           414 => x"81",
           415 => x"81",
           416 => x"81",
           417 => x"81",
           418 => x"81",
           419 => x"81",
           420 => x"81",
           421 => x"b0",
           422 => x"cb",
           423 => x"e4",
           424 => x"cb",
           425 => x"96",
           426 => x"b0",
           427 => x"90",
           428 => x"b0",
           429 => x"2d",
           430 => x"08",
           431 => x"04",
           432 => x"0c",
           433 => x"81",
           434 => x"81",
           435 => x"81",
           436 => x"94",
           437 => x"cb",
           438 => x"e4",
           439 => x"cb",
           440 => x"b7",
           441 => x"b0",
           442 => x"90",
           443 => x"b0",
           444 => x"b8",
           445 => x"b0",
           446 => x"90",
           447 => x"a4",
           448 => x"a8",
           449 => x"80",
           450 => x"05",
           451 => x"0b",
           452 => x"04",
           453 => x"81",
           454 => x"3c",
           455 => x"b0",
           456 => x"cb",
           457 => x"3d",
           458 => x"81",
           459 => x"8c",
           460 => x"81",
           461 => x"88",
           462 => x"80",
           463 => x"cb",
           464 => x"81",
           465 => x"54",
           466 => x"81",
           467 => x"04",
           468 => x"08",
           469 => x"b0",
           470 => x"0d",
           471 => x"cb",
           472 => x"05",
           473 => x"cb",
           474 => x"05",
           475 => x"3f",
           476 => x"08",
           477 => x"a4",
           478 => x"3d",
           479 => x"b0",
           480 => x"cb",
           481 => x"81",
           482 => x"fd",
           483 => x"0b",
           484 => x"08",
           485 => x"80",
           486 => x"b0",
           487 => x"0c",
           488 => x"08",
           489 => x"81",
           490 => x"88",
           491 => x"b9",
           492 => x"b0",
           493 => x"08",
           494 => x"38",
           495 => x"cb",
           496 => x"05",
           497 => x"38",
           498 => x"08",
           499 => x"10",
           500 => x"08",
           501 => x"81",
           502 => x"fc",
           503 => x"81",
           504 => x"fc",
           505 => x"b8",
           506 => x"b0",
           507 => x"08",
           508 => x"e1",
           509 => x"b0",
           510 => x"08",
           511 => x"08",
           512 => x"26",
           513 => x"cb",
           514 => x"05",
           515 => x"b0",
           516 => x"08",
           517 => x"b0",
           518 => x"0c",
           519 => x"08",
           520 => x"81",
           521 => x"fc",
           522 => x"81",
           523 => x"f8",
           524 => x"cb",
           525 => x"05",
           526 => x"81",
           527 => x"fc",
           528 => x"cb",
           529 => x"05",
           530 => x"81",
           531 => x"8c",
           532 => x"95",
           533 => x"b0",
           534 => x"08",
           535 => x"38",
           536 => x"08",
           537 => x"70",
           538 => x"08",
           539 => x"51",
           540 => x"cb",
           541 => x"05",
           542 => x"cb",
           543 => x"05",
           544 => x"cb",
           545 => x"05",
           546 => x"a4",
           547 => x"0d",
           548 => x"0c",
           549 => x"0d",
           550 => x"02",
           551 => x"05",
           552 => x"53",
           553 => x"27",
           554 => x"83",
           555 => x"80",
           556 => x"ff",
           557 => x"ff",
           558 => x"73",
           559 => x"05",
           560 => x"12",
           561 => x"2e",
           562 => x"ef",
           563 => x"cb",
           564 => x"3d",
           565 => x"74",
           566 => x"07",
           567 => x"2b",
           568 => x"51",
           569 => x"a5",
           570 => x"70",
           571 => x"0c",
           572 => x"84",
           573 => x"72",
           574 => x"05",
           575 => x"71",
           576 => x"53",
           577 => x"52",
           578 => x"dd",
           579 => x"27",
           580 => x"71",
           581 => x"53",
           582 => x"52",
           583 => x"f2",
           584 => x"ff",
           585 => x"3d",
           586 => x"70",
           587 => x"06",
           588 => x"70",
           589 => x"73",
           590 => x"56",
           591 => x"08",
           592 => x"38",
           593 => x"52",
           594 => x"81",
           595 => x"54",
           596 => x"9d",
           597 => x"55",
           598 => x"09",
           599 => x"38",
           600 => x"14",
           601 => x"81",
           602 => x"56",
           603 => x"e5",
           604 => x"55",
           605 => x"06",
           606 => x"06",
           607 => x"81",
           608 => x"52",
           609 => x"0d",
           610 => x"70",
           611 => x"ff",
           612 => x"f8",
           613 => x"80",
           614 => x"51",
           615 => x"84",
           616 => x"71",
           617 => x"54",
           618 => x"2e",
           619 => x"75",
           620 => x"94",
           621 => x"81",
           622 => x"87",
           623 => x"fe",
           624 => x"52",
           625 => x"88",
           626 => x"86",
           627 => x"a4",
           628 => x"06",
           629 => x"14",
           630 => x"80",
           631 => x"71",
           632 => x"0c",
           633 => x"04",
           634 => x"77",
           635 => x"53",
           636 => x"80",
           637 => x"38",
           638 => x"70",
           639 => x"81",
           640 => x"81",
           641 => x"39",
           642 => x"39",
           643 => x"80",
           644 => x"81",
           645 => x"55",
           646 => x"2e",
           647 => x"55",
           648 => x"84",
           649 => x"38",
           650 => x"06",
           651 => x"2e",
           652 => x"88",
           653 => x"70",
           654 => x"34",
           655 => x"71",
           656 => x"cb",
           657 => x"3d",
           658 => x"3d",
           659 => x"72",
           660 => x"91",
           661 => x"fc",
           662 => x"51",
           663 => x"81",
           664 => x"85",
           665 => x"83",
           666 => x"72",
           667 => x"0c",
           668 => x"04",
           669 => x"76",
           670 => x"ff",
           671 => x"81",
           672 => x"26",
           673 => x"83",
           674 => x"05",
           675 => x"70",
           676 => x"8a",
           677 => x"33",
           678 => x"70",
           679 => x"fe",
           680 => x"33",
           681 => x"70",
           682 => x"f2",
           683 => x"33",
           684 => x"70",
           685 => x"e6",
           686 => x"22",
           687 => x"74",
           688 => x"80",
           689 => x"13",
           690 => x"52",
           691 => x"26",
           692 => x"81",
           693 => x"98",
           694 => x"22",
           695 => x"bc",
           696 => x"33",
           697 => x"b8",
           698 => x"33",
           699 => x"b4",
           700 => x"33",
           701 => x"b0",
           702 => x"33",
           703 => x"ac",
           704 => x"33",
           705 => x"a8",
           706 => x"c0",
           707 => x"73",
           708 => x"a0",
           709 => x"87",
           710 => x"0c",
           711 => x"81",
           712 => x"86",
           713 => x"f3",
           714 => x"5b",
           715 => x"9c",
           716 => x"0c",
           717 => x"bc",
           718 => x"7b",
           719 => x"98",
           720 => x"79",
           721 => x"87",
           722 => x"08",
           723 => x"1c",
           724 => x"98",
           725 => x"79",
           726 => x"87",
           727 => x"08",
           728 => x"1c",
           729 => x"98",
           730 => x"79",
           731 => x"87",
           732 => x"08",
           733 => x"1c",
           734 => x"98",
           735 => x"79",
           736 => x"80",
           737 => x"83",
           738 => x"59",
           739 => x"ff",
           740 => x"1b",
           741 => x"1b",
           742 => x"1b",
           743 => x"1b",
           744 => x"1b",
           745 => x"83",
           746 => x"52",
           747 => x"51",
           748 => x"8f",
           749 => x"ff",
           750 => x"8f",
           751 => x"30",
           752 => x"51",
           753 => x"0b",
           754 => x"8c",
           755 => x"0d",
           756 => x"0d",
           757 => x"81",
           758 => x"70",
           759 => x"57",
           760 => x"c0",
           761 => x"74",
           762 => x"38",
           763 => x"94",
           764 => x"70",
           765 => x"81",
           766 => x"52",
           767 => x"8c",
           768 => x"2a",
           769 => x"51",
           770 => x"38",
           771 => x"70",
           772 => x"51",
           773 => x"8d",
           774 => x"2a",
           775 => x"51",
           776 => x"be",
           777 => x"ff",
           778 => x"c0",
           779 => x"70",
           780 => x"38",
           781 => x"90",
           782 => x"0c",
           783 => x"a4",
           784 => x"0d",
           785 => x"0d",
           786 => x"33",
           787 => x"c8",
           788 => x"81",
           789 => x"55",
           790 => x"94",
           791 => x"80",
           792 => x"87",
           793 => x"51",
           794 => x"96",
           795 => x"06",
           796 => x"70",
           797 => x"38",
           798 => x"70",
           799 => x"51",
           800 => x"72",
           801 => x"81",
           802 => x"70",
           803 => x"38",
           804 => x"70",
           805 => x"51",
           806 => x"38",
           807 => x"06",
           808 => x"94",
           809 => x"80",
           810 => x"87",
           811 => x"52",
           812 => x"87",
           813 => x"f9",
           814 => x"54",
           815 => x"70",
           816 => x"53",
           817 => x"77",
           818 => x"38",
           819 => x"06",
           820 => x"0b",
           821 => x"33",
           822 => x"06",
           823 => x"58",
           824 => x"84",
           825 => x"2e",
           826 => x"c0",
           827 => x"70",
           828 => x"2a",
           829 => x"53",
           830 => x"80",
           831 => x"71",
           832 => x"81",
           833 => x"70",
           834 => x"81",
           835 => x"06",
           836 => x"80",
           837 => x"71",
           838 => x"81",
           839 => x"70",
           840 => x"74",
           841 => x"51",
           842 => x"80",
           843 => x"2e",
           844 => x"c0",
           845 => x"77",
           846 => x"17",
           847 => x"81",
           848 => x"53",
           849 => x"84",
           850 => x"cb",
           851 => x"3d",
           852 => x"3d",
           853 => x"81",
           854 => x"70",
           855 => x"54",
           856 => x"94",
           857 => x"80",
           858 => x"87",
           859 => x"51",
           860 => x"82",
           861 => x"06",
           862 => x"70",
           863 => x"38",
           864 => x"06",
           865 => x"94",
           866 => x"80",
           867 => x"87",
           868 => x"52",
           869 => x"81",
           870 => x"cb",
           871 => x"84",
           872 => x"fe",
           873 => x"0b",
           874 => x"33",
           875 => x"06",
           876 => x"c0",
           877 => x"70",
           878 => x"38",
           879 => x"94",
           880 => x"70",
           881 => x"81",
           882 => x"51",
           883 => x"80",
           884 => x"72",
           885 => x"51",
           886 => x"80",
           887 => x"2e",
           888 => x"c0",
           889 => x"71",
           890 => x"2b",
           891 => x"51",
           892 => x"81",
           893 => x"84",
           894 => x"ff",
           895 => x"c0",
           896 => x"70",
           897 => x"06",
           898 => x"80",
           899 => x"38",
           900 => x"9c",
           901 => x"90",
           902 => x"9e",
           903 => x"c8",
           904 => x"c0",
           905 => x"81",
           906 => x"87",
           907 => x"08",
           908 => x"0c",
           909 => x"94",
           910 => x"a0",
           911 => x"9e",
           912 => x"c8",
           913 => x"c0",
           914 => x"81",
           915 => x"87",
           916 => x"08",
           917 => x"0c",
           918 => x"ac",
           919 => x"b0",
           920 => x"9e",
           921 => x"70",
           922 => x"23",
           923 => x"84",
           924 => x"b8",
           925 => x"81",
           926 => x"80",
           927 => x"9e",
           928 => x"a0",
           929 => x"52",
           930 => x"2e",
           931 => x"52",
           932 => x"bd",
           933 => x"87",
           934 => x"08",
           935 => x"80",
           936 => x"52",
           937 => x"83",
           938 => x"71",
           939 => x"34",
           940 => x"c0",
           941 => x"70",
           942 => x"06",
           943 => x"70",
           944 => x"38",
           945 => x"81",
           946 => x"80",
           947 => x"9e",
           948 => x"90",
           949 => x"52",
           950 => x"2e",
           951 => x"52",
           952 => x"c0",
           953 => x"87",
           954 => x"08",
           955 => x"06",
           956 => x"70",
           957 => x"38",
           958 => x"81",
           959 => x"80",
           960 => x"9e",
           961 => x"84",
           962 => x"52",
           963 => x"2e",
           964 => x"52",
           965 => x"c2",
           966 => x"87",
           967 => x"08",
           968 => x"06",
           969 => x"70",
           970 => x"38",
           971 => x"81",
           972 => x"80",
           973 => x"9e",
           974 => x"81",
           975 => x"52",
           976 => x"2e",
           977 => x"52",
           978 => x"c4",
           979 => x"9e",
           980 => x"80",
           981 => x"86",
           982 => x"51",
           983 => x"c5",
           984 => x"87",
           985 => x"08",
           986 => x"51",
           987 => x"80",
           988 => x"81",
           989 => x"c8",
           990 => x"0b",
           991 => x"88",
           992 => x"06",
           993 => x"70",
           994 => x"38",
           995 => x"81",
           996 => x"87",
           997 => x"08",
           998 => x"51",
           999 => x"c8",
          1000 => x"3d",
          1001 => x"3d",
          1002 => x"f0",
          1003 => x"3f",
          1004 => x"33",
          1005 => x"2e",
          1006 => x"b6",
          1007 => x"92",
          1008 => x"98",
          1009 => x"3f",
          1010 => x"33",
          1011 => x"2e",
          1012 => x"c8",
          1013 => x"81",
          1014 => x"52",
          1015 => x"51",
          1016 => x"81",
          1017 => x"54",
          1018 => x"92",
          1019 => x"9c",
          1020 => x"c8",
          1021 => x"81",
          1022 => x"89",
          1023 => x"c8",
          1024 => x"73",
          1025 => x"c8",
          1026 => x"73",
          1027 => x"38",
          1028 => x"08",
          1029 => x"a0",
          1030 => x"b6",
          1031 => x"96",
          1032 => x"c1",
          1033 => x"80",
          1034 => x"81",
          1035 => x"83",
          1036 => x"c8",
          1037 => x"73",
          1038 => x"38",
          1039 => x"51",
          1040 => x"81",
          1041 => x"54",
          1042 => x"88",
          1043 => x"b8",
          1044 => x"3f",
          1045 => x"33",
          1046 => x"2e",
          1047 => x"c8",
          1048 => x"81",
          1049 => x"88",
          1050 => x"c8",
          1051 => x"73",
          1052 => x"38",
          1053 => x"51",
          1054 => x"81",
          1055 => x"54",
          1056 => x"8d",
          1057 => x"c8",
          1058 => x"b8",
          1059 => x"a6",
          1060 => x"9c",
          1061 => x"3f",
          1062 => x"08",
          1063 => x"a8",
          1064 => x"3f",
          1065 => x"08",
          1066 => x"d0",
          1067 => x"3f",
          1068 => x"08",
          1069 => x"f8",
          1070 => x"3f",
          1071 => x"22",
          1072 => x"a0",
          1073 => x"3f",
          1074 => x"08",
          1075 => x"c8",
          1076 => x"3f",
          1077 => x"04",
          1078 => x"02",
          1079 => x"ff",
          1080 => x"84",
          1081 => x"71",
          1082 => x"0b",
          1083 => x"05",
          1084 => x"04",
          1085 => x"51",
          1086 => x"b9",
          1087 => x"39",
          1088 => x"51",
          1089 => x"ba",
          1090 => x"39",
          1091 => x"51",
          1092 => x"ba",
          1093 => x"9f",
          1094 => x"0d",
          1095 => x"80",
          1096 => x"0b",
          1097 => x"84",
          1098 => x"3d",
          1099 => x"96",
          1100 => x"52",
          1101 => x"0c",
          1102 => x"70",
          1103 => x"0c",
          1104 => x"3d",
          1105 => x"3d",
          1106 => x"96",
          1107 => x"81",
          1108 => x"52",
          1109 => x"73",
          1110 => x"c8",
          1111 => x"70",
          1112 => x"0c",
          1113 => x"83",
          1114 => x"81",
          1115 => x"87",
          1116 => x"0c",
          1117 => x"0d",
          1118 => x"33",
          1119 => x"2e",
          1120 => x"85",
          1121 => x"ed",
          1122 => x"bc",
          1123 => x"80",
          1124 => x"72",
          1125 => x"cb",
          1126 => x"05",
          1127 => x"0c",
          1128 => x"cb",
          1129 => x"71",
          1130 => x"38",
          1131 => x"2d",
          1132 => x"04",
          1133 => x"02",
          1134 => x"81",
          1135 => x"76",
          1136 => x"0c",
          1137 => x"ad",
          1138 => x"cb",
          1139 => x"3d",
          1140 => x"3d",
          1141 => x"73",
          1142 => x"ff",
          1143 => x"71",
          1144 => x"38",
          1145 => x"06",
          1146 => x"54",
          1147 => x"e7",
          1148 => x"0d",
          1149 => x"0d",
          1150 => x"b4",
          1151 => x"cb",
          1152 => x"54",
          1153 => x"81",
          1154 => x"53",
          1155 => x"8e",
          1156 => x"ff",
          1157 => x"14",
          1158 => x"3f",
          1159 => x"81",
          1160 => x"86",
          1161 => x"ec",
          1162 => x"68",
          1163 => x"70",
          1164 => x"33",
          1165 => x"2e",
          1166 => x"75",
          1167 => x"81",
          1168 => x"38",
          1169 => x"70",
          1170 => x"33",
          1171 => x"75",
          1172 => x"81",
          1173 => x"81",
          1174 => x"75",
          1175 => x"81",
          1176 => x"82",
          1177 => x"81",
          1178 => x"56",
          1179 => x"09",
          1180 => x"38",
          1181 => x"71",
          1182 => x"81",
          1183 => x"59",
          1184 => x"9d",
          1185 => x"53",
          1186 => x"95",
          1187 => x"29",
          1188 => x"76",
          1189 => x"79",
          1190 => x"5b",
          1191 => x"e5",
          1192 => x"ec",
          1193 => x"70",
          1194 => x"25",
          1195 => x"32",
          1196 => x"72",
          1197 => x"73",
          1198 => x"58",
          1199 => x"73",
          1200 => x"38",
          1201 => x"79",
          1202 => x"5b",
          1203 => x"75",
          1204 => x"de",
          1205 => x"80",
          1206 => x"89",
          1207 => x"70",
          1208 => x"55",
          1209 => x"cf",
          1210 => x"38",
          1211 => x"24",
          1212 => x"80",
          1213 => x"8e",
          1214 => x"c3",
          1215 => x"73",
          1216 => x"81",
          1217 => x"99",
          1218 => x"c4",
          1219 => x"38",
          1220 => x"73",
          1221 => x"81",
          1222 => x"80",
          1223 => x"38",
          1224 => x"2e",
          1225 => x"f9",
          1226 => x"d8",
          1227 => x"38",
          1228 => x"77",
          1229 => x"08",
          1230 => x"80",
          1231 => x"55",
          1232 => x"8d",
          1233 => x"70",
          1234 => x"51",
          1235 => x"f5",
          1236 => x"2a",
          1237 => x"74",
          1238 => x"53",
          1239 => x"8f",
          1240 => x"fc",
          1241 => x"81",
          1242 => x"80",
          1243 => x"73",
          1244 => x"3f",
          1245 => x"56",
          1246 => x"27",
          1247 => x"a0",
          1248 => x"3f",
          1249 => x"84",
          1250 => x"33",
          1251 => x"93",
          1252 => x"95",
          1253 => x"91",
          1254 => x"8d",
          1255 => x"89",
          1256 => x"fb",
          1257 => x"86",
          1258 => x"2a",
          1259 => x"51",
          1260 => x"2e",
          1261 => x"84",
          1262 => x"86",
          1263 => x"78",
          1264 => x"08",
          1265 => x"32",
          1266 => x"72",
          1267 => x"51",
          1268 => x"74",
          1269 => x"38",
          1270 => x"88",
          1271 => x"7a",
          1272 => x"55",
          1273 => x"3d",
          1274 => x"52",
          1275 => x"e0",
          1276 => x"a4",
          1277 => x"06",
          1278 => x"52",
          1279 => x"3f",
          1280 => x"08",
          1281 => x"27",
          1282 => x"14",
          1283 => x"f8",
          1284 => x"87",
          1285 => x"81",
          1286 => x"b0",
          1287 => x"7d",
          1288 => x"5f",
          1289 => x"75",
          1290 => x"07",
          1291 => x"54",
          1292 => x"26",
          1293 => x"ff",
          1294 => x"84",
          1295 => x"06",
          1296 => x"80",
          1297 => x"96",
          1298 => x"e0",
          1299 => x"73",
          1300 => x"57",
          1301 => x"06",
          1302 => x"54",
          1303 => x"a0",
          1304 => x"2a",
          1305 => x"54",
          1306 => x"38",
          1307 => x"76",
          1308 => x"38",
          1309 => x"fd",
          1310 => x"06",
          1311 => x"38",
          1312 => x"56",
          1313 => x"26",
          1314 => x"3d",
          1315 => x"05",
          1316 => x"ff",
          1317 => x"53",
          1318 => x"d9",
          1319 => x"38",
          1320 => x"56",
          1321 => x"27",
          1322 => x"a0",
          1323 => x"3f",
          1324 => x"3d",
          1325 => x"3d",
          1326 => x"70",
          1327 => x"52",
          1328 => x"73",
          1329 => x"3f",
          1330 => x"04",
          1331 => x"74",
          1332 => x"0c",
          1333 => x"05",
          1334 => x"fa",
          1335 => x"cb",
          1336 => x"80",
          1337 => x"0b",
          1338 => x"0c",
          1339 => x"04",
          1340 => x"81",
          1341 => x"76",
          1342 => x"0c",
          1343 => x"05",
          1344 => x"53",
          1345 => x"72",
          1346 => x"0c",
          1347 => x"04",
          1348 => x"77",
          1349 => x"b8",
          1350 => x"54",
          1351 => x"54",
          1352 => x"80",
          1353 => x"cb",
          1354 => x"71",
          1355 => x"a4",
          1356 => x"06",
          1357 => x"2e",
          1358 => x"72",
          1359 => x"38",
          1360 => x"70",
          1361 => x"25",
          1362 => x"73",
          1363 => x"38",
          1364 => x"86",
          1365 => x"54",
          1366 => x"73",
          1367 => x"ff",
          1368 => x"72",
          1369 => x"74",
          1370 => x"72",
          1371 => x"54",
          1372 => x"81",
          1373 => x"39",
          1374 => x"80",
          1375 => x"51",
          1376 => x"81",
          1377 => x"cb",
          1378 => x"3d",
          1379 => x"3d",
          1380 => x"b8",
          1381 => x"cb",
          1382 => x"53",
          1383 => x"fe",
          1384 => x"81",
          1385 => x"84",
          1386 => x"f8",
          1387 => x"7c",
          1388 => x"70",
          1389 => x"75",
          1390 => x"55",
          1391 => x"2e",
          1392 => x"87",
          1393 => x"76",
          1394 => x"73",
          1395 => x"81",
          1396 => x"81",
          1397 => x"77",
          1398 => x"70",
          1399 => x"58",
          1400 => x"09",
          1401 => x"c2",
          1402 => x"81",
          1403 => x"75",
          1404 => x"55",
          1405 => x"e2",
          1406 => x"90",
          1407 => x"f8",
          1408 => x"8f",
          1409 => x"81",
          1410 => x"75",
          1411 => x"55",
          1412 => x"81",
          1413 => x"27",
          1414 => x"d0",
          1415 => x"55",
          1416 => x"73",
          1417 => x"80",
          1418 => x"14",
          1419 => x"72",
          1420 => x"e0",
          1421 => x"80",
          1422 => x"39",
          1423 => x"55",
          1424 => x"80",
          1425 => x"e0",
          1426 => x"38",
          1427 => x"81",
          1428 => x"53",
          1429 => x"81",
          1430 => x"53",
          1431 => x"8e",
          1432 => x"70",
          1433 => x"55",
          1434 => x"27",
          1435 => x"77",
          1436 => x"74",
          1437 => x"76",
          1438 => x"77",
          1439 => x"70",
          1440 => x"55",
          1441 => x"77",
          1442 => x"38",
          1443 => x"74",
          1444 => x"55",
          1445 => x"a4",
          1446 => x"0d",
          1447 => x"0d",
          1448 => x"56",
          1449 => x"0c",
          1450 => x"70",
          1451 => x"73",
          1452 => x"81",
          1453 => x"81",
          1454 => x"ed",
          1455 => x"2e",
          1456 => x"8e",
          1457 => x"08",
          1458 => x"76",
          1459 => x"56",
          1460 => x"b0",
          1461 => x"06",
          1462 => x"75",
          1463 => x"76",
          1464 => x"70",
          1465 => x"73",
          1466 => x"8b",
          1467 => x"73",
          1468 => x"85",
          1469 => x"82",
          1470 => x"76",
          1471 => x"70",
          1472 => x"ac",
          1473 => x"a0",
          1474 => x"fa",
          1475 => x"53",
          1476 => x"57",
          1477 => x"98",
          1478 => x"39",
          1479 => x"80",
          1480 => x"26",
          1481 => x"86",
          1482 => x"80",
          1483 => x"57",
          1484 => x"74",
          1485 => x"38",
          1486 => x"27",
          1487 => x"14",
          1488 => x"06",
          1489 => x"14",
          1490 => x"06",
          1491 => x"74",
          1492 => x"f9",
          1493 => x"ff",
          1494 => x"89",
          1495 => x"38",
          1496 => x"c5",
          1497 => x"29",
          1498 => x"81",
          1499 => x"76",
          1500 => x"56",
          1501 => x"ba",
          1502 => x"2e",
          1503 => x"30",
          1504 => x"0c",
          1505 => x"81",
          1506 => x"8a",
          1507 => x"ff",
          1508 => x"8f",
          1509 => x"81",
          1510 => x"26",
          1511 => x"c8",
          1512 => x"52",
          1513 => x"a4",
          1514 => x"0d",
          1515 => x"0d",
          1516 => x"33",
          1517 => x"9f",
          1518 => x"53",
          1519 => x"81",
          1520 => x"38",
          1521 => x"87",
          1522 => x"11",
          1523 => x"54",
          1524 => x"84",
          1525 => x"54",
          1526 => x"87",
          1527 => x"11",
          1528 => x"0c",
          1529 => x"c0",
          1530 => x"70",
          1531 => x"70",
          1532 => x"51",
          1533 => x"8a",
          1534 => x"98",
          1535 => x"70",
          1536 => x"08",
          1537 => x"06",
          1538 => x"38",
          1539 => x"8c",
          1540 => x"80",
          1541 => x"71",
          1542 => x"14",
          1543 => x"d0",
          1544 => x"70",
          1545 => x"0c",
          1546 => x"04",
          1547 => x"60",
          1548 => x"8c",
          1549 => x"33",
          1550 => x"5b",
          1551 => x"5a",
          1552 => x"81",
          1553 => x"81",
          1554 => x"52",
          1555 => x"38",
          1556 => x"84",
          1557 => x"92",
          1558 => x"c0",
          1559 => x"87",
          1560 => x"13",
          1561 => x"57",
          1562 => x"0b",
          1563 => x"8c",
          1564 => x"0c",
          1565 => x"75",
          1566 => x"2a",
          1567 => x"51",
          1568 => x"80",
          1569 => x"7b",
          1570 => x"7b",
          1571 => x"5d",
          1572 => x"59",
          1573 => x"06",
          1574 => x"73",
          1575 => x"81",
          1576 => x"ff",
          1577 => x"72",
          1578 => x"38",
          1579 => x"8c",
          1580 => x"c3",
          1581 => x"98",
          1582 => x"71",
          1583 => x"38",
          1584 => x"2e",
          1585 => x"76",
          1586 => x"92",
          1587 => x"72",
          1588 => x"06",
          1589 => x"f7",
          1590 => x"5a",
          1591 => x"80",
          1592 => x"70",
          1593 => x"5a",
          1594 => x"80",
          1595 => x"73",
          1596 => x"06",
          1597 => x"38",
          1598 => x"fe",
          1599 => x"fc",
          1600 => x"52",
          1601 => x"83",
          1602 => x"71",
          1603 => x"cb",
          1604 => x"3d",
          1605 => x"3d",
          1606 => x"64",
          1607 => x"bf",
          1608 => x"40",
          1609 => x"59",
          1610 => x"58",
          1611 => x"81",
          1612 => x"81",
          1613 => x"52",
          1614 => x"09",
          1615 => x"b1",
          1616 => x"84",
          1617 => x"92",
          1618 => x"c0",
          1619 => x"87",
          1620 => x"13",
          1621 => x"56",
          1622 => x"87",
          1623 => x"0c",
          1624 => x"82",
          1625 => x"58",
          1626 => x"84",
          1627 => x"06",
          1628 => x"71",
          1629 => x"38",
          1630 => x"05",
          1631 => x"0c",
          1632 => x"73",
          1633 => x"81",
          1634 => x"71",
          1635 => x"38",
          1636 => x"8c",
          1637 => x"d0",
          1638 => x"98",
          1639 => x"71",
          1640 => x"38",
          1641 => x"2e",
          1642 => x"76",
          1643 => x"92",
          1644 => x"72",
          1645 => x"06",
          1646 => x"f7",
          1647 => x"59",
          1648 => x"1a",
          1649 => x"06",
          1650 => x"59",
          1651 => x"80",
          1652 => x"73",
          1653 => x"06",
          1654 => x"38",
          1655 => x"fe",
          1656 => x"fc",
          1657 => x"52",
          1658 => x"83",
          1659 => x"71",
          1660 => x"cb",
          1661 => x"3d",
          1662 => x"3d",
          1663 => x"84",
          1664 => x"33",
          1665 => x"b7",
          1666 => x"54",
          1667 => x"fa",
          1668 => x"cb",
          1669 => x"06",
          1670 => x"72",
          1671 => x"85",
          1672 => x"98",
          1673 => x"56",
          1674 => x"80",
          1675 => x"76",
          1676 => x"74",
          1677 => x"c0",
          1678 => x"54",
          1679 => x"2e",
          1680 => x"d4",
          1681 => x"2e",
          1682 => x"80",
          1683 => x"08",
          1684 => x"70",
          1685 => x"51",
          1686 => x"2e",
          1687 => x"c0",
          1688 => x"52",
          1689 => x"87",
          1690 => x"08",
          1691 => x"38",
          1692 => x"87",
          1693 => x"14",
          1694 => x"70",
          1695 => x"52",
          1696 => x"96",
          1697 => x"92",
          1698 => x"0a",
          1699 => x"39",
          1700 => x"0c",
          1701 => x"39",
          1702 => x"54",
          1703 => x"a4",
          1704 => x"0d",
          1705 => x"0d",
          1706 => x"33",
          1707 => x"88",
          1708 => x"cb",
          1709 => x"51",
          1710 => x"04",
          1711 => x"75",
          1712 => x"82",
          1713 => x"90",
          1714 => x"2b",
          1715 => x"33",
          1716 => x"88",
          1717 => x"71",
          1718 => x"a4",
          1719 => x"54",
          1720 => x"85",
          1721 => x"ff",
          1722 => x"02",
          1723 => x"05",
          1724 => x"70",
          1725 => x"05",
          1726 => x"88",
          1727 => x"72",
          1728 => x"0d",
          1729 => x"0d",
          1730 => x"52",
          1731 => x"81",
          1732 => x"70",
          1733 => x"70",
          1734 => x"05",
          1735 => x"88",
          1736 => x"72",
          1737 => x"54",
          1738 => x"2a",
          1739 => x"34",
          1740 => x"04",
          1741 => x"76",
          1742 => x"54",
          1743 => x"2e",
          1744 => x"70",
          1745 => x"33",
          1746 => x"05",
          1747 => x"11",
          1748 => x"84",
          1749 => x"fe",
          1750 => x"77",
          1751 => x"53",
          1752 => x"81",
          1753 => x"ff",
          1754 => x"f4",
          1755 => x"0d",
          1756 => x"0d",
          1757 => x"56",
          1758 => x"70",
          1759 => x"33",
          1760 => x"05",
          1761 => x"71",
          1762 => x"56",
          1763 => x"72",
          1764 => x"38",
          1765 => x"e2",
          1766 => x"cb",
          1767 => x"3d",
          1768 => x"3d",
          1769 => x"54",
          1770 => x"71",
          1771 => x"38",
          1772 => x"70",
          1773 => x"f3",
          1774 => x"81",
          1775 => x"84",
          1776 => x"80",
          1777 => x"a4",
          1778 => x"0b",
          1779 => x"0c",
          1780 => x"0d",
          1781 => x"0b",
          1782 => x"56",
          1783 => x"2e",
          1784 => x"81",
          1785 => x"08",
          1786 => x"70",
          1787 => x"33",
          1788 => x"a2",
          1789 => x"a4",
          1790 => x"09",
          1791 => x"38",
          1792 => x"08",
          1793 => x"b0",
          1794 => x"a4",
          1795 => x"9c",
          1796 => x"56",
          1797 => x"27",
          1798 => x"16",
          1799 => x"82",
          1800 => x"06",
          1801 => x"54",
          1802 => x"78",
          1803 => x"33",
          1804 => x"3f",
          1805 => x"5a",
          1806 => x"a4",
          1807 => x"0d",
          1808 => x"0d",
          1809 => x"56",
          1810 => x"b0",
          1811 => x"af",
          1812 => x"fe",
          1813 => x"cb",
          1814 => x"81",
          1815 => x"9f",
          1816 => x"74",
          1817 => x"52",
          1818 => x"51",
          1819 => x"81",
          1820 => x"80",
          1821 => x"ff",
          1822 => x"74",
          1823 => x"76",
          1824 => x"0c",
          1825 => x"04",
          1826 => x"7a",
          1827 => x"fe",
          1828 => x"cb",
          1829 => x"81",
          1830 => x"81",
          1831 => x"33",
          1832 => x"2e",
          1833 => x"80",
          1834 => x"17",
          1835 => x"81",
          1836 => x"06",
          1837 => x"84",
          1838 => x"cb",
          1839 => x"b4",
          1840 => x"56",
          1841 => x"82",
          1842 => x"84",
          1843 => x"fc",
          1844 => x"8b",
          1845 => x"52",
          1846 => x"a9",
          1847 => x"85",
          1848 => x"84",
          1849 => x"fc",
          1850 => x"17",
          1851 => x"9c",
          1852 => x"91",
          1853 => x"08",
          1854 => x"17",
          1855 => x"3f",
          1856 => x"81",
          1857 => x"19",
          1858 => x"53",
          1859 => x"17",
          1860 => x"82",
          1861 => x"18",
          1862 => x"80",
          1863 => x"33",
          1864 => x"3f",
          1865 => x"08",
          1866 => x"38",
          1867 => x"81",
          1868 => x"8a",
          1869 => x"fb",
          1870 => x"fe",
          1871 => x"08",
          1872 => x"56",
          1873 => x"74",
          1874 => x"38",
          1875 => x"75",
          1876 => x"16",
          1877 => x"53",
          1878 => x"a4",
          1879 => x"0d",
          1880 => x"0d",
          1881 => x"08",
          1882 => x"81",
          1883 => x"df",
          1884 => x"15",
          1885 => x"d7",
          1886 => x"33",
          1887 => x"82",
          1888 => x"38",
          1889 => x"89",
          1890 => x"2e",
          1891 => x"bf",
          1892 => x"2e",
          1893 => x"81",
          1894 => x"81",
          1895 => x"89",
          1896 => x"08",
          1897 => x"52",
          1898 => x"3f",
          1899 => x"08",
          1900 => x"74",
          1901 => x"14",
          1902 => x"81",
          1903 => x"2a",
          1904 => x"05",
          1905 => x"57",
          1906 => x"f5",
          1907 => x"a4",
          1908 => x"38",
          1909 => x"06",
          1910 => x"33",
          1911 => x"78",
          1912 => x"06",
          1913 => x"5c",
          1914 => x"53",
          1915 => x"38",
          1916 => x"06",
          1917 => x"39",
          1918 => x"a4",
          1919 => x"52",
          1920 => x"bd",
          1921 => x"a4",
          1922 => x"38",
          1923 => x"fe",
          1924 => x"b4",
          1925 => x"8d",
          1926 => x"a4",
          1927 => x"ff",
          1928 => x"39",
          1929 => x"a4",
          1930 => x"52",
          1931 => x"91",
          1932 => x"a4",
          1933 => x"76",
          1934 => x"fc",
          1935 => x"b4",
          1936 => x"f8",
          1937 => x"a4",
          1938 => x"06",
          1939 => x"81",
          1940 => x"cb",
          1941 => x"3d",
          1942 => x"3d",
          1943 => x"7e",
          1944 => x"82",
          1945 => x"27",
          1946 => x"76",
          1947 => x"27",
          1948 => x"75",
          1949 => x"79",
          1950 => x"38",
          1951 => x"89",
          1952 => x"2e",
          1953 => x"80",
          1954 => x"2e",
          1955 => x"81",
          1956 => x"81",
          1957 => x"89",
          1958 => x"08",
          1959 => x"52",
          1960 => x"3f",
          1961 => x"08",
          1962 => x"a4",
          1963 => x"38",
          1964 => x"06",
          1965 => x"81",
          1966 => x"06",
          1967 => x"77",
          1968 => x"2e",
          1969 => x"84",
          1970 => x"06",
          1971 => x"06",
          1972 => x"53",
          1973 => x"81",
          1974 => x"34",
          1975 => x"a4",
          1976 => x"52",
          1977 => x"d9",
          1978 => x"a4",
          1979 => x"cb",
          1980 => x"94",
          1981 => x"ff",
          1982 => x"05",
          1983 => x"54",
          1984 => x"38",
          1985 => x"74",
          1986 => x"06",
          1987 => x"07",
          1988 => x"74",
          1989 => x"39",
          1990 => x"a4",
          1991 => x"52",
          1992 => x"9d",
          1993 => x"a4",
          1994 => x"cb",
          1995 => x"d8",
          1996 => x"ff",
          1997 => x"76",
          1998 => x"06",
          1999 => x"05",
          2000 => x"3f",
          2001 => x"87",
          2002 => x"08",
          2003 => x"51",
          2004 => x"81",
          2005 => x"59",
          2006 => x"08",
          2007 => x"f0",
          2008 => x"82",
          2009 => x"06",
          2010 => x"05",
          2011 => x"54",
          2012 => x"3f",
          2013 => x"08",
          2014 => x"74",
          2015 => x"51",
          2016 => x"81",
          2017 => x"34",
          2018 => x"a4",
          2019 => x"0d",
          2020 => x"0d",
          2021 => x"72",
          2022 => x"56",
          2023 => x"27",
          2024 => x"98",
          2025 => x"9d",
          2026 => x"2e",
          2027 => x"53",
          2028 => x"51",
          2029 => x"81",
          2030 => x"54",
          2031 => x"08",
          2032 => x"93",
          2033 => x"80",
          2034 => x"54",
          2035 => x"81",
          2036 => x"54",
          2037 => x"74",
          2038 => x"fb",
          2039 => x"cb",
          2040 => x"81",
          2041 => x"80",
          2042 => x"38",
          2043 => x"08",
          2044 => x"38",
          2045 => x"08",
          2046 => x"38",
          2047 => x"52",
          2048 => x"d6",
          2049 => x"a4",
          2050 => x"98",
          2051 => x"11",
          2052 => x"57",
          2053 => x"74",
          2054 => x"81",
          2055 => x"0c",
          2056 => x"81",
          2057 => x"84",
          2058 => x"55",
          2059 => x"ff",
          2060 => x"54",
          2061 => x"a4",
          2062 => x"0d",
          2063 => x"0d",
          2064 => x"08",
          2065 => x"79",
          2066 => x"17",
          2067 => x"80",
          2068 => x"98",
          2069 => x"26",
          2070 => x"58",
          2071 => x"52",
          2072 => x"fd",
          2073 => x"74",
          2074 => x"08",
          2075 => x"38",
          2076 => x"08",
          2077 => x"a4",
          2078 => x"82",
          2079 => x"17",
          2080 => x"a4",
          2081 => x"c7",
          2082 => x"90",
          2083 => x"56",
          2084 => x"2e",
          2085 => x"77",
          2086 => x"81",
          2087 => x"38",
          2088 => x"98",
          2089 => x"26",
          2090 => x"56",
          2091 => x"51",
          2092 => x"80",
          2093 => x"a4",
          2094 => x"09",
          2095 => x"38",
          2096 => x"08",
          2097 => x"a4",
          2098 => x"30",
          2099 => x"80",
          2100 => x"07",
          2101 => x"08",
          2102 => x"55",
          2103 => x"ef",
          2104 => x"a4",
          2105 => x"95",
          2106 => x"08",
          2107 => x"27",
          2108 => x"98",
          2109 => x"89",
          2110 => x"85",
          2111 => x"db",
          2112 => x"81",
          2113 => x"17",
          2114 => x"89",
          2115 => x"75",
          2116 => x"ac",
          2117 => x"7a",
          2118 => x"3f",
          2119 => x"08",
          2120 => x"38",
          2121 => x"cb",
          2122 => x"2e",
          2123 => x"86",
          2124 => x"a4",
          2125 => x"cb",
          2126 => x"70",
          2127 => x"07",
          2128 => x"7c",
          2129 => x"55",
          2130 => x"f8",
          2131 => x"2e",
          2132 => x"ff",
          2133 => x"55",
          2134 => x"ff",
          2135 => x"76",
          2136 => x"3f",
          2137 => x"08",
          2138 => x"08",
          2139 => x"cb",
          2140 => x"80",
          2141 => x"55",
          2142 => x"94",
          2143 => x"2e",
          2144 => x"53",
          2145 => x"51",
          2146 => x"81",
          2147 => x"55",
          2148 => x"75",
          2149 => x"98",
          2150 => x"05",
          2151 => x"56",
          2152 => x"26",
          2153 => x"15",
          2154 => x"84",
          2155 => x"07",
          2156 => x"18",
          2157 => x"ff",
          2158 => x"2e",
          2159 => x"39",
          2160 => x"39",
          2161 => x"08",
          2162 => x"81",
          2163 => x"74",
          2164 => x"0c",
          2165 => x"04",
          2166 => x"7a",
          2167 => x"f3",
          2168 => x"cb",
          2169 => x"81",
          2170 => x"a4",
          2171 => x"38",
          2172 => x"51",
          2173 => x"81",
          2174 => x"81",
          2175 => x"b0",
          2176 => x"84",
          2177 => x"52",
          2178 => x"52",
          2179 => x"3f",
          2180 => x"39",
          2181 => x"8a",
          2182 => x"75",
          2183 => x"38",
          2184 => x"19",
          2185 => x"81",
          2186 => x"ed",
          2187 => x"cb",
          2188 => x"2e",
          2189 => x"15",
          2190 => x"70",
          2191 => x"07",
          2192 => x"53",
          2193 => x"75",
          2194 => x"0c",
          2195 => x"04",
          2196 => x"7a",
          2197 => x"58",
          2198 => x"f0",
          2199 => x"80",
          2200 => x"9f",
          2201 => x"80",
          2202 => x"90",
          2203 => x"17",
          2204 => x"aa",
          2205 => x"53",
          2206 => x"88",
          2207 => x"08",
          2208 => x"38",
          2209 => x"53",
          2210 => x"17",
          2211 => x"72",
          2212 => x"fe",
          2213 => x"08",
          2214 => x"80",
          2215 => x"16",
          2216 => x"2b",
          2217 => x"75",
          2218 => x"73",
          2219 => x"f5",
          2220 => x"cb",
          2221 => x"81",
          2222 => x"ff",
          2223 => x"81",
          2224 => x"a4",
          2225 => x"38",
          2226 => x"81",
          2227 => x"26",
          2228 => x"58",
          2229 => x"73",
          2230 => x"39",
          2231 => x"51",
          2232 => x"81",
          2233 => x"98",
          2234 => x"94",
          2235 => x"17",
          2236 => x"58",
          2237 => x"9a",
          2238 => x"81",
          2239 => x"74",
          2240 => x"98",
          2241 => x"83",
          2242 => x"b4",
          2243 => x"0c",
          2244 => x"81",
          2245 => x"8a",
          2246 => x"f8",
          2247 => x"70",
          2248 => x"08",
          2249 => x"57",
          2250 => x"0a",
          2251 => x"38",
          2252 => x"15",
          2253 => x"08",
          2254 => x"72",
          2255 => x"cb",
          2256 => x"ff",
          2257 => x"81",
          2258 => x"13",
          2259 => x"94",
          2260 => x"74",
          2261 => x"85",
          2262 => x"22",
          2263 => x"73",
          2264 => x"38",
          2265 => x"8a",
          2266 => x"05",
          2267 => x"06",
          2268 => x"8a",
          2269 => x"73",
          2270 => x"3f",
          2271 => x"08",
          2272 => x"81",
          2273 => x"a4",
          2274 => x"ff",
          2275 => x"81",
          2276 => x"ff",
          2277 => x"38",
          2278 => x"81",
          2279 => x"26",
          2280 => x"7b",
          2281 => x"98",
          2282 => x"55",
          2283 => x"94",
          2284 => x"73",
          2285 => x"3f",
          2286 => x"08",
          2287 => x"81",
          2288 => x"80",
          2289 => x"38",
          2290 => x"cb",
          2291 => x"2e",
          2292 => x"55",
          2293 => x"08",
          2294 => x"38",
          2295 => x"08",
          2296 => x"fb",
          2297 => x"cb",
          2298 => x"38",
          2299 => x"0c",
          2300 => x"51",
          2301 => x"81",
          2302 => x"98",
          2303 => x"90",
          2304 => x"16",
          2305 => x"15",
          2306 => x"74",
          2307 => x"0c",
          2308 => x"04",
          2309 => x"7b",
          2310 => x"5b",
          2311 => x"52",
          2312 => x"ac",
          2313 => x"a4",
          2314 => x"cb",
          2315 => x"ec",
          2316 => x"a4",
          2317 => x"17",
          2318 => x"51",
          2319 => x"81",
          2320 => x"54",
          2321 => x"08",
          2322 => x"81",
          2323 => x"9c",
          2324 => x"33",
          2325 => x"72",
          2326 => x"09",
          2327 => x"38",
          2328 => x"cb",
          2329 => x"72",
          2330 => x"55",
          2331 => x"53",
          2332 => x"8e",
          2333 => x"56",
          2334 => x"09",
          2335 => x"38",
          2336 => x"cb",
          2337 => x"81",
          2338 => x"fd",
          2339 => x"cb",
          2340 => x"81",
          2341 => x"80",
          2342 => x"38",
          2343 => x"09",
          2344 => x"38",
          2345 => x"81",
          2346 => x"8b",
          2347 => x"fd",
          2348 => x"9a",
          2349 => x"eb",
          2350 => x"cb",
          2351 => x"ff",
          2352 => x"70",
          2353 => x"53",
          2354 => x"09",
          2355 => x"38",
          2356 => x"eb",
          2357 => x"cb",
          2358 => x"2b",
          2359 => x"72",
          2360 => x"0c",
          2361 => x"04",
          2362 => x"77",
          2363 => x"ff",
          2364 => x"9a",
          2365 => x"55",
          2366 => x"76",
          2367 => x"53",
          2368 => x"09",
          2369 => x"38",
          2370 => x"52",
          2371 => x"eb",
          2372 => x"3d",
          2373 => x"3d",
          2374 => x"5b",
          2375 => x"08",
          2376 => x"15",
          2377 => x"81",
          2378 => x"15",
          2379 => x"51",
          2380 => x"81",
          2381 => x"58",
          2382 => x"08",
          2383 => x"9c",
          2384 => x"33",
          2385 => x"86",
          2386 => x"80",
          2387 => x"13",
          2388 => x"06",
          2389 => x"06",
          2390 => x"72",
          2391 => x"81",
          2392 => x"53",
          2393 => x"2e",
          2394 => x"53",
          2395 => x"a9",
          2396 => x"74",
          2397 => x"72",
          2398 => x"38",
          2399 => x"99",
          2400 => x"a4",
          2401 => x"06",
          2402 => x"88",
          2403 => x"06",
          2404 => x"54",
          2405 => x"a0",
          2406 => x"74",
          2407 => x"3f",
          2408 => x"08",
          2409 => x"a4",
          2410 => x"98",
          2411 => x"fa",
          2412 => x"80",
          2413 => x"0c",
          2414 => x"a4",
          2415 => x"0d",
          2416 => x"0d",
          2417 => x"57",
          2418 => x"73",
          2419 => x"3f",
          2420 => x"08",
          2421 => x"a4",
          2422 => x"98",
          2423 => x"75",
          2424 => x"3f",
          2425 => x"08",
          2426 => x"a4",
          2427 => x"a0",
          2428 => x"a4",
          2429 => x"14",
          2430 => x"db",
          2431 => x"a0",
          2432 => x"14",
          2433 => x"ac",
          2434 => x"83",
          2435 => x"81",
          2436 => x"87",
          2437 => x"fd",
          2438 => x"70",
          2439 => x"08",
          2440 => x"55",
          2441 => x"3f",
          2442 => x"08",
          2443 => x"13",
          2444 => x"73",
          2445 => x"83",
          2446 => x"3d",
          2447 => x"3d",
          2448 => x"57",
          2449 => x"89",
          2450 => x"17",
          2451 => x"81",
          2452 => x"70",
          2453 => x"55",
          2454 => x"08",
          2455 => x"81",
          2456 => x"52",
          2457 => x"a8",
          2458 => x"2e",
          2459 => x"84",
          2460 => x"52",
          2461 => x"09",
          2462 => x"38",
          2463 => x"81",
          2464 => x"81",
          2465 => x"73",
          2466 => x"55",
          2467 => x"55",
          2468 => x"c5",
          2469 => x"88",
          2470 => x"0b",
          2471 => x"9c",
          2472 => x"8b",
          2473 => x"17",
          2474 => x"08",
          2475 => x"52",
          2476 => x"81",
          2477 => x"76",
          2478 => x"51",
          2479 => x"81",
          2480 => x"86",
          2481 => x"12",
          2482 => x"3f",
          2483 => x"08",
          2484 => x"88",
          2485 => x"f3",
          2486 => x"70",
          2487 => x"80",
          2488 => x"51",
          2489 => x"af",
          2490 => x"81",
          2491 => x"dc",
          2492 => x"74",
          2493 => x"38",
          2494 => x"88",
          2495 => x"39",
          2496 => x"80",
          2497 => x"56",
          2498 => x"af",
          2499 => x"06",
          2500 => x"56",
          2501 => x"32",
          2502 => x"80",
          2503 => x"51",
          2504 => x"dc",
          2505 => x"1c",
          2506 => x"33",
          2507 => x"9f",
          2508 => x"ff",
          2509 => x"1c",
          2510 => x"7a",
          2511 => x"3f",
          2512 => x"08",
          2513 => x"39",
          2514 => x"a0",
          2515 => x"5e",
          2516 => x"52",
          2517 => x"ff",
          2518 => x"59",
          2519 => x"33",
          2520 => x"ae",
          2521 => x"06",
          2522 => x"78",
          2523 => x"81",
          2524 => x"32",
          2525 => x"9f",
          2526 => x"26",
          2527 => x"53",
          2528 => x"73",
          2529 => x"17",
          2530 => x"34",
          2531 => x"db",
          2532 => x"32",
          2533 => x"9f",
          2534 => x"54",
          2535 => x"2e",
          2536 => x"80",
          2537 => x"75",
          2538 => x"bd",
          2539 => x"7e",
          2540 => x"a0",
          2541 => x"bd",
          2542 => x"82",
          2543 => x"18",
          2544 => x"1a",
          2545 => x"a0",
          2546 => x"fc",
          2547 => x"32",
          2548 => x"80",
          2549 => x"30",
          2550 => x"71",
          2551 => x"51",
          2552 => x"55",
          2553 => x"ac",
          2554 => x"81",
          2555 => x"78",
          2556 => x"51",
          2557 => x"af",
          2558 => x"06",
          2559 => x"55",
          2560 => x"32",
          2561 => x"80",
          2562 => x"51",
          2563 => x"db",
          2564 => x"39",
          2565 => x"09",
          2566 => x"38",
          2567 => x"7c",
          2568 => x"54",
          2569 => x"a2",
          2570 => x"32",
          2571 => x"ae",
          2572 => x"72",
          2573 => x"9f",
          2574 => x"51",
          2575 => x"74",
          2576 => x"88",
          2577 => x"fe",
          2578 => x"98",
          2579 => x"80",
          2580 => x"75",
          2581 => x"81",
          2582 => x"33",
          2583 => x"51",
          2584 => x"81",
          2585 => x"80",
          2586 => x"78",
          2587 => x"81",
          2588 => x"5a",
          2589 => x"d2",
          2590 => x"a4",
          2591 => x"80",
          2592 => x"1c",
          2593 => x"27",
          2594 => x"79",
          2595 => x"74",
          2596 => x"7a",
          2597 => x"74",
          2598 => x"39",
          2599 => x"ba",
          2600 => x"fe",
          2601 => x"a4",
          2602 => x"ff",
          2603 => x"73",
          2604 => x"38",
          2605 => x"81",
          2606 => x"54",
          2607 => x"75",
          2608 => x"17",
          2609 => x"39",
          2610 => x"0c",
          2611 => x"99",
          2612 => x"54",
          2613 => x"2e",
          2614 => x"84",
          2615 => x"34",
          2616 => x"76",
          2617 => x"8b",
          2618 => x"81",
          2619 => x"56",
          2620 => x"80",
          2621 => x"1b",
          2622 => x"08",
          2623 => x"51",
          2624 => x"81",
          2625 => x"56",
          2626 => x"08",
          2627 => x"98",
          2628 => x"76",
          2629 => x"3f",
          2630 => x"08",
          2631 => x"a4",
          2632 => x"38",
          2633 => x"70",
          2634 => x"73",
          2635 => x"be",
          2636 => x"33",
          2637 => x"73",
          2638 => x"8b",
          2639 => x"83",
          2640 => x"06",
          2641 => x"73",
          2642 => x"53",
          2643 => x"51",
          2644 => x"81",
          2645 => x"80",
          2646 => x"75",
          2647 => x"f3",
          2648 => x"9f",
          2649 => x"1c",
          2650 => x"74",
          2651 => x"38",
          2652 => x"09",
          2653 => x"e7",
          2654 => x"2a",
          2655 => x"77",
          2656 => x"51",
          2657 => x"2e",
          2658 => x"81",
          2659 => x"80",
          2660 => x"38",
          2661 => x"ab",
          2662 => x"55",
          2663 => x"75",
          2664 => x"73",
          2665 => x"55",
          2666 => x"82",
          2667 => x"06",
          2668 => x"ab",
          2669 => x"33",
          2670 => x"70",
          2671 => x"55",
          2672 => x"2e",
          2673 => x"1b",
          2674 => x"06",
          2675 => x"52",
          2676 => x"db",
          2677 => x"a4",
          2678 => x"0c",
          2679 => x"74",
          2680 => x"0c",
          2681 => x"04",
          2682 => x"7c",
          2683 => x"08",
          2684 => x"55",
          2685 => x"59",
          2686 => x"81",
          2687 => x"70",
          2688 => x"33",
          2689 => x"52",
          2690 => x"2e",
          2691 => x"ee",
          2692 => x"2e",
          2693 => x"81",
          2694 => x"33",
          2695 => x"81",
          2696 => x"52",
          2697 => x"26",
          2698 => x"14",
          2699 => x"06",
          2700 => x"52",
          2701 => x"80",
          2702 => x"0b",
          2703 => x"59",
          2704 => x"7a",
          2705 => x"70",
          2706 => x"33",
          2707 => x"05",
          2708 => x"9f",
          2709 => x"53",
          2710 => x"89",
          2711 => x"70",
          2712 => x"54",
          2713 => x"12",
          2714 => x"26",
          2715 => x"12",
          2716 => x"06",
          2717 => x"30",
          2718 => x"51",
          2719 => x"2e",
          2720 => x"85",
          2721 => x"be",
          2722 => x"74",
          2723 => x"30",
          2724 => x"9f",
          2725 => x"2a",
          2726 => x"54",
          2727 => x"2e",
          2728 => x"15",
          2729 => x"55",
          2730 => x"ff",
          2731 => x"39",
          2732 => x"86",
          2733 => x"7c",
          2734 => x"51",
          2735 => x"cb",
          2736 => x"70",
          2737 => x"0c",
          2738 => x"04",
          2739 => x"78",
          2740 => x"83",
          2741 => x"0b",
          2742 => x"79",
          2743 => x"e2",
          2744 => x"55",
          2745 => x"08",
          2746 => x"84",
          2747 => x"df",
          2748 => x"cb",
          2749 => x"ff",
          2750 => x"83",
          2751 => x"d4",
          2752 => x"81",
          2753 => x"38",
          2754 => x"17",
          2755 => x"74",
          2756 => x"09",
          2757 => x"38",
          2758 => x"81",
          2759 => x"30",
          2760 => x"79",
          2761 => x"54",
          2762 => x"74",
          2763 => x"09",
          2764 => x"38",
          2765 => x"ba",
          2766 => x"ea",
          2767 => x"b1",
          2768 => x"a4",
          2769 => x"cb",
          2770 => x"2e",
          2771 => x"53",
          2772 => x"52",
          2773 => x"51",
          2774 => x"81",
          2775 => x"55",
          2776 => x"08",
          2777 => x"38",
          2778 => x"81",
          2779 => x"88",
          2780 => x"f2",
          2781 => x"02",
          2782 => x"cb",
          2783 => x"55",
          2784 => x"60",
          2785 => x"3f",
          2786 => x"08",
          2787 => x"80",
          2788 => x"a4",
          2789 => x"fc",
          2790 => x"a4",
          2791 => x"81",
          2792 => x"70",
          2793 => x"8c",
          2794 => x"2e",
          2795 => x"73",
          2796 => x"81",
          2797 => x"33",
          2798 => x"80",
          2799 => x"81",
          2800 => x"d7",
          2801 => x"cb",
          2802 => x"ff",
          2803 => x"06",
          2804 => x"98",
          2805 => x"2e",
          2806 => x"74",
          2807 => x"81",
          2808 => x"8a",
          2809 => x"ac",
          2810 => x"39",
          2811 => x"77",
          2812 => x"81",
          2813 => x"33",
          2814 => x"3f",
          2815 => x"08",
          2816 => x"70",
          2817 => x"55",
          2818 => x"86",
          2819 => x"80",
          2820 => x"74",
          2821 => x"81",
          2822 => x"8a",
          2823 => x"f4",
          2824 => x"53",
          2825 => x"fd",
          2826 => x"cb",
          2827 => x"ff",
          2828 => x"82",
          2829 => x"06",
          2830 => x"8c",
          2831 => x"58",
          2832 => x"f6",
          2833 => x"58",
          2834 => x"2e",
          2835 => x"fa",
          2836 => x"e8",
          2837 => x"a4",
          2838 => x"78",
          2839 => x"5a",
          2840 => x"90",
          2841 => x"75",
          2842 => x"38",
          2843 => x"3d",
          2844 => x"70",
          2845 => x"08",
          2846 => x"7a",
          2847 => x"38",
          2848 => x"51",
          2849 => x"81",
          2850 => x"81",
          2851 => x"81",
          2852 => x"38",
          2853 => x"83",
          2854 => x"38",
          2855 => x"84",
          2856 => x"38",
          2857 => x"81",
          2858 => x"38",
          2859 => x"db",
          2860 => x"cb",
          2861 => x"ff",
          2862 => x"72",
          2863 => x"09",
          2864 => x"d0",
          2865 => x"14",
          2866 => x"3f",
          2867 => x"08",
          2868 => x"06",
          2869 => x"38",
          2870 => x"51",
          2871 => x"81",
          2872 => x"58",
          2873 => x"0c",
          2874 => x"33",
          2875 => x"80",
          2876 => x"ff",
          2877 => x"ff",
          2878 => x"55",
          2879 => x"81",
          2880 => x"38",
          2881 => x"06",
          2882 => x"80",
          2883 => x"52",
          2884 => x"8a",
          2885 => x"80",
          2886 => x"ff",
          2887 => x"53",
          2888 => x"86",
          2889 => x"83",
          2890 => x"c5",
          2891 => x"f5",
          2892 => x"a4",
          2893 => x"cb",
          2894 => x"15",
          2895 => x"06",
          2896 => x"76",
          2897 => x"80",
          2898 => x"da",
          2899 => x"cb",
          2900 => x"ff",
          2901 => x"74",
          2902 => x"d4",
          2903 => x"dc",
          2904 => x"a4",
          2905 => x"c2",
          2906 => x"b9",
          2907 => x"a4",
          2908 => x"ff",
          2909 => x"56",
          2910 => x"83",
          2911 => x"14",
          2912 => x"71",
          2913 => x"5a",
          2914 => x"26",
          2915 => x"8a",
          2916 => x"74",
          2917 => x"ff",
          2918 => x"81",
          2919 => x"55",
          2920 => x"08",
          2921 => x"ec",
          2922 => x"a4",
          2923 => x"ff",
          2924 => x"83",
          2925 => x"74",
          2926 => x"26",
          2927 => x"57",
          2928 => x"26",
          2929 => x"57",
          2930 => x"56",
          2931 => x"82",
          2932 => x"15",
          2933 => x"0c",
          2934 => x"0c",
          2935 => x"a4",
          2936 => x"1d",
          2937 => x"54",
          2938 => x"2e",
          2939 => x"af",
          2940 => x"14",
          2941 => x"3f",
          2942 => x"08",
          2943 => x"06",
          2944 => x"72",
          2945 => x"79",
          2946 => x"80",
          2947 => x"d9",
          2948 => x"cb",
          2949 => x"15",
          2950 => x"2b",
          2951 => x"8d",
          2952 => x"2e",
          2953 => x"77",
          2954 => x"0c",
          2955 => x"76",
          2956 => x"38",
          2957 => x"70",
          2958 => x"81",
          2959 => x"53",
          2960 => x"89",
          2961 => x"56",
          2962 => x"08",
          2963 => x"38",
          2964 => x"15",
          2965 => x"8c",
          2966 => x"80",
          2967 => x"34",
          2968 => x"09",
          2969 => x"92",
          2970 => x"14",
          2971 => x"3f",
          2972 => x"08",
          2973 => x"06",
          2974 => x"2e",
          2975 => x"80",
          2976 => x"1b",
          2977 => x"db",
          2978 => x"cb",
          2979 => x"ea",
          2980 => x"a4",
          2981 => x"34",
          2982 => x"51",
          2983 => x"81",
          2984 => x"83",
          2985 => x"53",
          2986 => x"d5",
          2987 => x"06",
          2988 => x"b4",
          2989 => x"84",
          2990 => x"a4",
          2991 => x"85",
          2992 => x"09",
          2993 => x"38",
          2994 => x"51",
          2995 => x"81",
          2996 => x"86",
          2997 => x"f2",
          2998 => x"06",
          2999 => x"9c",
          3000 => x"d8",
          3001 => x"a4",
          3002 => x"0c",
          3003 => x"51",
          3004 => x"81",
          3005 => x"8c",
          3006 => x"74",
          3007 => x"d0",
          3008 => x"53",
          3009 => x"d0",
          3010 => x"15",
          3011 => x"94",
          3012 => x"56",
          3013 => x"a4",
          3014 => x"0d",
          3015 => x"0d",
          3016 => x"55",
          3017 => x"b9",
          3018 => x"53",
          3019 => x"b1",
          3020 => x"52",
          3021 => x"a9",
          3022 => x"22",
          3023 => x"57",
          3024 => x"2e",
          3025 => x"99",
          3026 => x"33",
          3027 => x"3f",
          3028 => x"08",
          3029 => x"71",
          3030 => x"74",
          3031 => x"83",
          3032 => x"78",
          3033 => x"52",
          3034 => x"a4",
          3035 => x"0d",
          3036 => x"0d",
          3037 => x"33",
          3038 => x"3d",
          3039 => x"56",
          3040 => x"8b",
          3041 => x"81",
          3042 => x"24",
          3043 => x"cb",
          3044 => x"29",
          3045 => x"05",
          3046 => x"55",
          3047 => x"84",
          3048 => x"34",
          3049 => x"80",
          3050 => x"80",
          3051 => x"75",
          3052 => x"75",
          3053 => x"38",
          3054 => x"3d",
          3055 => x"05",
          3056 => x"3f",
          3057 => x"08",
          3058 => x"cb",
          3059 => x"3d",
          3060 => x"3d",
          3061 => x"84",
          3062 => x"05",
          3063 => x"89",
          3064 => x"2e",
          3065 => x"77",
          3066 => x"54",
          3067 => x"05",
          3068 => x"84",
          3069 => x"f6",
          3070 => x"cb",
          3071 => x"81",
          3072 => x"84",
          3073 => x"5c",
          3074 => x"3d",
          3075 => x"ed",
          3076 => x"cb",
          3077 => x"81",
          3078 => x"92",
          3079 => x"d7",
          3080 => x"98",
          3081 => x"73",
          3082 => x"38",
          3083 => x"9c",
          3084 => x"80",
          3085 => x"38",
          3086 => x"95",
          3087 => x"2e",
          3088 => x"aa",
          3089 => x"ea",
          3090 => x"cb",
          3091 => x"9e",
          3092 => x"05",
          3093 => x"54",
          3094 => x"38",
          3095 => x"70",
          3096 => x"54",
          3097 => x"8e",
          3098 => x"83",
          3099 => x"88",
          3100 => x"83",
          3101 => x"83",
          3102 => x"06",
          3103 => x"80",
          3104 => x"38",
          3105 => x"51",
          3106 => x"81",
          3107 => x"56",
          3108 => x"0a",
          3109 => x"05",
          3110 => x"3f",
          3111 => x"0b",
          3112 => x"80",
          3113 => x"7a",
          3114 => x"3f",
          3115 => x"9c",
          3116 => x"d1",
          3117 => x"81",
          3118 => x"34",
          3119 => x"80",
          3120 => x"b0",
          3121 => x"54",
          3122 => x"52",
          3123 => x"05",
          3124 => x"3f",
          3125 => x"08",
          3126 => x"a4",
          3127 => x"38",
          3128 => x"82",
          3129 => x"b2",
          3130 => x"84",
          3131 => x"06",
          3132 => x"73",
          3133 => x"38",
          3134 => x"ad",
          3135 => x"2a",
          3136 => x"51",
          3137 => x"2e",
          3138 => x"81",
          3139 => x"80",
          3140 => x"87",
          3141 => x"39",
          3142 => x"51",
          3143 => x"81",
          3144 => x"7b",
          3145 => x"12",
          3146 => x"81",
          3147 => x"81",
          3148 => x"83",
          3149 => x"06",
          3150 => x"80",
          3151 => x"77",
          3152 => x"58",
          3153 => x"08",
          3154 => x"63",
          3155 => x"63",
          3156 => x"57",
          3157 => x"81",
          3158 => x"81",
          3159 => x"88",
          3160 => x"9c",
          3161 => x"d2",
          3162 => x"cb",
          3163 => x"cb",
          3164 => x"1b",
          3165 => x"0c",
          3166 => x"22",
          3167 => x"77",
          3168 => x"80",
          3169 => x"34",
          3170 => x"1a",
          3171 => x"94",
          3172 => x"85",
          3173 => x"06",
          3174 => x"80",
          3175 => x"38",
          3176 => x"08",
          3177 => x"84",
          3178 => x"a4",
          3179 => x"0c",
          3180 => x"70",
          3181 => x"52",
          3182 => x"39",
          3183 => x"51",
          3184 => x"81",
          3185 => x"57",
          3186 => x"08",
          3187 => x"38",
          3188 => x"cb",
          3189 => x"2e",
          3190 => x"83",
          3191 => x"75",
          3192 => x"74",
          3193 => x"07",
          3194 => x"54",
          3195 => x"8a",
          3196 => x"75",
          3197 => x"73",
          3198 => x"98",
          3199 => x"a9",
          3200 => x"ff",
          3201 => x"80",
          3202 => x"76",
          3203 => x"d6",
          3204 => x"cb",
          3205 => x"38",
          3206 => x"39",
          3207 => x"81",
          3208 => x"05",
          3209 => x"84",
          3210 => x"0c",
          3211 => x"81",
          3212 => x"97",
          3213 => x"f2",
          3214 => x"63",
          3215 => x"40",
          3216 => x"7e",
          3217 => x"fc",
          3218 => x"51",
          3219 => x"81",
          3220 => x"55",
          3221 => x"08",
          3222 => x"19",
          3223 => x"80",
          3224 => x"74",
          3225 => x"39",
          3226 => x"81",
          3227 => x"56",
          3228 => x"82",
          3229 => x"39",
          3230 => x"1a",
          3231 => x"82",
          3232 => x"0b",
          3233 => x"81",
          3234 => x"39",
          3235 => x"94",
          3236 => x"55",
          3237 => x"83",
          3238 => x"7b",
          3239 => x"89",
          3240 => x"08",
          3241 => x"06",
          3242 => x"81",
          3243 => x"8a",
          3244 => x"05",
          3245 => x"06",
          3246 => x"a8",
          3247 => x"38",
          3248 => x"55",
          3249 => x"19",
          3250 => x"51",
          3251 => x"81",
          3252 => x"55",
          3253 => x"ff",
          3254 => x"ff",
          3255 => x"38",
          3256 => x"0c",
          3257 => x"52",
          3258 => x"cb",
          3259 => x"a4",
          3260 => x"ff",
          3261 => x"cb",
          3262 => x"7c",
          3263 => x"57",
          3264 => x"80",
          3265 => x"1a",
          3266 => x"22",
          3267 => x"75",
          3268 => x"38",
          3269 => x"58",
          3270 => x"53",
          3271 => x"1b",
          3272 => x"88",
          3273 => x"a4",
          3274 => x"38",
          3275 => x"33",
          3276 => x"80",
          3277 => x"b0",
          3278 => x"31",
          3279 => x"27",
          3280 => x"80",
          3281 => x"52",
          3282 => x"77",
          3283 => x"7d",
          3284 => x"e0",
          3285 => x"2b",
          3286 => x"76",
          3287 => x"94",
          3288 => x"ff",
          3289 => x"71",
          3290 => x"7b",
          3291 => x"38",
          3292 => x"19",
          3293 => x"51",
          3294 => x"81",
          3295 => x"fe",
          3296 => x"53",
          3297 => x"83",
          3298 => x"b4",
          3299 => x"51",
          3300 => x"7b",
          3301 => x"08",
          3302 => x"76",
          3303 => x"08",
          3304 => x"0c",
          3305 => x"f3",
          3306 => x"75",
          3307 => x"0c",
          3308 => x"04",
          3309 => x"60",
          3310 => x"40",
          3311 => x"80",
          3312 => x"3d",
          3313 => x"77",
          3314 => x"3f",
          3315 => x"08",
          3316 => x"a4",
          3317 => x"91",
          3318 => x"74",
          3319 => x"38",
          3320 => x"b8",
          3321 => x"33",
          3322 => x"70",
          3323 => x"56",
          3324 => x"74",
          3325 => x"a4",
          3326 => x"82",
          3327 => x"34",
          3328 => x"98",
          3329 => x"91",
          3330 => x"56",
          3331 => x"94",
          3332 => x"11",
          3333 => x"76",
          3334 => x"75",
          3335 => x"80",
          3336 => x"38",
          3337 => x"70",
          3338 => x"56",
          3339 => x"fd",
          3340 => x"11",
          3341 => x"77",
          3342 => x"5c",
          3343 => x"38",
          3344 => x"88",
          3345 => x"74",
          3346 => x"52",
          3347 => x"18",
          3348 => x"51",
          3349 => x"81",
          3350 => x"55",
          3351 => x"08",
          3352 => x"ab",
          3353 => x"2e",
          3354 => x"74",
          3355 => x"95",
          3356 => x"19",
          3357 => x"08",
          3358 => x"88",
          3359 => x"55",
          3360 => x"9c",
          3361 => x"09",
          3362 => x"38",
          3363 => x"c1",
          3364 => x"a4",
          3365 => x"38",
          3366 => x"52",
          3367 => x"97",
          3368 => x"a4",
          3369 => x"fe",
          3370 => x"cb",
          3371 => x"7c",
          3372 => x"57",
          3373 => x"80",
          3374 => x"1b",
          3375 => x"22",
          3376 => x"75",
          3377 => x"38",
          3378 => x"59",
          3379 => x"53",
          3380 => x"1a",
          3381 => x"be",
          3382 => x"a4",
          3383 => x"38",
          3384 => x"08",
          3385 => x"56",
          3386 => x"9b",
          3387 => x"53",
          3388 => x"77",
          3389 => x"7d",
          3390 => x"16",
          3391 => x"3f",
          3392 => x"0b",
          3393 => x"78",
          3394 => x"80",
          3395 => x"18",
          3396 => x"08",
          3397 => x"7e",
          3398 => x"3f",
          3399 => x"08",
          3400 => x"7e",
          3401 => x"0c",
          3402 => x"19",
          3403 => x"08",
          3404 => x"84",
          3405 => x"57",
          3406 => x"27",
          3407 => x"56",
          3408 => x"52",
          3409 => x"f9",
          3410 => x"a4",
          3411 => x"38",
          3412 => x"52",
          3413 => x"83",
          3414 => x"b4",
          3415 => x"d4",
          3416 => x"81",
          3417 => x"34",
          3418 => x"7e",
          3419 => x"0c",
          3420 => x"1a",
          3421 => x"94",
          3422 => x"1b",
          3423 => x"5e",
          3424 => x"27",
          3425 => x"55",
          3426 => x"0c",
          3427 => x"90",
          3428 => x"c0",
          3429 => x"90",
          3430 => x"56",
          3431 => x"a4",
          3432 => x"0d",
          3433 => x"0d",
          3434 => x"fc",
          3435 => x"52",
          3436 => x"3f",
          3437 => x"08",
          3438 => x"a4",
          3439 => x"38",
          3440 => x"70",
          3441 => x"81",
          3442 => x"55",
          3443 => x"80",
          3444 => x"16",
          3445 => x"51",
          3446 => x"81",
          3447 => x"57",
          3448 => x"08",
          3449 => x"a4",
          3450 => x"11",
          3451 => x"55",
          3452 => x"16",
          3453 => x"08",
          3454 => x"75",
          3455 => x"e8",
          3456 => x"08",
          3457 => x"51",
          3458 => x"82",
          3459 => x"52",
          3460 => x"c9",
          3461 => x"52",
          3462 => x"c9",
          3463 => x"54",
          3464 => x"15",
          3465 => x"cc",
          3466 => x"cb",
          3467 => x"17",
          3468 => x"06",
          3469 => x"90",
          3470 => x"81",
          3471 => x"8a",
          3472 => x"fc",
          3473 => x"70",
          3474 => x"d9",
          3475 => x"a4",
          3476 => x"cb",
          3477 => x"38",
          3478 => x"05",
          3479 => x"f1",
          3480 => x"cb",
          3481 => x"81",
          3482 => x"87",
          3483 => x"a4",
          3484 => x"72",
          3485 => x"0c",
          3486 => x"04",
          3487 => x"84",
          3488 => x"e4",
          3489 => x"80",
          3490 => x"a4",
          3491 => x"38",
          3492 => x"08",
          3493 => x"34",
          3494 => x"81",
          3495 => x"83",
          3496 => x"ef",
          3497 => x"53",
          3498 => x"05",
          3499 => x"51",
          3500 => x"81",
          3501 => x"55",
          3502 => x"08",
          3503 => x"76",
          3504 => x"93",
          3505 => x"51",
          3506 => x"81",
          3507 => x"55",
          3508 => x"08",
          3509 => x"80",
          3510 => x"70",
          3511 => x"56",
          3512 => x"89",
          3513 => x"94",
          3514 => x"b2",
          3515 => x"05",
          3516 => x"2a",
          3517 => x"51",
          3518 => x"80",
          3519 => x"76",
          3520 => x"52",
          3521 => x"3f",
          3522 => x"08",
          3523 => x"8e",
          3524 => x"a4",
          3525 => x"09",
          3526 => x"38",
          3527 => x"81",
          3528 => x"93",
          3529 => x"e4",
          3530 => x"6f",
          3531 => x"7a",
          3532 => x"9e",
          3533 => x"05",
          3534 => x"51",
          3535 => x"81",
          3536 => x"57",
          3537 => x"08",
          3538 => x"7b",
          3539 => x"94",
          3540 => x"55",
          3541 => x"73",
          3542 => x"ed",
          3543 => x"93",
          3544 => x"55",
          3545 => x"81",
          3546 => x"57",
          3547 => x"08",
          3548 => x"68",
          3549 => x"c9",
          3550 => x"cb",
          3551 => x"81",
          3552 => x"82",
          3553 => x"52",
          3554 => x"a3",
          3555 => x"a4",
          3556 => x"52",
          3557 => x"b8",
          3558 => x"a4",
          3559 => x"cb",
          3560 => x"a2",
          3561 => x"74",
          3562 => x"3f",
          3563 => x"08",
          3564 => x"a4",
          3565 => x"69",
          3566 => x"d9",
          3567 => x"81",
          3568 => x"2e",
          3569 => x"52",
          3570 => x"cf",
          3571 => x"a4",
          3572 => x"cb",
          3573 => x"2e",
          3574 => x"84",
          3575 => x"06",
          3576 => x"57",
          3577 => x"76",
          3578 => x"9e",
          3579 => x"05",
          3580 => x"dc",
          3581 => x"90",
          3582 => x"81",
          3583 => x"56",
          3584 => x"80",
          3585 => x"02",
          3586 => x"81",
          3587 => x"70",
          3588 => x"56",
          3589 => x"81",
          3590 => x"78",
          3591 => x"38",
          3592 => x"99",
          3593 => x"81",
          3594 => x"18",
          3595 => x"18",
          3596 => x"58",
          3597 => x"33",
          3598 => x"ee",
          3599 => x"6f",
          3600 => x"af",
          3601 => x"8d",
          3602 => x"2e",
          3603 => x"8a",
          3604 => x"6f",
          3605 => x"af",
          3606 => x"0b",
          3607 => x"33",
          3608 => x"81",
          3609 => x"70",
          3610 => x"52",
          3611 => x"56",
          3612 => x"8d",
          3613 => x"70",
          3614 => x"51",
          3615 => x"f5",
          3616 => x"54",
          3617 => x"a7",
          3618 => x"74",
          3619 => x"38",
          3620 => x"73",
          3621 => x"81",
          3622 => x"81",
          3623 => x"39",
          3624 => x"81",
          3625 => x"74",
          3626 => x"81",
          3627 => x"91",
          3628 => x"6e",
          3629 => x"59",
          3630 => x"7a",
          3631 => x"5c",
          3632 => x"26",
          3633 => x"7a",
          3634 => x"cb",
          3635 => x"3d",
          3636 => x"3d",
          3637 => x"8d",
          3638 => x"54",
          3639 => x"55",
          3640 => x"81",
          3641 => x"53",
          3642 => x"08",
          3643 => x"91",
          3644 => x"72",
          3645 => x"8c",
          3646 => x"73",
          3647 => x"38",
          3648 => x"70",
          3649 => x"81",
          3650 => x"57",
          3651 => x"73",
          3652 => x"08",
          3653 => x"94",
          3654 => x"75",
          3655 => x"97",
          3656 => x"11",
          3657 => x"2b",
          3658 => x"73",
          3659 => x"38",
          3660 => x"16",
          3661 => x"e5",
          3662 => x"a4",
          3663 => x"78",
          3664 => x"55",
          3665 => x"d5",
          3666 => x"a4",
          3667 => x"96",
          3668 => x"70",
          3669 => x"94",
          3670 => x"71",
          3671 => x"08",
          3672 => x"53",
          3673 => x"15",
          3674 => x"a6",
          3675 => x"74",
          3676 => x"3f",
          3677 => x"08",
          3678 => x"a4",
          3679 => x"81",
          3680 => x"cb",
          3681 => x"2e",
          3682 => x"81",
          3683 => x"88",
          3684 => x"98",
          3685 => x"80",
          3686 => x"38",
          3687 => x"80",
          3688 => x"77",
          3689 => x"08",
          3690 => x"0c",
          3691 => x"70",
          3692 => x"81",
          3693 => x"5a",
          3694 => x"2e",
          3695 => x"52",
          3696 => x"f9",
          3697 => x"a4",
          3698 => x"cb",
          3699 => x"38",
          3700 => x"08",
          3701 => x"73",
          3702 => x"c7",
          3703 => x"cb",
          3704 => x"73",
          3705 => x"38",
          3706 => x"af",
          3707 => x"73",
          3708 => x"27",
          3709 => x"98",
          3710 => x"a0",
          3711 => x"08",
          3712 => x"0c",
          3713 => x"06",
          3714 => x"2e",
          3715 => x"52",
          3716 => x"a3",
          3717 => x"a4",
          3718 => x"82",
          3719 => x"34",
          3720 => x"c4",
          3721 => x"91",
          3722 => x"53",
          3723 => x"89",
          3724 => x"a4",
          3725 => x"94",
          3726 => x"8c",
          3727 => x"27",
          3728 => x"8c",
          3729 => x"15",
          3730 => x"07",
          3731 => x"16",
          3732 => x"ff",
          3733 => x"80",
          3734 => x"77",
          3735 => x"2e",
          3736 => x"9c",
          3737 => x"53",
          3738 => x"a4",
          3739 => x"0d",
          3740 => x"0d",
          3741 => x"54",
          3742 => x"81",
          3743 => x"53",
          3744 => x"05",
          3745 => x"84",
          3746 => x"e7",
          3747 => x"a4",
          3748 => x"cb",
          3749 => x"ea",
          3750 => x"0c",
          3751 => x"51",
          3752 => x"81",
          3753 => x"55",
          3754 => x"08",
          3755 => x"ab",
          3756 => x"98",
          3757 => x"80",
          3758 => x"38",
          3759 => x"70",
          3760 => x"81",
          3761 => x"57",
          3762 => x"ad",
          3763 => x"08",
          3764 => x"d3",
          3765 => x"cb",
          3766 => x"17",
          3767 => x"86",
          3768 => x"17",
          3769 => x"75",
          3770 => x"3f",
          3771 => x"08",
          3772 => x"2e",
          3773 => x"85",
          3774 => x"86",
          3775 => x"2e",
          3776 => x"76",
          3777 => x"73",
          3778 => x"0c",
          3779 => x"04",
          3780 => x"76",
          3781 => x"05",
          3782 => x"53",
          3783 => x"81",
          3784 => x"87",
          3785 => x"a4",
          3786 => x"86",
          3787 => x"fb",
          3788 => x"79",
          3789 => x"05",
          3790 => x"56",
          3791 => x"3f",
          3792 => x"08",
          3793 => x"a4",
          3794 => x"38",
          3795 => x"81",
          3796 => x"52",
          3797 => x"f8",
          3798 => x"a4",
          3799 => x"ca",
          3800 => x"a4",
          3801 => x"51",
          3802 => x"81",
          3803 => x"53",
          3804 => x"08",
          3805 => x"81",
          3806 => x"80",
          3807 => x"81",
          3808 => x"a6",
          3809 => x"73",
          3810 => x"3f",
          3811 => x"51",
          3812 => x"81",
          3813 => x"84",
          3814 => x"70",
          3815 => x"2c",
          3816 => x"a4",
          3817 => x"51",
          3818 => x"81",
          3819 => x"87",
          3820 => x"ee",
          3821 => x"57",
          3822 => x"3d",
          3823 => x"3d",
          3824 => x"af",
          3825 => x"a4",
          3826 => x"cb",
          3827 => x"38",
          3828 => x"51",
          3829 => x"81",
          3830 => x"55",
          3831 => x"08",
          3832 => x"80",
          3833 => x"70",
          3834 => x"58",
          3835 => x"85",
          3836 => x"8d",
          3837 => x"2e",
          3838 => x"52",
          3839 => x"be",
          3840 => x"cb",
          3841 => x"3d",
          3842 => x"3d",
          3843 => x"55",
          3844 => x"92",
          3845 => x"52",
          3846 => x"de",
          3847 => x"cb",
          3848 => x"81",
          3849 => x"82",
          3850 => x"74",
          3851 => x"98",
          3852 => x"11",
          3853 => x"59",
          3854 => x"75",
          3855 => x"38",
          3856 => x"81",
          3857 => x"5b",
          3858 => x"82",
          3859 => x"39",
          3860 => x"08",
          3861 => x"59",
          3862 => x"09",
          3863 => x"38",
          3864 => x"57",
          3865 => x"3d",
          3866 => x"c1",
          3867 => x"cb",
          3868 => x"2e",
          3869 => x"cb",
          3870 => x"2e",
          3871 => x"cb",
          3872 => x"70",
          3873 => x"08",
          3874 => x"7a",
          3875 => x"7f",
          3876 => x"54",
          3877 => x"77",
          3878 => x"80",
          3879 => x"15",
          3880 => x"a4",
          3881 => x"75",
          3882 => x"52",
          3883 => x"52",
          3884 => x"8d",
          3885 => x"a4",
          3886 => x"cb",
          3887 => x"d6",
          3888 => x"33",
          3889 => x"1a",
          3890 => x"54",
          3891 => x"09",
          3892 => x"38",
          3893 => x"ff",
          3894 => x"81",
          3895 => x"83",
          3896 => x"70",
          3897 => x"25",
          3898 => x"59",
          3899 => x"9b",
          3900 => x"51",
          3901 => x"3f",
          3902 => x"08",
          3903 => x"70",
          3904 => x"25",
          3905 => x"59",
          3906 => x"75",
          3907 => x"7a",
          3908 => x"ff",
          3909 => x"7c",
          3910 => x"90",
          3911 => x"11",
          3912 => x"56",
          3913 => x"15",
          3914 => x"cb",
          3915 => x"3d",
          3916 => x"3d",
          3917 => x"3d",
          3918 => x"70",
          3919 => x"dd",
          3920 => x"a4",
          3921 => x"cb",
          3922 => x"a8",
          3923 => x"33",
          3924 => x"a0",
          3925 => x"33",
          3926 => x"70",
          3927 => x"55",
          3928 => x"73",
          3929 => x"8e",
          3930 => x"08",
          3931 => x"18",
          3932 => x"80",
          3933 => x"38",
          3934 => x"08",
          3935 => x"08",
          3936 => x"c4",
          3937 => x"cb",
          3938 => x"88",
          3939 => x"80",
          3940 => x"17",
          3941 => x"51",
          3942 => x"3f",
          3943 => x"08",
          3944 => x"81",
          3945 => x"81",
          3946 => x"a4",
          3947 => x"09",
          3948 => x"38",
          3949 => x"39",
          3950 => x"77",
          3951 => x"a4",
          3952 => x"08",
          3953 => x"98",
          3954 => x"81",
          3955 => x"52",
          3956 => x"bd",
          3957 => x"a4",
          3958 => x"17",
          3959 => x"0c",
          3960 => x"80",
          3961 => x"73",
          3962 => x"75",
          3963 => x"38",
          3964 => x"34",
          3965 => x"81",
          3966 => x"89",
          3967 => x"e2",
          3968 => x"53",
          3969 => x"a4",
          3970 => x"3d",
          3971 => x"3f",
          3972 => x"08",
          3973 => x"a4",
          3974 => x"38",
          3975 => x"3d",
          3976 => x"3d",
          3977 => x"d1",
          3978 => x"cb",
          3979 => x"81",
          3980 => x"81",
          3981 => x"80",
          3982 => x"70",
          3983 => x"81",
          3984 => x"56",
          3985 => x"81",
          3986 => x"98",
          3987 => x"74",
          3988 => x"38",
          3989 => x"05",
          3990 => x"06",
          3991 => x"55",
          3992 => x"38",
          3993 => x"51",
          3994 => x"81",
          3995 => x"74",
          3996 => x"81",
          3997 => x"56",
          3998 => x"80",
          3999 => x"54",
          4000 => x"08",
          4001 => x"2e",
          4002 => x"73",
          4003 => x"a4",
          4004 => x"52",
          4005 => x"52",
          4006 => x"3f",
          4007 => x"08",
          4008 => x"a4",
          4009 => x"38",
          4010 => x"08",
          4011 => x"cc",
          4012 => x"cb",
          4013 => x"81",
          4014 => x"86",
          4015 => x"80",
          4016 => x"cb",
          4017 => x"2e",
          4018 => x"cb",
          4019 => x"c0",
          4020 => x"ce",
          4021 => x"cb",
          4022 => x"cb",
          4023 => x"70",
          4024 => x"08",
          4025 => x"51",
          4026 => x"80",
          4027 => x"73",
          4028 => x"38",
          4029 => x"52",
          4030 => x"95",
          4031 => x"a4",
          4032 => x"8c",
          4033 => x"ff",
          4034 => x"81",
          4035 => x"55",
          4036 => x"a4",
          4037 => x"0d",
          4038 => x"0d",
          4039 => x"3d",
          4040 => x"9a",
          4041 => x"cb",
          4042 => x"a4",
          4043 => x"cb",
          4044 => x"b0",
          4045 => x"69",
          4046 => x"70",
          4047 => x"97",
          4048 => x"a4",
          4049 => x"cb",
          4050 => x"38",
          4051 => x"94",
          4052 => x"a4",
          4053 => x"09",
          4054 => x"88",
          4055 => x"df",
          4056 => x"85",
          4057 => x"51",
          4058 => x"74",
          4059 => x"78",
          4060 => x"8a",
          4061 => x"57",
          4062 => x"81",
          4063 => x"75",
          4064 => x"cb",
          4065 => x"38",
          4066 => x"cb",
          4067 => x"2e",
          4068 => x"83",
          4069 => x"81",
          4070 => x"ff",
          4071 => x"06",
          4072 => x"54",
          4073 => x"73",
          4074 => x"81",
          4075 => x"52",
          4076 => x"a4",
          4077 => x"a4",
          4078 => x"cb",
          4079 => x"9a",
          4080 => x"a0",
          4081 => x"51",
          4082 => x"3f",
          4083 => x"0b",
          4084 => x"78",
          4085 => x"bf",
          4086 => x"88",
          4087 => x"80",
          4088 => x"ff",
          4089 => x"75",
          4090 => x"11",
          4091 => x"f8",
          4092 => x"78",
          4093 => x"80",
          4094 => x"ff",
          4095 => x"78",
          4096 => x"80",
          4097 => x"7f",
          4098 => x"d4",
          4099 => x"c9",
          4100 => x"54",
          4101 => x"15",
          4102 => x"cb",
          4103 => x"cb",
          4104 => x"81",
          4105 => x"b2",
          4106 => x"b2",
          4107 => x"96",
          4108 => x"b5",
          4109 => x"53",
          4110 => x"51",
          4111 => x"64",
          4112 => x"8b",
          4113 => x"54",
          4114 => x"15",
          4115 => x"ff",
          4116 => x"81",
          4117 => x"54",
          4118 => x"53",
          4119 => x"51",
          4120 => x"3f",
          4121 => x"a4",
          4122 => x"0d",
          4123 => x"0d",
          4124 => x"05",
          4125 => x"3f",
          4126 => x"3d",
          4127 => x"52",
          4128 => x"d5",
          4129 => x"cb",
          4130 => x"81",
          4131 => x"82",
          4132 => x"4d",
          4133 => x"52",
          4134 => x"52",
          4135 => x"3f",
          4136 => x"08",
          4137 => x"a4",
          4138 => x"38",
          4139 => x"05",
          4140 => x"06",
          4141 => x"73",
          4142 => x"a0",
          4143 => x"08",
          4144 => x"ff",
          4145 => x"ff",
          4146 => x"ac",
          4147 => x"92",
          4148 => x"54",
          4149 => x"3f",
          4150 => x"52",
          4151 => x"f7",
          4152 => x"a4",
          4153 => x"cb",
          4154 => x"38",
          4155 => x"09",
          4156 => x"38",
          4157 => x"08",
          4158 => x"88",
          4159 => x"39",
          4160 => x"08",
          4161 => x"81",
          4162 => x"38",
          4163 => x"b1",
          4164 => x"a4",
          4165 => x"cb",
          4166 => x"c8",
          4167 => x"93",
          4168 => x"ff",
          4169 => x"8d",
          4170 => x"b4",
          4171 => x"af",
          4172 => x"17",
          4173 => x"33",
          4174 => x"70",
          4175 => x"55",
          4176 => x"38",
          4177 => x"54",
          4178 => x"34",
          4179 => x"0b",
          4180 => x"8b",
          4181 => x"84",
          4182 => x"06",
          4183 => x"73",
          4184 => x"e5",
          4185 => x"2e",
          4186 => x"75",
          4187 => x"c6",
          4188 => x"cb",
          4189 => x"78",
          4190 => x"bb",
          4191 => x"81",
          4192 => x"80",
          4193 => x"38",
          4194 => x"08",
          4195 => x"ff",
          4196 => x"81",
          4197 => x"79",
          4198 => x"58",
          4199 => x"cb",
          4200 => x"c0",
          4201 => x"33",
          4202 => x"2e",
          4203 => x"99",
          4204 => x"75",
          4205 => x"c6",
          4206 => x"54",
          4207 => x"15",
          4208 => x"81",
          4209 => x"9c",
          4210 => x"c8",
          4211 => x"cb",
          4212 => x"81",
          4213 => x"8c",
          4214 => x"ff",
          4215 => x"81",
          4216 => x"55",
          4217 => x"a4",
          4218 => x"0d",
          4219 => x"0d",
          4220 => x"05",
          4221 => x"05",
          4222 => x"33",
          4223 => x"53",
          4224 => x"05",
          4225 => x"51",
          4226 => x"81",
          4227 => x"55",
          4228 => x"08",
          4229 => x"78",
          4230 => x"95",
          4231 => x"51",
          4232 => x"81",
          4233 => x"55",
          4234 => x"08",
          4235 => x"80",
          4236 => x"81",
          4237 => x"86",
          4238 => x"38",
          4239 => x"61",
          4240 => x"12",
          4241 => x"7a",
          4242 => x"51",
          4243 => x"74",
          4244 => x"78",
          4245 => x"83",
          4246 => x"51",
          4247 => x"3f",
          4248 => x"08",
          4249 => x"cb",
          4250 => x"3d",
          4251 => x"3d",
          4252 => x"82",
          4253 => x"d0",
          4254 => x"3d",
          4255 => x"3f",
          4256 => x"08",
          4257 => x"a4",
          4258 => x"38",
          4259 => x"52",
          4260 => x"05",
          4261 => x"3f",
          4262 => x"08",
          4263 => x"a4",
          4264 => x"02",
          4265 => x"33",
          4266 => x"54",
          4267 => x"a6",
          4268 => x"22",
          4269 => x"71",
          4270 => x"53",
          4271 => x"51",
          4272 => x"3f",
          4273 => x"0b",
          4274 => x"76",
          4275 => x"b8",
          4276 => x"a4",
          4277 => x"81",
          4278 => x"93",
          4279 => x"ea",
          4280 => x"6b",
          4281 => x"53",
          4282 => x"05",
          4283 => x"51",
          4284 => x"81",
          4285 => x"81",
          4286 => x"30",
          4287 => x"a4",
          4288 => x"25",
          4289 => x"79",
          4290 => x"85",
          4291 => x"75",
          4292 => x"73",
          4293 => x"f9",
          4294 => x"80",
          4295 => x"8d",
          4296 => x"54",
          4297 => x"3f",
          4298 => x"08",
          4299 => x"a4",
          4300 => x"38",
          4301 => x"51",
          4302 => x"81",
          4303 => x"57",
          4304 => x"08",
          4305 => x"cb",
          4306 => x"cb",
          4307 => x"5b",
          4308 => x"18",
          4309 => x"18",
          4310 => x"74",
          4311 => x"81",
          4312 => x"78",
          4313 => x"8b",
          4314 => x"54",
          4315 => x"75",
          4316 => x"38",
          4317 => x"1b",
          4318 => x"55",
          4319 => x"2e",
          4320 => x"39",
          4321 => x"09",
          4322 => x"38",
          4323 => x"80",
          4324 => x"70",
          4325 => x"25",
          4326 => x"80",
          4327 => x"38",
          4328 => x"bc",
          4329 => x"11",
          4330 => x"ff",
          4331 => x"81",
          4332 => x"57",
          4333 => x"08",
          4334 => x"70",
          4335 => x"80",
          4336 => x"83",
          4337 => x"80",
          4338 => x"84",
          4339 => x"a7",
          4340 => x"b4",
          4341 => x"ad",
          4342 => x"cb",
          4343 => x"0c",
          4344 => x"a4",
          4345 => x"0d",
          4346 => x"0d",
          4347 => x"3d",
          4348 => x"52",
          4349 => x"ce",
          4350 => x"cb",
          4351 => x"cb",
          4352 => x"54",
          4353 => x"08",
          4354 => x"8b",
          4355 => x"8b",
          4356 => x"59",
          4357 => x"3f",
          4358 => x"33",
          4359 => x"06",
          4360 => x"57",
          4361 => x"81",
          4362 => x"58",
          4363 => x"06",
          4364 => x"4e",
          4365 => x"ff",
          4366 => x"81",
          4367 => x"80",
          4368 => x"6c",
          4369 => x"53",
          4370 => x"ae",
          4371 => x"cb",
          4372 => x"2e",
          4373 => x"88",
          4374 => x"6d",
          4375 => x"55",
          4376 => x"cb",
          4377 => x"ff",
          4378 => x"83",
          4379 => x"51",
          4380 => x"26",
          4381 => x"15",
          4382 => x"ff",
          4383 => x"80",
          4384 => x"87",
          4385 => x"80",
          4386 => x"74",
          4387 => x"38",
          4388 => x"bc",
          4389 => x"ae",
          4390 => x"cb",
          4391 => x"38",
          4392 => x"27",
          4393 => x"89",
          4394 => x"8b",
          4395 => x"27",
          4396 => x"55",
          4397 => x"81",
          4398 => x"8f",
          4399 => x"2a",
          4400 => x"70",
          4401 => x"34",
          4402 => x"74",
          4403 => x"05",
          4404 => x"17",
          4405 => x"70",
          4406 => x"52",
          4407 => x"73",
          4408 => x"c8",
          4409 => x"33",
          4410 => x"73",
          4411 => x"81",
          4412 => x"80",
          4413 => x"02",
          4414 => x"76",
          4415 => x"51",
          4416 => x"2e",
          4417 => x"87",
          4418 => x"57",
          4419 => x"79",
          4420 => x"80",
          4421 => x"70",
          4422 => x"ba",
          4423 => x"cb",
          4424 => x"81",
          4425 => x"80",
          4426 => x"52",
          4427 => x"bf",
          4428 => x"cb",
          4429 => x"81",
          4430 => x"8d",
          4431 => x"c4",
          4432 => x"e5",
          4433 => x"c6",
          4434 => x"a4",
          4435 => x"09",
          4436 => x"cc",
          4437 => x"76",
          4438 => x"c4",
          4439 => x"74",
          4440 => x"b0",
          4441 => x"a4",
          4442 => x"cb",
          4443 => x"38",
          4444 => x"cb",
          4445 => x"67",
          4446 => x"db",
          4447 => x"88",
          4448 => x"34",
          4449 => x"52",
          4450 => x"ab",
          4451 => x"54",
          4452 => x"15",
          4453 => x"ff",
          4454 => x"81",
          4455 => x"54",
          4456 => x"81",
          4457 => x"9c",
          4458 => x"f2",
          4459 => x"62",
          4460 => x"80",
          4461 => x"93",
          4462 => x"55",
          4463 => x"5e",
          4464 => x"3f",
          4465 => x"08",
          4466 => x"a4",
          4467 => x"38",
          4468 => x"58",
          4469 => x"38",
          4470 => x"97",
          4471 => x"08",
          4472 => x"38",
          4473 => x"70",
          4474 => x"81",
          4475 => x"55",
          4476 => x"87",
          4477 => x"39",
          4478 => x"90",
          4479 => x"82",
          4480 => x"8a",
          4481 => x"89",
          4482 => x"7f",
          4483 => x"56",
          4484 => x"3f",
          4485 => x"06",
          4486 => x"72",
          4487 => x"81",
          4488 => x"05",
          4489 => x"7c",
          4490 => x"55",
          4491 => x"27",
          4492 => x"16",
          4493 => x"83",
          4494 => x"76",
          4495 => x"80",
          4496 => x"79",
          4497 => x"99",
          4498 => x"7f",
          4499 => x"14",
          4500 => x"83",
          4501 => x"81",
          4502 => x"81",
          4503 => x"38",
          4504 => x"08",
          4505 => x"95",
          4506 => x"a4",
          4507 => x"81",
          4508 => x"7b",
          4509 => x"06",
          4510 => x"39",
          4511 => x"56",
          4512 => x"09",
          4513 => x"b9",
          4514 => x"80",
          4515 => x"80",
          4516 => x"78",
          4517 => x"7a",
          4518 => x"38",
          4519 => x"73",
          4520 => x"81",
          4521 => x"ff",
          4522 => x"74",
          4523 => x"ff",
          4524 => x"81",
          4525 => x"58",
          4526 => x"08",
          4527 => x"74",
          4528 => x"16",
          4529 => x"73",
          4530 => x"39",
          4531 => x"7e",
          4532 => x"0c",
          4533 => x"2e",
          4534 => x"88",
          4535 => x"8c",
          4536 => x"1a",
          4537 => x"07",
          4538 => x"1b",
          4539 => x"08",
          4540 => x"16",
          4541 => x"75",
          4542 => x"38",
          4543 => x"90",
          4544 => x"15",
          4545 => x"54",
          4546 => x"34",
          4547 => x"81",
          4548 => x"90",
          4549 => x"e9",
          4550 => x"6d",
          4551 => x"80",
          4552 => x"9d",
          4553 => x"5c",
          4554 => x"3f",
          4555 => x"0b",
          4556 => x"08",
          4557 => x"38",
          4558 => x"08",
          4559 => x"cb",
          4560 => x"08",
          4561 => x"80",
          4562 => x"80",
          4563 => x"cb",
          4564 => x"ff",
          4565 => x"52",
          4566 => x"a0",
          4567 => x"cb",
          4568 => x"ff",
          4569 => x"06",
          4570 => x"56",
          4571 => x"38",
          4572 => x"70",
          4573 => x"55",
          4574 => x"8b",
          4575 => x"3d",
          4576 => x"83",
          4577 => x"ff",
          4578 => x"81",
          4579 => x"99",
          4580 => x"74",
          4581 => x"38",
          4582 => x"80",
          4583 => x"ff",
          4584 => x"55",
          4585 => x"83",
          4586 => x"78",
          4587 => x"38",
          4588 => x"26",
          4589 => x"81",
          4590 => x"8b",
          4591 => x"79",
          4592 => x"80",
          4593 => x"93",
          4594 => x"39",
          4595 => x"6e",
          4596 => x"89",
          4597 => x"48",
          4598 => x"83",
          4599 => x"61",
          4600 => x"25",
          4601 => x"55",
          4602 => x"8a",
          4603 => x"3d",
          4604 => x"81",
          4605 => x"ff",
          4606 => x"81",
          4607 => x"a4",
          4608 => x"38",
          4609 => x"70",
          4610 => x"cb",
          4611 => x"56",
          4612 => x"38",
          4613 => x"55",
          4614 => x"75",
          4615 => x"38",
          4616 => x"70",
          4617 => x"ff",
          4618 => x"83",
          4619 => x"78",
          4620 => x"89",
          4621 => x"81",
          4622 => x"06",
          4623 => x"80",
          4624 => x"77",
          4625 => x"74",
          4626 => x"8d",
          4627 => x"06",
          4628 => x"2e",
          4629 => x"77",
          4630 => x"93",
          4631 => x"74",
          4632 => x"cb",
          4633 => x"7d",
          4634 => x"81",
          4635 => x"38",
          4636 => x"66",
          4637 => x"81",
          4638 => x"a4",
          4639 => x"74",
          4640 => x"38",
          4641 => x"98",
          4642 => x"a4",
          4643 => x"82",
          4644 => x"57",
          4645 => x"80",
          4646 => x"76",
          4647 => x"38",
          4648 => x"51",
          4649 => x"3f",
          4650 => x"08",
          4651 => x"87",
          4652 => x"2a",
          4653 => x"5c",
          4654 => x"cb",
          4655 => x"80",
          4656 => x"44",
          4657 => x"0a",
          4658 => x"ec",
          4659 => x"39",
          4660 => x"66",
          4661 => x"81",
          4662 => x"94",
          4663 => x"74",
          4664 => x"38",
          4665 => x"98",
          4666 => x"94",
          4667 => x"82",
          4668 => x"57",
          4669 => x"80",
          4670 => x"76",
          4671 => x"38",
          4672 => x"51",
          4673 => x"3f",
          4674 => x"08",
          4675 => x"57",
          4676 => x"08",
          4677 => x"96",
          4678 => x"81",
          4679 => x"10",
          4680 => x"08",
          4681 => x"72",
          4682 => x"59",
          4683 => x"ff",
          4684 => x"5d",
          4685 => x"44",
          4686 => x"11",
          4687 => x"70",
          4688 => x"71",
          4689 => x"06",
          4690 => x"52",
          4691 => x"40",
          4692 => x"09",
          4693 => x"38",
          4694 => x"18",
          4695 => x"39",
          4696 => x"79",
          4697 => x"70",
          4698 => x"58",
          4699 => x"76",
          4700 => x"38",
          4701 => x"7d",
          4702 => x"70",
          4703 => x"55",
          4704 => x"3f",
          4705 => x"08",
          4706 => x"2e",
          4707 => x"9b",
          4708 => x"a4",
          4709 => x"f5",
          4710 => x"38",
          4711 => x"38",
          4712 => x"59",
          4713 => x"38",
          4714 => x"7d",
          4715 => x"81",
          4716 => x"38",
          4717 => x"0b",
          4718 => x"08",
          4719 => x"78",
          4720 => x"1a",
          4721 => x"c0",
          4722 => x"74",
          4723 => x"39",
          4724 => x"55",
          4725 => x"8f",
          4726 => x"fd",
          4727 => x"cb",
          4728 => x"f5",
          4729 => x"78",
          4730 => x"79",
          4731 => x"80",
          4732 => x"f1",
          4733 => x"39",
          4734 => x"81",
          4735 => x"06",
          4736 => x"55",
          4737 => x"27",
          4738 => x"81",
          4739 => x"56",
          4740 => x"38",
          4741 => x"80",
          4742 => x"ff",
          4743 => x"8b",
          4744 => x"bc",
          4745 => x"ff",
          4746 => x"84",
          4747 => x"1b",
          4748 => x"b3",
          4749 => x"1c",
          4750 => x"ff",
          4751 => x"8e",
          4752 => x"a1",
          4753 => x"0b",
          4754 => x"7d",
          4755 => x"30",
          4756 => x"84",
          4757 => x"51",
          4758 => x"51",
          4759 => x"3f",
          4760 => x"83",
          4761 => x"90",
          4762 => x"ff",
          4763 => x"93",
          4764 => x"a0",
          4765 => x"39",
          4766 => x"1b",
          4767 => x"85",
          4768 => x"95",
          4769 => x"52",
          4770 => x"ff",
          4771 => x"81",
          4772 => x"1b",
          4773 => x"cf",
          4774 => x"9c",
          4775 => x"a0",
          4776 => x"83",
          4777 => x"06",
          4778 => x"82",
          4779 => x"52",
          4780 => x"51",
          4781 => x"3f",
          4782 => x"1b",
          4783 => x"c5",
          4784 => x"ac",
          4785 => x"a0",
          4786 => x"52",
          4787 => x"ff",
          4788 => x"86",
          4789 => x"51",
          4790 => x"3f",
          4791 => x"80",
          4792 => x"a9",
          4793 => x"1c",
          4794 => x"81",
          4795 => x"80",
          4796 => x"ae",
          4797 => x"b2",
          4798 => x"1b",
          4799 => x"85",
          4800 => x"ff",
          4801 => x"96",
          4802 => x"9f",
          4803 => x"80",
          4804 => x"34",
          4805 => x"1c",
          4806 => x"81",
          4807 => x"ab",
          4808 => x"a0",
          4809 => x"d4",
          4810 => x"fe",
          4811 => x"59",
          4812 => x"3f",
          4813 => x"53",
          4814 => x"51",
          4815 => x"3f",
          4816 => x"cb",
          4817 => x"e7",
          4818 => x"2e",
          4819 => x"80",
          4820 => x"54",
          4821 => x"53",
          4822 => x"51",
          4823 => x"3f",
          4824 => x"80",
          4825 => x"ff",
          4826 => x"84",
          4827 => x"d2",
          4828 => x"ff",
          4829 => x"86",
          4830 => x"f2",
          4831 => x"1b",
          4832 => x"81",
          4833 => x"52",
          4834 => x"51",
          4835 => x"3f",
          4836 => x"ec",
          4837 => x"9e",
          4838 => x"d4",
          4839 => x"51",
          4840 => x"3f",
          4841 => x"87",
          4842 => x"52",
          4843 => x"9a",
          4844 => x"54",
          4845 => x"7a",
          4846 => x"ff",
          4847 => x"65",
          4848 => x"7a",
          4849 => x"8f",
          4850 => x"80",
          4851 => x"2e",
          4852 => x"9a",
          4853 => x"7a",
          4854 => x"a9",
          4855 => x"84",
          4856 => x"9e",
          4857 => x"0a",
          4858 => x"51",
          4859 => x"ff",
          4860 => x"7d",
          4861 => x"38",
          4862 => x"52",
          4863 => x"9e",
          4864 => x"55",
          4865 => x"62",
          4866 => x"74",
          4867 => x"75",
          4868 => x"7e",
          4869 => x"fe",
          4870 => x"a4",
          4871 => x"38",
          4872 => x"81",
          4873 => x"52",
          4874 => x"9e",
          4875 => x"16",
          4876 => x"56",
          4877 => x"38",
          4878 => x"77",
          4879 => x"8d",
          4880 => x"7d",
          4881 => x"38",
          4882 => x"57",
          4883 => x"83",
          4884 => x"76",
          4885 => x"7a",
          4886 => x"ff",
          4887 => x"81",
          4888 => x"81",
          4889 => x"16",
          4890 => x"56",
          4891 => x"38",
          4892 => x"83",
          4893 => x"86",
          4894 => x"ff",
          4895 => x"38",
          4896 => x"82",
          4897 => x"81",
          4898 => x"06",
          4899 => x"fe",
          4900 => x"53",
          4901 => x"51",
          4902 => x"3f",
          4903 => x"52",
          4904 => x"9c",
          4905 => x"be",
          4906 => x"75",
          4907 => x"81",
          4908 => x"0b",
          4909 => x"77",
          4910 => x"75",
          4911 => x"60",
          4912 => x"80",
          4913 => x"75",
          4914 => x"d1",
          4915 => x"85",
          4916 => x"cb",
          4917 => x"2a",
          4918 => x"75",
          4919 => x"81",
          4920 => x"87",
          4921 => x"52",
          4922 => x"51",
          4923 => x"3f",
          4924 => x"ca",
          4925 => x"9c",
          4926 => x"54",
          4927 => x"52",
          4928 => x"98",
          4929 => x"56",
          4930 => x"08",
          4931 => x"53",
          4932 => x"51",
          4933 => x"3f",
          4934 => x"cb",
          4935 => x"38",
          4936 => x"56",
          4937 => x"56",
          4938 => x"cb",
          4939 => x"75",
          4940 => x"0c",
          4941 => x"04",
          4942 => x"73",
          4943 => x"26",
          4944 => x"71",
          4945 => x"b5",
          4946 => x"71",
          4947 => x"bd",
          4948 => x"80",
          4949 => x"c8",
          4950 => x"39",
          4951 => x"51",
          4952 => x"81",
          4953 => x"80",
          4954 => x"be",
          4955 => x"e4",
          4956 => x"90",
          4957 => x"39",
          4958 => x"51",
          4959 => x"81",
          4960 => x"80",
          4961 => x"be",
          4962 => x"c8",
          4963 => x"e4",
          4964 => x"39",
          4965 => x"51",
          4966 => x"bf",
          4967 => x"39",
          4968 => x"51",
          4969 => x"bf",
          4970 => x"39",
          4971 => x"51",
          4972 => x"c0",
          4973 => x"39",
          4974 => x"51",
          4975 => x"c0",
          4976 => x"39",
          4977 => x"51",
          4978 => x"c0",
          4979 => x"39",
          4980 => x"51",
          4981 => x"3f",
          4982 => x"04",
          4983 => x"77",
          4984 => x"74",
          4985 => x"8a",
          4986 => x"75",
          4987 => x"51",
          4988 => x"e8",
          4989 => x"fe",
          4990 => x"81",
          4991 => x"52",
          4992 => x"f2",
          4993 => x"cb",
          4994 => x"79",
          4995 => x"81",
          4996 => x"ff",
          4997 => x"87",
          4998 => x"f5",
          4999 => x"7f",
          5000 => x"05",
          5001 => x"33",
          5002 => x"66",
          5003 => x"5a",
          5004 => x"78",
          5005 => x"a8",
          5006 => x"fa",
          5007 => x"b0",
          5008 => x"8e",
          5009 => x"74",
          5010 => x"fc",
          5011 => x"2e",
          5012 => x"a0",
          5013 => x"80",
          5014 => x"16",
          5015 => x"27",
          5016 => x"22",
          5017 => x"b4",
          5018 => x"ca",
          5019 => x"81",
          5020 => x"ff",
          5021 => x"82",
          5022 => x"c3",
          5023 => x"53",
          5024 => x"8e",
          5025 => x"52",
          5026 => x"51",
          5027 => x"3f",
          5028 => x"c1",
          5029 => x"86",
          5030 => x"15",
          5031 => x"74",
          5032 => x"78",
          5033 => x"72",
          5034 => x"c1",
          5035 => x"8c",
          5036 => x"39",
          5037 => x"51",
          5038 => x"3f",
          5039 => x"a0",
          5040 => x"8d",
          5041 => x"39",
          5042 => x"51",
          5043 => x"3f",
          5044 => x"77",
          5045 => x"74",
          5046 => x"79",
          5047 => x"55",
          5048 => x"27",
          5049 => x"80",
          5050 => x"73",
          5051 => x"85",
          5052 => x"83",
          5053 => x"fe",
          5054 => x"81",
          5055 => x"39",
          5056 => x"51",
          5057 => x"3f",
          5058 => x"1a",
          5059 => x"fd",
          5060 => x"cb",
          5061 => x"2b",
          5062 => x"51",
          5063 => x"2e",
          5064 => x"a5",
          5065 => x"fb",
          5066 => x"a4",
          5067 => x"70",
          5068 => x"a0",
          5069 => x"70",
          5070 => x"2a",
          5071 => x"51",
          5072 => x"2e",
          5073 => x"dd",
          5074 => x"2e",
          5075 => x"85",
          5076 => x"8c",
          5077 => x"53",
          5078 => x"fd",
          5079 => x"53",
          5080 => x"a4",
          5081 => x"0d",
          5082 => x"0d",
          5083 => x"05",
          5084 => x"33",
          5085 => x"70",
          5086 => x"25",
          5087 => x"74",
          5088 => x"51",
          5089 => x"56",
          5090 => x"80",
          5091 => x"53",
          5092 => x"3d",
          5093 => x"c0",
          5094 => x"cb",
          5095 => x"81",
          5096 => x"b8",
          5097 => x"a4",
          5098 => x"98",
          5099 => x"cb",
          5100 => x"96",
          5101 => x"54",
          5102 => x"77",
          5103 => x"c4",
          5104 => x"cb",
          5105 => x"81",
          5106 => x"90",
          5107 => x"74",
          5108 => x"38",
          5109 => x"19",
          5110 => x"39",
          5111 => x"05",
          5112 => x"3f",
          5113 => x"77",
          5114 => x"51",
          5115 => x"2e",
          5116 => x"80",
          5117 => x"81",
          5118 => x"87",
          5119 => x"08",
          5120 => x"fb",
          5121 => x"57",
          5122 => x"a4",
          5123 => x"0d",
          5124 => x"0d",
          5125 => x"05",
          5126 => x"57",
          5127 => x"80",
          5128 => x"79",
          5129 => x"3f",
          5130 => x"08",
          5131 => x"80",
          5132 => x"75",
          5133 => x"38",
          5134 => x"55",
          5135 => x"cb",
          5136 => x"52",
          5137 => x"2d",
          5138 => x"08",
          5139 => x"77",
          5140 => x"cb",
          5141 => x"3d",
          5142 => x"3d",
          5143 => x"05",
          5144 => x"e4",
          5145 => x"ec",
          5146 => x"88",
          5147 => x"c8",
          5148 => x"ff",
          5149 => x"81",
          5150 => x"81",
          5151 => x"81",
          5152 => x"52",
          5153 => x"51",
          5154 => x"3f",
          5155 => x"85",
          5156 => x"92",
          5157 => x"0d",
          5158 => x"0d",
          5159 => x"80",
          5160 => x"80",
          5161 => x"51",
          5162 => x"3f",
          5163 => x"51",
          5164 => x"3f",
          5165 => x"f5",
          5166 => x"81",
          5167 => x"06",
          5168 => x"80",
          5169 => x"81",
          5170 => x"eb",
          5171 => x"c4",
          5172 => x"e3",
          5173 => x"fe",
          5174 => x"72",
          5175 => x"81",
          5176 => x"71",
          5177 => x"38",
          5178 => x"f5",
          5179 => x"c2",
          5180 => x"f7",
          5181 => x"51",
          5182 => x"3f",
          5183 => x"70",
          5184 => x"52",
          5185 => x"95",
          5186 => x"fe",
          5187 => x"81",
          5188 => x"fe",
          5189 => x"80",
          5190 => x"9b",
          5191 => x"2a",
          5192 => x"51",
          5193 => x"2e",
          5194 => x"51",
          5195 => x"3f",
          5196 => x"51",
          5197 => x"3f",
          5198 => x"f4",
          5199 => x"85",
          5200 => x"06",
          5201 => x"80",
          5202 => x"81",
          5203 => x"e7",
          5204 => x"90",
          5205 => x"df",
          5206 => x"fe",
          5207 => x"72",
          5208 => x"81",
          5209 => x"71",
          5210 => x"38",
          5211 => x"f4",
          5212 => x"c3",
          5213 => x"f6",
          5214 => x"51",
          5215 => x"3f",
          5216 => x"70",
          5217 => x"52",
          5218 => x"95",
          5219 => x"fe",
          5220 => x"81",
          5221 => x"fe",
          5222 => x"80",
          5223 => x"97",
          5224 => x"2a",
          5225 => x"51",
          5226 => x"2e",
          5227 => x"51",
          5228 => x"3f",
          5229 => x"51",
          5230 => x"3f",
          5231 => x"f3",
          5232 => x"ff",
          5233 => x"3d",
          5234 => x"3d",
          5235 => x"08",
          5236 => x"57",
          5237 => x"80",
          5238 => x"39",
          5239 => x"85",
          5240 => x"80",
          5241 => x"14",
          5242 => x"33",
          5243 => x"06",
          5244 => x"74",
          5245 => x"38",
          5246 => x"80",
          5247 => x"72",
          5248 => x"81",
          5249 => x"72",
          5250 => x"81",
          5251 => x"80",
          5252 => x"05",
          5253 => x"56",
          5254 => x"81",
          5255 => x"77",
          5256 => x"08",
          5257 => x"ed",
          5258 => x"cb",
          5259 => x"38",
          5260 => x"53",
          5261 => x"ff",
          5262 => x"16",
          5263 => x"06",
          5264 => x"76",
          5265 => x"ff",
          5266 => x"cb",
          5267 => x"3d",
          5268 => x"3d",
          5269 => x"71",
          5270 => x"0c",
          5271 => x"52",
          5272 => x"8a",
          5273 => x"cb",
          5274 => x"ff",
          5275 => x"7c",
          5276 => x"06",
          5277 => x"c4",
          5278 => x"3d",
          5279 => x"ff",
          5280 => x"7b",
          5281 => x"81",
          5282 => x"ff",
          5283 => x"81",
          5284 => x"7c",
          5285 => x"81",
          5286 => x"8e",
          5287 => x"70",
          5288 => x"c4",
          5289 => x"fe",
          5290 => x"3d",
          5291 => x"80",
          5292 => x"52",
          5293 => x"eb",
          5294 => x"f8",
          5295 => x"ff",
          5296 => x"b7",
          5297 => x"05",
          5298 => x"3f",
          5299 => x"08",
          5300 => x"90",
          5301 => x"78",
          5302 => x"8a",
          5303 => x"80",
          5304 => x"dc",
          5305 => x"2e",
          5306 => x"78",
          5307 => x"38",
          5308 => x"81",
          5309 => x"82",
          5310 => x"78",
          5311 => x"a2",
          5312 => x"39",
          5313 => x"82",
          5314 => x"94",
          5315 => x"38",
          5316 => x"78",
          5317 => x"85",
          5318 => x"80",
          5319 => x"38",
          5320 => x"83",
          5321 => x"bc",
          5322 => x"38",
          5323 => x"78",
          5324 => x"86",
          5325 => x"80",
          5326 => x"8c",
          5327 => x"39",
          5328 => x"2e",
          5329 => x"78",
          5330 => x"a9",
          5331 => x"d1",
          5332 => x"38",
          5333 => x"24",
          5334 => x"80",
          5335 => x"c4",
          5336 => x"39",
          5337 => x"2e",
          5338 => x"78",
          5339 => x"8a",
          5340 => x"97",
          5341 => x"83",
          5342 => x"38",
          5343 => x"24",
          5344 => x"80",
          5345 => x"9d",
          5346 => x"82",
          5347 => x"38",
          5348 => x"78",
          5349 => x"8b",
          5350 => x"81",
          5351 => x"82",
          5352 => x"39",
          5353 => x"f4",
          5354 => x"f8",
          5355 => x"83",
          5356 => x"cb",
          5357 => x"38",
          5358 => x"51",
          5359 => x"b7",
          5360 => x"11",
          5361 => x"05",
          5362 => x"df",
          5363 => x"a4",
          5364 => x"88",
          5365 => x"25",
          5366 => x"43",
          5367 => x"05",
          5368 => x"80",
          5369 => x"51",
          5370 => x"3f",
          5371 => x"08",
          5372 => x"59",
          5373 => x"81",
          5374 => x"fe",
          5375 => x"81",
          5376 => x"39",
          5377 => x"51",
          5378 => x"b7",
          5379 => x"11",
          5380 => x"05",
          5381 => x"93",
          5382 => x"a4",
          5383 => x"fd",
          5384 => x"53",
          5385 => x"80",
          5386 => x"51",
          5387 => x"3f",
          5388 => x"08",
          5389 => x"84",
          5390 => x"39",
          5391 => x"f4",
          5392 => x"f8",
          5393 => x"82",
          5394 => x"cb",
          5395 => x"2e",
          5396 => x"89",
          5397 => x"38",
          5398 => x"f0",
          5399 => x"f8",
          5400 => x"82",
          5401 => x"cb",
          5402 => x"38",
          5403 => x"08",
          5404 => x"81",
          5405 => x"79",
          5406 => x"d0",
          5407 => x"cb",
          5408 => x"79",
          5409 => x"b4",
          5410 => x"d4",
          5411 => x"b5",
          5412 => x"cb",
          5413 => x"93",
          5414 => x"dc",
          5415 => x"b2",
          5416 => x"fb",
          5417 => x"3d",
          5418 => x"51",
          5419 => x"3f",
          5420 => x"08",
          5421 => x"f8",
          5422 => x"fe",
          5423 => x"81",
          5424 => x"a4",
          5425 => x"51",
          5426 => x"80",
          5427 => x"3d",
          5428 => x"51",
          5429 => x"3f",
          5430 => x"08",
          5431 => x"f8",
          5432 => x"fe",
          5433 => x"81",
          5434 => x"b8",
          5435 => x"05",
          5436 => x"ea",
          5437 => x"cb",
          5438 => x"3d",
          5439 => x"52",
          5440 => x"c6",
          5441 => x"90",
          5442 => x"d8",
          5443 => x"80",
          5444 => x"a4",
          5445 => x"06",
          5446 => x"79",
          5447 => x"f5",
          5448 => x"cb",
          5449 => x"2e",
          5450 => x"81",
          5451 => x"51",
          5452 => x"fa",
          5453 => x"3d",
          5454 => x"53",
          5455 => x"51",
          5456 => x"3f",
          5457 => x"08",
          5458 => x"d6",
          5459 => x"fe",
          5460 => x"fe",
          5461 => x"ff",
          5462 => x"81",
          5463 => x"80",
          5464 => x"38",
          5465 => x"ec",
          5466 => x"f8",
          5467 => x"80",
          5468 => x"cb",
          5469 => x"38",
          5470 => x"08",
          5471 => x"90",
          5472 => x"ce",
          5473 => x"5c",
          5474 => x"27",
          5475 => x"59",
          5476 => x"84",
          5477 => x"7a",
          5478 => x"38",
          5479 => x"51",
          5480 => x"b7",
          5481 => x"11",
          5482 => x"05",
          5483 => x"fb",
          5484 => x"a4",
          5485 => x"38",
          5486 => x"33",
          5487 => x"2e",
          5488 => x"c8",
          5489 => x"b3",
          5490 => x"be",
          5491 => x"80",
          5492 => x"81",
          5493 => x"44",
          5494 => x"c8",
          5495 => x"78",
          5496 => x"c8",
          5497 => x"78",
          5498 => x"38",
          5499 => x"08",
          5500 => x"81",
          5501 => x"fc",
          5502 => x"b7",
          5503 => x"11",
          5504 => x"05",
          5505 => x"a3",
          5506 => x"a4",
          5507 => x"38",
          5508 => x"33",
          5509 => x"2e",
          5510 => x"c8",
          5511 => x"b2",
          5512 => x"be",
          5513 => x"80",
          5514 => x"81",
          5515 => x"43",
          5516 => x"c8",
          5517 => x"78",
          5518 => x"c8",
          5519 => x"78",
          5520 => x"38",
          5521 => x"08",
          5522 => x"81",
          5523 => x"88",
          5524 => x"3d",
          5525 => x"53",
          5526 => x"51",
          5527 => x"3f",
          5528 => x"08",
          5529 => x"38",
          5530 => x"59",
          5531 => x"83",
          5532 => x"79",
          5533 => x"38",
          5534 => x"88",
          5535 => x"2e",
          5536 => x"42",
          5537 => x"51",
          5538 => x"3f",
          5539 => x"54",
          5540 => x"52",
          5541 => x"83",
          5542 => x"ac",
          5543 => x"39",
          5544 => x"f4",
          5545 => x"f8",
          5546 => x"fd",
          5547 => x"cb",
          5548 => x"2e",
          5549 => x"b7",
          5550 => x"11",
          5551 => x"05",
          5552 => x"e7",
          5553 => x"a4",
          5554 => x"a5",
          5555 => x"02",
          5556 => x"33",
          5557 => x"81",
          5558 => x"3d",
          5559 => x"53",
          5560 => x"51",
          5561 => x"3f",
          5562 => x"08",
          5563 => x"b2",
          5564 => x"33",
          5565 => x"c5",
          5566 => x"fb",
          5567 => x"f8",
          5568 => x"fe",
          5569 => x"79",
          5570 => x"59",
          5571 => x"f7",
          5572 => x"79",
          5573 => x"b7",
          5574 => x"11",
          5575 => x"05",
          5576 => x"87",
          5577 => x"a4",
          5578 => x"91",
          5579 => x"02",
          5580 => x"33",
          5581 => x"81",
          5582 => x"b5",
          5583 => x"c4",
          5584 => x"8e",
          5585 => x"39",
          5586 => x"e8",
          5587 => x"f8",
          5588 => x"fe",
          5589 => x"cb",
          5590 => x"2e",
          5591 => x"b7",
          5592 => x"11",
          5593 => x"05",
          5594 => x"b1",
          5595 => x"a4",
          5596 => x"a6",
          5597 => x"02",
          5598 => x"79",
          5599 => x"5b",
          5600 => x"b7",
          5601 => x"11",
          5602 => x"05",
          5603 => x"8d",
          5604 => x"a4",
          5605 => x"f6",
          5606 => x"70",
          5607 => x"81",
          5608 => x"fe",
          5609 => x"80",
          5610 => x"51",
          5611 => x"3f",
          5612 => x"33",
          5613 => x"2e",
          5614 => x"78",
          5615 => x"38",
          5616 => x"41",
          5617 => x"3d",
          5618 => x"53",
          5619 => x"51",
          5620 => x"3f",
          5621 => x"08",
          5622 => x"38",
          5623 => x"be",
          5624 => x"70",
          5625 => x"23",
          5626 => x"ae",
          5627 => x"c4",
          5628 => x"de",
          5629 => x"39",
          5630 => x"e8",
          5631 => x"f8",
          5632 => x"fd",
          5633 => x"cb",
          5634 => x"2e",
          5635 => x"b7",
          5636 => x"11",
          5637 => x"05",
          5638 => x"81",
          5639 => x"a4",
          5640 => x"a1",
          5641 => x"71",
          5642 => x"84",
          5643 => x"3d",
          5644 => x"53",
          5645 => x"51",
          5646 => x"3f",
          5647 => x"08",
          5648 => x"de",
          5649 => x"08",
          5650 => x"c5",
          5651 => x"f8",
          5652 => x"f8",
          5653 => x"fe",
          5654 => x"79",
          5655 => x"59",
          5656 => x"f4",
          5657 => x"79",
          5658 => x"b7",
          5659 => x"11",
          5660 => x"05",
          5661 => x"a5",
          5662 => x"a4",
          5663 => x"99",
          5664 => x"60",
          5665 => x"d8",
          5666 => x"aa",
          5667 => x"71",
          5668 => x"84",
          5669 => x"ad",
          5670 => x"c4",
          5671 => x"b2",
          5672 => x"39",
          5673 => x"51",
          5674 => x"3f",
          5675 => x"f1",
          5676 => x"ee",
          5677 => x"fc",
          5678 => x"96",
          5679 => x"fe",
          5680 => x"f3",
          5681 => x"80",
          5682 => x"c0",
          5683 => x"84",
          5684 => x"87",
          5685 => x"0c",
          5686 => x"51",
          5687 => x"3f",
          5688 => x"81",
          5689 => x"fe",
          5690 => x"8c",
          5691 => x"87",
          5692 => x"0c",
          5693 => x"0b",
          5694 => x"94",
          5695 => x"39",
          5696 => x"f4",
          5697 => x"f8",
          5698 => x"f9",
          5699 => x"cb",
          5700 => x"2e",
          5701 => x"63",
          5702 => x"bc",
          5703 => x"96",
          5704 => x"78",
          5705 => x"fe",
          5706 => x"fe",
          5707 => x"fe",
          5708 => x"81",
          5709 => x"80",
          5710 => x"38",
          5711 => x"c6",
          5712 => x"f6",
          5713 => x"59",
          5714 => x"cb",
          5715 => x"81",
          5716 => x"80",
          5717 => x"38",
          5718 => x"08",
          5719 => x"f4",
          5720 => x"d2",
          5721 => x"39",
          5722 => x"51",
          5723 => x"3f",
          5724 => x"3f",
          5725 => x"81",
          5726 => x"fe",
          5727 => x"80",
          5728 => x"39",
          5729 => x"3f",
          5730 => x"64",
          5731 => x"59",
          5732 => x"f2",
          5733 => x"80",
          5734 => x"38",
          5735 => x"80",
          5736 => x"3d",
          5737 => x"51",
          5738 => x"3f",
          5739 => x"56",
          5740 => x"08",
          5741 => x"c4",
          5742 => x"81",
          5743 => x"a3",
          5744 => x"5a",
          5745 => x"3f",
          5746 => x"58",
          5747 => x"57",
          5748 => x"81",
          5749 => x"05",
          5750 => x"81",
          5751 => x"81",
          5752 => x"79",
          5753 => x"3f",
          5754 => x"08",
          5755 => x"32",
          5756 => x"07",
          5757 => x"38",
          5758 => x"09",
          5759 => x"a2",
          5760 => x"d8",
          5761 => x"ae",
          5762 => x"39",
          5763 => x"80",
          5764 => x"d8",
          5765 => x"8d",
          5766 => x"c0",
          5767 => x"b6",
          5768 => x"0b",
          5769 => x"9c",
          5770 => x"83",
          5771 => x"94",
          5772 => x"80",
          5773 => x"c0",
          5774 => x"97",
          5775 => x"cb",
          5776 => x"d2",
          5777 => x"b8",
          5778 => x"af",
          5779 => x"d2",
          5780 => x"e8",
          5781 => x"df",
          5782 => x"f4",
          5783 => x"f2",
          5784 => x"99",
          5785 => x"b5",
          5786 => x"eb",
          5787 => x"e2",
          5788 => x"00",
          5789 => x"f4",
          5790 => x"fa",
          5791 => x"00",
          5792 => x"06",
          5793 => x"0c",
          5794 => x"ca",
          5795 => x"4e",
          5796 => x"55",
          5797 => x"5c",
          5798 => x"63",
          5799 => x"6a",
          5800 => x"71",
          5801 => x"78",
          5802 => x"7f",
          5803 => x"86",
          5804 => x"8d",
          5805 => x"94",
          5806 => x"9a",
          5807 => x"a0",
          5808 => x"a6",
          5809 => x"ac",
          5810 => x"b2",
          5811 => x"b8",
          5812 => x"be",
          5813 => x"c4",
          5814 => x"25",
          5815 => x"64",
          5816 => x"3a",
          5817 => x"25",
          5818 => x"64",
          5819 => x"00",
          5820 => x"20",
          5821 => x"66",
          5822 => x"72",
          5823 => x"6f",
          5824 => x"00",
          5825 => x"72",
          5826 => x"53",
          5827 => x"63",
          5828 => x"69",
          5829 => x"00",
          5830 => x"65",
          5831 => x"65",
          5832 => x"6d",
          5833 => x"6d",
          5834 => x"65",
          5835 => x"00",
          5836 => x"20",
          5837 => x"4e",
          5838 => x"41",
          5839 => x"53",
          5840 => x"74",
          5841 => x"38",
          5842 => x"53",
          5843 => x"3d",
          5844 => x"58",
          5845 => x"00",
          5846 => x"20",
          5847 => x"4d",
          5848 => x"74",
          5849 => x"3d",
          5850 => x"58",
          5851 => x"69",
          5852 => x"25",
          5853 => x"29",
          5854 => x"00",
          5855 => x"20",
          5856 => x"20",
          5857 => x"61",
          5858 => x"25",
          5859 => x"2c",
          5860 => x"7a",
          5861 => x"30",
          5862 => x"2e",
          5863 => x"00",
          5864 => x"20",
          5865 => x"54",
          5866 => x"00",
          5867 => x"20",
          5868 => x"0a",
          5869 => x"00",
          5870 => x"20",
          5871 => x"0a",
          5872 => x"00",
          5873 => x"20",
          5874 => x"43",
          5875 => x"20",
          5876 => x"76",
          5877 => x"73",
          5878 => x"32",
          5879 => x"0a",
          5880 => x"00",
          5881 => x"20",
          5882 => x"45",
          5883 => x"50",
          5884 => x"4f",
          5885 => x"4f",
          5886 => x"52",
          5887 => x"00",
          5888 => x"20",
          5889 => x"45",
          5890 => x"28",
          5891 => x"65",
          5892 => x"25",
          5893 => x"29",
          5894 => x"00",
          5895 => x"72",
          5896 => x"65",
          5897 => x"00",
          5898 => x"20",
          5899 => x"20",
          5900 => x"65",
          5901 => x"65",
          5902 => x"72",
          5903 => x"64",
          5904 => x"73",
          5905 => x"25",
          5906 => x"0a",
          5907 => x"00",
          5908 => x"20",
          5909 => x"20",
          5910 => x"6f",
          5911 => x"53",
          5912 => x"74",
          5913 => x"64",
          5914 => x"73",
          5915 => x"25",
          5916 => x"0a",
          5917 => x"00",
          5918 => x"20",
          5919 => x"63",
          5920 => x"74",
          5921 => x"20",
          5922 => x"72",
          5923 => x"20",
          5924 => x"20",
          5925 => x"25",
          5926 => x"0a",
          5927 => x"00",
          5928 => x"20",
          5929 => x"20",
          5930 => x"20",
          5931 => x"20",
          5932 => x"20",
          5933 => x"20",
          5934 => x"20",
          5935 => x"25",
          5936 => x"0a",
          5937 => x"00",
          5938 => x"20",
          5939 => x"74",
          5940 => x"43",
          5941 => x"6b",
          5942 => x"65",
          5943 => x"20",
          5944 => x"20",
          5945 => x"25",
          5946 => x"0a",
          5947 => x"00",
          5948 => x"6c",
          5949 => x"00",
          5950 => x"69",
          5951 => x"00",
          5952 => x"78",
          5953 => x"00",
          5954 => x"00",
          5955 => x"6d",
          5956 => x"00",
          5957 => x"6e",
          5958 => x"00",
          5959 => x"00",
          5960 => x"2c",
          5961 => x"3d",
          5962 => x"5d",
          5963 => x"00",
          5964 => x"00",
          5965 => x"33",
          5966 => x"00",
          5967 => x"4d",
          5968 => x"53",
          5969 => x"00",
          5970 => x"4e",
          5971 => x"20",
          5972 => x"46",
          5973 => x"32",
          5974 => x"00",
          5975 => x"4e",
          5976 => x"20",
          5977 => x"46",
          5978 => x"20",
          5979 => x"00",
          5980 => x"1c",
          5981 => x"00",
          5982 => x"00",
          5983 => x"00",
          5984 => x"41",
          5985 => x"80",
          5986 => x"49",
          5987 => x"8f",
          5988 => x"4f",
          5989 => x"55",
          5990 => x"9b",
          5991 => x"9f",
          5992 => x"55",
          5993 => x"a7",
          5994 => x"ab",
          5995 => x"af",
          5996 => x"b3",
          5997 => x"b7",
          5998 => x"bb",
          5999 => x"bf",
          6000 => x"c3",
          6001 => x"c7",
          6002 => x"cb",
          6003 => x"cf",
          6004 => x"d3",
          6005 => x"d7",
          6006 => x"db",
          6007 => x"df",
          6008 => x"e3",
          6009 => x"e7",
          6010 => x"eb",
          6011 => x"ef",
          6012 => x"f3",
          6013 => x"f7",
          6014 => x"fb",
          6015 => x"ff",
          6016 => x"3b",
          6017 => x"2f",
          6018 => x"3a",
          6019 => x"7c",
          6020 => x"00",
          6021 => x"04",
          6022 => x"40",
          6023 => x"00",
          6024 => x"00",
          6025 => x"02",
          6026 => x"08",
          6027 => x"20",
          6028 => x"00",
          6029 => x"69",
          6030 => x"00",
          6031 => x"63",
          6032 => x"00",
          6033 => x"69",
          6034 => x"00",
          6035 => x"61",
          6036 => x"00",
          6037 => x"65",
          6038 => x"00",
          6039 => x"65",
          6040 => x"00",
          6041 => x"6d",
          6042 => x"00",
          6043 => x"73",
          6044 => x"00",
          6045 => x"00",
          6046 => x"00",
          6047 => x"00",
          6048 => x"00",
          6049 => x"00",
          6050 => x"00",
          6051 => x"00",
          6052 => x"6c",
          6053 => x"00",
          6054 => x"00",
          6055 => x"74",
          6056 => x"00",
          6057 => x"65",
          6058 => x"00",
          6059 => x"6f",
          6060 => x"00",
          6061 => x"74",
          6062 => x"00",
          6063 => x"6b",
          6064 => x"72",
          6065 => x"00",
          6066 => x"65",
          6067 => x"6c",
          6068 => x"72",
          6069 => x"0a",
          6070 => x"00",
          6071 => x"6b",
          6072 => x"74",
          6073 => x"61",
          6074 => x"0a",
          6075 => x"00",
          6076 => x"66",
          6077 => x"20",
          6078 => x"6e",
          6079 => x"00",
          6080 => x"70",
          6081 => x"20",
          6082 => x"6e",
          6083 => x"00",
          6084 => x"61",
          6085 => x"20",
          6086 => x"65",
          6087 => x"65",
          6088 => x"00",
          6089 => x"65",
          6090 => x"64",
          6091 => x"65",
          6092 => x"00",
          6093 => x"65",
          6094 => x"72",
          6095 => x"79",
          6096 => x"69",
          6097 => x"2e",
          6098 => x"00",
          6099 => x"65",
          6100 => x"6e",
          6101 => x"20",
          6102 => x"61",
          6103 => x"2e",
          6104 => x"00",
          6105 => x"69",
          6106 => x"72",
          6107 => x"20",
          6108 => x"74",
          6109 => x"65",
          6110 => x"00",
          6111 => x"76",
          6112 => x"75",
          6113 => x"72",
          6114 => x"20",
          6115 => x"61",
          6116 => x"2e",
          6117 => x"00",
          6118 => x"6b",
          6119 => x"74",
          6120 => x"61",
          6121 => x"64",
          6122 => x"00",
          6123 => x"63",
          6124 => x"61",
          6125 => x"6c",
          6126 => x"69",
          6127 => x"79",
          6128 => x"6d",
          6129 => x"75",
          6130 => x"6f",
          6131 => x"69",
          6132 => x"0a",
          6133 => x"00",
          6134 => x"6d",
          6135 => x"61",
          6136 => x"74",
          6137 => x"0a",
          6138 => x"00",
          6139 => x"65",
          6140 => x"2c",
          6141 => x"65",
          6142 => x"69",
          6143 => x"63",
          6144 => x"65",
          6145 => x"64",
          6146 => x"00",
          6147 => x"65",
          6148 => x"20",
          6149 => x"6b",
          6150 => x"0a",
          6151 => x"00",
          6152 => x"75",
          6153 => x"63",
          6154 => x"74",
          6155 => x"6d",
          6156 => x"2e",
          6157 => x"00",
          6158 => x"20",
          6159 => x"79",
          6160 => x"65",
          6161 => x"69",
          6162 => x"2e",
          6163 => x"00",
          6164 => x"61",
          6165 => x"65",
          6166 => x"69",
          6167 => x"72",
          6168 => x"74",
          6169 => x"00",
          6170 => x"63",
          6171 => x"2e",
          6172 => x"00",
          6173 => x"6e",
          6174 => x"20",
          6175 => x"6f",
          6176 => x"00",
          6177 => x"75",
          6178 => x"74",
          6179 => x"25",
          6180 => x"74",
          6181 => x"75",
          6182 => x"74",
          6183 => x"73",
          6184 => x"0a",
          6185 => x"00",
          6186 => x"58",
          6187 => x"00",
          6188 => x"00",
          6189 => x"58",
          6190 => x"00",
          6191 => x"20",
          6192 => x"20",
          6193 => x"00",
          6194 => x"58",
          6195 => x"00",
          6196 => x"00",
          6197 => x"00",
          6198 => x"00",
          6199 => x"64",
          6200 => x"00",
          6201 => x"54",
          6202 => x"00",
          6203 => x"20",
          6204 => x"28",
          6205 => x"00",
          6206 => x"30",
          6207 => x"30",
          6208 => x"00",
          6209 => x"33",
          6210 => x"00",
          6211 => x"55",
          6212 => x"65",
          6213 => x"30",
          6214 => x"20",
          6215 => x"25",
          6216 => x"2a",
          6217 => x"00",
          6218 => x"54",
          6219 => x"6e",
          6220 => x"72",
          6221 => x"20",
          6222 => x"64",
          6223 => x"0a",
          6224 => x"00",
          6225 => x"65",
          6226 => x"6e",
          6227 => x"72",
          6228 => x"0a",
          6229 => x"00",
          6230 => x"20",
          6231 => x"65",
          6232 => x"70",
          6233 => x"00",
          6234 => x"54",
          6235 => x"44",
          6236 => x"74",
          6237 => x"75",
          6238 => x"00",
          6239 => x"54",
          6240 => x"52",
          6241 => x"74",
          6242 => x"75",
          6243 => x"00",
          6244 => x"54",
          6245 => x"58",
          6246 => x"74",
          6247 => x"75",
          6248 => x"00",
          6249 => x"54",
          6250 => x"58",
          6251 => x"74",
          6252 => x"75",
          6253 => x"00",
          6254 => x"54",
          6255 => x"58",
          6256 => x"74",
          6257 => x"75",
          6258 => x"00",
          6259 => x"54",
          6260 => x"58",
          6261 => x"74",
          6262 => x"75",
          6263 => x"00",
          6264 => x"74",
          6265 => x"20",
          6266 => x"74",
          6267 => x"72",
          6268 => x"0a",
          6269 => x"00",
          6270 => x"62",
          6271 => x"67",
          6272 => x"6d",
          6273 => x"2e",
          6274 => x"00",
          6275 => x"00",
          6276 => x"6c",
          6277 => x"74",
          6278 => x"6e",
          6279 => x"61",
          6280 => x"65",
          6281 => x"20",
          6282 => x"64",
          6283 => x"20",
          6284 => x"61",
          6285 => x"69",
          6286 => x"20",
          6287 => x"75",
          6288 => x"79",
          6289 => x"00",
          6290 => x"00",
          6291 => x"20",
          6292 => x"6b",
          6293 => x"21",
          6294 => x"00",
          6295 => x"74",
          6296 => x"69",
          6297 => x"2e",
          6298 => x"00",
          6299 => x"6c",
          6300 => x"74",
          6301 => x"6e",
          6302 => x"61",
          6303 => x"65",
          6304 => x"00",
          6305 => x"25",
          6306 => x"00",
          6307 => x"00",
          6308 => x"61",
          6309 => x"67",
          6310 => x"00",
          6311 => x"70",
          6312 => x"6d",
          6313 => x"0a",
          6314 => x"00",
          6315 => x"6d",
          6316 => x"74",
          6317 => x"00",
          6318 => x"58",
          6319 => x"32",
          6320 => x"00",
          6321 => x"0a",
          6322 => x"00",
          6323 => x"58",
          6324 => x"34",
          6325 => x"00",
          6326 => x"58",
          6327 => x"38",
          6328 => x"00",
          6329 => x"61",
          6330 => x"6e",
          6331 => x"6e",
          6332 => x"72",
          6333 => x"73",
          6334 => x"00",
          6335 => x"62",
          6336 => x"67",
          6337 => x"74",
          6338 => x"75",
          6339 => x"0a",
          6340 => x"00",
          6341 => x"61",
          6342 => x"64",
          6343 => x"72",
          6344 => x"69",
          6345 => x"00",
          6346 => x"62",
          6347 => x"67",
          6348 => x"72",
          6349 => x"69",
          6350 => x"00",
          6351 => x"63",
          6352 => x"6e",
          6353 => x"6f",
          6354 => x"40",
          6355 => x"38",
          6356 => x"2e",
          6357 => x"00",
          6358 => x"6c",
          6359 => x"20",
          6360 => x"65",
          6361 => x"25",
          6362 => x"20",
          6363 => x"0a",
          6364 => x"00",
          6365 => x"6c",
          6366 => x"74",
          6367 => x"65",
          6368 => x"6f",
          6369 => x"28",
          6370 => x"2e",
          6371 => x"00",
          6372 => x"74",
          6373 => x"69",
          6374 => x"61",
          6375 => x"69",
          6376 => x"69",
          6377 => x"2e",
          6378 => x"00",
          6379 => x"64",
          6380 => x"62",
          6381 => x"69",
          6382 => x"2e",
          6383 => x"00",
          6384 => x"00",
          6385 => x"00",
          6386 => x"5c",
          6387 => x"25",
          6388 => x"73",
          6389 => x"00",
          6390 => x"20",
          6391 => x"6d",
          6392 => x"2e",
          6393 => x"00",
          6394 => x"6e",
          6395 => x"2e",
          6396 => x"00",
          6397 => x"62",
          6398 => x"67",
          6399 => x"74",
          6400 => x"75",
          6401 => x"2e",
          6402 => x"00",
          6403 => x"00",
          6404 => x"00",
          6405 => x"ff",
          6406 => x"00",
          6407 => x"ff",
          6408 => x"00",
          6409 => x"ff",
          6410 => x"00",
          6411 => x"00",
          6412 => x"00",
          6413 => x"00",
          6414 => x"00",
          6415 => x"01",
          6416 => x"01",
          6417 => x"01",
          6418 => x"00",
          6419 => x"00",
          6420 => x"00",
          6421 => x"34",
          6422 => x"00",
          6423 => x"00",
          6424 => x"00",
          6425 => x"3c",
          6426 => x"00",
          6427 => x"00",
          6428 => x"00",
          6429 => x"44",
          6430 => x"00",
          6431 => x"00",
          6432 => x"00",
          6433 => x"4c",
          6434 => x"00",
          6435 => x"00",
          6436 => x"00",
          6437 => x"54",
          6438 => x"00",
          6439 => x"00",
          6440 => x"00",
          6441 => x"5c",
          6442 => x"00",
          6443 => x"00",
          6444 => x"00",
          6445 => x"64",
          6446 => x"00",
          6447 => x"00",
          6448 => x"00",
          6449 => x"6c",
          6450 => x"00",
          6451 => x"00",
          6452 => x"00",
          6453 => x"74",
          6454 => x"00",
          6455 => x"00",
          6456 => x"00",
          6457 => x"78",
          6458 => x"00",
          6459 => x"00",
          6460 => x"00",
          6461 => x"7c",
          6462 => x"00",
          6463 => x"00",
          6464 => x"00",
          6465 => x"80",
          6466 => x"00",
          6467 => x"00",
          6468 => x"00",
          6469 => x"84",
          6470 => x"00",
          6471 => x"00",
          6472 => x"00",
          6473 => x"88",
          6474 => x"00",
          6475 => x"00",
          6476 => x"00",
          6477 => x"8c",
          6478 => x"00",
          6479 => x"00",
          6480 => x"00",
          6481 => x"90",
          6482 => x"00",
          6483 => x"00",
          6484 => x"00",
          6485 => x"98",
          6486 => x"00",
          6487 => x"00",
          6488 => x"00",
          6489 => x"9c",
          6490 => x"00",
          6491 => x"00",
          6492 => x"00",
          6493 => x"a4",
          6494 => x"00",
          6495 => x"00",
          6496 => x"00",
          6497 => x"ac",
          6498 => x"00",
          6499 => x"00",
          6500 => x"00",
          6501 => x"b4",
          6502 => x"00",
          6503 => x"00",
          6504 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"fd",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"0b",
            10 => x"84",
            11 => x"0b",
            12 => x"0b",
            13 => x"a2",
            14 => x"0b",
            15 => x"0b",
            16 => x"c0",
            17 => x"0b",
            18 => x"0b",
            19 => x"de",
            20 => x"0b",
            21 => x"0b",
            22 => x"fc",
            23 => x"0b",
            24 => x"0b",
            25 => x"9a",
            26 => x"0b",
            27 => x"0b",
            28 => x"b8",
            29 => x"0b",
            30 => x"0b",
            31 => x"d6",
            32 => x"0b",
            33 => x"0b",
            34 => x"f4",
            35 => x"0b",
            36 => x"0b",
            37 => x"93",
            38 => x"0b",
            39 => x"0b",
            40 => x"b3",
            41 => x"0b",
            42 => x"0b",
            43 => x"d3",
            44 => x"0b",
            45 => x"0b",
            46 => x"f3",
            47 => x"0b",
            48 => x"0b",
            49 => x"93",
            50 => x"0b",
            51 => x"0b",
            52 => x"b3",
            53 => x"0b",
            54 => x"0b",
            55 => x"d3",
            56 => x"0b",
            57 => x"0b",
            58 => x"f3",
            59 => x"0b",
            60 => x"0b",
            61 => x"93",
            62 => x"0b",
            63 => x"0b",
            64 => x"b3",
            65 => x"0b",
            66 => x"0b",
            67 => x"d3",
            68 => x"0b",
            69 => x"0b",
            70 => x"f3",
            71 => x"0b",
            72 => x"0b",
            73 => x"93",
            74 => x"0b",
            75 => x"0b",
            76 => x"b1",
            77 => x"0b",
            78 => x"0b",
            79 => x"cf",
            80 => x"0b",
            81 => x"0b",
            82 => x"ed",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"00",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"00",
           137 => x"00",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"00",
           145 => x"00",
           146 => x"00",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"00",
           153 => x"00",
           154 => x"00",
           155 => x"00",
           156 => x"00",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"00",
           161 => x"00",
           162 => x"00",
           163 => x"00",
           164 => x"00",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"00",
           169 => x"00",
           170 => x"00",
           171 => x"00",
           172 => x"00",
           173 => x"00",
           174 => x"00",
           175 => x"00",
           176 => x"00",
           177 => x"00",
           178 => x"00",
           179 => x"00",
           180 => x"00",
           181 => x"00",
           182 => x"00",
           183 => x"00",
           184 => x"00",
           185 => x"00",
           186 => x"00",
           187 => x"00",
           188 => x"00",
           189 => x"00",
           190 => x"00",
           191 => x"00",
           192 => x"00",
           193 => x"00",
           194 => x"00",
           195 => x"00",
           196 => x"00",
           197 => x"00",
           198 => x"00",
           199 => x"00",
           200 => x"00",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"00",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"00",
           233 => x"00",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"00",
           249 => x"00",
           250 => x"00",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"80",
           257 => x"b0",
           258 => x"2d",
           259 => x"08",
           260 => x"04",
           261 => x"0c",
           262 => x"81",
           263 => x"81",
           264 => x"81",
           265 => x"a3",
           266 => x"cb",
           267 => x"e4",
           268 => x"cb",
           269 => x"d2",
           270 => x"b0",
           271 => x"90",
           272 => x"b0",
           273 => x"2d",
           274 => x"08",
           275 => x"04",
           276 => x"0c",
           277 => x"81",
           278 => x"81",
           279 => x"81",
           280 => x"a3",
           281 => x"cb",
           282 => x"e4",
           283 => x"cb",
           284 => x"ab",
           285 => x"b0",
           286 => x"90",
           287 => x"b0",
           288 => x"2d",
           289 => x"08",
           290 => x"04",
           291 => x"0c",
           292 => x"81",
           293 => x"81",
           294 => x"81",
           295 => x"a9",
           296 => x"cb",
           297 => x"e4",
           298 => x"cb",
           299 => x"f0",
           300 => x"b0",
           301 => x"90",
           302 => x"b0",
           303 => x"2d",
           304 => x"08",
           305 => x"04",
           306 => x"0c",
           307 => x"81",
           308 => x"81",
           309 => x"81",
           310 => x"93",
           311 => x"cb",
           312 => x"e4",
           313 => x"cb",
           314 => x"f4",
           315 => x"b0",
           316 => x"90",
           317 => x"b0",
           318 => x"2d",
           319 => x"08",
           320 => x"04",
           321 => x"0c",
           322 => x"2d",
           323 => x"08",
           324 => x"04",
           325 => x"0c",
           326 => x"2d",
           327 => x"08",
           328 => x"04",
           329 => x"0c",
           330 => x"2d",
           331 => x"08",
           332 => x"04",
           333 => x"0c",
           334 => x"2d",
           335 => x"08",
           336 => x"04",
           337 => x"0c",
           338 => x"2d",
           339 => x"08",
           340 => x"04",
           341 => x"0c",
           342 => x"2d",
           343 => x"08",
           344 => x"04",
           345 => x"0c",
           346 => x"2d",
           347 => x"08",
           348 => x"04",
           349 => x"0c",
           350 => x"2d",
           351 => x"08",
           352 => x"04",
           353 => x"0c",
           354 => x"2d",
           355 => x"08",
           356 => x"04",
           357 => x"0c",
           358 => x"2d",
           359 => x"08",
           360 => x"04",
           361 => x"0c",
           362 => x"2d",
           363 => x"08",
           364 => x"04",
           365 => x"0c",
           366 => x"2d",
           367 => x"08",
           368 => x"04",
           369 => x"0c",
           370 => x"2d",
           371 => x"08",
           372 => x"04",
           373 => x"0c",
           374 => x"2d",
           375 => x"08",
           376 => x"04",
           377 => x"0c",
           378 => x"2d",
           379 => x"08",
           380 => x"04",
           381 => x"0c",
           382 => x"2d",
           383 => x"08",
           384 => x"04",
           385 => x"0c",
           386 => x"2d",
           387 => x"08",
           388 => x"04",
           389 => x"0c",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"2d",
           407 => x"08",
           408 => x"04",
           409 => x"0c",
           410 => x"2d",
           411 => x"08",
           412 => x"04",
           413 => x"0c",
           414 => x"2d",
           415 => x"08",
           416 => x"04",
           417 => x"0c",
           418 => x"2d",
           419 => x"08",
           420 => x"04",
           421 => x"0c",
           422 => x"81",
           423 => x"81",
           424 => x"81",
           425 => x"b2",
           426 => x"cb",
           427 => x"e4",
           428 => x"cb",
           429 => x"fa",
           430 => x"b0",
           431 => x"90",
           432 => x"b0",
           433 => x"2d",
           434 => x"08",
           435 => x"04",
           436 => x"0c",
           437 => x"81",
           438 => x"81",
           439 => x"81",
           440 => x"97",
           441 => x"cb",
           442 => x"e4",
           443 => x"cb",
           444 => x"9a",
           445 => x"cb",
           446 => x"e4",
           447 => x"cb",
           448 => x"e2",
           449 => x"38",
           450 => x"84",
           451 => x"0b",
           452 => x"80",
           453 => x"51",
           454 => x"04",
           455 => x"cb",
           456 => x"81",
           457 => x"fd",
           458 => x"53",
           459 => x"08",
           460 => x"52",
           461 => x"08",
           462 => x"51",
           463 => x"81",
           464 => x"70",
           465 => x"0c",
           466 => x"0d",
           467 => x"0c",
           468 => x"b0",
           469 => x"cb",
           470 => x"3d",
           471 => x"81",
           472 => x"8c",
           473 => x"81",
           474 => x"88",
           475 => x"93",
           476 => x"a4",
           477 => x"cb",
           478 => x"85",
           479 => x"cb",
           480 => x"81",
           481 => x"02",
           482 => x"0c",
           483 => x"81",
           484 => x"b0",
           485 => x"0c",
           486 => x"cb",
           487 => x"05",
           488 => x"b0",
           489 => x"08",
           490 => x"08",
           491 => x"27",
           492 => x"cb",
           493 => x"05",
           494 => x"ae",
           495 => x"81",
           496 => x"8c",
           497 => x"a2",
           498 => x"b0",
           499 => x"08",
           500 => x"b0",
           501 => x"0c",
           502 => x"08",
           503 => x"10",
           504 => x"08",
           505 => x"ff",
           506 => x"cb",
           507 => x"05",
           508 => x"80",
           509 => x"cb",
           510 => x"05",
           511 => x"b0",
           512 => x"08",
           513 => x"81",
           514 => x"88",
           515 => x"cb",
           516 => x"05",
           517 => x"cb",
           518 => x"05",
           519 => x"b0",
           520 => x"08",
           521 => x"08",
           522 => x"07",
           523 => x"08",
           524 => x"81",
           525 => x"fc",
           526 => x"2a",
           527 => x"08",
           528 => x"81",
           529 => x"8c",
           530 => x"2a",
           531 => x"08",
           532 => x"ff",
           533 => x"cb",
           534 => x"05",
           535 => x"93",
           536 => x"b0",
           537 => x"08",
           538 => x"b0",
           539 => x"0c",
           540 => x"81",
           541 => x"f8",
           542 => x"81",
           543 => x"f4",
           544 => x"81",
           545 => x"f4",
           546 => x"cb",
           547 => x"3d",
           548 => x"b0",
           549 => x"3d",
           550 => x"71",
           551 => x"9f",
           552 => x"55",
           553 => x"72",
           554 => x"74",
           555 => x"70",
           556 => x"38",
           557 => x"71",
           558 => x"38",
           559 => x"81",
           560 => x"ff",
           561 => x"ff",
           562 => x"06",
           563 => x"81",
           564 => x"86",
           565 => x"74",
           566 => x"75",
           567 => x"90",
           568 => x"54",
           569 => x"27",
           570 => x"71",
           571 => x"53",
           572 => x"70",
           573 => x"0c",
           574 => x"84",
           575 => x"72",
           576 => x"05",
           577 => x"12",
           578 => x"26",
           579 => x"72",
           580 => x"72",
           581 => x"05",
           582 => x"12",
           583 => x"26",
           584 => x"53",
           585 => x"fb",
           586 => x"79",
           587 => x"83",
           588 => x"52",
           589 => x"71",
           590 => x"54",
           591 => x"73",
           592 => x"c6",
           593 => x"54",
           594 => x"70",
           595 => x"52",
           596 => x"2e",
           597 => x"33",
           598 => x"2e",
           599 => x"95",
           600 => x"81",
           601 => x"70",
           602 => x"54",
           603 => x"70",
           604 => x"33",
           605 => x"ff",
           606 => x"ff",
           607 => x"31",
           608 => x"0c",
           609 => x"3d",
           610 => x"09",
           611 => x"fd",
           612 => x"70",
           613 => x"81",
           614 => x"51",
           615 => x"38",
           616 => x"16",
           617 => x"56",
           618 => x"08",
           619 => x"73",
           620 => x"ff",
           621 => x"0b",
           622 => x"0c",
           623 => x"04",
           624 => x"80",
           625 => x"71",
           626 => x"87",
           627 => x"cb",
           628 => x"ff",
           629 => x"ff",
           630 => x"72",
           631 => x"38",
           632 => x"a4",
           633 => x"0d",
           634 => x"0d",
           635 => x"70",
           636 => x"71",
           637 => x"ca",
           638 => x"51",
           639 => x"09",
           640 => x"38",
           641 => x"f1",
           642 => x"84",
           643 => x"53",
           644 => x"70",
           645 => x"53",
           646 => x"a0",
           647 => x"81",
           648 => x"2e",
           649 => x"e5",
           650 => x"ff",
           651 => x"a0",
           652 => x"06",
           653 => x"73",
           654 => x"55",
           655 => x"0c",
           656 => x"81",
           657 => x"87",
           658 => x"fc",
           659 => x"53",
           660 => x"2e",
           661 => x"3d",
           662 => x"72",
           663 => x"3f",
           664 => x"08",
           665 => x"53",
           666 => x"53",
           667 => x"a4",
           668 => x"0d",
           669 => x"0d",
           670 => x"33",
           671 => x"53",
           672 => x"8b",
           673 => x"38",
           674 => x"ff",
           675 => x"52",
           676 => x"81",
           677 => x"13",
           678 => x"52",
           679 => x"80",
           680 => x"13",
           681 => x"52",
           682 => x"80",
           683 => x"13",
           684 => x"52",
           685 => x"80",
           686 => x"13",
           687 => x"52",
           688 => x"26",
           689 => x"8a",
           690 => x"87",
           691 => x"e7",
           692 => x"38",
           693 => x"c0",
           694 => x"72",
           695 => x"98",
           696 => x"13",
           697 => x"98",
           698 => x"13",
           699 => x"98",
           700 => x"13",
           701 => x"98",
           702 => x"13",
           703 => x"98",
           704 => x"13",
           705 => x"98",
           706 => x"87",
           707 => x"0c",
           708 => x"98",
           709 => x"0b",
           710 => x"9c",
           711 => x"71",
           712 => x"0c",
           713 => x"04",
           714 => x"7f",
           715 => x"98",
           716 => x"7d",
           717 => x"98",
           718 => x"7d",
           719 => x"c0",
           720 => x"5a",
           721 => x"34",
           722 => x"b4",
           723 => x"83",
           724 => x"c0",
           725 => x"5a",
           726 => x"34",
           727 => x"ac",
           728 => x"85",
           729 => x"c0",
           730 => x"5a",
           731 => x"34",
           732 => x"a4",
           733 => x"88",
           734 => x"c0",
           735 => x"5a",
           736 => x"23",
           737 => x"79",
           738 => x"06",
           739 => x"ff",
           740 => x"86",
           741 => x"85",
           742 => x"84",
           743 => x"83",
           744 => x"82",
           745 => x"7d",
           746 => x"06",
           747 => x"d8",
           748 => x"3f",
           749 => x"04",
           750 => x"02",
           751 => x"70",
           752 => x"2a",
           753 => x"70",
           754 => x"c8",
           755 => x"3d",
           756 => x"3d",
           757 => x"0b",
           758 => x"33",
           759 => x"06",
           760 => x"87",
           761 => x"51",
           762 => x"86",
           763 => x"94",
           764 => x"08",
           765 => x"70",
           766 => x"54",
           767 => x"2e",
           768 => x"91",
           769 => x"06",
           770 => x"d7",
           771 => x"32",
           772 => x"51",
           773 => x"2e",
           774 => x"93",
           775 => x"06",
           776 => x"ff",
           777 => x"81",
           778 => x"87",
           779 => x"52",
           780 => x"86",
           781 => x"94",
           782 => x"72",
           783 => x"cb",
           784 => x"3d",
           785 => x"3d",
           786 => x"05",
           787 => x"81",
           788 => x"70",
           789 => x"57",
           790 => x"c0",
           791 => x"74",
           792 => x"38",
           793 => x"94",
           794 => x"70",
           795 => x"81",
           796 => x"52",
           797 => x"8c",
           798 => x"2a",
           799 => x"51",
           800 => x"38",
           801 => x"70",
           802 => x"51",
           803 => x"8d",
           804 => x"2a",
           805 => x"51",
           806 => x"be",
           807 => x"ff",
           808 => x"c0",
           809 => x"70",
           810 => x"38",
           811 => x"90",
           812 => x"0c",
           813 => x"04",
           814 => x"79",
           815 => x"33",
           816 => x"06",
           817 => x"70",
           818 => x"fe",
           819 => x"ff",
           820 => x"0b",
           821 => x"8c",
           822 => x"ff",
           823 => x"55",
           824 => x"94",
           825 => x"80",
           826 => x"87",
           827 => x"51",
           828 => x"96",
           829 => x"06",
           830 => x"70",
           831 => x"38",
           832 => x"70",
           833 => x"51",
           834 => x"72",
           835 => x"81",
           836 => x"70",
           837 => x"38",
           838 => x"70",
           839 => x"51",
           840 => x"38",
           841 => x"06",
           842 => x"94",
           843 => x"80",
           844 => x"87",
           845 => x"52",
           846 => x"81",
           847 => x"70",
           848 => x"53",
           849 => x"ff",
           850 => x"81",
           851 => x"89",
           852 => x"fe",
           853 => x"0b",
           854 => x"33",
           855 => x"06",
           856 => x"c0",
           857 => x"72",
           858 => x"38",
           859 => x"94",
           860 => x"70",
           861 => x"81",
           862 => x"51",
           863 => x"e2",
           864 => x"ff",
           865 => x"c0",
           866 => x"70",
           867 => x"38",
           868 => x"90",
           869 => x"70",
           870 => x"81",
           871 => x"51",
           872 => x"04",
           873 => x"0b",
           874 => x"8c",
           875 => x"ff",
           876 => x"87",
           877 => x"52",
           878 => x"86",
           879 => x"94",
           880 => x"08",
           881 => x"70",
           882 => x"51",
           883 => x"70",
           884 => x"38",
           885 => x"06",
           886 => x"94",
           887 => x"80",
           888 => x"87",
           889 => x"52",
           890 => x"98",
           891 => x"2c",
           892 => x"71",
           893 => x"0c",
           894 => x"04",
           895 => x"87",
           896 => x"08",
           897 => x"8a",
           898 => x"70",
           899 => x"93",
           900 => x"9e",
           901 => x"c8",
           902 => x"c0",
           903 => x"81",
           904 => x"87",
           905 => x"08",
           906 => x"0c",
           907 => x"90",
           908 => x"9c",
           909 => x"9e",
           910 => x"c8",
           911 => x"c0",
           912 => x"81",
           913 => x"87",
           914 => x"08",
           915 => x"0c",
           916 => x"a8",
           917 => x"ac",
           918 => x"9e",
           919 => x"c8",
           920 => x"c0",
           921 => x"51",
           922 => x"b4",
           923 => x"9e",
           924 => x"c8",
           925 => x"0b",
           926 => x"34",
           927 => x"c0",
           928 => x"70",
           929 => x"51",
           930 => x"80",
           931 => x"81",
           932 => x"c8",
           933 => x"0b",
           934 => x"88",
           935 => x"80",
           936 => x"52",
           937 => x"2e",
           938 => x"52",
           939 => x"be",
           940 => x"87",
           941 => x"08",
           942 => x"80",
           943 => x"52",
           944 => x"83",
           945 => x"71",
           946 => x"34",
           947 => x"c0",
           948 => x"70",
           949 => x"51",
           950 => x"80",
           951 => x"81",
           952 => x"c8",
           953 => x"0b",
           954 => x"88",
           955 => x"80",
           956 => x"52",
           957 => x"83",
           958 => x"71",
           959 => x"34",
           960 => x"c0",
           961 => x"70",
           962 => x"51",
           963 => x"80",
           964 => x"81",
           965 => x"c8",
           966 => x"0b",
           967 => x"88",
           968 => x"80",
           969 => x"52",
           970 => x"83",
           971 => x"71",
           972 => x"34",
           973 => x"c0",
           974 => x"70",
           975 => x"51",
           976 => x"80",
           977 => x"81",
           978 => x"c8",
           979 => x"c0",
           980 => x"70",
           981 => x"70",
           982 => x"51",
           983 => x"c8",
           984 => x"0b",
           985 => x"88",
           986 => x"06",
           987 => x"70",
           988 => x"38",
           989 => x"81",
           990 => x"80",
           991 => x"9e",
           992 => x"88",
           993 => x"52",
           994 => x"83",
           995 => x"71",
           996 => x"34",
           997 => x"88",
           998 => x"06",
           999 => x"81",
          1000 => x"83",
          1001 => x"fd",
          1002 => x"b5",
          1003 => x"a3",
          1004 => x"bc",
          1005 => x"80",
          1006 => x"81",
          1007 => x"84",
          1008 => x"b6",
          1009 => x"8b",
          1010 => x"bd",
          1011 => x"80",
          1012 => x"81",
          1013 => x"53",
          1014 => x"08",
          1015 => x"b0",
          1016 => x"3f",
          1017 => x"33",
          1018 => x"2e",
          1019 => x"c8",
          1020 => x"81",
          1021 => x"52",
          1022 => x"51",
          1023 => x"81",
          1024 => x"54",
          1025 => x"81",
          1026 => x"54",
          1027 => x"92",
          1028 => x"a4",
          1029 => x"c8",
          1030 => x"81",
          1031 => x"89",
          1032 => x"c8",
          1033 => x"73",
          1034 => x"38",
          1035 => x"51",
          1036 => x"81",
          1037 => x"54",
          1038 => x"88",
          1039 => x"ac",
          1040 => x"3f",
          1041 => x"33",
          1042 => x"2e",
          1043 => x"b7",
          1044 => x"ff",
          1045 => x"c4",
          1046 => x"80",
          1047 => x"81",
          1048 => x"52",
          1049 => x"51",
          1050 => x"81",
          1051 => x"54",
          1052 => x"88",
          1053 => x"e4",
          1054 => x"3f",
          1055 => x"33",
          1056 => x"2e",
          1057 => x"c8",
          1058 => x"81",
          1059 => x"88",
          1060 => x"b8",
          1061 => x"bb",
          1062 => x"a8",
          1063 => x"b8",
          1064 => x"93",
          1065 => x"ac",
          1066 => x"b8",
          1067 => x"87",
          1068 => x"b0",
          1069 => x"b8",
          1070 => x"fb",
          1071 => x"b4",
          1072 => x"b9",
          1073 => x"ef",
          1074 => x"b8",
          1075 => x"b9",
          1076 => x"e3",
          1077 => x"0d",
          1078 => x"0d",
          1079 => x"33",
          1080 => x"71",
          1081 => x"38",
          1082 => x"0b",
          1083 => x"f4",
          1084 => x"08",
          1085 => x"f0",
          1086 => x"81",
          1087 => x"97",
          1088 => x"80",
          1089 => x"81",
          1090 => x"8b",
          1091 => x"8c",
          1092 => x"81",
          1093 => x"f7",
          1094 => x"3d",
          1095 => x"88",
          1096 => x"80",
          1097 => x"96",
          1098 => x"ff",
          1099 => x"c0",
          1100 => x"08",
          1101 => x"72",
          1102 => x"07",
          1103 => x"cc",
          1104 => x"83",
          1105 => x"ff",
          1106 => x"c0",
          1107 => x"08",
          1108 => x"0c",
          1109 => x"0c",
          1110 => x"81",
          1111 => x"06",
          1112 => x"cc",
          1113 => x"51",
          1114 => x"04",
          1115 => x"08",
          1116 => x"84",
          1117 => x"3d",
          1118 => x"05",
          1119 => x"8a",
          1120 => x"06",
          1121 => x"51",
          1122 => x"cb",
          1123 => x"71",
          1124 => x"38",
          1125 => x"81",
          1126 => x"81",
          1127 => x"bc",
          1128 => x"81",
          1129 => x"52",
          1130 => x"85",
          1131 => x"71",
          1132 => x"0d",
          1133 => x"0d",
          1134 => x"33",
          1135 => x"08",
          1136 => x"b4",
          1137 => x"ff",
          1138 => x"81",
          1139 => x"84",
          1140 => x"fd",
          1141 => x"54",
          1142 => x"81",
          1143 => x"53",
          1144 => x"8e",
          1145 => x"ff",
          1146 => x"14",
          1147 => x"3f",
          1148 => x"3d",
          1149 => x"3d",
          1150 => x"cb",
          1151 => x"81",
          1152 => x"56",
          1153 => x"70",
          1154 => x"53",
          1155 => x"2e",
          1156 => x"81",
          1157 => x"81",
          1158 => x"da",
          1159 => x"74",
          1160 => x"0c",
          1161 => x"04",
          1162 => x"66",
          1163 => x"78",
          1164 => x"5a",
          1165 => x"80",
          1166 => x"38",
          1167 => x"09",
          1168 => x"de",
          1169 => x"7a",
          1170 => x"5c",
          1171 => x"5b",
          1172 => x"09",
          1173 => x"38",
          1174 => x"39",
          1175 => x"09",
          1176 => x"38",
          1177 => x"70",
          1178 => x"33",
          1179 => x"2e",
          1180 => x"92",
          1181 => x"19",
          1182 => x"70",
          1183 => x"33",
          1184 => x"53",
          1185 => x"16",
          1186 => x"26",
          1187 => x"88",
          1188 => x"05",
          1189 => x"05",
          1190 => x"05",
          1191 => x"5b",
          1192 => x"80",
          1193 => x"30",
          1194 => x"80",
          1195 => x"cc",
          1196 => x"70",
          1197 => x"25",
          1198 => x"54",
          1199 => x"53",
          1200 => x"8c",
          1201 => x"07",
          1202 => x"05",
          1203 => x"5a",
          1204 => x"83",
          1205 => x"54",
          1206 => x"27",
          1207 => x"16",
          1208 => x"06",
          1209 => x"80",
          1210 => x"aa",
          1211 => x"cf",
          1212 => x"73",
          1213 => x"81",
          1214 => x"80",
          1215 => x"38",
          1216 => x"2e",
          1217 => x"81",
          1218 => x"80",
          1219 => x"8a",
          1220 => x"39",
          1221 => x"2e",
          1222 => x"73",
          1223 => x"8a",
          1224 => x"d3",
          1225 => x"80",
          1226 => x"80",
          1227 => x"ee",
          1228 => x"39",
          1229 => x"71",
          1230 => x"53",
          1231 => x"54",
          1232 => x"2e",
          1233 => x"15",
          1234 => x"33",
          1235 => x"72",
          1236 => x"81",
          1237 => x"39",
          1238 => x"56",
          1239 => x"27",
          1240 => x"51",
          1241 => x"75",
          1242 => x"72",
          1243 => x"38",
          1244 => x"df",
          1245 => x"16",
          1246 => x"7b",
          1247 => x"38",
          1248 => x"f2",
          1249 => x"77",
          1250 => x"12",
          1251 => x"53",
          1252 => x"5c",
          1253 => x"5c",
          1254 => x"5c",
          1255 => x"5c",
          1256 => x"51",
          1257 => x"fd",
          1258 => x"82",
          1259 => x"06",
          1260 => x"80",
          1261 => x"77",
          1262 => x"53",
          1263 => x"18",
          1264 => x"72",
          1265 => x"c4",
          1266 => x"70",
          1267 => x"25",
          1268 => x"55",
          1269 => x"8d",
          1270 => x"2e",
          1271 => x"30",
          1272 => x"5b",
          1273 => x"8f",
          1274 => x"7b",
          1275 => x"e6",
          1276 => x"cb",
          1277 => x"ff",
          1278 => x"75",
          1279 => x"9e",
          1280 => x"a4",
          1281 => x"74",
          1282 => x"a7",
          1283 => x"80",
          1284 => x"38",
          1285 => x"72",
          1286 => x"54",
          1287 => x"72",
          1288 => x"05",
          1289 => x"17",
          1290 => x"77",
          1291 => x"51",
          1292 => x"9f",
          1293 => x"72",
          1294 => x"79",
          1295 => x"81",
          1296 => x"72",
          1297 => x"38",
          1298 => x"05",
          1299 => x"ad",
          1300 => x"17",
          1301 => x"81",
          1302 => x"b0",
          1303 => x"38",
          1304 => x"81",
          1305 => x"06",
          1306 => x"9f",
          1307 => x"55",
          1308 => x"97",
          1309 => x"f9",
          1310 => x"81",
          1311 => x"8b",
          1312 => x"16",
          1313 => x"73",
          1314 => x"96",
          1315 => x"e0",
          1316 => x"17",
          1317 => x"33",
          1318 => x"f9",
          1319 => x"f2",
          1320 => x"16",
          1321 => x"7b",
          1322 => x"38",
          1323 => x"c6",
          1324 => x"96",
          1325 => x"fd",
          1326 => x"3d",
          1327 => x"05",
          1328 => x"52",
          1329 => x"e0",
          1330 => x"0d",
          1331 => x"0d",
          1332 => x"bc",
          1333 => x"88",
          1334 => x"51",
          1335 => x"81",
          1336 => x"53",
          1337 => x"80",
          1338 => x"bc",
          1339 => x"0d",
          1340 => x"0d",
          1341 => x"08",
          1342 => x"b4",
          1343 => x"88",
          1344 => x"52",
          1345 => x"3f",
          1346 => x"b4",
          1347 => x"0d",
          1348 => x"0d",
          1349 => x"cb",
          1350 => x"56",
          1351 => x"80",
          1352 => x"2e",
          1353 => x"81",
          1354 => x"52",
          1355 => x"cb",
          1356 => x"ff",
          1357 => x"80",
          1358 => x"38",
          1359 => x"b9",
          1360 => x"32",
          1361 => x"80",
          1362 => x"52",
          1363 => x"8b",
          1364 => x"2e",
          1365 => x"14",
          1366 => x"9f",
          1367 => x"38",
          1368 => x"73",
          1369 => x"38",
          1370 => x"72",
          1371 => x"14",
          1372 => x"f8",
          1373 => x"af",
          1374 => x"52",
          1375 => x"8a",
          1376 => x"3f",
          1377 => x"81",
          1378 => x"87",
          1379 => x"fe",
          1380 => x"cb",
          1381 => x"81",
          1382 => x"77",
          1383 => x"53",
          1384 => x"72",
          1385 => x"0c",
          1386 => x"04",
          1387 => x"7a",
          1388 => x"80",
          1389 => x"58",
          1390 => x"33",
          1391 => x"a0",
          1392 => x"06",
          1393 => x"13",
          1394 => x"39",
          1395 => x"09",
          1396 => x"38",
          1397 => x"11",
          1398 => x"08",
          1399 => x"54",
          1400 => x"2e",
          1401 => x"80",
          1402 => x"08",
          1403 => x"0c",
          1404 => x"33",
          1405 => x"80",
          1406 => x"38",
          1407 => x"80",
          1408 => x"38",
          1409 => x"57",
          1410 => x"0c",
          1411 => x"33",
          1412 => x"39",
          1413 => x"74",
          1414 => x"38",
          1415 => x"80",
          1416 => x"89",
          1417 => x"38",
          1418 => x"d0",
          1419 => x"55",
          1420 => x"80",
          1421 => x"39",
          1422 => x"d9",
          1423 => x"80",
          1424 => x"27",
          1425 => x"80",
          1426 => x"89",
          1427 => x"70",
          1428 => x"55",
          1429 => x"70",
          1430 => x"55",
          1431 => x"27",
          1432 => x"14",
          1433 => x"06",
          1434 => x"74",
          1435 => x"73",
          1436 => x"38",
          1437 => x"14",
          1438 => x"05",
          1439 => x"08",
          1440 => x"54",
          1441 => x"39",
          1442 => x"84",
          1443 => x"55",
          1444 => x"81",
          1445 => x"cb",
          1446 => x"3d",
          1447 => x"3d",
          1448 => x"5a",
          1449 => x"7a",
          1450 => x"08",
          1451 => x"53",
          1452 => x"09",
          1453 => x"38",
          1454 => x"0c",
          1455 => x"ad",
          1456 => x"06",
          1457 => x"76",
          1458 => x"0c",
          1459 => x"33",
          1460 => x"73",
          1461 => x"81",
          1462 => x"38",
          1463 => x"05",
          1464 => x"08",
          1465 => x"53",
          1466 => x"2e",
          1467 => x"57",
          1468 => x"2e",
          1469 => x"39",
          1470 => x"13",
          1471 => x"08",
          1472 => x"53",
          1473 => x"55",
          1474 => x"80",
          1475 => x"14",
          1476 => x"88",
          1477 => x"27",
          1478 => x"eb",
          1479 => x"53",
          1480 => x"89",
          1481 => x"38",
          1482 => x"55",
          1483 => x"8a",
          1484 => x"a0",
          1485 => x"c2",
          1486 => x"74",
          1487 => x"e0",
          1488 => x"ff",
          1489 => x"d0",
          1490 => x"ff",
          1491 => x"90",
          1492 => x"38",
          1493 => x"81",
          1494 => x"53",
          1495 => x"ca",
          1496 => x"27",
          1497 => x"77",
          1498 => x"08",
          1499 => x"0c",
          1500 => x"33",
          1501 => x"ff",
          1502 => x"80",
          1503 => x"74",
          1504 => x"79",
          1505 => x"74",
          1506 => x"0c",
          1507 => x"04",
          1508 => x"02",
          1509 => x"51",
          1510 => x"72",
          1511 => x"81",
          1512 => x"33",
          1513 => x"cb",
          1514 => x"3d",
          1515 => x"3d",
          1516 => x"05",
          1517 => x"05",
          1518 => x"56",
          1519 => x"72",
          1520 => x"e0",
          1521 => x"2b",
          1522 => x"8c",
          1523 => x"88",
          1524 => x"2e",
          1525 => x"88",
          1526 => x"0c",
          1527 => x"8c",
          1528 => x"71",
          1529 => x"87",
          1530 => x"0c",
          1531 => x"08",
          1532 => x"51",
          1533 => x"2e",
          1534 => x"c0",
          1535 => x"51",
          1536 => x"71",
          1537 => x"80",
          1538 => x"92",
          1539 => x"98",
          1540 => x"70",
          1541 => x"38",
          1542 => x"d0",
          1543 => x"c8",
          1544 => x"51",
          1545 => x"a4",
          1546 => x"0d",
          1547 => x"0d",
          1548 => x"02",
          1549 => x"05",
          1550 => x"58",
          1551 => x"52",
          1552 => x"3f",
          1553 => x"08",
          1554 => x"54",
          1555 => x"be",
          1556 => x"75",
          1557 => x"c0",
          1558 => x"87",
          1559 => x"12",
          1560 => x"84",
          1561 => x"40",
          1562 => x"85",
          1563 => x"98",
          1564 => x"7d",
          1565 => x"0c",
          1566 => x"85",
          1567 => x"06",
          1568 => x"71",
          1569 => x"38",
          1570 => x"71",
          1571 => x"05",
          1572 => x"19",
          1573 => x"a2",
          1574 => x"71",
          1575 => x"38",
          1576 => x"83",
          1577 => x"38",
          1578 => x"8a",
          1579 => x"98",
          1580 => x"71",
          1581 => x"c0",
          1582 => x"52",
          1583 => x"87",
          1584 => x"80",
          1585 => x"81",
          1586 => x"c0",
          1587 => x"53",
          1588 => x"82",
          1589 => x"71",
          1590 => x"1a",
          1591 => x"84",
          1592 => x"19",
          1593 => x"06",
          1594 => x"79",
          1595 => x"38",
          1596 => x"80",
          1597 => x"87",
          1598 => x"26",
          1599 => x"73",
          1600 => x"06",
          1601 => x"2e",
          1602 => x"52",
          1603 => x"81",
          1604 => x"8f",
          1605 => x"f3",
          1606 => x"62",
          1607 => x"05",
          1608 => x"57",
          1609 => x"83",
          1610 => x"52",
          1611 => x"3f",
          1612 => x"08",
          1613 => x"54",
          1614 => x"2e",
          1615 => x"81",
          1616 => x"74",
          1617 => x"c0",
          1618 => x"87",
          1619 => x"12",
          1620 => x"84",
          1621 => x"5f",
          1622 => x"0b",
          1623 => x"8c",
          1624 => x"0c",
          1625 => x"80",
          1626 => x"70",
          1627 => x"81",
          1628 => x"54",
          1629 => x"8c",
          1630 => x"81",
          1631 => x"7c",
          1632 => x"58",
          1633 => x"70",
          1634 => x"52",
          1635 => x"8a",
          1636 => x"98",
          1637 => x"71",
          1638 => x"c0",
          1639 => x"52",
          1640 => x"87",
          1641 => x"80",
          1642 => x"81",
          1643 => x"c0",
          1644 => x"53",
          1645 => x"82",
          1646 => x"71",
          1647 => x"19",
          1648 => x"81",
          1649 => x"ff",
          1650 => x"19",
          1651 => x"78",
          1652 => x"38",
          1653 => x"80",
          1654 => x"87",
          1655 => x"26",
          1656 => x"73",
          1657 => x"06",
          1658 => x"2e",
          1659 => x"52",
          1660 => x"81",
          1661 => x"8f",
          1662 => x"f6",
          1663 => x"02",
          1664 => x"05",
          1665 => x"05",
          1666 => x"71",
          1667 => x"57",
          1668 => x"81",
          1669 => x"81",
          1670 => x"54",
          1671 => x"38",
          1672 => x"c0",
          1673 => x"81",
          1674 => x"2e",
          1675 => x"71",
          1676 => x"38",
          1677 => x"87",
          1678 => x"11",
          1679 => x"80",
          1680 => x"80",
          1681 => x"83",
          1682 => x"38",
          1683 => x"72",
          1684 => x"2a",
          1685 => x"51",
          1686 => x"80",
          1687 => x"87",
          1688 => x"08",
          1689 => x"38",
          1690 => x"8c",
          1691 => x"96",
          1692 => x"0c",
          1693 => x"8c",
          1694 => x"08",
          1695 => x"51",
          1696 => x"38",
          1697 => x"56",
          1698 => x"80",
          1699 => x"85",
          1700 => x"77",
          1701 => x"83",
          1702 => x"75",
          1703 => x"cb",
          1704 => x"3d",
          1705 => x"3d",
          1706 => x"11",
          1707 => x"71",
          1708 => x"81",
          1709 => x"53",
          1710 => x"0d",
          1711 => x"0d",
          1712 => x"33",
          1713 => x"71",
          1714 => x"88",
          1715 => x"14",
          1716 => x"07",
          1717 => x"33",
          1718 => x"cb",
          1719 => x"53",
          1720 => x"52",
          1721 => x"04",
          1722 => x"73",
          1723 => x"92",
          1724 => x"52",
          1725 => x"81",
          1726 => x"70",
          1727 => x"70",
          1728 => x"3d",
          1729 => x"3d",
          1730 => x"52",
          1731 => x"70",
          1732 => x"34",
          1733 => x"51",
          1734 => x"81",
          1735 => x"70",
          1736 => x"70",
          1737 => x"05",
          1738 => x"88",
          1739 => x"72",
          1740 => x"0d",
          1741 => x"0d",
          1742 => x"54",
          1743 => x"80",
          1744 => x"71",
          1745 => x"53",
          1746 => x"81",
          1747 => x"ff",
          1748 => x"39",
          1749 => x"04",
          1750 => x"75",
          1751 => x"52",
          1752 => x"70",
          1753 => x"34",
          1754 => x"70",
          1755 => x"3d",
          1756 => x"3d",
          1757 => x"79",
          1758 => x"74",
          1759 => x"56",
          1760 => x"81",
          1761 => x"71",
          1762 => x"16",
          1763 => x"52",
          1764 => x"86",
          1765 => x"2e",
          1766 => x"81",
          1767 => x"86",
          1768 => x"fe",
          1769 => x"76",
          1770 => x"39",
          1771 => x"8a",
          1772 => x"51",
          1773 => x"71",
          1774 => x"33",
          1775 => x"0c",
          1776 => x"04",
          1777 => x"cb",
          1778 => x"80",
          1779 => x"a4",
          1780 => x"3d",
          1781 => x"80",
          1782 => x"33",
          1783 => x"7a",
          1784 => x"38",
          1785 => x"16",
          1786 => x"16",
          1787 => x"17",
          1788 => x"fa",
          1789 => x"cb",
          1790 => x"2e",
          1791 => x"b7",
          1792 => x"a4",
          1793 => x"34",
          1794 => x"70",
          1795 => x"31",
          1796 => x"59",
          1797 => x"77",
          1798 => x"82",
          1799 => x"74",
          1800 => x"81",
          1801 => x"81",
          1802 => x"53",
          1803 => x"16",
          1804 => x"e3",
          1805 => x"81",
          1806 => x"cb",
          1807 => x"3d",
          1808 => x"3d",
          1809 => x"56",
          1810 => x"74",
          1811 => x"2e",
          1812 => x"51",
          1813 => x"81",
          1814 => x"57",
          1815 => x"08",
          1816 => x"54",
          1817 => x"16",
          1818 => x"33",
          1819 => x"3f",
          1820 => x"08",
          1821 => x"38",
          1822 => x"57",
          1823 => x"0c",
          1824 => x"a4",
          1825 => x"0d",
          1826 => x"0d",
          1827 => x"57",
          1828 => x"81",
          1829 => x"58",
          1830 => x"08",
          1831 => x"76",
          1832 => x"83",
          1833 => x"06",
          1834 => x"84",
          1835 => x"78",
          1836 => x"81",
          1837 => x"38",
          1838 => x"81",
          1839 => x"52",
          1840 => x"52",
          1841 => x"3f",
          1842 => x"52",
          1843 => x"51",
          1844 => x"84",
          1845 => x"d2",
          1846 => x"fc",
          1847 => x"8a",
          1848 => x"52",
          1849 => x"51",
          1850 => x"90",
          1851 => x"84",
          1852 => x"fc",
          1853 => x"17",
          1854 => x"a0",
          1855 => x"86",
          1856 => x"08",
          1857 => x"b0",
          1858 => x"55",
          1859 => x"81",
          1860 => x"f8",
          1861 => x"84",
          1862 => x"53",
          1863 => x"17",
          1864 => x"d7",
          1865 => x"a4",
          1866 => x"83",
          1867 => x"77",
          1868 => x"0c",
          1869 => x"04",
          1870 => x"77",
          1871 => x"12",
          1872 => x"55",
          1873 => x"56",
          1874 => x"8d",
          1875 => x"22",
          1876 => x"ac",
          1877 => x"57",
          1878 => x"cb",
          1879 => x"3d",
          1880 => x"3d",
          1881 => x"70",
          1882 => x"57",
          1883 => x"81",
          1884 => x"98",
          1885 => x"81",
          1886 => x"74",
          1887 => x"72",
          1888 => x"f5",
          1889 => x"24",
          1890 => x"81",
          1891 => x"81",
          1892 => x"83",
          1893 => x"38",
          1894 => x"76",
          1895 => x"70",
          1896 => x"16",
          1897 => x"74",
          1898 => x"96",
          1899 => x"a4",
          1900 => x"38",
          1901 => x"06",
          1902 => x"33",
          1903 => x"89",
          1904 => x"08",
          1905 => x"54",
          1906 => x"fc",
          1907 => x"cb",
          1908 => x"fe",
          1909 => x"ff",
          1910 => x"11",
          1911 => x"2b",
          1912 => x"81",
          1913 => x"2a",
          1914 => x"51",
          1915 => x"e2",
          1916 => x"ff",
          1917 => x"da",
          1918 => x"2a",
          1919 => x"05",
          1920 => x"fc",
          1921 => x"cb",
          1922 => x"c6",
          1923 => x"83",
          1924 => x"05",
          1925 => x"f9",
          1926 => x"cb",
          1927 => x"ff",
          1928 => x"ae",
          1929 => x"2a",
          1930 => x"05",
          1931 => x"fc",
          1932 => x"cb",
          1933 => x"38",
          1934 => x"83",
          1935 => x"05",
          1936 => x"f8",
          1937 => x"cb",
          1938 => x"0a",
          1939 => x"39",
          1940 => x"81",
          1941 => x"89",
          1942 => x"f8",
          1943 => x"7c",
          1944 => x"56",
          1945 => x"77",
          1946 => x"38",
          1947 => x"08",
          1948 => x"38",
          1949 => x"72",
          1950 => x"9d",
          1951 => x"24",
          1952 => x"81",
          1953 => x"82",
          1954 => x"83",
          1955 => x"38",
          1956 => x"76",
          1957 => x"70",
          1958 => x"18",
          1959 => x"76",
          1960 => x"9e",
          1961 => x"a4",
          1962 => x"cb",
          1963 => x"d9",
          1964 => x"ff",
          1965 => x"05",
          1966 => x"81",
          1967 => x"54",
          1968 => x"80",
          1969 => x"77",
          1970 => x"f0",
          1971 => x"8f",
          1972 => x"51",
          1973 => x"34",
          1974 => x"17",
          1975 => x"2a",
          1976 => x"05",
          1977 => x"fa",
          1978 => x"cb",
          1979 => x"81",
          1980 => x"81",
          1981 => x"83",
          1982 => x"b4",
          1983 => x"2a",
          1984 => x"8f",
          1985 => x"2a",
          1986 => x"f0",
          1987 => x"06",
          1988 => x"72",
          1989 => x"ec",
          1990 => x"2a",
          1991 => x"05",
          1992 => x"fa",
          1993 => x"cb",
          1994 => x"81",
          1995 => x"80",
          1996 => x"83",
          1997 => x"52",
          1998 => x"fe",
          1999 => x"b4",
          2000 => x"a4",
          2001 => x"76",
          2002 => x"17",
          2003 => x"75",
          2004 => x"3f",
          2005 => x"08",
          2006 => x"a4",
          2007 => x"77",
          2008 => x"77",
          2009 => x"fc",
          2010 => x"b4",
          2011 => x"51",
          2012 => x"c9",
          2013 => x"a4",
          2014 => x"06",
          2015 => x"72",
          2016 => x"3f",
          2017 => x"17",
          2018 => x"cb",
          2019 => x"3d",
          2020 => x"3d",
          2021 => x"7e",
          2022 => x"56",
          2023 => x"75",
          2024 => x"74",
          2025 => x"27",
          2026 => x"80",
          2027 => x"ff",
          2028 => x"75",
          2029 => x"3f",
          2030 => x"08",
          2031 => x"a4",
          2032 => x"38",
          2033 => x"54",
          2034 => x"81",
          2035 => x"39",
          2036 => x"08",
          2037 => x"39",
          2038 => x"51",
          2039 => x"81",
          2040 => x"58",
          2041 => x"08",
          2042 => x"c7",
          2043 => x"a4",
          2044 => x"d2",
          2045 => x"a4",
          2046 => x"cf",
          2047 => x"74",
          2048 => x"fc",
          2049 => x"cb",
          2050 => x"38",
          2051 => x"fe",
          2052 => x"08",
          2053 => x"74",
          2054 => x"38",
          2055 => x"17",
          2056 => x"33",
          2057 => x"73",
          2058 => x"77",
          2059 => x"26",
          2060 => x"80",
          2061 => x"cb",
          2062 => x"3d",
          2063 => x"3d",
          2064 => x"71",
          2065 => x"5b",
          2066 => x"8c",
          2067 => x"77",
          2068 => x"38",
          2069 => x"78",
          2070 => x"81",
          2071 => x"79",
          2072 => x"f9",
          2073 => x"55",
          2074 => x"a4",
          2075 => x"e0",
          2076 => x"a4",
          2077 => x"cb",
          2078 => x"2e",
          2079 => x"98",
          2080 => x"cb",
          2081 => x"82",
          2082 => x"58",
          2083 => x"70",
          2084 => x"80",
          2085 => x"38",
          2086 => x"09",
          2087 => x"e2",
          2088 => x"56",
          2089 => x"76",
          2090 => x"82",
          2091 => x"7a",
          2092 => x"3f",
          2093 => x"cb",
          2094 => x"2e",
          2095 => x"86",
          2096 => x"a4",
          2097 => x"cb",
          2098 => x"70",
          2099 => x"07",
          2100 => x"7c",
          2101 => x"a4",
          2102 => x"51",
          2103 => x"81",
          2104 => x"cb",
          2105 => x"2e",
          2106 => x"17",
          2107 => x"74",
          2108 => x"73",
          2109 => x"27",
          2110 => x"58",
          2111 => x"80",
          2112 => x"56",
          2113 => x"98",
          2114 => x"26",
          2115 => x"56",
          2116 => x"81",
          2117 => x"52",
          2118 => x"c6",
          2119 => x"a4",
          2120 => x"b8",
          2121 => x"81",
          2122 => x"81",
          2123 => x"06",
          2124 => x"cb",
          2125 => x"81",
          2126 => x"09",
          2127 => x"72",
          2128 => x"70",
          2129 => x"51",
          2130 => x"80",
          2131 => x"78",
          2132 => x"06",
          2133 => x"73",
          2134 => x"39",
          2135 => x"52",
          2136 => x"f7",
          2137 => x"a4",
          2138 => x"a4",
          2139 => x"81",
          2140 => x"07",
          2141 => x"55",
          2142 => x"2e",
          2143 => x"80",
          2144 => x"75",
          2145 => x"76",
          2146 => x"3f",
          2147 => x"08",
          2148 => x"38",
          2149 => x"0c",
          2150 => x"fe",
          2151 => x"08",
          2152 => x"74",
          2153 => x"ff",
          2154 => x"0c",
          2155 => x"81",
          2156 => x"84",
          2157 => x"39",
          2158 => x"81",
          2159 => x"8c",
          2160 => x"8c",
          2161 => x"a4",
          2162 => x"39",
          2163 => x"55",
          2164 => x"a4",
          2165 => x"0d",
          2166 => x"0d",
          2167 => x"55",
          2168 => x"81",
          2169 => x"58",
          2170 => x"cb",
          2171 => x"d8",
          2172 => x"74",
          2173 => x"3f",
          2174 => x"08",
          2175 => x"08",
          2176 => x"59",
          2177 => x"77",
          2178 => x"70",
          2179 => x"c8",
          2180 => x"84",
          2181 => x"56",
          2182 => x"58",
          2183 => x"97",
          2184 => x"75",
          2185 => x"52",
          2186 => x"51",
          2187 => x"81",
          2188 => x"80",
          2189 => x"8a",
          2190 => x"32",
          2191 => x"72",
          2192 => x"2a",
          2193 => x"56",
          2194 => x"a4",
          2195 => x"0d",
          2196 => x"0d",
          2197 => x"08",
          2198 => x"74",
          2199 => x"26",
          2200 => x"74",
          2201 => x"72",
          2202 => x"74",
          2203 => x"88",
          2204 => x"73",
          2205 => x"33",
          2206 => x"27",
          2207 => x"16",
          2208 => x"9b",
          2209 => x"2a",
          2210 => x"88",
          2211 => x"58",
          2212 => x"80",
          2213 => x"16",
          2214 => x"0c",
          2215 => x"8a",
          2216 => x"89",
          2217 => x"72",
          2218 => x"38",
          2219 => x"51",
          2220 => x"81",
          2221 => x"54",
          2222 => x"08",
          2223 => x"38",
          2224 => x"cb",
          2225 => x"8b",
          2226 => x"08",
          2227 => x"08",
          2228 => x"82",
          2229 => x"74",
          2230 => x"cb",
          2231 => x"75",
          2232 => x"3f",
          2233 => x"08",
          2234 => x"73",
          2235 => x"98",
          2236 => x"82",
          2237 => x"2e",
          2238 => x"39",
          2239 => x"39",
          2240 => x"13",
          2241 => x"74",
          2242 => x"16",
          2243 => x"18",
          2244 => x"77",
          2245 => x"0c",
          2246 => x"04",
          2247 => x"7a",
          2248 => x"12",
          2249 => x"59",
          2250 => x"80",
          2251 => x"86",
          2252 => x"98",
          2253 => x"14",
          2254 => x"55",
          2255 => x"81",
          2256 => x"83",
          2257 => x"77",
          2258 => x"81",
          2259 => x"0c",
          2260 => x"55",
          2261 => x"76",
          2262 => x"17",
          2263 => x"74",
          2264 => x"9b",
          2265 => x"39",
          2266 => x"ff",
          2267 => x"2a",
          2268 => x"81",
          2269 => x"52",
          2270 => x"e6",
          2271 => x"a4",
          2272 => x"55",
          2273 => x"cb",
          2274 => x"80",
          2275 => x"55",
          2276 => x"08",
          2277 => x"f4",
          2278 => x"08",
          2279 => x"08",
          2280 => x"38",
          2281 => x"77",
          2282 => x"84",
          2283 => x"39",
          2284 => x"52",
          2285 => x"86",
          2286 => x"a4",
          2287 => x"55",
          2288 => x"08",
          2289 => x"c4",
          2290 => x"81",
          2291 => x"81",
          2292 => x"81",
          2293 => x"a4",
          2294 => x"b0",
          2295 => x"a4",
          2296 => x"51",
          2297 => x"81",
          2298 => x"a0",
          2299 => x"15",
          2300 => x"75",
          2301 => x"3f",
          2302 => x"08",
          2303 => x"76",
          2304 => x"77",
          2305 => x"9c",
          2306 => x"55",
          2307 => x"a4",
          2308 => x"0d",
          2309 => x"0d",
          2310 => x"08",
          2311 => x"80",
          2312 => x"fc",
          2313 => x"cb",
          2314 => x"81",
          2315 => x"80",
          2316 => x"cb",
          2317 => x"98",
          2318 => x"78",
          2319 => x"3f",
          2320 => x"08",
          2321 => x"a4",
          2322 => x"38",
          2323 => x"08",
          2324 => x"70",
          2325 => x"58",
          2326 => x"2e",
          2327 => x"83",
          2328 => x"81",
          2329 => x"55",
          2330 => x"81",
          2331 => x"07",
          2332 => x"2e",
          2333 => x"16",
          2334 => x"2e",
          2335 => x"88",
          2336 => x"81",
          2337 => x"56",
          2338 => x"51",
          2339 => x"81",
          2340 => x"54",
          2341 => x"08",
          2342 => x"9b",
          2343 => x"2e",
          2344 => x"83",
          2345 => x"73",
          2346 => x"0c",
          2347 => x"04",
          2348 => x"76",
          2349 => x"54",
          2350 => x"81",
          2351 => x"83",
          2352 => x"76",
          2353 => x"53",
          2354 => x"2e",
          2355 => x"90",
          2356 => x"51",
          2357 => x"81",
          2358 => x"90",
          2359 => x"53",
          2360 => x"a4",
          2361 => x"0d",
          2362 => x"0d",
          2363 => x"83",
          2364 => x"54",
          2365 => x"55",
          2366 => x"3f",
          2367 => x"51",
          2368 => x"2e",
          2369 => x"8b",
          2370 => x"2a",
          2371 => x"51",
          2372 => x"86",
          2373 => x"f7",
          2374 => x"7d",
          2375 => x"75",
          2376 => x"98",
          2377 => x"2e",
          2378 => x"98",
          2379 => x"78",
          2380 => x"3f",
          2381 => x"08",
          2382 => x"a4",
          2383 => x"38",
          2384 => x"70",
          2385 => x"73",
          2386 => x"58",
          2387 => x"8b",
          2388 => x"bf",
          2389 => x"ff",
          2390 => x"53",
          2391 => x"34",
          2392 => x"08",
          2393 => x"e5",
          2394 => x"81",
          2395 => x"2e",
          2396 => x"70",
          2397 => x"57",
          2398 => x"9e",
          2399 => x"2e",
          2400 => x"cb",
          2401 => x"df",
          2402 => x"72",
          2403 => x"81",
          2404 => x"76",
          2405 => x"2e",
          2406 => x"52",
          2407 => x"fc",
          2408 => x"a4",
          2409 => x"cb",
          2410 => x"38",
          2411 => x"fe",
          2412 => x"39",
          2413 => x"16",
          2414 => x"cb",
          2415 => x"3d",
          2416 => x"3d",
          2417 => x"08",
          2418 => x"52",
          2419 => x"c5",
          2420 => x"a4",
          2421 => x"cb",
          2422 => x"38",
          2423 => x"52",
          2424 => x"de",
          2425 => x"a4",
          2426 => x"cb",
          2427 => x"38",
          2428 => x"cb",
          2429 => x"9c",
          2430 => x"ea",
          2431 => x"53",
          2432 => x"9c",
          2433 => x"ea",
          2434 => x"0b",
          2435 => x"74",
          2436 => x"0c",
          2437 => x"04",
          2438 => x"75",
          2439 => x"12",
          2440 => x"53",
          2441 => x"9a",
          2442 => x"a4",
          2443 => x"9c",
          2444 => x"e5",
          2445 => x"0b",
          2446 => x"85",
          2447 => x"fa",
          2448 => x"7a",
          2449 => x"0b",
          2450 => x"98",
          2451 => x"2e",
          2452 => x"80",
          2453 => x"55",
          2454 => x"17",
          2455 => x"33",
          2456 => x"51",
          2457 => x"2e",
          2458 => x"85",
          2459 => x"06",
          2460 => x"e5",
          2461 => x"2e",
          2462 => x"8b",
          2463 => x"70",
          2464 => x"34",
          2465 => x"71",
          2466 => x"05",
          2467 => x"15",
          2468 => x"27",
          2469 => x"15",
          2470 => x"80",
          2471 => x"34",
          2472 => x"52",
          2473 => x"88",
          2474 => x"17",
          2475 => x"52",
          2476 => x"3f",
          2477 => x"08",
          2478 => x"12",
          2479 => x"3f",
          2480 => x"08",
          2481 => x"98",
          2482 => x"da",
          2483 => x"a4",
          2484 => x"23",
          2485 => x"04",
          2486 => x"7f",
          2487 => x"5b",
          2488 => x"33",
          2489 => x"73",
          2490 => x"38",
          2491 => x"80",
          2492 => x"38",
          2493 => x"8c",
          2494 => x"08",
          2495 => x"aa",
          2496 => x"41",
          2497 => x"33",
          2498 => x"73",
          2499 => x"81",
          2500 => x"81",
          2501 => x"dc",
          2502 => x"70",
          2503 => x"07",
          2504 => x"73",
          2505 => x"88",
          2506 => x"70",
          2507 => x"73",
          2508 => x"38",
          2509 => x"ab",
          2510 => x"52",
          2511 => x"91",
          2512 => x"a4",
          2513 => x"98",
          2514 => x"61",
          2515 => x"5a",
          2516 => x"a0",
          2517 => x"e7",
          2518 => x"70",
          2519 => x"79",
          2520 => x"73",
          2521 => x"81",
          2522 => x"38",
          2523 => x"33",
          2524 => x"ae",
          2525 => x"70",
          2526 => x"82",
          2527 => x"51",
          2528 => x"54",
          2529 => x"79",
          2530 => x"74",
          2531 => x"57",
          2532 => x"af",
          2533 => x"70",
          2534 => x"51",
          2535 => x"dc",
          2536 => x"73",
          2537 => x"38",
          2538 => x"82",
          2539 => x"19",
          2540 => x"54",
          2541 => x"82",
          2542 => x"54",
          2543 => x"78",
          2544 => x"81",
          2545 => x"54",
          2546 => x"81",
          2547 => x"af",
          2548 => x"77",
          2549 => x"70",
          2550 => x"25",
          2551 => x"07",
          2552 => x"51",
          2553 => x"2e",
          2554 => x"39",
          2555 => x"80",
          2556 => x"33",
          2557 => x"73",
          2558 => x"81",
          2559 => x"81",
          2560 => x"dc",
          2561 => x"70",
          2562 => x"07",
          2563 => x"73",
          2564 => x"b5",
          2565 => x"2e",
          2566 => x"83",
          2567 => x"76",
          2568 => x"07",
          2569 => x"2e",
          2570 => x"8b",
          2571 => x"77",
          2572 => x"30",
          2573 => x"71",
          2574 => x"53",
          2575 => x"55",
          2576 => x"38",
          2577 => x"5c",
          2578 => x"75",
          2579 => x"73",
          2580 => x"38",
          2581 => x"06",
          2582 => x"11",
          2583 => x"75",
          2584 => x"3f",
          2585 => x"08",
          2586 => x"38",
          2587 => x"33",
          2588 => x"54",
          2589 => x"e6",
          2590 => x"cb",
          2591 => x"2e",
          2592 => x"ff",
          2593 => x"74",
          2594 => x"38",
          2595 => x"75",
          2596 => x"17",
          2597 => x"57",
          2598 => x"a7",
          2599 => x"81",
          2600 => x"e5",
          2601 => x"cb",
          2602 => x"38",
          2603 => x"54",
          2604 => x"89",
          2605 => x"70",
          2606 => x"57",
          2607 => x"54",
          2608 => x"81",
          2609 => x"f7",
          2610 => x"7e",
          2611 => x"2e",
          2612 => x"33",
          2613 => x"e5",
          2614 => x"06",
          2615 => x"7a",
          2616 => x"a0",
          2617 => x"38",
          2618 => x"55",
          2619 => x"84",
          2620 => x"39",
          2621 => x"8b",
          2622 => x"7b",
          2623 => x"7a",
          2624 => x"3f",
          2625 => x"08",
          2626 => x"a4",
          2627 => x"38",
          2628 => x"52",
          2629 => x"aa",
          2630 => x"a4",
          2631 => x"cb",
          2632 => x"c2",
          2633 => x"08",
          2634 => x"55",
          2635 => x"ff",
          2636 => x"15",
          2637 => x"54",
          2638 => x"34",
          2639 => x"70",
          2640 => x"81",
          2641 => x"58",
          2642 => x"8b",
          2643 => x"74",
          2644 => x"3f",
          2645 => x"08",
          2646 => x"38",
          2647 => x"51",
          2648 => x"ff",
          2649 => x"ab",
          2650 => x"55",
          2651 => x"bb",
          2652 => x"2e",
          2653 => x"80",
          2654 => x"85",
          2655 => x"06",
          2656 => x"58",
          2657 => x"80",
          2658 => x"75",
          2659 => x"73",
          2660 => x"b5",
          2661 => x"0b",
          2662 => x"80",
          2663 => x"39",
          2664 => x"54",
          2665 => x"85",
          2666 => x"75",
          2667 => x"81",
          2668 => x"73",
          2669 => x"1b",
          2670 => x"2a",
          2671 => x"51",
          2672 => x"80",
          2673 => x"90",
          2674 => x"ff",
          2675 => x"05",
          2676 => x"f5",
          2677 => x"cb",
          2678 => x"1c",
          2679 => x"39",
          2680 => x"a4",
          2681 => x"0d",
          2682 => x"0d",
          2683 => x"7b",
          2684 => x"73",
          2685 => x"55",
          2686 => x"2e",
          2687 => x"75",
          2688 => x"57",
          2689 => x"26",
          2690 => x"ba",
          2691 => x"70",
          2692 => x"ba",
          2693 => x"06",
          2694 => x"73",
          2695 => x"70",
          2696 => x"51",
          2697 => x"89",
          2698 => x"82",
          2699 => x"ff",
          2700 => x"56",
          2701 => x"2e",
          2702 => x"80",
          2703 => x"f0",
          2704 => x"08",
          2705 => x"76",
          2706 => x"58",
          2707 => x"81",
          2708 => x"ff",
          2709 => x"53",
          2710 => x"26",
          2711 => x"13",
          2712 => x"06",
          2713 => x"9f",
          2714 => x"99",
          2715 => x"e0",
          2716 => x"ff",
          2717 => x"72",
          2718 => x"2a",
          2719 => x"72",
          2720 => x"06",
          2721 => x"ff",
          2722 => x"30",
          2723 => x"70",
          2724 => x"07",
          2725 => x"9f",
          2726 => x"54",
          2727 => x"80",
          2728 => x"81",
          2729 => x"59",
          2730 => x"25",
          2731 => x"8b",
          2732 => x"24",
          2733 => x"76",
          2734 => x"78",
          2735 => x"81",
          2736 => x"51",
          2737 => x"a4",
          2738 => x"0d",
          2739 => x"0d",
          2740 => x"0b",
          2741 => x"ff",
          2742 => x"0c",
          2743 => x"51",
          2744 => x"84",
          2745 => x"a4",
          2746 => x"38",
          2747 => x"51",
          2748 => x"81",
          2749 => x"83",
          2750 => x"54",
          2751 => x"82",
          2752 => x"09",
          2753 => x"e3",
          2754 => x"b4",
          2755 => x"57",
          2756 => x"2e",
          2757 => x"83",
          2758 => x"74",
          2759 => x"70",
          2760 => x"25",
          2761 => x"51",
          2762 => x"38",
          2763 => x"2e",
          2764 => x"b5",
          2765 => x"81",
          2766 => x"80",
          2767 => x"e0",
          2768 => x"cb",
          2769 => x"81",
          2770 => x"80",
          2771 => x"85",
          2772 => x"b4",
          2773 => x"16",
          2774 => x"3f",
          2775 => x"08",
          2776 => x"a4",
          2777 => x"83",
          2778 => x"74",
          2779 => x"0c",
          2780 => x"04",
          2781 => x"61",
          2782 => x"80",
          2783 => x"58",
          2784 => x"0c",
          2785 => x"e1",
          2786 => x"a4",
          2787 => x"56",
          2788 => x"cb",
          2789 => x"86",
          2790 => x"cb",
          2791 => x"29",
          2792 => x"05",
          2793 => x"53",
          2794 => x"80",
          2795 => x"38",
          2796 => x"76",
          2797 => x"74",
          2798 => x"72",
          2799 => x"38",
          2800 => x"51",
          2801 => x"81",
          2802 => x"81",
          2803 => x"81",
          2804 => x"72",
          2805 => x"80",
          2806 => x"38",
          2807 => x"70",
          2808 => x"53",
          2809 => x"86",
          2810 => x"a7",
          2811 => x"34",
          2812 => x"34",
          2813 => x"14",
          2814 => x"b2",
          2815 => x"a4",
          2816 => x"06",
          2817 => x"54",
          2818 => x"72",
          2819 => x"76",
          2820 => x"38",
          2821 => x"70",
          2822 => x"53",
          2823 => x"85",
          2824 => x"70",
          2825 => x"5b",
          2826 => x"81",
          2827 => x"81",
          2828 => x"76",
          2829 => x"81",
          2830 => x"38",
          2831 => x"56",
          2832 => x"83",
          2833 => x"70",
          2834 => x"80",
          2835 => x"83",
          2836 => x"dc",
          2837 => x"cb",
          2838 => x"76",
          2839 => x"05",
          2840 => x"16",
          2841 => x"56",
          2842 => x"d7",
          2843 => x"8d",
          2844 => x"72",
          2845 => x"54",
          2846 => x"57",
          2847 => x"95",
          2848 => x"73",
          2849 => x"3f",
          2850 => x"08",
          2851 => x"57",
          2852 => x"89",
          2853 => x"56",
          2854 => x"d7",
          2855 => x"76",
          2856 => x"f1",
          2857 => x"76",
          2858 => x"e9",
          2859 => x"51",
          2860 => x"81",
          2861 => x"83",
          2862 => x"53",
          2863 => x"2e",
          2864 => x"84",
          2865 => x"ca",
          2866 => x"da",
          2867 => x"a4",
          2868 => x"ff",
          2869 => x"8d",
          2870 => x"14",
          2871 => x"3f",
          2872 => x"08",
          2873 => x"15",
          2874 => x"14",
          2875 => x"34",
          2876 => x"33",
          2877 => x"81",
          2878 => x"54",
          2879 => x"72",
          2880 => x"91",
          2881 => x"ff",
          2882 => x"29",
          2883 => x"33",
          2884 => x"72",
          2885 => x"72",
          2886 => x"38",
          2887 => x"06",
          2888 => x"2e",
          2889 => x"56",
          2890 => x"80",
          2891 => x"da",
          2892 => x"cb",
          2893 => x"81",
          2894 => x"88",
          2895 => x"8f",
          2896 => x"56",
          2897 => x"38",
          2898 => x"51",
          2899 => x"81",
          2900 => x"83",
          2901 => x"55",
          2902 => x"80",
          2903 => x"da",
          2904 => x"cb",
          2905 => x"80",
          2906 => x"da",
          2907 => x"cb",
          2908 => x"ff",
          2909 => x"8d",
          2910 => x"2e",
          2911 => x"88",
          2912 => x"14",
          2913 => x"05",
          2914 => x"75",
          2915 => x"38",
          2916 => x"52",
          2917 => x"51",
          2918 => x"3f",
          2919 => x"08",
          2920 => x"a4",
          2921 => x"82",
          2922 => x"cb",
          2923 => x"ff",
          2924 => x"26",
          2925 => x"57",
          2926 => x"f5",
          2927 => x"82",
          2928 => x"f5",
          2929 => x"81",
          2930 => x"8d",
          2931 => x"2e",
          2932 => x"82",
          2933 => x"16",
          2934 => x"16",
          2935 => x"70",
          2936 => x"7a",
          2937 => x"0c",
          2938 => x"83",
          2939 => x"06",
          2940 => x"de",
          2941 => x"ae",
          2942 => x"a4",
          2943 => x"ff",
          2944 => x"56",
          2945 => x"38",
          2946 => x"38",
          2947 => x"51",
          2948 => x"81",
          2949 => x"a8",
          2950 => x"82",
          2951 => x"39",
          2952 => x"80",
          2953 => x"38",
          2954 => x"15",
          2955 => x"53",
          2956 => x"8d",
          2957 => x"15",
          2958 => x"76",
          2959 => x"51",
          2960 => x"13",
          2961 => x"8d",
          2962 => x"15",
          2963 => x"c5",
          2964 => x"90",
          2965 => x"0b",
          2966 => x"ff",
          2967 => x"15",
          2968 => x"2e",
          2969 => x"81",
          2970 => x"e4",
          2971 => x"b6",
          2972 => x"a4",
          2973 => x"ff",
          2974 => x"81",
          2975 => x"06",
          2976 => x"81",
          2977 => x"51",
          2978 => x"81",
          2979 => x"80",
          2980 => x"cb",
          2981 => x"15",
          2982 => x"14",
          2983 => x"3f",
          2984 => x"08",
          2985 => x"06",
          2986 => x"d4",
          2987 => x"81",
          2988 => x"38",
          2989 => x"d8",
          2990 => x"cb",
          2991 => x"8b",
          2992 => x"2e",
          2993 => x"b3",
          2994 => x"14",
          2995 => x"3f",
          2996 => x"08",
          2997 => x"e4",
          2998 => x"81",
          2999 => x"84",
          3000 => x"d7",
          3001 => x"cb",
          3002 => x"15",
          3003 => x"14",
          3004 => x"3f",
          3005 => x"08",
          3006 => x"76",
          3007 => x"cb",
          3008 => x"05",
          3009 => x"cb",
          3010 => x"86",
          3011 => x"0b",
          3012 => x"80",
          3013 => x"cb",
          3014 => x"3d",
          3015 => x"3d",
          3016 => x"89",
          3017 => x"2e",
          3018 => x"08",
          3019 => x"2e",
          3020 => x"33",
          3021 => x"2e",
          3022 => x"13",
          3023 => x"22",
          3024 => x"76",
          3025 => x"06",
          3026 => x"13",
          3027 => x"c0",
          3028 => x"a4",
          3029 => x"52",
          3030 => x"71",
          3031 => x"55",
          3032 => x"53",
          3033 => x"0c",
          3034 => x"cb",
          3035 => x"3d",
          3036 => x"3d",
          3037 => x"05",
          3038 => x"89",
          3039 => x"52",
          3040 => x"3f",
          3041 => x"0b",
          3042 => x"08",
          3043 => x"81",
          3044 => x"84",
          3045 => x"c0",
          3046 => x"55",
          3047 => x"2e",
          3048 => x"74",
          3049 => x"73",
          3050 => x"38",
          3051 => x"78",
          3052 => x"54",
          3053 => x"92",
          3054 => x"89",
          3055 => x"84",
          3056 => x"b0",
          3057 => x"a4",
          3058 => x"81",
          3059 => x"88",
          3060 => x"eb",
          3061 => x"02",
          3062 => x"e7",
          3063 => x"59",
          3064 => x"80",
          3065 => x"38",
          3066 => x"70",
          3067 => x"d0",
          3068 => x"3d",
          3069 => x"58",
          3070 => x"81",
          3071 => x"55",
          3072 => x"08",
          3073 => x"7a",
          3074 => x"8c",
          3075 => x"56",
          3076 => x"81",
          3077 => x"55",
          3078 => x"08",
          3079 => x"80",
          3080 => x"70",
          3081 => x"57",
          3082 => x"83",
          3083 => x"77",
          3084 => x"73",
          3085 => x"ab",
          3086 => x"2e",
          3087 => x"84",
          3088 => x"06",
          3089 => x"51",
          3090 => x"81",
          3091 => x"55",
          3092 => x"b2",
          3093 => x"06",
          3094 => x"b8",
          3095 => x"2a",
          3096 => x"51",
          3097 => x"2e",
          3098 => x"55",
          3099 => x"77",
          3100 => x"74",
          3101 => x"77",
          3102 => x"81",
          3103 => x"73",
          3104 => x"af",
          3105 => x"7a",
          3106 => x"3f",
          3107 => x"08",
          3108 => x"b2",
          3109 => x"8e",
          3110 => x"ea",
          3111 => x"a0",
          3112 => x"34",
          3113 => x"52",
          3114 => x"bd",
          3115 => x"62",
          3116 => x"d4",
          3117 => x"54",
          3118 => x"15",
          3119 => x"2e",
          3120 => x"7a",
          3121 => x"51",
          3122 => x"75",
          3123 => x"d4",
          3124 => x"be",
          3125 => x"a4",
          3126 => x"cb",
          3127 => x"ca",
          3128 => x"74",
          3129 => x"02",
          3130 => x"70",
          3131 => x"81",
          3132 => x"56",
          3133 => x"86",
          3134 => x"82",
          3135 => x"81",
          3136 => x"06",
          3137 => x"80",
          3138 => x"75",
          3139 => x"73",
          3140 => x"38",
          3141 => x"92",
          3142 => x"7a",
          3143 => x"3f",
          3144 => x"08",
          3145 => x"8c",
          3146 => x"55",
          3147 => x"08",
          3148 => x"77",
          3149 => x"81",
          3150 => x"73",
          3151 => x"38",
          3152 => x"07",
          3153 => x"11",
          3154 => x"0c",
          3155 => x"0c",
          3156 => x"52",
          3157 => x"3f",
          3158 => x"08",
          3159 => x"08",
          3160 => x"63",
          3161 => x"5a",
          3162 => x"81",
          3163 => x"81",
          3164 => x"8c",
          3165 => x"7a",
          3166 => x"17",
          3167 => x"23",
          3168 => x"34",
          3169 => x"1a",
          3170 => x"9c",
          3171 => x"0b",
          3172 => x"77",
          3173 => x"81",
          3174 => x"73",
          3175 => x"8d",
          3176 => x"a4",
          3177 => x"81",
          3178 => x"cb",
          3179 => x"1a",
          3180 => x"22",
          3181 => x"7b",
          3182 => x"a8",
          3183 => x"78",
          3184 => x"3f",
          3185 => x"08",
          3186 => x"a4",
          3187 => x"83",
          3188 => x"81",
          3189 => x"ff",
          3190 => x"06",
          3191 => x"55",
          3192 => x"56",
          3193 => x"76",
          3194 => x"51",
          3195 => x"27",
          3196 => x"70",
          3197 => x"5a",
          3198 => x"76",
          3199 => x"74",
          3200 => x"83",
          3201 => x"73",
          3202 => x"38",
          3203 => x"51",
          3204 => x"81",
          3205 => x"85",
          3206 => x"8e",
          3207 => x"2a",
          3208 => x"08",
          3209 => x"0c",
          3210 => x"79",
          3211 => x"73",
          3212 => x"0c",
          3213 => x"04",
          3214 => x"60",
          3215 => x"40",
          3216 => x"80",
          3217 => x"3d",
          3218 => x"78",
          3219 => x"3f",
          3220 => x"08",
          3221 => x"a4",
          3222 => x"91",
          3223 => x"74",
          3224 => x"38",
          3225 => x"c4",
          3226 => x"33",
          3227 => x"87",
          3228 => x"2e",
          3229 => x"95",
          3230 => x"91",
          3231 => x"56",
          3232 => x"81",
          3233 => x"34",
          3234 => x"a0",
          3235 => x"08",
          3236 => x"31",
          3237 => x"27",
          3238 => x"5c",
          3239 => x"82",
          3240 => x"19",
          3241 => x"ff",
          3242 => x"74",
          3243 => x"7e",
          3244 => x"ff",
          3245 => x"2a",
          3246 => x"79",
          3247 => x"87",
          3248 => x"08",
          3249 => x"98",
          3250 => x"78",
          3251 => x"3f",
          3252 => x"08",
          3253 => x"27",
          3254 => x"74",
          3255 => x"a3",
          3256 => x"1a",
          3257 => x"08",
          3258 => x"d4",
          3259 => x"cb",
          3260 => x"2e",
          3261 => x"81",
          3262 => x"1a",
          3263 => x"59",
          3264 => x"2e",
          3265 => x"77",
          3266 => x"11",
          3267 => x"55",
          3268 => x"85",
          3269 => x"31",
          3270 => x"76",
          3271 => x"81",
          3272 => x"ca",
          3273 => x"cb",
          3274 => x"d7",
          3275 => x"11",
          3276 => x"74",
          3277 => x"38",
          3278 => x"77",
          3279 => x"78",
          3280 => x"84",
          3281 => x"16",
          3282 => x"08",
          3283 => x"2b",
          3284 => x"cf",
          3285 => x"89",
          3286 => x"39",
          3287 => x"0c",
          3288 => x"83",
          3289 => x"80",
          3290 => x"55",
          3291 => x"83",
          3292 => x"9c",
          3293 => x"7e",
          3294 => x"3f",
          3295 => x"08",
          3296 => x"75",
          3297 => x"08",
          3298 => x"1f",
          3299 => x"7c",
          3300 => x"3f",
          3301 => x"7e",
          3302 => x"0c",
          3303 => x"1b",
          3304 => x"1c",
          3305 => x"fd",
          3306 => x"56",
          3307 => x"a4",
          3308 => x"0d",
          3309 => x"0d",
          3310 => x"64",
          3311 => x"58",
          3312 => x"90",
          3313 => x"52",
          3314 => x"d2",
          3315 => x"a4",
          3316 => x"cb",
          3317 => x"38",
          3318 => x"55",
          3319 => x"86",
          3320 => x"83",
          3321 => x"18",
          3322 => x"2a",
          3323 => x"51",
          3324 => x"56",
          3325 => x"83",
          3326 => x"39",
          3327 => x"19",
          3328 => x"83",
          3329 => x"0b",
          3330 => x"81",
          3331 => x"39",
          3332 => x"7c",
          3333 => x"74",
          3334 => x"38",
          3335 => x"7b",
          3336 => x"ec",
          3337 => x"08",
          3338 => x"06",
          3339 => x"81",
          3340 => x"8a",
          3341 => x"05",
          3342 => x"06",
          3343 => x"bf",
          3344 => x"38",
          3345 => x"55",
          3346 => x"7a",
          3347 => x"98",
          3348 => x"77",
          3349 => x"3f",
          3350 => x"08",
          3351 => x"a4",
          3352 => x"82",
          3353 => x"81",
          3354 => x"38",
          3355 => x"ff",
          3356 => x"98",
          3357 => x"18",
          3358 => x"74",
          3359 => x"7e",
          3360 => x"08",
          3361 => x"2e",
          3362 => x"8d",
          3363 => x"ce",
          3364 => x"cb",
          3365 => x"ee",
          3366 => x"08",
          3367 => x"d1",
          3368 => x"cb",
          3369 => x"2e",
          3370 => x"81",
          3371 => x"1b",
          3372 => x"5a",
          3373 => x"2e",
          3374 => x"78",
          3375 => x"11",
          3376 => x"55",
          3377 => x"85",
          3378 => x"31",
          3379 => x"76",
          3380 => x"81",
          3381 => x"c8",
          3382 => x"cb",
          3383 => x"a6",
          3384 => x"11",
          3385 => x"56",
          3386 => x"27",
          3387 => x"80",
          3388 => x"08",
          3389 => x"2b",
          3390 => x"b4",
          3391 => x"b5",
          3392 => x"80",
          3393 => x"34",
          3394 => x"56",
          3395 => x"8c",
          3396 => x"19",
          3397 => x"38",
          3398 => x"b6",
          3399 => x"a4",
          3400 => x"38",
          3401 => x"12",
          3402 => x"9c",
          3403 => x"18",
          3404 => x"06",
          3405 => x"31",
          3406 => x"76",
          3407 => x"7b",
          3408 => x"08",
          3409 => x"cd",
          3410 => x"cb",
          3411 => x"b6",
          3412 => x"7c",
          3413 => x"08",
          3414 => x"1f",
          3415 => x"cb",
          3416 => x"55",
          3417 => x"16",
          3418 => x"31",
          3419 => x"7f",
          3420 => x"94",
          3421 => x"70",
          3422 => x"8c",
          3423 => x"58",
          3424 => x"76",
          3425 => x"75",
          3426 => x"19",
          3427 => x"39",
          3428 => x"80",
          3429 => x"74",
          3430 => x"80",
          3431 => x"cb",
          3432 => x"3d",
          3433 => x"3d",
          3434 => x"3d",
          3435 => x"70",
          3436 => x"ea",
          3437 => x"a4",
          3438 => x"cb",
          3439 => x"fb",
          3440 => x"33",
          3441 => x"70",
          3442 => x"55",
          3443 => x"2e",
          3444 => x"a0",
          3445 => x"78",
          3446 => x"3f",
          3447 => x"08",
          3448 => x"a4",
          3449 => x"38",
          3450 => x"8b",
          3451 => x"07",
          3452 => x"8b",
          3453 => x"16",
          3454 => x"52",
          3455 => x"dd",
          3456 => x"16",
          3457 => x"15",
          3458 => x"3f",
          3459 => x"0a",
          3460 => x"51",
          3461 => x"76",
          3462 => x"51",
          3463 => x"78",
          3464 => x"83",
          3465 => x"51",
          3466 => x"81",
          3467 => x"90",
          3468 => x"bf",
          3469 => x"73",
          3470 => x"76",
          3471 => x"0c",
          3472 => x"04",
          3473 => x"76",
          3474 => x"fe",
          3475 => x"cb",
          3476 => x"81",
          3477 => x"9c",
          3478 => x"fc",
          3479 => x"51",
          3480 => x"81",
          3481 => x"53",
          3482 => x"08",
          3483 => x"cb",
          3484 => x"0c",
          3485 => x"a4",
          3486 => x"0d",
          3487 => x"0d",
          3488 => x"e6",
          3489 => x"52",
          3490 => x"cb",
          3491 => x"8b",
          3492 => x"a4",
          3493 => x"d4",
          3494 => x"71",
          3495 => x"0c",
          3496 => x"04",
          3497 => x"80",
          3498 => x"d0",
          3499 => x"3d",
          3500 => x"3f",
          3501 => x"08",
          3502 => x"a4",
          3503 => x"38",
          3504 => x"52",
          3505 => x"05",
          3506 => x"3f",
          3507 => x"08",
          3508 => x"a4",
          3509 => x"02",
          3510 => x"33",
          3511 => x"55",
          3512 => x"25",
          3513 => x"7a",
          3514 => x"54",
          3515 => x"a2",
          3516 => x"84",
          3517 => x"06",
          3518 => x"73",
          3519 => x"38",
          3520 => x"70",
          3521 => x"a8",
          3522 => x"a4",
          3523 => x"0c",
          3524 => x"cb",
          3525 => x"2e",
          3526 => x"83",
          3527 => x"74",
          3528 => x"0c",
          3529 => x"04",
          3530 => x"6f",
          3531 => x"80",
          3532 => x"53",
          3533 => x"b8",
          3534 => x"3d",
          3535 => x"3f",
          3536 => x"08",
          3537 => x"a4",
          3538 => x"38",
          3539 => x"7c",
          3540 => x"47",
          3541 => x"54",
          3542 => x"81",
          3543 => x"52",
          3544 => x"52",
          3545 => x"3f",
          3546 => x"08",
          3547 => x"a4",
          3548 => x"38",
          3549 => x"51",
          3550 => x"81",
          3551 => x"57",
          3552 => x"08",
          3553 => x"69",
          3554 => x"da",
          3555 => x"cb",
          3556 => x"76",
          3557 => x"d5",
          3558 => x"cb",
          3559 => x"81",
          3560 => x"82",
          3561 => x"52",
          3562 => x"eb",
          3563 => x"a4",
          3564 => x"cb",
          3565 => x"38",
          3566 => x"51",
          3567 => x"73",
          3568 => x"08",
          3569 => x"76",
          3570 => x"d6",
          3571 => x"cb",
          3572 => x"81",
          3573 => x"80",
          3574 => x"76",
          3575 => x"81",
          3576 => x"82",
          3577 => x"39",
          3578 => x"38",
          3579 => x"bc",
          3580 => x"51",
          3581 => x"76",
          3582 => x"11",
          3583 => x"51",
          3584 => x"73",
          3585 => x"38",
          3586 => x"55",
          3587 => x"16",
          3588 => x"56",
          3589 => x"38",
          3590 => x"73",
          3591 => x"90",
          3592 => x"2e",
          3593 => x"16",
          3594 => x"ff",
          3595 => x"ff",
          3596 => x"58",
          3597 => x"74",
          3598 => x"75",
          3599 => x"18",
          3600 => x"58",
          3601 => x"fe",
          3602 => x"7b",
          3603 => x"06",
          3604 => x"18",
          3605 => x"58",
          3606 => x"80",
          3607 => x"d4",
          3608 => x"29",
          3609 => x"05",
          3610 => x"33",
          3611 => x"56",
          3612 => x"2e",
          3613 => x"16",
          3614 => x"33",
          3615 => x"73",
          3616 => x"16",
          3617 => x"26",
          3618 => x"55",
          3619 => x"91",
          3620 => x"54",
          3621 => x"70",
          3622 => x"34",
          3623 => x"ec",
          3624 => x"70",
          3625 => x"34",
          3626 => x"09",
          3627 => x"38",
          3628 => x"39",
          3629 => x"19",
          3630 => x"33",
          3631 => x"05",
          3632 => x"78",
          3633 => x"80",
          3634 => x"81",
          3635 => x"9e",
          3636 => x"f7",
          3637 => x"7d",
          3638 => x"05",
          3639 => x"57",
          3640 => x"3f",
          3641 => x"08",
          3642 => x"a4",
          3643 => x"38",
          3644 => x"53",
          3645 => x"38",
          3646 => x"54",
          3647 => x"92",
          3648 => x"33",
          3649 => x"70",
          3650 => x"54",
          3651 => x"38",
          3652 => x"15",
          3653 => x"70",
          3654 => x"58",
          3655 => x"82",
          3656 => x"8a",
          3657 => x"89",
          3658 => x"53",
          3659 => x"b7",
          3660 => x"ff",
          3661 => x"9b",
          3662 => x"cb",
          3663 => x"15",
          3664 => x"53",
          3665 => x"9b",
          3666 => x"cb",
          3667 => x"26",
          3668 => x"30",
          3669 => x"70",
          3670 => x"77",
          3671 => x"18",
          3672 => x"51",
          3673 => x"88",
          3674 => x"73",
          3675 => x"52",
          3676 => x"ca",
          3677 => x"a4",
          3678 => x"cb",
          3679 => x"2e",
          3680 => x"81",
          3681 => x"ff",
          3682 => x"38",
          3683 => x"08",
          3684 => x"73",
          3685 => x"73",
          3686 => x"9c",
          3687 => x"27",
          3688 => x"75",
          3689 => x"16",
          3690 => x"17",
          3691 => x"33",
          3692 => x"70",
          3693 => x"55",
          3694 => x"80",
          3695 => x"73",
          3696 => x"cc",
          3697 => x"cb",
          3698 => x"81",
          3699 => x"94",
          3700 => x"a4",
          3701 => x"39",
          3702 => x"51",
          3703 => x"81",
          3704 => x"54",
          3705 => x"be",
          3706 => x"27",
          3707 => x"53",
          3708 => x"08",
          3709 => x"73",
          3710 => x"ff",
          3711 => x"15",
          3712 => x"16",
          3713 => x"ff",
          3714 => x"80",
          3715 => x"73",
          3716 => x"c6",
          3717 => x"cb",
          3718 => x"38",
          3719 => x"16",
          3720 => x"80",
          3721 => x"0b",
          3722 => x"81",
          3723 => x"75",
          3724 => x"cb",
          3725 => x"58",
          3726 => x"54",
          3727 => x"74",
          3728 => x"73",
          3729 => x"90",
          3730 => x"c0",
          3731 => x"90",
          3732 => x"83",
          3733 => x"72",
          3734 => x"38",
          3735 => x"08",
          3736 => x"77",
          3737 => x"80",
          3738 => x"cb",
          3739 => x"3d",
          3740 => x"3d",
          3741 => x"89",
          3742 => x"2e",
          3743 => x"80",
          3744 => x"fc",
          3745 => x"3d",
          3746 => x"e1",
          3747 => x"cb",
          3748 => x"81",
          3749 => x"80",
          3750 => x"76",
          3751 => x"75",
          3752 => x"3f",
          3753 => x"08",
          3754 => x"a4",
          3755 => x"38",
          3756 => x"70",
          3757 => x"57",
          3758 => x"a2",
          3759 => x"33",
          3760 => x"70",
          3761 => x"55",
          3762 => x"2e",
          3763 => x"16",
          3764 => x"51",
          3765 => x"81",
          3766 => x"88",
          3767 => x"54",
          3768 => x"84",
          3769 => x"52",
          3770 => x"e5",
          3771 => x"a4",
          3772 => x"84",
          3773 => x"06",
          3774 => x"55",
          3775 => x"80",
          3776 => x"80",
          3777 => x"54",
          3778 => x"a4",
          3779 => x"0d",
          3780 => x"0d",
          3781 => x"fc",
          3782 => x"52",
          3783 => x"3f",
          3784 => x"08",
          3785 => x"cb",
          3786 => x"0c",
          3787 => x"04",
          3788 => x"77",
          3789 => x"fc",
          3790 => x"53",
          3791 => x"de",
          3792 => x"a4",
          3793 => x"cb",
          3794 => x"df",
          3795 => x"38",
          3796 => x"08",
          3797 => x"cd",
          3798 => x"cb",
          3799 => x"80",
          3800 => x"cb",
          3801 => x"73",
          3802 => x"3f",
          3803 => x"08",
          3804 => x"a4",
          3805 => x"09",
          3806 => x"38",
          3807 => x"39",
          3808 => x"08",
          3809 => x"52",
          3810 => x"b3",
          3811 => x"73",
          3812 => x"3f",
          3813 => x"08",
          3814 => x"30",
          3815 => x"9f",
          3816 => x"cb",
          3817 => x"51",
          3818 => x"72",
          3819 => x"0c",
          3820 => x"04",
          3821 => x"65",
          3822 => x"89",
          3823 => x"96",
          3824 => x"df",
          3825 => x"cb",
          3826 => x"81",
          3827 => x"b2",
          3828 => x"75",
          3829 => x"3f",
          3830 => x"08",
          3831 => x"a4",
          3832 => x"02",
          3833 => x"33",
          3834 => x"55",
          3835 => x"25",
          3836 => x"55",
          3837 => x"80",
          3838 => x"76",
          3839 => x"d4",
          3840 => x"81",
          3841 => x"94",
          3842 => x"f0",
          3843 => x"65",
          3844 => x"53",
          3845 => x"05",
          3846 => x"51",
          3847 => x"81",
          3848 => x"5b",
          3849 => x"08",
          3850 => x"7c",
          3851 => x"08",
          3852 => x"fe",
          3853 => x"08",
          3854 => x"55",
          3855 => x"91",
          3856 => x"0c",
          3857 => x"81",
          3858 => x"39",
          3859 => x"c7",
          3860 => x"a4",
          3861 => x"55",
          3862 => x"2e",
          3863 => x"bf",
          3864 => x"5f",
          3865 => x"92",
          3866 => x"51",
          3867 => x"81",
          3868 => x"ff",
          3869 => x"81",
          3870 => x"81",
          3871 => x"81",
          3872 => x"30",
          3873 => x"a4",
          3874 => x"25",
          3875 => x"19",
          3876 => x"5a",
          3877 => x"08",
          3878 => x"38",
          3879 => x"a4",
          3880 => x"cb",
          3881 => x"58",
          3882 => x"77",
          3883 => x"7d",
          3884 => x"bf",
          3885 => x"cb",
          3886 => x"81",
          3887 => x"80",
          3888 => x"70",
          3889 => x"ff",
          3890 => x"56",
          3891 => x"2e",
          3892 => x"9e",
          3893 => x"51",
          3894 => x"3f",
          3895 => x"08",
          3896 => x"06",
          3897 => x"80",
          3898 => x"19",
          3899 => x"54",
          3900 => x"14",
          3901 => x"c5",
          3902 => x"a4",
          3903 => x"06",
          3904 => x"80",
          3905 => x"19",
          3906 => x"54",
          3907 => x"06",
          3908 => x"79",
          3909 => x"78",
          3910 => x"79",
          3911 => x"84",
          3912 => x"07",
          3913 => x"84",
          3914 => x"81",
          3915 => x"92",
          3916 => x"f9",
          3917 => x"8a",
          3918 => x"53",
          3919 => x"e3",
          3920 => x"cb",
          3921 => x"81",
          3922 => x"81",
          3923 => x"17",
          3924 => x"81",
          3925 => x"17",
          3926 => x"2a",
          3927 => x"51",
          3928 => x"55",
          3929 => x"81",
          3930 => x"17",
          3931 => x"8c",
          3932 => x"81",
          3933 => x"9b",
          3934 => x"a4",
          3935 => x"17",
          3936 => x"51",
          3937 => x"81",
          3938 => x"74",
          3939 => x"56",
          3940 => x"98",
          3941 => x"76",
          3942 => x"c6",
          3943 => x"a4",
          3944 => x"09",
          3945 => x"38",
          3946 => x"cb",
          3947 => x"2e",
          3948 => x"85",
          3949 => x"a3",
          3950 => x"38",
          3951 => x"cb",
          3952 => x"15",
          3953 => x"38",
          3954 => x"53",
          3955 => x"08",
          3956 => x"c3",
          3957 => x"cb",
          3958 => x"94",
          3959 => x"18",
          3960 => x"33",
          3961 => x"54",
          3962 => x"34",
          3963 => x"85",
          3964 => x"18",
          3965 => x"74",
          3966 => x"0c",
          3967 => x"04",
          3968 => x"82",
          3969 => x"ff",
          3970 => x"a1",
          3971 => x"e4",
          3972 => x"a4",
          3973 => x"cb",
          3974 => x"f5",
          3975 => x"a1",
          3976 => x"95",
          3977 => x"58",
          3978 => x"81",
          3979 => x"55",
          3980 => x"08",
          3981 => x"02",
          3982 => x"33",
          3983 => x"70",
          3984 => x"55",
          3985 => x"73",
          3986 => x"75",
          3987 => x"80",
          3988 => x"bd",
          3989 => x"d6",
          3990 => x"81",
          3991 => x"87",
          3992 => x"ad",
          3993 => x"78",
          3994 => x"3f",
          3995 => x"08",
          3996 => x"70",
          3997 => x"55",
          3998 => x"2e",
          3999 => x"78",
          4000 => x"a4",
          4001 => x"08",
          4002 => x"38",
          4003 => x"cb",
          4004 => x"76",
          4005 => x"70",
          4006 => x"b5",
          4007 => x"a4",
          4008 => x"cb",
          4009 => x"e9",
          4010 => x"a4",
          4011 => x"51",
          4012 => x"81",
          4013 => x"55",
          4014 => x"08",
          4015 => x"55",
          4016 => x"81",
          4017 => x"84",
          4018 => x"81",
          4019 => x"80",
          4020 => x"51",
          4021 => x"81",
          4022 => x"81",
          4023 => x"30",
          4024 => x"a4",
          4025 => x"25",
          4026 => x"75",
          4027 => x"38",
          4028 => x"8f",
          4029 => x"75",
          4030 => x"c1",
          4031 => x"cb",
          4032 => x"74",
          4033 => x"51",
          4034 => x"3f",
          4035 => x"08",
          4036 => x"cb",
          4037 => x"3d",
          4038 => x"3d",
          4039 => x"99",
          4040 => x"52",
          4041 => x"d8",
          4042 => x"cb",
          4043 => x"81",
          4044 => x"82",
          4045 => x"5e",
          4046 => x"3d",
          4047 => x"cf",
          4048 => x"cb",
          4049 => x"81",
          4050 => x"86",
          4051 => x"82",
          4052 => x"cb",
          4053 => x"2e",
          4054 => x"82",
          4055 => x"80",
          4056 => x"70",
          4057 => x"06",
          4058 => x"54",
          4059 => x"38",
          4060 => x"52",
          4061 => x"52",
          4062 => x"3f",
          4063 => x"08",
          4064 => x"81",
          4065 => x"83",
          4066 => x"81",
          4067 => x"81",
          4068 => x"06",
          4069 => x"54",
          4070 => x"08",
          4071 => x"81",
          4072 => x"81",
          4073 => x"39",
          4074 => x"38",
          4075 => x"08",
          4076 => x"c4",
          4077 => x"cb",
          4078 => x"81",
          4079 => x"81",
          4080 => x"53",
          4081 => x"19",
          4082 => x"8c",
          4083 => x"ae",
          4084 => x"34",
          4085 => x"0b",
          4086 => x"82",
          4087 => x"52",
          4088 => x"51",
          4089 => x"3f",
          4090 => x"b4",
          4091 => x"c9",
          4092 => x"53",
          4093 => x"53",
          4094 => x"51",
          4095 => x"3f",
          4096 => x"0b",
          4097 => x"34",
          4098 => x"80",
          4099 => x"51",
          4100 => x"78",
          4101 => x"83",
          4102 => x"51",
          4103 => x"81",
          4104 => x"54",
          4105 => x"08",
          4106 => x"88",
          4107 => x"64",
          4108 => x"ff",
          4109 => x"75",
          4110 => x"78",
          4111 => x"3f",
          4112 => x"0b",
          4113 => x"78",
          4114 => x"83",
          4115 => x"51",
          4116 => x"3f",
          4117 => x"08",
          4118 => x"80",
          4119 => x"76",
          4120 => x"ae",
          4121 => x"cb",
          4122 => x"3d",
          4123 => x"3d",
          4124 => x"84",
          4125 => x"f1",
          4126 => x"a8",
          4127 => x"05",
          4128 => x"51",
          4129 => x"81",
          4130 => x"55",
          4131 => x"08",
          4132 => x"78",
          4133 => x"08",
          4134 => x"70",
          4135 => x"b8",
          4136 => x"a4",
          4137 => x"cb",
          4138 => x"b9",
          4139 => x"9b",
          4140 => x"a0",
          4141 => x"55",
          4142 => x"38",
          4143 => x"3d",
          4144 => x"3d",
          4145 => x"51",
          4146 => x"3f",
          4147 => x"52",
          4148 => x"52",
          4149 => x"dd",
          4150 => x"08",
          4151 => x"cb",
          4152 => x"cb",
          4153 => x"81",
          4154 => x"95",
          4155 => x"2e",
          4156 => x"88",
          4157 => x"3d",
          4158 => x"38",
          4159 => x"e5",
          4160 => x"a4",
          4161 => x"09",
          4162 => x"b8",
          4163 => x"c9",
          4164 => x"cb",
          4165 => x"81",
          4166 => x"81",
          4167 => x"56",
          4168 => x"3d",
          4169 => x"52",
          4170 => x"ff",
          4171 => x"02",
          4172 => x"8b",
          4173 => x"16",
          4174 => x"2a",
          4175 => x"51",
          4176 => x"89",
          4177 => x"07",
          4178 => x"17",
          4179 => x"81",
          4180 => x"34",
          4181 => x"70",
          4182 => x"81",
          4183 => x"55",
          4184 => x"80",
          4185 => x"64",
          4186 => x"38",
          4187 => x"51",
          4188 => x"81",
          4189 => x"52",
          4190 => x"b7",
          4191 => x"55",
          4192 => x"08",
          4193 => x"dd",
          4194 => x"a4",
          4195 => x"51",
          4196 => x"3f",
          4197 => x"08",
          4198 => x"11",
          4199 => x"81",
          4200 => x"80",
          4201 => x"16",
          4202 => x"ae",
          4203 => x"06",
          4204 => x"53",
          4205 => x"51",
          4206 => x"78",
          4207 => x"83",
          4208 => x"39",
          4209 => x"08",
          4210 => x"51",
          4211 => x"81",
          4212 => x"55",
          4213 => x"08",
          4214 => x"51",
          4215 => x"3f",
          4216 => x"08",
          4217 => x"cb",
          4218 => x"3d",
          4219 => x"3d",
          4220 => x"db",
          4221 => x"84",
          4222 => x"05",
          4223 => x"82",
          4224 => x"d0",
          4225 => x"3d",
          4226 => x"3f",
          4227 => x"08",
          4228 => x"a4",
          4229 => x"38",
          4230 => x"52",
          4231 => x"05",
          4232 => x"3f",
          4233 => x"08",
          4234 => x"a4",
          4235 => x"02",
          4236 => x"33",
          4237 => x"54",
          4238 => x"aa",
          4239 => x"06",
          4240 => x"8b",
          4241 => x"06",
          4242 => x"07",
          4243 => x"56",
          4244 => x"34",
          4245 => x"0b",
          4246 => x"78",
          4247 => x"a9",
          4248 => x"a4",
          4249 => x"81",
          4250 => x"95",
          4251 => x"ef",
          4252 => x"56",
          4253 => x"3d",
          4254 => x"94",
          4255 => x"f4",
          4256 => x"a4",
          4257 => x"cb",
          4258 => x"cb",
          4259 => x"63",
          4260 => x"d4",
          4261 => x"c0",
          4262 => x"a4",
          4263 => x"cb",
          4264 => x"38",
          4265 => x"05",
          4266 => x"06",
          4267 => x"73",
          4268 => x"16",
          4269 => x"22",
          4270 => x"07",
          4271 => x"1f",
          4272 => x"c2",
          4273 => x"81",
          4274 => x"34",
          4275 => x"b3",
          4276 => x"cb",
          4277 => x"74",
          4278 => x"0c",
          4279 => x"04",
          4280 => x"69",
          4281 => x"80",
          4282 => x"d0",
          4283 => x"3d",
          4284 => x"3f",
          4285 => x"08",
          4286 => x"08",
          4287 => x"cb",
          4288 => x"80",
          4289 => x"57",
          4290 => x"81",
          4291 => x"70",
          4292 => x"55",
          4293 => x"80",
          4294 => x"5d",
          4295 => x"52",
          4296 => x"52",
          4297 => x"a9",
          4298 => x"a4",
          4299 => x"cb",
          4300 => x"d1",
          4301 => x"73",
          4302 => x"3f",
          4303 => x"08",
          4304 => x"a4",
          4305 => x"81",
          4306 => x"81",
          4307 => x"65",
          4308 => x"78",
          4309 => x"7b",
          4310 => x"55",
          4311 => x"34",
          4312 => x"8a",
          4313 => x"38",
          4314 => x"1a",
          4315 => x"34",
          4316 => x"9e",
          4317 => x"70",
          4318 => x"51",
          4319 => x"a0",
          4320 => x"8e",
          4321 => x"2e",
          4322 => x"86",
          4323 => x"34",
          4324 => x"30",
          4325 => x"80",
          4326 => x"7a",
          4327 => x"c1",
          4328 => x"2e",
          4329 => x"a0",
          4330 => x"51",
          4331 => x"3f",
          4332 => x"08",
          4333 => x"a4",
          4334 => x"7b",
          4335 => x"55",
          4336 => x"73",
          4337 => x"38",
          4338 => x"73",
          4339 => x"38",
          4340 => x"15",
          4341 => x"ff",
          4342 => x"81",
          4343 => x"7b",
          4344 => x"cb",
          4345 => x"3d",
          4346 => x"3d",
          4347 => x"9c",
          4348 => x"05",
          4349 => x"51",
          4350 => x"81",
          4351 => x"81",
          4352 => x"56",
          4353 => x"a4",
          4354 => x"38",
          4355 => x"52",
          4356 => x"52",
          4357 => x"c0",
          4358 => x"70",
          4359 => x"ff",
          4360 => x"55",
          4361 => x"27",
          4362 => x"78",
          4363 => x"ff",
          4364 => x"05",
          4365 => x"55",
          4366 => x"3f",
          4367 => x"08",
          4368 => x"38",
          4369 => x"70",
          4370 => x"ff",
          4371 => x"81",
          4372 => x"80",
          4373 => x"74",
          4374 => x"07",
          4375 => x"4e",
          4376 => x"81",
          4377 => x"55",
          4378 => x"70",
          4379 => x"06",
          4380 => x"99",
          4381 => x"e0",
          4382 => x"ff",
          4383 => x"54",
          4384 => x"27",
          4385 => x"ba",
          4386 => x"55",
          4387 => x"a3",
          4388 => x"81",
          4389 => x"ff",
          4390 => x"81",
          4391 => x"93",
          4392 => x"75",
          4393 => x"76",
          4394 => x"38",
          4395 => x"77",
          4396 => x"86",
          4397 => x"39",
          4398 => x"27",
          4399 => x"88",
          4400 => x"78",
          4401 => x"5a",
          4402 => x"57",
          4403 => x"81",
          4404 => x"81",
          4405 => x"33",
          4406 => x"06",
          4407 => x"57",
          4408 => x"fe",
          4409 => x"3d",
          4410 => x"55",
          4411 => x"2e",
          4412 => x"76",
          4413 => x"38",
          4414 => x"55",
          4415 => x"33",
          4416 => x"a0",
          4417 => x"06",
          4418 => x"17",
          4419 => x"38",
          4420 => x"43",
          4421 => x"3d",
          4422 => x"ff",
          4423 => x"81",
          4424 => x"54",
          4425 => x"08",
          4426 => x"81",
          4427 => x"ff",
          4428 => x"81",
          4429 => x"54",
          4430 => x"08",
          4431 => x"80",
          4432 => x"54",
          4433 => x"80",
          4434 => x"cb",
          4435 => x"2e",
          4436 => x"80",
          4437 => x"54",
          4438 => x"80",
          4439 => x"52",
          4440 => x"bd",
          4441 => x"cb",
          4442 => x"81",
          4443 => x"b1",
          4444 => x"81",
          4445 => x"52",
          4446 => x"ab",
          4447 => x"54",
          4448 => x"15",
          4449 => x"78",
          4450 => x"ff",
          4451 => x"79",
          4452 => x"83",
          4453 => x"51",
          4454 => x"3f",
          4455 => x"08",
          4456 => x"74",
          4457 => x"0c",
          4458 => x"04",
          4459 => x"60",
          4460 => x"05",
          4461 => x"33",
          4462 => x"05",
          4463 => x"40",
          4464 => x"da",
          4465 => x"a4",
          4466 => x"cb",
          4467 => x"bd",
          4468 => x"33",
          4469 => x"b5",
          4470 => x"2e",
          4471 => x"1a",
          4472 => x"90",
          4473 => x"33",
          4474 => x"70",
          4475 => x"55",
          4476 => x"38",
          4477 => x"97",
          4478 => x"82",
          4479 => x"58",
          4480 => x"7e",
          4481 => x"70",
          4482 => x"55",
          4483 => x"56",
          4484 => x"8a",
          4485 => x"7d",
          4486 => x"70",
          4487 => x"2a",
          4488 => x"08",
          4489 => x"08",
          4490 => x"5d",
          4491 => x"77",
          4492 => x"98",
          4493 => x"26",
          4494 => x"57",
          4495 => x"59",
          4496 => x"52",
          4497 => x"ae",
          4498 => x"15",
          4499 => x"98",
          4500 => x"26",
          4501 => x"55",
          4502 => x"08",
          4503 => x"99",
          4504 => x"a4",
          4505 => x"ff",
          4506 => x"cb",
          4507 => x"38",
          4508 => x"75",
          4509 => x"81",
          4510 => x"93",
          4511 => x"80",
          4512 => x"2e",
          4513 => x"ff",
          4514 => x"58",
          4515 => x"7d",
          4516 => x"38",
          4517 => x"55",
          4518 => x"b4",
          4519 => x"56",
          4520 => x"09",
          4521 => x"38",
          4522 => x"53",
          4523 => x"51",
          4524 => x"3f",
          4525 => x"08",
          4526 => x"a4",
          4527 => x"38",
          4528 => x"ff",
          4529 => x"5c",
          4530 => x"84",
          4531 => x"5c",
          4532 => x"12",
          4533 => x"80",
          4534 => x"78",
          4535 => x"7c",
          4536 => x"90",
          4537 => x"c0",
          4538 => x"90",
          4539 => x"15",
          4540 => x"90",
          4541 => x"54",
          4542 => x"91",
          4543 => x"31",
          4544 => x"84",
          4545 => x"07",
          4546 => x"16",
          4547 => x"73",
          4548 => x"0c",
          4549 => x"04",
          4550 => x"6b",
          4551 => x"05",
          4552 => x"33",
          4553 => x"5a",
          4554 => x"bd",
          4555 => x"80",
          4556 => x"a4",
          4557 => x"f8",
          4558 => x"a4",
          4559 => x"81",
          4560 => x"70",
          4561 => x"74",
          4562 => x"38",
          4563 => x"81",
          4564 => x"81",
          4565 => x"81",
          4566 => x"ff",
          4567 => x"81",
          4568 => x"81",
          4569 => x"81",
          4570 => x"83",
          4571 => x"c0",
          4572 => x"2a",
          4573 => x"51",
          4574 => x"74",
          4575 => x"99",
          4576 => x"53",
          4577 => x"51",
          4578 => x"3f",
          4579 => x"08",
          4580 => x"55",
          4581 => x"92",
          4582 => x"80",
          4583 => x"38",
          4584 => x"06",
          4585 => x"2e",
          4586 => x"48",
          4587 => x"87",
          4588 => x"79",
          4589 => x"78",
          4590 => x"26",
          4591 => x"19",
          4592 => x"74",
          4593 => x"38",
          4594 => x"e4",
          4595 => x"2a",
          4596 => x"70",
          4597 => x"59",
          4598 => x"7a",
          4599 => x"56",
          4600 => x"80",
          4601 => x"51",
          4602 => x"74",
          4603 => x"99",
          4604 => x"53",
          4605 => x"51",
          4606 => x"3f",
          4607 => x"cb",
          4608 => x"ac",
          4609 => x"2a",
          4610 => x"81",
          4611 => x"43",
          4612 => x"83",
          4613 => x"66",
          4614 => x"60",
          4615 => x"90",
          4616 => x"31",
          4617 => x"80",
          4618 => x"8a",
          4619 => x"56",
          4620 => x"26",
          4621 => x"77",
          4622 => x"81",
          4623 => x"74",
          4624 => x"38",
          4625 => x"55",
          4626 => x"83",
          4627 => x"81",
          4628 => x"80",
          4629 => x"38",
          4630 => x"55",
          4631 => x"5e",
          4632 => x"89",
          4633 => x"5a",
          4634 => x"09",
          4635 => x"e1",
          4636 => x"38",
          4637 => x"57",
          4638 => x"bc",
          4639 => x"5a",
          4640 => x"9d",
          4641 => x"26",
          4642 => x"bc",
          4643 => x"10",
          4644 => x"22",
          4645 => x"74",
          4646 => x"38",
          4647 => x"ee",
          4648 => x"66",
          4649 => x"f6",
          4650 => x"a4",
          4651 => x"84",
          4652 => x"89",
          4653 => x"a0",
          4654 => x"81",
          4655 => x"fc",
          4656 => x"56",
          4657 => x"f0",
          4658 => x"80",
          4659 => x"d3",
          4660 => x"38",
          4661 => x"57",
          4662 => x"bc",
          4663 => x"5a",
          4664 => x"9d",
          4665 => x"26",
          4666 => x"bc",
          4667 => x"10",
          4668 => x"22",
          4669 => x"74",
          4670 => x"38",
          4671 => x"ee",
          4672 => x"66",
          4673 => x"96",
          4674 => x"a4",
          4675 => x"05",
          4676 => x"a4",
          4677 => x"26",
          4678 => x"0b",
          4679 => x"08",
          4680 => x"a4",
          4681 => x"11",
          4682 => x"05",
          4683 => x"83",
          4684 => x"2a",
          4685 => x"a0",
          4686 => x"7d",
          4687 => x"69",
          4688 => x"05",
          4689 => x"72",
          4690 => x"5c",
          4691 => x"59",
          4692 => x"2e",
          4693 => x"89",
          4694 => x"60",
          4695 => x"84",
          4696 => x"5d",
          4697 => x"18",
          4698 => x"68",
          4699 => x"74",
          4700 => x"af",
          4701 => x"31",
          4702 => x"53",
          4703 => x"52",
          4704 => x"9a",
          4705 => x"a4",
          4706 => x"83",
          4707 => x"06",
          4708 => x"cb",
          4709 => x"ff",
          4710 => x"dd",
          4711 => x"83",
          4712 => x"2a",
          4713 => x"be",
          4714 => x"39",
          4715 => x"09",
          4716 => x"c5",
          4717 => x"f5",
          4718 => x"a4",
          4719 => x"38",
          4720 => x"79",
          4721 => x"80",
          4722 => x"38",
          4723 => x"96",
          4724 => x"06",
          4725 => x"2e",
          4726 => x"5e",
          4727 => x"81",
          4728 => x"9f",
          4729 => x"38",
          4730 => x"38",
          4731 => x"81",
          4732 => x"fc",
          4733 => x"ab",
          4734 => x"7d",
          4735 => x"81",
          4736 => x"7d",
          4737 => x"78",
          4738 => x"74",
          4739 => x"8e",
          4740 => x"9c",
          4741 => x"53",
          4742 => x"51",
          4743 => x"3f",
          4744 => x"ba",
          4745 => x"51",
          4746 => x"3f",
          4747 => x"8b",
          4748 => x"a1",
          4749 => x"8d",
          4750 => x"83",
          4751 => x"52",
          4752 => x"ff",
          4753 => x"81",
          4754 => x"34",
          4755 => x"70",
          4756 => x"2a",
          4757 => x"54",
          4758 => x"1b",
          4759 => x"88",
          4760 => x"74",
          4761 => x"26",
          4762 => x"83",
          4763 => x"52",
          4764 => x"ff",
          4765 => x"8a",
          4766 => x"a0",
          4767 => x"a1",
          4768 => x"0b",
          4769 => x"bf",
          4770 => x"51",
          4771 => x"3f",
          4772 => x"9a",
          4773 => x"a0",
          4774 => x"52",
          4775 => x"ff",
          4776 => x"7d",
          4777 => x"81",
          4778 => x"38",
          4779 => x"0a",
          4780 => x"1b",
          4781 => x"ce",
          4782 => x"a4",
          4783 => x"a0",
          4784 => x"52",
          4785 => x"ff",
          4786 => x"81",
          4787 => x"51",
          4788 => x"3f",
          4789 => x"1b",
          4790 => x"8c",
          4791 => x"0b",
          4792 => x"34",
          4793 => x"c2",
          4794 => x"53",
          4795 => x"52",
          4796 => x"51",
          4797 => x"88",
          4798 => x"a7",
          4799 => x"a0",
          4800 => x"83",
          4801 => x"52",
          4802 => x"ff",
          4803 => x"ff",
          4804 => x"1c",
          4805 => x"a6",
          4806 => x"53",
          4807 => x"52",
          4808 => x"ff",
          4809 => x"82",
          4810 => x"83",
          4811 => x"52",
          4812 => x"b4",
          4813 => x"60",
          4814 => x"7e",
          4815 => x"d7",
          4816 => x"81",
          4817 => x"83",
          4818 => x"83",
          4819 => x"06",
          4820 => x"75",
          4821 => x"05",
          4822 => x"7e",
          4823 => x"b7",
          4824 => x"53",
          4825 => x"51",
          4826 => x"3f",
          4827 => x"a4",
          4828 => x"51",
          4829 => x"3f",
          4830 => x"e4",
          4831 => x"e4",
          4832 => x"9f",
          4833 => x"18",
          4834 => x"1b",
          4835 => x"f6",
          4836 => x"83",
          4837 => x"ff",
          4838 => x"82",
          4839 => x"78",
          4840 => x"c4",
          4841 => x"60",
          4842 => x"7a",
          4843 => x"ff",
          4844 => x"75",
          4845 => x"53",
          4846 => x"51",
          4847 => x"3f",
          4848 => x"52",
          4849 => x"9f",
          4850 => x"56",
          4851 => x"83",
          4852 => x"06",
          4853 => x"52",
          4854 => x"9e",
          4855 => x"52",
          4856 => x"ff",
          4857 => x"f0",
          4858 => x"1b",
          4859 => x"87",
          4860 => x"55",
          4861 => x"83",
          4862 => x"74",
          4863 => x"ff",
          4864 => x"7c",
          4865 => x"74",
          4866 => x"38",
          4867 => x"54",
          4868 => x"52",
          4869 => x"99",
          4870 => x"cb",
          4871 => x"87",
          4872 => x"53",
          4873 => x"08",
          4874 => x"ff",
          4875 => x"76",
          4876 => x"31",
          4877 => x"cd",
          4878 => x"58",
          4879 => x"ff",
          4880 => x"55",
          4881 => x"83",
          4882 => x"61",
          4883 => x"26",
          4884 => x"57",
          4885 => x"53",
          4886 => x"51",
          4887 => x"3f",
          4888 => x"08",
          4889 => x"76",
          4890 => x"31",
          4891 => x"db",
          4892 => x"7d",
          4893 => x"38",
          4894 => x"83",
          4895 => x"8a",
          4896 => x"7d",
          4897 => x"38",
          4898 => x"81",
          4899 => x"80",
          4900 => x"80",
          4901 => x"7a",
          4902 => x"bc",
          4903 => x"d5",
          4904 => x"ff",
          4905 => x"83",
          4906 => x"77",
          4907 => x"0b",
          4908 => x"81",
          4909 => x"34",
          4910 => x"34",
          4911 => x"34",
          4912 => x"56",
          4913 => x"52",
          4914 => x"f4",
          4915 => x"0b",
          4916 => x"81",
          4917 => x"82",
          4918 => x"56",
          4919 => x"34",
          4920 => x"08",
          4921 => x"60",
          4922 => x"1b",
          4923 => x"96",
          4924 => x"83",
          4925 => x"ff",
          4926 => x"81",
          4927 => x"7a",
          4928 => x"ff",
          4929 => x"81",
          4930 => x"a4",
          4931 => x"80",
          4932 => x"7e",
          4933 => x"e3",
          4934 => x"81",
          4935 => x"90",
          4936 => x"8e",
          4937 => x"81",
          4938 => x"81",
          4939 => x"56",
          4940 => x"a4",
          4941 => x"0d",
          4942 => x"0d",
          4943 => x"93",
          4944 => x"38",
          4945 => x"81",
          4946 => x"52",
          4947 => x"81",
          4948 => x"81",
          4949 => x"bd",
          4950 => x"f9",
          4951 => x"dc",
          4952 => x"39",
          4953 => x"51",
          4954 => x"81",
          4955 => x"80",
          4956 => x"be",
          4957 => x"dd",
          4958 => x"a4",
          4959 => x"39",
          4960 => x"51",
          4961 => x"81",
          4962 => x"80",
          4963 => x"be",
          4964 => x"c1",
          4965 => x"fc",
          4966 => x"81",
          4967 => x"b5",
          4968 => x"ac",
          4969 => x"81",
          4970 => x"a9",
          4971 => x"ec",
          4972 => x"81",
          4973 => x"9d",
          4974 => x"a0",
          4975 => x"81",
          4976 => x"91",
          4977 => x"d0",
          4978 => x"81",
          4979 => x"85",
          4980 => x"f4",
          4981 => x"fb",
          4982 => x"0d",
          4983 => x"0d",
          4984 => x"56",
          4985 => x"26",
          4986 => x"52",
          4987 => x"29",
          4988 => x"87",
          4989 => x"51",
          4990 => x"3f",
          4991 => x"08",
          4992 => x"fe",
          4993 => x"81",
          4994 => x"54",
          4995 => x"52",
          4996 => x"51",
          4997 => x"3f",
          4998 => x"04",
          4999 => x"7d",
          5000 => x"8c",
          5001 => x"05",
          5002 => x"15",
          5003 => x"5a",
          5004 => x"5c",
          5005 => x"c1",
          5006 => x"8c",
          5007 => x"c1",
          5008 => x"87",
          5009 => x"55",
          5010 => x"80",
          5011 => x"90",
          5012 => x"79",
          5013 => x"38",
          5014 => x"74",
          5015 => x"78",
          5016 => x"72",
          5017 => x"c1",
          5018 => x"8c",
          5019 => x"39",
          5020 => x"51",
          5021 => x"3f",
          5022 => x"80",
          5023 => x"16",
          5024 => x"27",
          5025 => x"08",
          5026 => x"a8",
          5027 => x"a7",
          5028 => x"81",
          5029 => x"ff",
          5030 => x"84",
          5031 => x"39",
          5032 => x"72",
          5033 => x"38",
          5034 => x"81",
          5035 => x"ff",
          5036 => x"89",
          5037 => x"d0",
          5038 => x"97",
          5039 => x"55",
          5040 => x"fa",
          5041 => x"80",
          5042 => x"d4",
          5043 => x"83",
          5044 => x"74",
          5045 => x"38",
          5046 => x"33",
          5047 => x"52",
          5048 => x"74",
          5049 => x"72",
          5050 => x"38",
          5051 => x"26",
          5052 => x"51",
          5053 => x"51",
          5054 => x"3f",
          5055 => x"d3",
          5056 => x"d8",
          5057 => x"cb",
          5058 => x"77",
          5059 => x"fe",
          5060 => x"81",
          5061 => x"98",
          5062 => x"2c",
          5063 => x"a0",
          5064 => x"06",
          5065 => x"fc",
          5066 => x"cb",
          5067 => x"2b",
          5068 => x"70",
          5069 => x"30",
          5070 => x"9f",
          5071 => x"56",
          5072 => x"9b",
          5073 => x"72",
          5074 => x"9b",
          5075 => x"06",
          5076 => x"53",
          5077 => x"1c",
          5078 => x"26",
          5079 => x"ff",
          5080 => x"cb",
          5081 => x"3d",
          5082 => x"3d",
          5083 => x"84",
          5084 => x"05",
          5085 => x"30",
          5086 => x"80",
          5087 => x"ff",
          5088 => x"51",
          5089 => x"5b",
          5090 => x"74",
          5091 => x"81",
          5092 => x"8c",
          5093 => x"57",
          5094 => x"81",
          5095 => x"56",
          5096 => x"08",
          5097 => x"cb",
          5098 => x"c0",
          5099 => x"81",
          5100 => x"59",
          5101 => x"05",
          5102 => x"53",
          5103 => x"51",
          5104 => x"81",
          5105 => x"56",
          5106 => x"08",
          5107 => x"55",
          5108 => x"89",
          5109 => x"75",
          5110 => x"d8",
          5111 => x"d8",
          5112 => x"e0",
          5113 => x"70",
          5114 => x"25",
          5115 => x"80",
          5116 => x"74",
          5117 => x"38",
          5118 => x"53",
          5119 => x"88",
          5120 => x"51",
          5121 => x"75",
          5122 => x"cb",
          5123 => x"3d",
          5124 => x"3d",
          5125 => x"84",
          5126 => x"33",
          5127 => x"57",
          5128 => x"52",
          5129 => x"c2",
          5130 => x"a4",
          5131 => x"75",
          5132 => x"38",
          5133 => x"98",
          5134 => x"60",
          5135 => x"81",
          5136 => x"7e",
          5137 => x"77",
          5138 => x"a4",
          5139 => x"39",
          5140 => x"81",
          5141 => x"89",
          5142 => x"fc",
          5143 => x"9b",
          5144 => x"c1",
          5145 => x"c1",
          5146 => x"ff",
          5147 => x"81",
          5148 => x"51",
          5149 => x"3f",
          5150 => x"54",
          5151 => x"53",
          5152 => x"33",
          5153 => x"8c",
          5154 => x"ab",
          5155 => x"2e",
          5156 => x"fe",
          5157 => x"3d",
          5158 => x"3d",
          5159 => x"96",
          5160 => x"ff",
          5161 => x"81",
          5162 => x"8c",
          5163 => x"a8",
          5164 => x"84",
          5165 => x"fe",
          5166 => x"72",
          5167 => x"81",
          5168 => x"71",
          5169 => x"38",
          5170 => x"f5",
          5171 => x"c2",
          5172 => x"f7",
          5173 => x"51",
          5174 => x"3f",
          5175 => x"70",
          5176 => x"52",
          5177 => x"95",
          5178 => x"fe",
          5179 => x"81",
          5180 => x"fe",
          5181 => x"80",
          5182 => x"bc",
          5183 => x"2a",
          5184 => x"51",
          5185 => x"2e",
          5186 => x"51",
          5187 => x"3f",
          5188 => x"51",
          5189 => x"3f",
          5190 => x"f5",
          5191 => x"84",
          5192 => x"06",
          5193 => x"80",
          5194 => x"81",
          5195 => x"88",
          5196 => x"fc",
          5197 => x"80",
          5198 => x"fe",
          5199 => x"72",
          5200 => x"81",
          5201 => x"71",
          5202 => x"38",
          5203 => x"f4",
          5204 => x"c3",
          5205 => x"f6",
          5206 => x"51",
          5207 => x"3f",
          5208 => x"70",
          5209 => x"52",
          5210 => x"95",
          5211 => x"fe",
          5212 => x"81",
          5213 => x"fe",
          5214 => x"80",
          5215 => x"b8",
          5216 => x"2a",
          5217 => x"51",
          5218 => x"2e",
          5219 => x"51",
          5220 => x"3f",
          5221 => x"51",
          5222 => x"3f",
          5223 => x"f4",
          5224 => x"88",
          5225 => x"06",
          5226 => x"80",
          5227 => x"81",
          5228 => x"84",
          5229 => x"cc",
          5230 => x"fc",
          5231 => x"fe",
          5232 => x"fe",
          5233 => x"84",
          5234 => x"fa",
          5235 => x"70",
          5236 => x"55",
          5237 => x"2e",
          5238 => x"8e",
          5239 => x"0c",
          5240 => x"53",
          5241 => x"81",
          5242 => x"74",
          5243 => x"ff",
          5244 => x"53",
          5245 => x"83",
          5246 => x"74",
          5247 => x"38",
          5248 => x"75",
          5249 => x"53",
          5250 => x"09",
          5251 => x"38",
          5252 => x"81",
          5253 => x"80",
          5254 => x"29",
          5255 => x"05",
          5256 => x"70",
          5257 => x"fe",
          5258 => x"81",
          5259 => x"8b",
          5260 => x"33",
          5261 => x"2e",
          5262 => x"81",
          5263 => x"ff",
          5264 => x"94",
          5265 => x"38",
          5266 => x"81",
          5267 => x"88",
          5268 => x"cb",
          5269 => x"70",
          5270 => x"a4",
          5271 => x"81",
          5272 => x"ff",
          5273 => x"81",
          5274 => x"81",
          5275 => x"78",
          5276 => x"81",
          5277 => x"81",
          5278 => x"99",
          5279 => x"59",
          5280 => x"3f",
          5281 => x"52",
          5282 => x"51",
          5283 => x"3f",
          5284 => x"08",
          5285 => x"38",
          5286 => x"51",
          5287 => x"81",
          5288 => x"81",
          5289 => x"fe",
          5290 => x"99",
          5291 => x"5a",
          5292 => x"80",
          5293 => x"fe",
          5294 => x"80",
          5295 => x"51",
          5296 => x"3f",
          5297 => x"f8",
          5298 => x"ff",
          5299 => x"a4",
          5300 => x"70",
          5301 => x"59",
          5302 => x"2e",
          5303 => x"78",
          5304 => x"80",
          5305 => x"ab",
          5306 => x"38",
          5307 => x"a4",
          5308 => x"2e",
          5309 => x"78",
          5310 => x"38",
          5311 => x"ff",
          5312 => x"88",
          5313 => x"2e",
          5314 => x"78",
          5315 => x"ad",
          5316 => x"39",
          5317 => x"2e",
          5318 => x"78",
          5319 => x"90",
          5320 => x"2e",
          5321 => x"78",
          5322 => x"8b",
          5323 => x"39",
          5324 => x"2e",
          5325 => x"78",
          5326 => x"88",
          5327 => x"cc",
          5328 => x"f8",
          5329 => x"38",
          5330 => x"24",
          5331 => x"80",
          5332 => x"e2",
          5333 => x"d1",
          5334 => x"78",
          5335 => x"8a",
          5336 => x"a8",
          5337 => x"d4",
          5338 => x"38",
          5339 => x"2e",
          5340 => x"8c",
          5341 => x"81",
          5342 => x"fc",
          5343 => x"83",
          5344 => x"78",
          5345 => x"8b",
          5346 => x"81",
          5347 => x"d9",
          5348 => x"39",
          5349 => x"2e",
          5350 => x"78",
          5351 => x"fe",
          5352 => x"e8",
          5353 => x"fe",
          5354 => x"fe",
          5355 => x"ff",
          5356 => x"81",
          5357 => x"88",
          5358 => x"cc",
          5359 => x"39",
          5360 => x"f0",
          5361 => x"f8",
          5362 => x"83",
          5363 => x"cb",
          5364 => x"2e",
          5365 => x"63",
          5366 => x"80",
          5367 => x"cb",
          5368 => x"02",
          5369 => x"33",
          5370 => x"c2",
          5371 => x"a4",
          5372 => x"06",
          5373 => x"38",
          5374 => x"51",
          5375 => x"3f",
          5376 => x"9f",
          5377 => x"ec",
          5378 => x"39",
          5379 => x"f4",
          5380 => x"f8",
          5381 => x"83",
          5382 => x"cb",
          5383 => x"2e",
          5384 => x"80",
          5385 => x"02",
          5386 => x"33",
          5387 => x"cb",
          5388 => x"a4",
          5389 => x"c5",
          5390 => x"a6",
          5391 => x"fe",
          5392 => x"fe",
          5393 => x"ff",
          5394 => x"81",
          5395 => x"80",
          5396 => x"63",
          5397 => x"cb",
          5398 => x"fe",
          5399 => x"fe",
          5400 => x"ff",
          5401 => x"81",
          5402 => x"86",
          5403 => x"a4",
          5404 => x"53",
          5405 => x"52",
          5406 => x"80",
          5407 => x"80",
          5408 => x"53",
          5409 => x"84",
          5410 => x"cc",
          5411 => x"ff",
          5412 => x"81",
          5413 => x"81",
          5414 => x"c4",
          5415 => x"fa",
          5416 => x"5c",
          5417 => x"b7",
          5418 => x"05",
          5419 => x"b9",
          5420 => x"a4",
          5421 => x"fe",
          5422 => x"5b",
          5423 => x"3f",
          5424 => x"cb",
          5425 => x"7a",
          5426 => x"3f",
          5427 => x"b7",
          5428 => x"05",
          5429 => x"91",
          5430 => x"a4",
          5431 => x"fe",
          5432 => x"5b",
          5433 => x"3f",
          5434 => x"08",
          5435 => x"f8",
          5436 => x"fe",
          5437 => x"81",
          5438 => x"b8",
          5439 => x"05",
          5440 => x"ea",
          5441 => x"c8",
          5442 => x"cb",
          5443 => x"56",
          5444 => x"cb",
          5445 => x"ff",
          5446 => x"53",
          5447 => x"51",
          5448 => x"81",
          5449 => x"80",
          5450 => x"38",
          5451 => x"08",
          5452 => x"3f",
          5453 => x"b7",
          5454 => x"11",
          5455 => x"05",
          5456 => x"e8",
          5457 => x"a4",
          5458 => x"fa",
          5459 => x"3d",
          5460 => x"53",
          5461 => x"51",
          5462 => x"3f",
          5463 => x"08",
          5464 => x"bf",
          5465 => x"fe",
          5466 => x"fe",
          5467 => x"ff",
          5468 => x"81",
          5469 => x"86",
          5470 => x"a4",
          5471 => x"c5",
          5472 => x"f8",
          5473 => x"63",
          5474 => x"7b",
          5475 => x"61",
          5476 => x"70",
          5477 => x"0c",
          5478 => x"f5",
          5479 => x"d8",
          5480 => x"39",
          5481 => x"f4",
          5482 => x"f8",
          5483 => x"ff",
          5484 => x"cb",
          5485 => x"c4",
          5486 => x"bd",
          5487 => x"80",
          5488 => x"81",
          5489 => x"44",
          5490 => x"c8",
          5491 => x"78",
          5492 => x"38",
          5493 => x"08",
          5494 => x"81",
          5495 => x"59",
          5496 => x"81",
          5497 => x"59",
          5498 => x"88",
          5499 => x"a0",
          5500 => x"39",
          5501 => x"08",
          5502 => x"44",
          5503 => x"f0",
          5504 => x"f8",
          5505 => x"ff",
          5506 => x"cb",
          5507 => x"c3",
          5508 => x"bd",
          5509 => x"80",
          5510 => x"81",
          5511 => x"43",
          5512 => x"c8",
          5513 => x"78",
          5514 => x"38",
          5515 => x"08",
          5516 => x"81",
          5517 => x"59",
          5518 => x"81",
          5519 => x"59",
          5520 => x"88",
          5521 => x"a4",
          5522 => x"39",
          5523 => x"08",
          5524 => x"b7",
          5525 => x"11",
          5526 => x"05",
          5527 => x"cc",
          5528 => x"a4",
          5529 => x"9b",
          5530 => x"5b",
          5531 => x"2e",
          5532 => x"59",
          5533 => x"8d",
          5534 => x"2e",
          5535 => x"a0",
          5536 => x"88",
          5537 => x"9c",
          5538 => x"c7",
          5539 => x"63",
          5540 => x"62",
          5541 => x"ef",
          5542 => x"c5",
          5543 => x"bd",
          5544 => x"fe",
          5545 => x"fe",
          5546 => x"fe",
          5547 => x"81",
          5548 => x"80",
          5549 => x"38",
          5550 => x"f0",
          5551 => x"f8",
          5552 => x"fd",
          5553 => x"cb",
          5554 => x"2e",
          5555 => x"59",
          5556 => x"05",
          5557 => x"63",
          5558 => x"b7",
          5559 => x"11",
          5560 => x"05",
          5561 => x"c4",
          5562 => x"a4",
          5563 => x"f7",
          5564 => x"70",
          5565 => x"81",
          5566 => x"fe",
          5567 => x"80",
          5568 => x"51",
          5569 => x"3f",
          5570 => x"33",
          5571 => x"2e",
          5572 => x"9f",
          5573 => x"38",
          5574 => x"f0",
          5575 => x"f8",
          5576 => x"fd",
          5577 => x"cb",
          5578 => x"2e",
          5579 => x"59",
          5580 => x"05",
          5581 => x"63",
          5582 => x"ff",
          5583 => x"c5",
          5584 => x"f5",
          5585 => x"aa",
          5586 => x"fe",
          5587 => x"fe",
          5588 => x"fe",
          5589 => x"81",
          5590 => x"80",
          5591 => x"38",
          5592 => x"e4",
          5593 => x"f8",
          5594 => x"fe",
          5595 => x"cb",
          5596 => x"2e",
          5597 => x"59",
          5598 => x"22",
          5599 => x"05",
          5600 => x"41",
          5601 => x"e4",
          5602 => x"f8",
          5603 => x"fe",
          5604 => x"cb",
          5605 => x"38",
          5606 => x"60",
          5607 => x"52",
          5608 => x"51",
          5609 => x"3f",
          5610 => x"79",
          5611 => x"e1",
          5612 => x"79",
          5613 => x"ae",
          5614 => x"38",
          5615 => x"87",
          5616 => x"05",
          5617 => x"b7",
          5618 => x"11",
          5619 => x"05",
          5620 => x"ca",
          5621 => x"a4",
          5622 => x"92",
          5623 => x"02",
          5624 => x"79",
          5625 => x"5b",
          5626 => x"ff",
          5627 => x"c5",
          5628 => x"f3",
          5629 => x"a3",
          5630 => x"fe",
          5631 => x"fe",
          5632 => x"fe",
          5633 => x"81",
          5634 => x"80",
          5635 => x"38",
          5636 => x"e4",
          5637 => x"f8",
          5638 => x"fd",
          5639 => x"cb",
          5640 => x"2e",
          5641 => x"60",
          5642 => x"60",
          5643 => x"b7",
          5644 => x"11",
          5645 => x"05",
          5646 => x"e2",
          5647 => x"a4",
          5648 => x"f4",
          5649 => x"70",
          5650 => x"81",
          5651 => x"fe",
          5652 => x"80",
          5653 => x"51",
          5654 => x"3f",
          5655 => x"33",
          5656 => x"2e",
          5657 => x"9f",
          5658 => x"38",
          5659 => x"e4",
          5660 => x"f8",
          5661 => x"fc",
          5662 => x"cb",
          5663 => x"2e",
          5664 => x"53",
          5665 => x"c5",
          5666 => x"f8",
          5667 => x"60",
          5668 => x"60",
          5669 => x"ff",
          5670 => x"c5",
          5671 => x"f2",
          5672 => x"a2",
          5673 => x"e4",
          5674 => x"a7",
          5675 => x"fe",
          5676 => x"f3",
          5677 => x"c5",
          5678 => x"f2",
          5679 => x"51",
          5680 => x"3f",
          5681 => x"84",
          5682 => x"87",
          5683 => x"0c",
          5684 => x"0b",
          5685 => x"94",
          5686 => x"94",
          5687 => x"f3",
          5688 => x"39",
          5689 => x"51",
          5690 => x"3f",
          5691 => x"0b",
          5692 => x"84",
          5693 => x"83",
          5694 => x"94",
          5695 => x"a3",
          5696 => x"fe",
          5697 => x"fe",
          5698 => x"fe",
          5699 => x"81",
          5700 => x"80",
          5701 => x"38",
          5702 => x"c6",
          5703 => x"f7",
          5704 => x"59",
          5705 => x"3d",
          5706 => x"53",
          5707 => x"51",
          5708 => x"3f",
          5709 => x"08",
          5710 => x"e7",
          5711 => x"81",
          5712 => x"fe",
          5713 => x"63",
          5714 => x"81",
          5715 => x"5e",
          5716 => x"08",
          5717 => x"cb",
          5718 => x"a4",
          5719 => x"c6",
          5720 => x"f6",
          5721 => x"bb",
          5722 => x"90",
          5723 => x"e3",
          5724 => x"8d",
          5725 => x"39",
          5726 => x"51",
          5727 => x"3f",
          5728 => x"a0",
          5729 => x"9f",
          5730 => x"39",
          5731 => x"51",
          5732 => x"2e",
          5733 => x"7b",
          5734 => x"d2",
          5735 => x"2e",
          5736 => x"b7",
          5737 => x"05",
          5738 => x"bd",
          5739 => x"c0",
          5740 => x"a4",
          5741 => x"c7",
          5742 => x"53",
          5743 => x"52",
          5744 => x"52",
          5745 => x"85",
          5746 => x"90",
          5747 => x"d8",
          5748 => x"64",
          5749 => x"81",
          5750 => x"54",
          5751 => x"53",
          5752 => x"52",
          5753 => x"aa",
          5754 => x"a4",
          5755 => x"81",
          5756 => x"32",
          5757 => x"8a",
          5758 => x"2e",
          5759 => x"f1",
          5760 => x"c7",
          5761 => x"f5",
          5762 => x"97",
          5763 => x"0d",
          5764 => x"cb",
          5765 => x"a0",
          5766 => x"87",
          5767 => x"0c",
          5768 => x"c8",
          5769 => x"94",
          5770 => x"80",
          5771 => x"c0",
          5772 => x"8c",
          5773 => x"87",
          5774 => x"0c",
          5775 => x"81",
          5776 => x"9a",
          5777 => x"cb",
          5778 => x"e7",
          5779 => x"ed",
          5780 => x"c7",
          5781 => x"e4",
          5782 => x"c7",
          5783 => x"ee",
          5784 => x"a1",
          5785 => x"ed",
          5786 => x"51",
          5787 => x"ef",
          5788 => x"04",
          5789 => x"10",
          5790 => x"10",
          5791 => x"11",
          5792 => x"11",
          5793 => x"11",
          5794 => x"4d",
          5795 => x"4d",
          5796 => x"4d",
          5797 => x"4d",
          5798 => x"4d",
          5799 => x"4d",
          5800 => x"4d",
          5801 => x"4d",
          5802 => x"4d",
          5803 => x"4d",
          5804 => x"4d",
          5805 => x"4d",
          5806 => x"4d",
          5807 => x"4d",
          5808 => x"4d",
          5809 => x"4d",
          5810 => x"4d",
          5811 => x"4d",
          5812 => x"4d",
          5813 => x"4d",
          5814 => x"2f",
          5815 => x"25",
          5816 => x"64",
          5817 => x"3a",
          5818 => x"25",
          5819 => x"0a",
          5820 => x"43",
          5821 => x"6e",
          5822 => x"75",
          5823 => x"69",
          5824 => x"00",
          5825 => x"66",
          5826 => x"20",
          5827 => x"20",
          5828 => x"66",
          5829 => x"00",
          5830 => x"44",
          5831 => x"63",
          5832 => x"69",
          5833 => x"65",
          5834 => x"74",
          5835 => x"0a",
          5836 => x"20",
          5837 => x"53",
          5838 => x"52",
          5839 => x"28",
          5840 => x"72",
          5841 => x"30",
          5842 => x"20",
          5843 => x"65",
          5844 => x"38",
          5845 => x"0a",
          5846 => x"20",
          5847 => x"41",
          5848 => x"53",
          5849 => x"74",
          5850 => x"38",
          5851 => x"53",
          5852 => x"3d",
          5853 => x"58",
          5854 => x"00",
          5855 => x"20",
          5856 => x"4d",
          5857 => x"74",
          5858 => x"3d",
          5859 => x"58",
          5860 => x"69",
          5861 => x"25",
          5862 => x"29",
          5863 => x"00",
          5864 => x"20",
          5865 => x"43",
          5866 => x"00",
          5867 => x"20",
          5868 => x"32",
          5869 => x"00",
          5870 => x"20",
          5871 => x"49",
          5872 => x"00",
          5873 => x"20",
          5874 => x"20",
          5875 => x"64",
          5876 => x"65",
          5877 => x"65",
          5878 => x"30",
          5879 => x"2e",
          5880 => x"00",
          5881 => x"20",
          5882 => x"54",
          5883 => x"55",
          5884 => x"43",
          5885 => x"52",
          5886 => x"45",
          5887 => x"00",
          5888 => x"20",
          5889 => x"4d",
          5890 => x"20",
          5891 => x"6d",
          5892 => x"3d",
          5893 => x"58",
          5894 => x"00",
          5895 => x"64",
          5896 => x"73",
          5897 => x"0a",
          5898 => x"20",
          5899 => x"55",
          5900 => x"73",
          5901 => x"56",
          5902 => x"6f",
          5903 => x"64",
          5904 => x"73",
          5905 => x"20",
          5906 => x"58",
          5907 => x"00",
          5908 => x"20",
          5909 => x"55",
          5910 => x"6d",
          5911 => x"20",
          5912 => x"72",
          5913 => x"64",
          5914 => x"73",
          5915 => x"20",
          5916 => x"58",
          5917 => x"00",
          5918 => x"20",
          5919 => x"61",
          5920 => x"53",
          5921 => x"74",
          5922 => x"64",
          5923 => x"73",
          5924 => x"20",
          5925 => x"20",
          5926 => x"58",
          5927 => x"00",
          5928 => x"20",
          5929 => x"55",
          5930 => x"20",
          5931 => x"20",
          5932 => x"20",
          5933 => x"20",
          5934 => x"20",
          5935 => x"20",
          5936 => x"58",
          5937 => x"00",
          5938 => x"20",
          5939 => x"73",
          5940 => x"20",
          5941 => x"63",
          5942 => x"72",
          5943 => x"20",
          5944 => x"20",
          5945 => x"20",
          5946 => x"58",
          5947 => x"00",
          5948 => x"61",
          5949 => x"00",
          5950 => x"64",
          5951 => x"00",
          5952 => x"65",
          5953 => x"00",
          5954 => x"4f",
          5955 => x"4f",
          5956 => x"00",
          5957 => x"6b",
          5958 => x"6e",
          5959 => x"00",
          5960 => x"2b",
          5961 => x"3c",
          5962 => x"5b",
          5963 => x"00",
          5964 => x"54",
          5965 => x"54",
          5966 => x"00",
          5967 => x"90",
          5968 => x"4f",
          5969 => x"30",
          5970 => x"20",
          5971 => x"45",
          5972 => x"20",
          5973 => x"33",
          5974 => x"20",
          5975 => x"20",
          5976 => x"45",
          5977 => x"20",
          5978 => x"20",
          5979 => x"20",
          5980 => x"5d",
          5981 => x"00",
          5982 => x"00",
          5983 => x"00",
          5984 => x"45",
          5985 => x"8f",
          5986 => x"45",
          5987 => x"8e",
          5988 => x"92",
          5989 => x"55",
          5990 => x"9a",
          5991 => x"9e",
          5992 => x"4f",
          5993 => x"a6",
          5994 => x"aa",
          5995 => x"ae",
          5996 => x"b2",
          5997 => x"b6",
          5998 => x"ba",
          5999 => x"be",
          6000 => x"c2",
          6001 => x"c6",
          6002 => x"ca",
          6003 => x"ce",
          6004 => x"d2",
          6005 => x"d6",
          6006 => x"da",
          6007 => x"de",
          6008 => x"e2",
          6009 => x"e6",
          6010 => x"ea",
          6011 => x"ee",
          6012 => x"f2",
          6013 => x"f6",
          6014 => x"fa",
          6015 => x"fe",
          6016 => x"2c",
          6017 => x"5d",
          6018 => x"2a",
          6019 => x"3f",
          6020 => x"00",
          6021 => x"00",
          6022 => x"00",
          6023 => x"02",
          6024 => x"00",
          6025 => x"00",
          6026 => x"00",
          6027 => x"00",
          6028 => x"00",
          6029 => x"6e",
          6030 => x"00",
          6031 => x"6f",
          6032 => x"00",
          6033 => x"6e",
          6034 => x"00",
          6035 => x"6f",
          6036 => x"00",
          6037 => x"78",
          6038 => x"00",
          6039 => x"6c",
          6040 => x"00",
          6041 => x"75",
          6042 => x"00",
          6043 => x"65",
          6044 => x"00",
          6045 => x"62",
          6046 => x"68",
          6047 => x"77",
          6048 => x"64",
          6049 => x"65",
          6050 => x"64",
          6051 => x"65",
          6052 => x"6c",
          6053 => x"00",
          6054 => x"70",
          6055 => x"73",
          6056 => x"74",
          6057 => x"73",
          6058 => x"00",
          6059 => x"66",
          6060 => x"00",
          6061 => x"73",
          6062 => x"00",
          6063 => x"73",
          6064 => x"72",
          6065 => x"0a",
          6066 => x"74",
          6067 => x"61",
          6068 => x"72",
          6069 => x"2e",
          6070 => x"00",
          6071 => x"73",
          6072 => x"6f",
          6073 => x"65",
          6074 => x"2e",
          6075 => x"00",
          6076 => x"20",
          6077 => x"65",
          6078 => x"75",
          6079 => x"0a",
          6080 => x"20",
          6081 => x"68",
          6082 => x"75",
          6083 => x"0a",
          6084 => x"76",
          6085 => x"64",
          6086 => x"6c",
          6087 => x"6d",
          6088 => x"00",
          6089 => x"63",
          6090 => x"20",
          6091 => x"69",
          6092 => x"0a",
          6093 => x"6c",
          6094 => x"6c",
          6095 => x"64",
          6096 => x"78",
          6097 => x"73",
          6098 => x"00",
          6099 => x"6c",
          6100 => x"61",
          6101 => x"65",
          6102 => x"76",
          6103 => x"64",
          6104 => x"00",
          6105 => x"20",
          6106 => x"77",
          6107 => x"65",
          6108 => x"6f",
          6109 => x"74",
          6110 => x"0a",
          6111 => x"69",
          6112 => x"6e",
          6113 => x"65",
          6114 => x"73",
          6115 => x"76",
          6116 => x"64",
          6117 => x"00",
          6118 => x"73",
          6119 => x"6f",
          6120 => x"6e",
          6121 => x"65",
          6122 => x"00",
          6123 => x"20",
          6124 => x"70",
          6125 => x"62",
          6126 => x"66",
          6127 => x"73",
          6128 => x"65",
          6129 => x"6f",
          6130 => x"20",
          6131 => x"64",
          6132 => x"2e",
          6133 => x"00",
          6134 => x"72",
          6135 => x"20",
          6136 => x"72",
          6137 => x"2e",
          6138 => x"00",
          6139 => x"6d",
          6140 => x"74",
          6141 => x"70",
          6142 => x"74",
          6143 => x"20",
          6144 => x"63",
          6145 => x"65",
          6146 => x"00",
          6147 => x"6c",
          6148 => x"73",
          6149 => x"63",
          6150 => x"2e",
          6151 => x"00",
          6152 => x"73",
          6153 => x"69",
          6154 => x"6e",
          6155 => x"65",
          6156 => x"79",
          6157 => x"00",
          6158 => x"6f",
          6159 => x"6e",
          6160 => x"70",
          6161 => x"66",
          6162 => x"73",
          6163 => x"00",
          6164 => x"72",
          6165 => x"74",
          6166 => x"20",
          6167 => x"6f",
          6168 => x"63",
          6169 => x"00",
          6170 => x"63",
          6171 => x"73",
          6172 => x"00",
          6173 => x"6b",
          6174 => x"6e",
          6175 => x"72",
          6176 => x"0a",
          6177 => x"6c",
          6178 => x"79",
          6179 => x"20",
          6180 => x"61",
          6181 => x"6c",
          6182 => x"79",
          6183 => x"2f",
          6184 => x"2e",
          6185 => x"00",
          6186 => x"38",
          6187 => x"00",
          6188 => x"20",
          6189 => x"34",
          6190 => x"00",
          6191 => x"20",
          6192 => x"20",
          6193 => x"00",
          6194 => x"32",
          6195 => x"00",
          6196 => x"00",
          6197 => x"00",
          6198 => x"0a",
          6199 => x"61",
          6200 => x"00",
          6201 => x"55",
          6202 => x"00",
          6203 => x"2a",
          6204 => x"20",
          6205 => x"00",
          6206 => x"2f",
          6207 => x"32",
          6208 => x"00",
          6209 => x"2e",
          6210 => x"00",
          6211 => x"50",
          6212 => x"72",
          6213 => x"25",
          6214 => x"29",
          6215 => x"20",
          6216 => x"2a",
          6217 => x"00",
          6218 => x"55",
          6219 => x"49",
          6220 => x"72",
          6221 => x"74",
          6222 => x"6e",
          6223 => x"72",
          6224 => x"00",
          6225 => x"6d",
          6226 => x"69",
          6227 => x"72",
          6228 => x"74",
          6229 => x"00",
          6230 => x"32",
          6231 => x"74",
          6232 => x"75",
          6233 => x"00",
          6234 => x"43",
          6235 => x"52",
          6236 => x"6e",
          6237 => x"72",
          6238 => x"0a",
          6239 => x"43",
          6240 => x"57",
          6241 => x"6e",
          6242 => x"72",
          6243 => x"0a",
          6244 => x"52",
          6245 => x"52",
          6246 => x"6e",
          6247 => x"72",
          6248 => x"0a",
          6249 => x"52",
          6250 => x"54",
          6251 => x"6e",
          6252 => x"72",
          6253 => x"0a",
          6254 => x"52",
          6255 => x"52",
          6256 => x"6e",
          6257 => x"72",
          6258 => x"0a",
          6259 => x"52",
          6260 => x"54",
          6261 => x"6e",
          6262 => x"72",
          6263 => x"0a",
          6264 => x"74",
          6265 => x"67",
          6266 => x"20",
          6267 => x"65",
          6268 => x"2e",
          6269 => x"00",
          6270 => x"61",
          6271 => x"6e",
          6272 => x"69",
          6273 => x"2e",
          6274 => x"00",
          6275 => x"00",
          6276 => x"69",
          6277 => x"20",
          6278 => x"69",
          6279 => x"69",
          6280 => x"73",
          6281 => x"64",
          6282 => x"72",
          6283 => x"2c",
          6284 => x"65",
          6285 => x"20",
          6286 => x"74",
          6287 => x"6e",
          6288 => x"6c",
          6289 => x"00",
          6290 => x"00",
          6291 => x"64",
          6292 => x"73",
          6293 => x"64",
          6294 => x"00",
          6295 => x"69",
          6296 => x"6c",
          6297 => x"64",
          6298 => x"00",
          6299 => x"69",
          6300 => x"20",
          6301 => x"69",
          6302 => x"69",
          6303 => x"73",
          6304 => x"00",
          6305 => x"3d",
          6306 => x"00",
          6307 => x"3a",
          6308 => x"65",
          6309 => x"6e",
          6310 => x"2e",
          6311 => x"6d",
          6312 => x"65",
          6313 => x"79",
          6314 => x"00",
          6315 => x"6f",
          6316 => x"65",
          6317 => x"0a",
          6318 => x"38",
          6319 => x"30",
          6320 => x"00",
          6321 => x"3f",
          6322 => x"00",
          6323 => x"38",
          6324 => x"30",
          6325 => x"00",
          6326 => x"38",
          6327 => x"30",
          6328 => x"00",
          6329 => x"73",
          6330 => x"69",
          6331 => x"69",
          6332 => x"72",
          6333 => x"74",
          6334 => x"00",
          6335 => x"61",
          6336 => x"6e",
          6337 => x"6e",
          6338 => x"72",
          6339 => x"73",
          6340 => x"00",
          6341 => x"73",
          6342 => x"65",
          6343 => x"61",
          6344 => x"66",
          6345 => x"0a",
          6346 => x"61",
          6347 => x"6e",
          6348 => x"61",
          6349 => x"66",
          6350 => x"0a",
          6351 => x"65",
          6352 => x"69",
          6353 => x"63",
          6354 => x"20",
          6355 => x"30",
          6356 => x"2e",
          6357 => x"00",
          6358 => x"6c",
          6359 => x"67",
          6360 => x"64",
          6361 => x"20",
          6362 => x"78",
          6363 => x"2e",
          6364 => x"00",
          6365 => x"6c",
          6366 => x"65",
          6367 => x"6e",
          6368 => x"63",
          6369 => x"20",
          6370 => x"29",
          6371 => x"00",
          6372 => x"73",
          6373 => x"74",
          6374 => x"20",
          6375 => x"6c",
          6376 => x"74",
          6377 => x"2e",
          6378 => x"00",
          6379 => x"6c",
          6380 => x"65",
          6381 => x"74",
          6382 => x"2e",
          6383 => x"00",
          6384 => x"55",
          6385 => x"6e",
          6386 => x"3a",
          6387 => x"5c",
          6388 => x"25",
          6389 => x"00",
          6390 => x"64",
          6391 => x"6d",
          6392 => x"64",
          6393 => x"00",
          6394 => x"6e",
          6395 => x"67",
          6396 => x"0a",
          6397 => x"61",
          6398 => x"6e",
          6399 => x"6e",
          6400 => x"72",
          6401 => x"73",
          6402 => x"0a",
          6403 => x"00",
          6404 => x"00",
          6405 => x"7f",
          6406 => x"00",
          6407 => x"7f",
          6408 => x"00",
          6409 => x"7f",
          6410 => x"00",
          6411 => x"00",
          6412 => x"78",
          6413 => x"00",
          6414 => x"e1",
          6415 => x"01",
          6416 => x"01",
          6417 => x"01",
          6418 => x"00",
          6419 => x"00",
          6420 => x"00",
          6421 => x"5e",
          6422 => x"01",
          6423 => x"00",
          6424 => x"00",
          6425 => x"5e",
          6426 => x"01",
          6427 => x"00",
          6428 => x"00",
          6429 => x"5e",
          6430 => x"03",
          6431 => x"00",
          6432 => x"00",
          6433 => x"5e",
          6434 => x"03",
          6435 => x"00",
          6436 => x"00",
          6437 => x"5e",
          6438 => x"03",
          6439 => x"00",
          6440 => x"00",
          6441 => x"5e",
          6442 => x"04",
          6443 => x"00",
          6444 => x"00",
          6445 => x"5e",
          6446 => x"04",
          6447 => x"00",
          6448 => x"00",
          6449 => x"5e",
          6450 => x"04",
          6451 => x"00",
          6452 => x"00",
          6453 => x"5e",
          6454 => x"04",
          6455 => x"00",
          6456 => x"00",
          6457 => x"5e",
          6458 => x"04",
          6459 => x"00",
          6460 => x"00",
          6461 => x"5e",
          6462 => x"04",
          6463 => x"00",
          6464 => x"00",
          6465 => x"5e",
          6466 => x"05",
          6467 => x"00",
          6468 => x"00",
          6469 => x"5e",
          6470 => x"05",
          6471 => x"00",
          6472 => x"00",
          6473 => x"5e",
          6474 => x"05",
          6475 => x"00",
          6476 => x"00",
          6477 => x"5e",
          6478 => x"05",
          6479 => x"00",
          6480 => x"00",
          6481 => x"5e",
          6482 => x"07",
          6483 => x"00",
          6484 => x"00",
          6485 => x"5e",
          6486 => x"07",
          6487 => x"00",
          6488 => x"00",
          6489 => x"5e",
          6490 => x"08",
          6491 => x"00",
          6492 => x"00",
          6493 => x"5e",
          6494 => x"08",
          6495 => x"00",
          6496 => x"00",
          6497 => x"5e",
          6498 => x"08",
          6499 => x"00",
          6500 => x"00",
          6501 => x"5e",
          6502 => x"08",
          6503 => x"00",
          6504 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"8d",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"04",
            10 => x"88",
            11 => x"0b",
            12 => x"04",
            13 => x"88",
            14 => x"0b",
            15 => x"04",
            16 => x"88",
            17 => x"0b",
            18 => x"04",
            19 => x"88",
            20 => x"0b",
            21 => x"04",
            22 => x"88",
            23 => x"0b",
            24 => x"04",
            25 => x"89",
            26 => x"0b",
            27 => x"04",
            28 => x"89",
            29 => x"0b",
            30 => x"04",
            31 => x"89",
            32 => x"0b",
            33 => x"04",
            34 => x"89",
            35 => x"0b",
            36 => x"04",
            37 => x"8a",
            38 => x"0b",
            39 => x"04",
            40 => x"8a",
            41 => x"0b",
            42 => x"04",
            43 => x"8a",
            44 => x"0b",
            45 => x"04",
            46 => x"8a",
            47 => x"0b",
            48 => x"04",
            49 => x"8b",
            50 => x"0b",
            51 => x"04",
            52 => x"8b",
            53 => x"0b",
            54 => x"04",
            55 => x"8b",
            56 => x"0b",
            57 => x"04",
            58 => x"8b",
            59 => x"0b",
            60 => x"04",
            61 => x"8c",
            62 => x"0b",
            63 => x"04",
            64 => x"8c",
            65 => x"0b",
            66 => x"04",
            67 => x"8c",
            68 => x"0b",
            69 => x"04",
            70 => x"8c",
            71 => x"0b",
            72 => x"04",
            73 => x"8d",
            74 => x"0b",
            75 => x"04",
            76 => x"8d",
            77 => x"0b",
            78 => x"04",
            79 => x"8d",
            80 => x"0b",
            81 => x"04",
            82 => x"8d",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"00",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"00",
           137 => x"00",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"00",
           145 => x"00",
           146 => x"00",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"00",
           153 => x"00",
           154 => x"00",
           155 => x"00",
           156 => x"00",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"00",
           161 => x"00",
           162 => x"00",
           163 => x"00",
           164 => x"00",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"00",
           169 => x"00",
           170 => x"00",
           171 => x"00",
           172 => x"00",
           173 => x"00",
           174 => x"00",
           175 => x"00",
           176 => x"00",
           177 => x"00",
           178 => x"00",
           179 => x"00",
           180 => x"00",
           181 => x"00",
           182 => x"00",
           183 => x"00",
           184 => x"00",
           185 => x"00",
           186 => x"00",
           187 => x"00",
           188 => x"00",
           189 => x"00",
           190 => x"00",
           191 => x"00",
           192 => x"00",
           193 => x"00",
           194 => x"00",
           195 => x"00",
           196 => x"00",
           197 => x"00",
           198 => x"00",
           199 => x"00",
           200 => x"00",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"00",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"00",
           233 => x"00",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"00",
           249 => x"00",
           250 => x"00",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"88",
           257 => x"cb",
           258 => x"c5",
           259 => x"b0",
           260 => x"90",
           261 => x"b0",
           262 => x"2d",
           263 => x"08",
           264 => x"04",
           265 => x"0c",
           266 => x"81",
           267 => x"81",
           268 => x"81",
           269 => x"a3",
           270 => x"cb",
           271 => x"e4",
           272 => x"cb",
           273 => x"90",
           274 => x"b0",
           275 => x"90",
           276 => x"b0",
           277 => x"2d",
           278 => x"08",
           279 => x"04",
           280 => x"0c",
           281 => x"81",
           282 => x"81",
           283 => x"81",
           284 => x"ab",
           285 => x"cb",
           286 => x"e4",
           287 => x"cb",
           288 => x"9d",
           289 => x"b0",
           290 => x"90",
           291 => x"b0",
           292 => x"2d",
           293 => x"08",
           294 => x"04",
           295 => x"0c",
           296 => x"81",
           297 => x"81",
           298 => x"81",
           299 => x"a9",
           300 => x"cb",
           301 => x"e4",
           302 => x"cb",
           303 => x"d2",
           304 => x"b0",
           305 => x"90",
           306 => x"b0",
           307 => x"2d",
           308 => x"08",
           309 => x"04",
           310 => x"0c",
           311 => x"81",
           312 => x"81",
           313 => x"81",
           314 => x"94",
           315 => x"cb",
           316 => x"e4",
           317 => x"cb",
           318 => x"a7",
           319 => x"b0",
           320 => x"90",
           321 => x"b0",
           322 => x"d2",
           323 => x"b0",
           324 => x"90",
           325 => x"b0",
           326 => x"c3",
           327 => x"b0",
           328 => x"90",
           329 => x"b0",
           330 => x"b7",
           331 => x"b0",
           332 => x"90",
           333 => x"b0",
           334 => x"b4",
           335 => x"b0",
           336 => x"90",
           337 => x"b0",
           338 => x"d2",
           339 => x"b0",
           340 => x"90",
           341 => x"b0",
           342 => x"b2",
           343 => x"b0",
           344 => x"90",
           345 => x"b0",
           346 => x"a5",
           347 => x"b0",
           348 => x"90",
           349 => x"b0",
           350 => x"f1",
           351 => x"b0",
           352 => x"90",
           353 => x"b0",
           354 => x"90",
           355 => x"b0",
           356 => x"90",
           357 => x"b0",
           358 => x"af",
           359 => x"b0",
           360 => x"90",
           361 => x"b0",
           362 => x"99",
           363 => x"b0",
           364 => x"90",
           365 => x"b0",
           366 => x"ff",
           367 => x"b0",
           368 => x"90",
           369 => x"b0",
           370 => x"ed",
           371 => x"b0",
           372 => x"90",
           373 => x"b0",
           374 => x"b3",
           375 => x"b0",
           376 => x"90",
           377 => x"b0",
           378 => x"ed",
           379 => x"b0",
           380 => x"90",
           381 => x"b0",
           382 => x"ee",
           383 => x"b0",
           384 => x"90",
           385 => x"b0",
           386 => x"a3",
           387 => x"b0",
           388 => x"90",
           389 => x"b0",
           390 => x"fc",
           391 => x"b0",
           392 => x"90",
           393 => x"b0",
           394 => x"a7",
           395 => x"b0",
           396 => x"90",
           397 => x"b0",
           398 => x"8a",
           399 => x"b0",
           400 => x"90",
           401 => x"b0",
           402 => x"df",
           403 => x"b0",
           404 => x"90",
           405 => x"b0",
           406 => x"e9",
           407 => x"b0",
           408 => x"90",
           409 => x"b0",
           410 => x"ab",
           411 => x"b0",
           412 => x"90",
           413 => x"b0",
           414 => x"f1",
           415 => x"b0",
           416 => x"90",
           417 => x"b0",
           418 => x"97",
           419 => x"b0",
           420 => x"90",
           421 => x"b0",
           422 => x"2d",
           423 => x"08",
           424 => x"04",
           425 => x"0c",
           426 => x"81",
           427 => x"81",
           428 => x"81",
           429 => x"b3",
           430 => x"cb",
           431 => x"e4",
           432 => x"cb",
           433 => x"e8",
           434 => x"b0",
           435 => x"90",
           436 => x"b0",
           437 => x"2d",
           438 => x"08",
           439 => x"04",
           440 => x"0c",
           441 => x"81",
           442 => x"81",
           443 => x"81",
           444 => x"81",
           445 => x"81",
           446 => x"81",
           447 => x"81",
           448 => x"81",
           449 => x"8e",
           450 => x"70",
           451 => x"0c",
           452 => x"8e",
           453 => x"80",
           454 => x"8c",
           455 => x"81",
           456 => x"02",
           457 => x"0c",
           458 => x"80",
           459 => x"b0",
           460 => x"08",
           461 => x"b0",
           462 => x"08",
           463 => x"3f",
           464 => x"08",
           465 => x"a4",
           466 => x"3d",
           467 => x"b0",
           468 => x"cb",
           469 => x"81",
           470 => x"fd",
           471 => x"53",
           472 => x"08",
           473 => x"52",
           474 => x"08",
           475 => x"51",
           476 => x"cb",
           477 => x"81",
           478 => x"54",
           479 => x"81",
           480 => x"04",
           481 => x"08",
           482 => x"b0",
           483 => x"0d",
           484 => x"cb",
           485 => x"05",
           486 => x"81",
           487 => x"f8",
           488 => x"cb",
           489 => x"05",
           490 => x"b0",
           491 => x"08",
           492 => x"81",
           493 => x"fc",
           494 => x"2e",
           495 => x"0b",
           496 => x"08",
           497 => x"24",
           498 => x"cb",
           499 => x"05",
           500 => x"cb",
           501 => x"05",
           502 => x"b0",
           503 => x"08",
           504 => x"b0",
           505 => x"0c",
           506 => x"81",
           507 => x"fc",
           508 => x"2e",
           509 => x"81",
           510 => x"8c",
           511 => x"cb",
           512 => x"05",
           513 => x"38",
           514 => x"08",
           515 => x"81",
           516 => x"8c",
           517 => x"81",
           518 => x"88",
           519 => x"cb",
           520 => x"05",
           521 => x"b0",
           522 => x"08",
           523 => x"b0",
           524 => x"0c",
           525 => x"08",
           526 => x"81",
           527 => x"b0",
           528 => x"0c",
           529 => x"08",
           530 => x"81",
           531 => x"b0",
           532 => x"0c",
           533 => x"81",
           534 => x"90",
           535 => x"2e",
           536 => x"cb",
           537 => x"05",
           538 => x"cb",
           539 => x"05",
           540 => x"39",
           541 => x"08",
           542 => x"70",
           543 => x"08",
           544 => x"51",
           545 => x"08",
           546 => x"81",
           547 => x"85",
           548 => x"cb",
           549 => x"fc",
           550 => x"79",
           551 => x"05",
           552 => x"57",
           553 => x"83",
           554 => x"38",
           555 => x"51",
           556 => x"a4",
           557 => x"52",
           558 => x"93",
           559 => x"70",
           560 => x"34",
           561 => x"71",
           562 => x"81",
           563 => x"74",
           564 => x"0c",
           565 => x"04",
           566 => x"2b",
           567 => x"71",
           568 => x"51",
           569 => x"72",
           570 => x"72",
           571 => x"05",
           572 => x"71",
           573 => x"53",
           574 => x"70",
           575 => x"0c",
           576 => x"84",
           577 => x"f0",
           578 => x"8f",
           579 => x"83",
           580 => x"38",
           581 => x"84",
           582 => x"fc",
           583 => x"83",
           584 => x"70",
           585 => x"39",
           586 => x"77",
           587 => x"07",
           588 => x"54",
           589 => x"38",
           590 => x"08",
           591 => x"71",
           592 => x"80",
           593 => x"75",
           594 => x"33",
           595 => x"06",
           596 => x"80",
           597 => x"72",
           598 => x"75",
           599 => x"06",
           600 => x"12",
           601 => x"33",
           602 => x"06",
           603 => x"52",
           604 => x"72",
           605 => x"81",
           606 => x"81",
           607 => x"71",
           608 => x"a4",
           609 => x"87",
           610 => x"71",
           611 => x"fb",
           612 => x"06",
           613 => x"82",
           614 => x"51",
           615 => x"97",
           616 => x"84",
           617 => x"54",
           618 => x"75",
           619 => x"38",
           620 => x"52",
           621 => x"80",
           622 => x"a4",
           623 => x"0d",
           624 => x"0d",
           625 => x"53",
           626 => x"52",
           627 => x"81",
           628 => x"81",
           629 => x"07",
           630 => x"52",
           631 => x"e8",
           632 => x"cb",
           633 => x"3d",
           634 => x"3d",
           635 => x"08",
           636 => x"56",
           637 => x"80",
           638 => x"33",
           639 => x"2e",
           640 => x"86",
           641 => x"52",
           642 => x"53",
           643 => x"13",
           644 => x"33",
           645 => x"06",
           646 => x"70",
           647 => x"38",
           648 => x"80",
           649 => x"74",
           650 => x"81",
           651 => x"70",
           652 => x"81",
           653 => x"80",
           654 => x"05",
           655 => x"76",
           656 => x"70",
           657 => x"0c",
           658 => x"04",
           659 => x"76",
           660 => x"80",
           661 => x"86",
           662 => x"52",
           663 => x"bf",
           664 => x"a4",
           665 => x"80",
           666 => x"74",
           667 => x"cb",
           668 => x"3d",
           669 => x"3d",
           670 => x"11",
           671 => x"52",
           672 => x"70",
           673 => x"98",
           674 => x"33",
           675 => x"82",
           676 => x"26",
           677 => x"84",
           678 => x"83",
           679 => x"26",
           680 => x"85",
           681 => x"84",
           682 => x"26",
           683 => x"86",
           684 => x"85",
           685 => x"26",
           686 => x"88",
           687 => x"86",
           688 => x"e7",
           689 => x"38",
           690 => x"54",
           691 => x"87",
           692 => x"cc",
           693 => x"87",
           694 => x"0c",
           695 => x"c0",
           696 => x"82",
           697 => x"c0",
           698 => x"83",
           699 => x"c0",
           700 => x"84",
           701 => x"c0",
           702 => x"85",
           703 => x"c0",
           704 => x"86",
           705 => x"c0",
           706 => x"74",
           707 => x"a4",
           708 => x"c0",
           709 => x"80",
           710 => x"98",
           711 => x"52",
           712 => x"a4",
           713 => x"0d",
           714 => x"0d",
           715 => x"c0",
           716 => x"81",
           717 => x"c0",
           718 => x"5e",
           719 => x"87",
           720 => x"08",
           721 => x"1c",
           722 => x"98",
           723 => x"79",
           724 => x"87",
           725 => x"08",
           726 => x"1c",
           727 => x"98",
           728 => x"79",
           729 => x"87",
           730 => x"08",
           731 => x"1c",
           732 => x"98",
           733 => x"7b",
           734 => x"87",
           735 => x"08",
           736 => x"1c",
           737 => x"0c",
           738 => x"ff",
           739 => x"83",
           740 => x"58",
           741 => x"57",
           742 => x"56",
           743 => x"55",
           744 => x"54",
           745 => x"53",
           746 => x"ff",
           747 => x"b5",
           748 => x"84",
           749 => x"0d",
           750 => x"0d",
           751 => x"33",
           752 => x"9f",
           753 => x"52",
           754 => x"81",
           755 => x"83",
           756 => x"fb",
           757 => x"0b",
           758 => x"8c",
           759 => x"ff",
           760 => x"56",
           761 => x"84",
           762 => x"2e",
           763 => x"c0",
           764 => x"70",
           765 => x"2a",
           766 => x"53",
           767 => x"80",
           768 => x"71",
           769 => x"81",
           770 => x"70",
           771 => x"81",
           772 => x"06",
           773 => x"80",
           774 => x"71",
           775 => x"81",
           776 => x"70",
           777 => x"73",
           778 => x"51",
           779 => x"80",
           780 => x"2e",
           781 => x"c0",
           782 => x"75",
           783 => x"81",
           784 => x"87",
           785 => x"fb",
           786 => x"9f",
           787 => x"0b",
           788 => x"33",
           789 => x"06",
           790 => x"87",
           791 => x"51",
           792 => x"86",
           793 => x"94",
           794 => x"08",
           795 => x"70",
           796 => x"54",
           797 => x"2e",
           798 => x"91",
           799 => x"06",
           800 => x"d7",
           801 => x"32",
           802 => x"51",
           803 => x"2e",
           804 => x"93",
           805 => x"06",
           806 => x"ff",
           807 => x"81",
           808 => x"87",
           809 => x"52",
           810 => x"86",
           811 => x"94",
           812 => x"72",
           813 => x"0d",
           814 => x"0d",
           815 => x"74",
           816 => x"ff",
           817 => x"57",
           818 => x"80",
           819 => x"81",
           820 => x"15",
           821 => x"c8",
           822 => x"81",
           823 => x"57",
           824 => x"c0",
           825 => x"75",
           826 => x"38",
           827 => x"94",
           828 => x"70",
           829 => x"81",
           830 => x"52",
           831 => x"8c",
           832 => x"2a",
           833 => x"51",
           834 => x"38",
           835 => x"70",
           836 => x"51",
           837 => x"8d",
           838 => x"2a",
           839 => x"51",
           840 => x"be",
           841 => x"ff",
           842 => x"c0",
           843 => x"70",
           844 => x"38",
           845 => x"90",
           846 => x"0c",
           847 => x"33",
           848 => x"06",
           849 => x"70",
           850 => x"76",
           851 => x"0c",
           852 => x"04",
           853 => x"0b",
           854 => x"8c",
           855 => x"ff",
           856 => x"87",
           857 => x"51",
           858 => x"86",
           859 => x"94",
           860 => x"08",
           861 => x"70",
           862 => x"51",
           863 => x"2e",
           864 => x"81",
           865 => x"87",
           866 => x"52",
           867 => x"86",
           868 => x"94",
           869 => x"08",
           870 => x"06",
           871 => x"0c",
           872 => x"0d",
           873 => x"0d",
           874 => x"c8",
           875 => x"81",
           876 => x"53",
           877 => x"84",
           878 => x"2e",
           879 => x"c0",
           880 => x"71",
           881 => x"2a",
           882 => x"51",
           883 => x"52",
           884 => x"a0",
           885 => x"ff",
           886 => x"c0",
           887 => x"70",
           888 => x"38",
           889 => x"90",
           890 => x"70",
           891 => x"98",
           892 => x"51",
           893 => x"a4",
           894 => x"0d",
           895 => x"0d",
           896 => x"80",
           897 => x"2a",
           898 => x"51",
           899 => x"83",
           900 => x"c0",
           901 => x"81",
           902 => x"87",
           903 => x"08",
           904 => x"0c",
           905 => x"8c",
           906 => x"98",
           907 => x"9e",
           908 => x"c8",
           909 => x"c0",
           910 => x"81",
           911 => x"87",
           912 => x"08",
           913 => x"0c",
           914 => x"a4",
           915 => x"a8",
           916 => x"9e",
           917 => x"c8",
           918 => x"c0",
           919 => x"81",
           920 => x"87",
           921 => x"08",
           922 => x"c8",
           923 => x"c0",
           924 => x"81",
           925 => x"81",
           926 => x"bc",
           927 => x"87",
           928 => x"08",
           929 => x"06",
           930 => x"70",
           931 => x"38",
           932 => x"81",
           933 => x"80",
           934 => x"9e",
           935 => x"81",
           936 => x"51",
           937 => x"80",
           938 => x"81",
           939 => x"c8",
           940 => x"0b",
           941 => x"88",
           942 => x"c0",
           943 => x"52",
           944 => x"2e",
           945 => x"52",
           946 => x"bf",
           947 => x"87",
           948 => x"08",
           949 => x"06",
           950 => x"70",
           951 => x"38",
           952 => x"81",
           953 => x"80",
           954 => x"9e",
           955 => x"88",
           956 => x"52",
           957 => x"2e",
           958 => x"52",
           959 => x"c1",
           960 => x"87",
           961 => x"08",
           962 => x"06",
           963 => x"70",
           964 => x"38",
           965 => x"81",
           966 => x"80",
           967 => x"9e",
           968 => x"82",
           969 => x"52",
           970 => x"2e",
           971 => x"52",
           972 => x"c3",
           973 => x"87",
           974 => x"08",
           975 => x"06",
           976 => x"70",
           977 => x"38",
           978 => x"81",
           979 => x"87",
           980 => x"08",
           981 => x"06",
           982 => x"51",
           983 => x"81",
           984 => x"80",
           985 => x"9e",
           986 => x"90",
           987 => x"52",
           988 => x"83",
           989 => x"71",
           990 => x"34",
           991 => x"c0",
           992 => x"70",
           993 => x"52",
           994 => x"2e",
           995 => x"52",
           996 => x"c7",
           997 => x"9e",
           998 => x"87",
           999 => x"70",
          1000 => x"34",
          1001 => x"04",
          1002 => x"81",
          1003 => x"84",
          1004 => x"c8",
          1005 => x"73",
          1006 => x"38",
          1007 => x"51",
          1008 => x"81",
          1009 => x"84",
          1010 => x"c8",
          1011 => x"73",
          1012 => x"38",
          1013 => x"08",
          1014 => x"90",
          1015 => x"b6",
          1016 => x"d4",
          1017 => x"be",
          1018 => x"80",
          1019 => x"81",
          1020 => x"53",
          1021 => x"08",
          1022 => x"d8",
          1023 => x"3f",
          1024 => x"33",
          1025 => x"38",
          1026 => x"33",
          1027 => x"2e",
          1028 => x"c8",
          1029 => x"81",
          1030 => x"52",
          1031 => x"51",
          1032 => x"81",
          1033 => x"54",
          1034 => x"88",
          1035 => x"a0",
          1036 => x"3f",
          1037 => x"33",
          1038 => x"2e",
          1039 => x"b7",
          1040 => x"90",
          1041 => x"c3",
          1042 => x"80",
          1043 => x"81",
          1044 => x"82",
          1045 => x"c8",
          1046 => x"73",
          1047 => x"38",
          1048 => x"33",
          1049 => x"c4",
          1050 => x"3f",
          1051 => x"33",
          1052 => x"2e",
          1053 => x"b7",
          1054 => x"d8",
          1055 => x"c7",
          1056 => x"80",
          1057 => x"81",
          1058 => x"52",
          1059 => x"51",
          1060 => x"81",
          1061 => x"82",
          1062 => x"c8",
          1063 => x"81",
          1064 => x"88",
          1065 => x"c8",
          1066 => x"81",
          1067 => x"88",
          1068 => x"c8",
          1069 => x"81",
          1070 => x"87",
          1071 => x"c8",
          1072 => x"81",
          1073 => x"87",
          1074 => x"c8",
          1075 => x"81",
          1076 => x"87",
          1077 => x"3d",
          1078 => x"3d",
          1079 => x"05",
          1080 => x"52",
          1081 => x"ac",
          1082 => x"29",
          1083 => x"b4",
          1084 => x"71",
          1085 => x"b9",
          1086 => x"39",
          1087 => x"51",
          1088 => x"ba",
          1089 => x"39",
          1090 => x"51",
          1091 => x"ba",
          1092 => x"39",
          1093 => x"51",
          1094 => x"84",
          1095 => x"71",
          1096 => x"04",
          1097 => x"c0",
          1098 => x"04",
          1099 => x"87",
          1100 => x"70",
          1101 => x"80",
          1102 => x"74",
          1103 => x"c8",
          1104 => x"0c",
          1105 => x"04",
          1106 => x"87",
          1107 => x"70",
          1108 => x"cc",
          1109 => x"72",
          1110 => x"70",
          1111 => x"08",
          1112 => x"c8",
          1113 => x"0c",
          1114 => x"0d",
          1115 => x"cc",
          1116 => x"96",
          1117 => x"fe",
          1118 => x"93",
          1119 => x"72",
          1120 => x"81",
          1121 => x"8d",
          1122 => x"81",
          1123 => x"52",
          1124 => x"90",
          1125 => x"34",
          1126 => x"08",
          1127 => x"cb",
          1128 => x"39",
          1129 => x"08",
          1130 => x"2e",
          1131 => x"51",
          1132 => x"3d",
          1133 => x"3d",
          1134 => x"05",
          1135 => x"b4",
          1136 => x"cb",
          1137 => x"51",
          1138 => x"72",
          1139 => x"0c",
          1140 => x"04",
          1141 => x"75",
          1142 => x"70",
          1143 => x"53",
          1144 => x"2e",
          1145 => x"81",
          1146 => x"81",
          1147 => x"87",
          1148 => x"85",
          1149 => x"fc",
          1150 => x"81",
          1151 => x"78",
          1152 => x"0c",
          1153 => x"33",
          1154 => x"06",
          1155 => x"80",
          1156 => x"72",
          1157 => x"51",
          1158 => x"fe",
          1159 => x"39",
          1160 => x"b4",
          1161 => x"0d",
          1162 => x"0d",
          1163 => x"59",
          1164 => x"05",
          1165 => x"75",
          1166 => x"f8",
          1167 => x"2e",
          1168 => x"82",
          1169 => x"70",
          1170 => x"05",
          1171 => x"5b",
          1172 => x"2e",
          1173 => x"85",
          1174 => x"8b",
          1175 => x"2e",
          1176 => x"8a",
          1177 => x"78",
          1178 => x"5a",
          1179 => x"aa",
          1180 => x"06",
          1181 => x"84",
          1182 => x"7b",
          1183 => x"5d",
          1184 => x"59",
          1185 => x"d0",
          1186 => x"89",
          1187 => x"7a",
          1188 => x"10",
          1189 => x"d0",
          1190 => x"81",
          1191 => x"57",
          1192 => x"75",
          1193 => x"70",
          1194 => x"07",
          1195 => x"80",
          1196 => x"30",
          1197 => x"80",
          1198 => x"53",
          1199 => x"55",
          1200 => x"2e",
          1201 => x"84",
          1202 => x"81",
          1203 => x"57",
          1204 => x"2e",
          1205 => x"75",
          1206 => x"76",
          1207 => x"e0",
          1208 => x"ff",
          1209 => x"73",
          1210 => x"81",
          1211 => x"80",
          1212 => x"38",
          1213 => x"2e",
          1214 => x"73",
          1215 => x"8b",
          1216 => x"c2",
          1217 => x"38",
          1218 => x"73",
          1219 => x"81",
          1220 => x"8f",
          1221 => x"d5",
          1222 => x"38",
          1223 => x"24",
          1224 => x"80",
          1225 => x"38",
          1226 => x"73",
          1227 => x"80",
          1228 => x"ef",
          1229 => x"19",
          1230 => x"59",
          1231 => x"33",
          1232 => x"75",
          1233 => x"81",
          1234 => x"70",
          1235 => x"55",
          1236 => x"79",
          1237 => x"90",
          1238 => x"16",
          1239 => x"7b",
          1240 => x"a0",
          1241 => x"3f",
          1242 => x"53",
          1243 => x"e9",
          1244 => x"fc",
          1245 => x"81",
          1246 => x"72",
          1247 => x"b0",
          1248 => x"fb",
          1249 => x"39",
          1250 => x"83",
          1251 => x"59",
          1252 => x"82",
          1253 => x"88",
          1254 => x"8a",
          1255 => x"90",
          1256 => x"75",
          1257 => x"3f",
          1258 => x"79",
          1259 => x"81",
          1260 => x"72",
          1261 => x"38",
          1262 => x"59",
          1263 => x"84",
          1264 => x"58",
          1265 => x"80",
          1266 => x"30",
          1267 => x"80",
          1268 => x"55",
          1269 => x"25",
          1270 => x"80",
          1271 => x"74",
          1272 => x"07",
          1273 => x"0b",
          1274 => x"57",
          1275 => x"51",
          1276 => x"81",
          1277 => x"81",
          1278 => x"53",
          1279 => x"e6",
          1280 => x"cb",
          1281 => x"89",
          1282 => x"38",
          1283 => x"75",
          1284 => x"84",
          1285 => x"53",
          1286 => x"06",
          1287 => x"53",
          1288 => x"81",
          1289 => x"81",
          1290 => x"70",
          1291 => x"2a",
          1292 => x"76",
          1293 => x"38",
          1294 => x"38",
          1295 => x"70",
          1296 => x"53",
          1297 => x"8e",
          1298 => x"77",
          1299 => x"53",
          1300 => x"81",
          1301 => x"7a",
          1302 => x"55",
          1303 => x"83",
          1304 => x"79",
          1305 => x"81",
          1306 => x"72",
          1307 => x"17",
          1308 => x"27",
          1309 => x"51",
          1310 => x"75",
          1311 => x"72",
          1312 => x"81",
          1313 => x"7a",
          1314 => x"38",
          1315 => x"05",
          1316 => x"ff",
          1317 => x"70",
          1318 => x"57",
          1319 => x"76",
          1320 => x"81",
          1321 => x"72",
          1322 => x"84",
          1323 => x"f9",
          1324 => x"39",
          1325 => x"04",
          1326 => x"86",
          1327 => x"84",
          1328 => x"55",
          1329 => x"fa",
          1330 => x"3d",
          1331 => x"3d",
          1332 => x"cb",
          1333 => x"3d",
          1334 => x"75",
          1335 => x"3f",
          1336 => x"08",
          1337 => x"34",
          1338 => x"cb",
          1339 => x"3d",
          1340 => x"3d",
          1341 => x"b4",
          1342 => x"cb",
          1343 => x"3d",
          1344 => x"77",
          1345 => x"a1",
          1346 => x"cb",
          1347 => x"3d",
          1348 => x"3d",
          1349 => x"81",
          1350 => x"70",
          1351 => x"55",
          1352 => x"80",
          1353 => x"38",
          1354 => x"08",
          1355 => x"81",
          1356 => x"81",
          1357 => x"72",
          1358 => x"cb",
          1359 => x"2e",
          1360 => x"88",
          1361 => x"70",
          1362 => x"51",
          1363 => x"2e",
          1364 => x"80",
          1365 => x"ff",
          1366 => x"39",
          1367 => x"c8",
          1368 => x"52",
          1369 => x"c0",
          1370 => x"52",
          1371 => x"81",
          1372 => x"51",
          1373 => x"ff",
          1374 => x"15",
          1375 => x"34",
          1376 => x"f3",
          1377 => x"72",
          1378 => x"0c",
          1379 => x"04",
          1380 => x"81",
          1381 => x"75",
          1382 => x"0c",
          1383 => x"52",
          1384 => x"3f",
          1385 => x"b8",
          1386 => x"0d",
          1387 => x"0d",
          1388 => x"56",
          1389 => x"0c",
          1390 => x"70",
          1391 => x"73",
          1392 => x"81",
          1393 => x"81",
          1394 => x"ed",
          1395 => x"2e",
          1396 => x"8e",
          1397 => x"08",
          1398 => x"76",
          1399 => x"56",
          1400 => x"b0",
          1401 => x"06",
          1402 => x"75",
          1403 => x"76",
          1404 => x"70",
          1405 => x"73",
          1406 => x"8b",
          1407 => x"73",
          1408 => x"85",
          1409 => x"82",
          1410 => x"76",
          1411 => x"70",
          1412 => x"ac",
          1413 => x"a0",
          1414 => x"fa",
          1415 => x"53",
          1416 => x"57",
          1417 => x"98",
          1418 => x"39",
          1419 => x"80",
          1420 => x"26",
          1421 => x"86",
          1422 => x"80",
          1423 => x"57",
          1424 => x"74",
          1425 => x"38",
          1426 => x"27",
          1427 => x"14",
          1428 => x"06",
          1429 => x"14",
          1430 => x"06",
          1431 => x"74",
          1432 => x"f9",
          1433 => x"ff",
          1434 => x"89",
          1435 => x"38",
          1436 => x"c5",
          1437 => x"29",
          1438 => x"81",
          1439 => x"76",
          1440 => x"56",
          1441 => x"ba",
          1442 => x"2e",
          1443 => x"30",
          1444 => x"0c",
          1445 => x"81",
          1446 => x"8a",
          1447 => x"f8",
          1448 => x"7c",
          1449 => x"70",
          1450 => x"75",
          1451 => x"55",
          1452 => x"2e",
          1453 => x"87",
          1454 => x"76",
          1455 => x"73",
          1456 => x"81",
          1457 => x"81",
          1458 => x"77",
          1459 => x"70",
          1460 => x"58",
          1461 => x"09",
          1462 => x"c2",
          1463 => x"81",
          1464 => x"75",
          1465 => x"55",
          1466 => x"e2",
          1467 => x"90",
          1468 => x"f8",
          1469 => x"8f",
          1470 => x"81",
          1471 => x"75",
          1472 => x"55",
          1473 => x"81",
          1474 => x"27",
          1475 => x"d0",
          1476 => x"55",
          1477 => x"73",
          1478 => x"80",
          1479 => x"14",
          1480 => x"72",
          1481 => x"e0",
          1482 => x"80",
          1483 => x"39",
          1484 => x"55",
          1485 => x"80",
          1486 => x"e0",
          1487 => x"38",
          1488 => x"81",
          1489 => x"53",
          1490 => x"81",
          1491 => x"53",
          1492 => x"8e",
          1493 => x"70",
          1494 => x"55",
          1495 => x"27",
          1496 => x"77",
          1497 => x"74",
          1498 => x"76",
          1499 => x"77",
          1500 => x"70",
          1501 => x"55",
          1502 => x"77",
          1503 => x"38",
          1504 => x"74",
          1505 => x"55",
          1506 => x"a4",
          1507 => x"0d",
          1508 => x"0d",
          1509 => x"33",
          1510 => x"70",
          1511 => x"38",
          1512 => x"11",
          1513 => x"81",
          1514 => x"83",
          1515 => x"fc",
          1516 => x"9b",
          1517 => x"84",
          1518 => x"33",
          1519 => x"51",
          1520 => x"80",
          1521 => x"84",
          1522 => x"92",
          1523 => x"51",
          1524 => x"80",
          1525 => x"81",
          1526 => x"72",
          1527 => x"92",
          1528 => x"81",
          1529 => x"0b",
          1530 => x"8c",
          1531 => x"71",
          1532 => x"06",
          1533 => x"80",
          1534 => x"87",
          1535 => x"08",
          1536 => x"38",
          1537 => x"80",
          1538 => x"71",
          1539 => x"c0",
          1540 => x"51",
          1541 => x"87",
          1542 => x"c8",
          1543 => x"81",
          1544 => x"33",
          1545 => x"cb",
          1546 => x"3d",
          1547 => x"3d",
          1548 => x"64",
          1549 => x"bf",
          1550 => x"40",
          1551 => x"74",
          1552 => x"cd",
          1553 => x"a4",
          1554 => x"7a",
          1555 => x"81",
          1556 => x"72",
          1557 => x"87",
          1558 => x"11",
          1559 => x"8c",
          1560 => x"92",
          1561 => x"5a",
          1562 => x"58",
          1563 => x"c0",
          1564 => x"76",
          1565 => x"76",
          1566 => x"70",
          1567 => x"81",
          1568 => x"54",
          1569 => x"8e",
          1570 => x"52",
          1571 => x"81",
          1572 => x"81",
          1573 => x"74",
          1574 => x"53",
          1575 => x"83",
          1576 => x"78",
          1577 => x"8f",
          1578 => x"2e",
          1579 => x"c0",
          1580 => x"52",
          1581 => x"87",
          1582 => x"08",
          1583 => x"2e",
          1584 => x"84",
          1585 => x"38",
          1586 => x"87",
          1587 => x"15",
          1588 => x"70",
          1589 => x"52",
          1590 => x"ff",
          1591 => x"39",
          1592 => x"81",
          1593 => x"ff",
          1594 => x"57",
          1595 => x"90",
          1596 => x"80",
          1597 => x"71",
          1598 => x"78",
          1599 => x"38",
          1600 => x"80",
          1601 => x"80",
          1602 => x"81",
          1603 => x"72",
          1604 => x"0c",
          1605 => x"04",
          1606 => x"60",
          1607 => x"8c",
          1608 => x"33",
          1609 => x"5b",
          1610 => x"74",
          1611 => x"e1",
          1612 => x"a4",
          1613 => x"79",
          1614 => x"78",
          1615 => x"06",
          1616 => x"77",
          1617 => x"87",
          1618 => x"11",
          1619 => x"8c",
          1620 => x"92",
          1621 => x"59",
          1622 => x"85",
          1623 => x"98",
          1624 => x"7d",
          1625 => x"0c",
          1626 => x"08",
          1627 => x"70",
          1628 => x"53",
          1629 => x"2e",
          1630 => x"70",
          1631 => x"33",
          1632 => x"18",
          1633 => x"2a",
          1634 => x"51",
          1635 => x"2e",
          1636 => x"c0",
          1637 => x"52",
          1638 => x"87",
          1639 => x"08",
          1640 => x"2e",
          1641 => x"84",
          1642 => x"38",
          1643 => x"87",
          1644 => x"15",
          1645 => x"70",
          1646 => x"52",
          1647 => x"ff",
          1648 => x"39",
          1649 => x"81",
          1650 => x"80",
          1651 => x"52",
          1652 => x"90",
          1653 => x"80",
          1654 => x"71",
          1655 => x"7a",
          1656 => x"38",
          1657 => x"80",
          1658 => x"80",
          1659 => x"81",
          1660 => x"72",
          1661 => x"0c",
          1662 => x"04",
          1663 => x"7e",
          1664 => x"b3",
          1665 => x"88",
          1666 => x"33",
          1667 => x"56",
          1668 => x"3f",
          1669 => x"08",
          1670 => x"83",
          1671 => x"fe",
          1672 => x"87",
          1673 => x"0c",
          1674 => x"76",
          1675 => x"38",
          1676 => x"93",
          1677 => x"2b",
          1678 => x"8c",
          1679 => x"71",
          1680 => x"38",
          1681 => x"71",
          1682 => x"c6",
          1683 => x"39",
          1684 => x"81",
          1685 => x"06",
          1686 => x"71",
          1687 => x"38",
          1688 => x"8c",
          1689 => x"e8",
          1690 => x"98",
          1691 => x"71",
          1692 => x"73",
          1693 => x"92",
          1694 => x"72",
          1695 => x"06",
          1696 => x"f7",
          1697 => x"80",
          1698 => x"88",
          1699 => x"0c",
          1700 => x"80",
          1701 => x"56",
          1702 => x"56",
          1703 => x"81",
          1704 => x"8c",
          1705 => x"fe",
          1706 => x"81",
          1707 => x"33",
          1708 => x"07",
          1709 => x"0c",
          1710 => x"3d",
          1711 => x"3d",
          1712 => x"11",
          1713 => x"33",
          1714 => x"71",
          1715 => x"81",
          1716 => x"72",
          1717 => x"75",
          1718 => x"81",
          1719 => x"52",
          1720 => x"54",
          1721 => x"0d",
          1722 => x"0d",
          1723 => x"05",
          1724 => x"52",
          1725 => x"70",
          1726 => x"34",
          1727 => x"51",
          1728 => x"83",
          1729 => x"ff",
          1730 => x"75",
          1731 => x"72",
          1732 => x"54",
          1733 => x"2a",
          1734 => x"70",
          1735 => x"34",
          1736 => x"51",
          1737 => x"81",
          1738 => x"70",
          1739 => x"70",
          1740 => x"3d",
          1741 => x"3d",
          1742 => x"77",
          1743 => x"70",
          1744 => x"38",
          1745 => x"05",
          1746 => x"70",
          1747 => x"34",
          1748 => x"eb",
          1749 => x"0d",
          1750 => x"0d",
          1751 => x"54",
          1752 => x"72",
          1753 => x"54",
          1754 => x"51",
          1755 => x"84",
          1756 => x"fc",
          1757 => x"77",
          1758 => x"53",
          1759 => x"05",
          1760 => x"70",
          1761 => x"33",
          1762 => x"ff",
          1763 => x"52",
          1764 => x"2e",
          1765 => x"80",
          1766 => x"71",
          1767 => x"0c",
          1768 => x"04",
          1769 => x"74",
          1770 => x"89",
          1771 => x"2e",
          1772 => x"11",
          1773 => x"52",
          1774 => x"70",
          1775 => x"a4",
          1776 => x"0d",
          1777 => x"81",
          1778 => x"04",
          1779 => x"cb",
          1780 => x"f7",
          1781 => x"56",
          1782 => x"17",
          1783 => x"74",
          1784 => x"d6",
          1785 => x"b0",
          1786 => x"b4",
          1787 => x"81",
          1788 => x"59",
          1789 => x"81",
          1790 => x"7a",
          1791 => x"06",
          1792 => x"cb",
          1793 => x"17",
          1794 => x"08",
          1795 => x"08",
          1796 => x"08",
          1797 => x"74",
          1798 => x"38",
          1799 => x"55",
          1800 => x"09",
          1801 => x"38",
          1802 => x"18",
          1803 => x"81",
          1804 => x"f9",
          1805 => x"39",
          1806 => x"81",
          1807 => x"8b",
          1808 => x"fa",
          1809 => x"7a",
          1810 => x"57",
          1811 => x"08",
          1812 => x"75",
          1813 => x"3f",
          1814 => x"08",
          1815 => x"a4",
          1816 => x"81",
          1817 => x"b4",
          1818 => x"16",
          1819 => x"be",
          1820 => x"a4",
          1821 => x"85",
          1822 => x"81",
          1823 => x"17",
          1824 => x"cb",
          1825 => x"3d",
          1826 => x"3d",
          1827 => x"52",
          1828 => x"3f",
          1829 => x"08",
          1830 => x"a4",
          1831 => x"38",
          1832 => x"74",
          1833 => x"81",
          1834 => x"38",
          1835 => x"59",
          1836 => x"09",
          1837 => x"e3",
          1838 => x"53",
          1839 => x"08",
          1840 => x"70",
          1841 => x"91",
          1842 => x"d5",
          1843 => x"17",
          1844 => x"3f",
          1845 => x"a4",
          1846 => x"51",
          1847 => x"86",
          1848 => x"f2",
          1849 => x"17",
          1850 => x"3f",
          1851 => x"52",
          1852 => x"51",
          1853 => x"8c",
          1854 => x"84",
          1855 => x"fc",
          1856 => x"17",
          1857 => x"70",
          1858 => x"79",
          1859 => x"52",
          1860 => x"51",
          1861 => x"77",
          1862 => x"80",
          1863 => x"81",
          1864 => x"f9",
          1865 => x"cb",
          1866 => x"2e",
          1867 => x"58",
          1868 => x"a4",
          1869 => x"0d",
          1870 => x"0d",
          1871 => x"98",
          1872 => x"05",
          1873 => x"80",
          1874 => x"27",
          1875 => x"14",
          1876 => x"29",
          1877 => x"05",
          1878 => x"81",
          1879 => x"87",
          1880 => x"f9",
          1881 => x"7a",
          1882 => x"54",
          1883 => x"27",
          1884 => x"76",
          1885 => x"27",
          1886 => x"ff",
          1887 => x"58",
          1888 => x"80",
          1889 => x"82",
          1890 => x"72",
          1891 => x"38",
          1892 => x"72",
          1893 => x"8e",
          1894 => x"39",
          1895 => x"17",
          1896 => x"a4",
          1897 => x"53",
          1898 => x"fd",
          1899 => x"cb",
          1900 => x"9f",
          1901 => x"ff",
          1902 => x"11",
          1903 => x"70",
          1904 => x"18",
          1905 => x"76",
          1906 => x"53",
          1907 => x"81",
          1908 => x"80",
          1909 => x"83",
          1910 => x"b4",
          1911 => x"88",
          1912 => x"79",
          1913 => x"84",
          1914 => x"58",
          1915 => x"80",
          1916 => x"9f",
          1917 => x"80",
          1918 => x"88",
          1919 => x"08",
          1920 => x"51",
          1921 => x"81",
          1922 => x"80",
          1923 => x"10",
          1924 => x"74",
          1925 => x"51",
          1926 => x"81",
          1927 => x"83",
          1928 => x"58",
          1929 => x"87",
          1930 => x"08",
          1931 => x"51",
          1932 => x"81",
          1933 => x"9b",
          1934 => x"2b",
          1935 => x"74",
          1936 => x"51",
          1937 => x"81",
          1938 => x"f0",
          1939 => x"83",
          1940 => x"77",
          1941 => x"0c",
          1942 => x"04",
          1943 => x"7a",
          1944 => x"58",
          1945 => x"81",
          1946 => x"9e",
          1947 => x"17",
          1948 => x"96",
          1949 => x"53",
          1950 => x"81",
          1951 => x"79",
          1952 => x"72",
          1953 => x"38",
          1954 => x"72",
          1955 => x"b8",
          1956 => x"39",
          1957 => x"17",
          1958 => x"a4",
          1959 => x"53",
          1960 => x"fb",
          1961 => x"cb",
          1962 => x"81",
          1963 => x"81",
          1964 => x"83",
          1965 => x"b4",
          1966 => x"78",
          1967 => x"56",
          1968 => x"76",
          1969 => x"38",
          1970 => x"9f",
          1971 => x"33",
          1972 => x"07",
          1973 => x"74",
          1974 => x"83",
          1975 => x"89",
          1976 => x"08",
          1977 => x"51",
          1978 => x"81",
          1979 => x"59",
          1980 => x"08",
          1981 => x"74",
          1982 => x"16",
          1983 => x"84",
          1984 => x"76",
          1985 => x"88",
          1986 => x"81",
          1987 => x"8f",
          1988 => x"53",
          1989 => x"80",
          1990 => x"88",
          1991 => x"08",
          1992 => x"51",
          1993 => x"81",
          1994 => x"59",
          1995 => x"08",
          1996 => x"77",
          1997 => x"06",
          1998 => x"83",
          1999 => x"05",
          2000 => x"f7",
          2001 => x"39",
          2002 => x"a4",
          2003 => x"52",
          2004 => x"ef",
          2005 => x"a4",
          2006 => x"cb",
          2007 => x"38",
          2008 => x"06",
          2009 => x"83",
          2010 => x"18",
          2011 => x"54",
          2012 => x"f6",
          2013 => x"cb",
          2014 => x"0a",
          2015 => x"52",
          2016 => x"83",
          2017 => x"83",
          2018 => x"81",
          2019 => x"8a",
          2020 => x"f8",
          2021 => x"7c",
          2022 => x"59",
          2023 => x"81",
          2024 => x"38",
          2025 => x"08",
          2026 => x"73",
          2027 => x"38",
          2028 => x"52",
          2029 => x"a4",
          2030 => x"a4",
          2031 => x"cb",
          2032 => x"f2",
          2033 => x"82",
          2034 => x"39",
          2035 => x"e6",
          2036 => x"a4",
          2037 => x"de",
          2038 => x"78",
          2039 => x"3f",
          2040 => x"08",
          2041 => x"a4",
          2042 => x"80",
          2043 => x"cb",
          2044 => x"2e",
          2045 => x"cb",
          2046 => x"2e",
          2047 => x"53",
          2048 => x"51",
          2049 => x"81",
          2050 => x"c5",
          2051 => x"08",
          2052 => x"18",
          2053 => x"57",
          2054 => x"90",
          2055 => x"90",
          2056 => x"16",
          2057 => x"54",
          2058 => x"34",
          2059 => x"78",
          2060 => x"38",
          2061 => x"81",
          2062 => x"8a",
          2063 => x"f6",
          2064 => x"7e",
          2065 => x"5b",
          2066 => x"38",
          2067 => x"58",
          2068 => x"88",
          2069 => x"08",
          2070 => x"38",
          2071 => x"39",
          2072 => x"51",
          2073 => x"81",
          2074 => x"cb",
          2075 => x"82",
          2076 => x"cb",
          2077 => x"81",
          2078 => x"ff",
          2079 => x"38",
          2080 => x"81",
          2081 => x"26",
          2082 => x"79",
          2083 => x"08",
          2084 => x"73",
          2085 => x"b9",
          2086 => x"2e",
          2087 => x"80",
          2088 => x"1a",
          2089 => x"08",
          2090 => x"38",
          2091 => x"52",
          2092 => x"af",
          2093 => x"81",
          2094 => x"81",
          2095 => x"06",
          2096 => x"cb",
          2097 => x"81",
          2098 => x"09",
          2099 => x"72",
          2100 => x"70",
          2101 => x"cb",
          2102 => x"51",
          2103 => x"73",
          2104 => x"81",
          2105 => x"80",
          2106 => x"8c",
          2107 => x"81",
          2108 => x"38",
          2109 => x"08",
          2110 => x"73",
          2111 => x"75",
          2112 => x"77",
          2113 => x"56",
          2114 => x"76",
          2115 => x"82",
          2116 => x"26",
          2117 => x"75",
          2118 => x"f8",
          2119 => x"cb",
          2120 => x"2e",
          2121 => x"59",
          2122 => x"08",
          2123 => x"81",
          2124 => x"81",
          2125 => x"59",
          2126 => x"08",
          2127 => x"70",
          2128 => x"25",
          2129 => x"51",
          2130 => x"73",
          2131 => x"75",
          2132 => x"81",
          2133 => x"38",
          2134 => x"f5",
          2135 => x"75",
          2136 => x"f9",
          2137 => x"cb",
          2138 => x"cb",
          2139 => x"70",
          2140 => x"08",
          2141 => x"51",
          2142 => x"80",
          2143 => x"73",
          2144 => x"38",
          2145 => x"52",
          2146 => x"d0",
          2147 => x"a4",
          2148 => x"a5",
          2149 => x"18",
          2150 => x"08",
          2151 => x"18",
          2152 => x"74",
          2153 => x"38",
          2154 => x"18",
          2155 => x"33",
          2156 => x"73",
          2157 => x"97",
          2158 => x"74",
          2159 => x"38",
          2160 => x"55",
          2161 => x"cb",
          2162 => x"85",
          2163 => x"75",
          2164 => x"cb",
          2165 => x"3d",
          2166 => x"3d",
          2167 => x"52",
          2168 => x"3f",
          2169 => x"08",
          2170 => x"81",
          2171 => x"80",
          2172 => x"52",
          2173 => x"c1",
          2174 => x"a4",
          2175 => x"a4",
          2176 => x"0c",
          2177 => x"53",
          2178 => x"15",
          2179 => x"f2",
          2180 => x"56",
          2181 => x"16",
          2182 => x"22",
          2183 => x"27",
          2184 => x"54",
          2185 => x"76",
          2186 => x"33",
          2187 => x"3f",
          2188 => x"08",
          2189 => x"38",
          2190 => x"76",
          2191 => x"70",
          2192 => x"9f",
          2193 => x"56",
          2194 => x"cb",
          2195 => x"3d",
          2196 => x"3d",
          2197 => x"71",
          2198 => x"57",
          2199 => x"0a",
          2200 => x"38",
          2201 => x"53",
          2202 => x"38",
          2203 => x"0c",
          2204 => x"54",
          2205 => x"75",
          2206 => x"73",
          2207 => x"a8",
          2208 => x"73",
          2209 => x"85",
          2210 => x"0b",
          2211 => x"5a",
          2212 => x"27",
          2213 => x"a8",
          2214 => x"18",
          2215 => x"39",
          2216 => x"70",
          2217 => x"58",
          2218 => x"b2",
          2219 => x"76",
          2220 => x"3f",
          2221 => x"08",
          2222 => x"a4",
          2223 => x"bd",
          2224 => x"81",
          2225 => x"27",
          2226 => x"16",
          2227 => x"a4",
          2228 => x"38",
          2229 => x"39",
          2230 => x"55",
          2231 => x"52",
          2232 => x"d5",
          2233 => x"a4",
          2234 => x"0c",
          2235 => x"0c",
          2236 => x"53",
          2237 => x"80",
          2238 => x"85",
          2239 => x"94",
          2240 => x"2a",
          2241 => x"0c",
          2242 => x"06",
          2243 => x"9c",
          2244 => x"58",
          2245 => x"a4",
          2246 => x"0d",
          2247 => x"0d",
          2248 => x"90",
          2249 => x"05",
          2250 => x"f0",
          2251 => x"27",
          2252 => x"0b",
          2253 => x"98",
          2254 => x"84",
          2255 => x"2e",
          2256 => x"76",
          2257 => x"58",
          2258 => x"38",
          2259 => x"15",
          2260 => x"08",
          2261 => x"38",
          2262 => x"88",
          2263 => x"53",
          2264 => x"81",
          2265 => x"c0",
          2266 => x"22",
          2267 => x"89",
          2268 => x"72",
          2269 => x"74",
          2270 => x"f3",
          2271 => x"cb",
          2272 => x"82",
          2273 => x"81",
          2274 => x"27",
          2275 => x"81",
          2276 => x"a4",
          2277 => x"80",
          2278 => x"16",
          2279 => x"a4",
          2280 => x"ca",
          2281 => x"38",
          2282 => x"0c",
          2283 => x"dd",
          2284 => x"08",
          2285 => x"f9",
          2286 => x"cb",
          2287 => x"87",
          2288 => x"a4",
          2289 => x"80",
          2290 => x"55",
          2291 => x"08",
          2292 => x"38",
          2293 => x"cb",
          2294 => x"2e",
          2295 => x"cb",
          2296 => x"75",
          2297 => x"3f",
          2298 => x"08",
          2299 => x"94",
          2300 => x"52",
          2301 => x"c1",
          2302 => x"a4",
          2303 => x"0c",
          2304 => x"0c",
          2305 => x"05",
          2306 => x"80",
          2307 => x"cb",
          2308 => x"3d",
          2309 => x"3d",
          2310 => x"71",
          2311 => x"57",
          2312 => x"51",
          2313 => x"81",
          2314 => x"54",
          2315 => x"08",
          2316 => x"81",
          2317 => x"56",
          2318 => x"52",
          2319 => x"83",
          2320 => x"a4",
          2321 => x"cb",
          2322 => x"d2",
          2323 => x"a4",
          2324 => x"08",
          2325 => x"54",
          2326 => x"e5",
          2327 => x"06",
          2328 => x"58",
          2329 => x"08",
          2330 => x"38",
          2331 => x"75",
          2332 => x"80",
          2333 => x"81",
          2334 => x"7a",
          2335 => x"06",
          2336 => x"39",
          2337 => x"08",
          2338 => x"76",
          2339 => x"3f",
          2340 => x"08",
          2341 => x"a4",
          2342 => x"ff",
          2343 => x"84",
          2344 => x"06",
          2345 => x"54",
          2346 => x"a4",
          2347 => x"0d",
          2348 => x"0d",
          2349 => x"52",
          2350 => x"3f",
          2351 => x"08",
          2352 => x"06",
          2353 => x"51",
          2354 => x"83",
          2355 => x"06",
          2356 => x"14",
          2357 => x"3f",
          2358 => x"08",
          2359 => x"07",
          2360 => x"cb",
          2361 => x"3d",
          2362 => x"3d",
          2363 => x"70",
          2364 => x"06",
          2365 => x"53",
          2366 => x"ed",
          2367 => x"33",
          2368 => x"83",
          2369 => x"06",
          2370 => x"90",
          2371 => x"15",
          2372 => x"3f",
          2373 => x"04",
          2374 => x"7b",
          2375 => x"84",
          2376 => x"58",
          2377 => x"80",
          2378 => x"38",
          2379 => x"52",
          2380 => x"8f",
          2381 => x"a4",
          2382 => x"cb",
          2383 => x"f5",
          2384 => x"08",
          2385 => x"53",
          2386 => x"84",
          2387 => x"39",
          2388 => x"70",
          2389 => x"81",
          2390 => x"51",
          2391 => x"16",
          2392 => x"a4",
          2393 => x"81",
          2394 => x"38",
          2395 => x"ae",
          2396 => x"81",
          2397 => x"54",
          2398 => x"2e",
          2399 => x"8f",
          2400 => x"81",
          2401 => x"76",
          2402 => x"54",
          2403 => x"09",
          2404 => x"38",
          2405 => x"7a",
          2406 => x"80",
          2407 => x"fa",
          2408 => x"cb",
          2409 => x"81",
          2410 => x"89",
          2411 => x"08",
          2412 => x"86",
          2413 => x"98",
          2414 => x"81",
          2415 => x"8b",
          2416 => x"fb",
          2417 => x"70",
          2418 => x"81",
          2419 => x"fc",
          2420 => x"cb",
          2421 => x"81",
          2422 => x"b4",
          2423 => x"08",
          2424 => x"ec",
          2425 => x"cb",
          2426 => x"81",
          2427 => x"a0",
          2428 => x"81",
          2429 => x"52",
          2430 => x"51",
          2431 => x"8b",
          2432 => x"52",
          2433 => x"51",
          2434 => x"81",
          2435 => x"34",
          2436 => x"a4",
          2437 => x"0d",
          2438 => x"0d",
          2439 => x"98",
          2440 => x"70",
          2441 => x"ec",
          2442 => x"cb",
          2443 => x"38",
          2444 => x"53",
          2445 => x"81",
          2446 => x"34",
          2447 => x"04",
          2448 => x"78",
          2449 => x"80",
          2450 => x"34",
          2451 => x"80",
          2452 => x"38",
          2453 => x"18",
          2454 => x"9c",
          2455 => x"70",
          2456 => x"56",
          2457 => x"a0",
          2458 => x"71",
          2459 => x"81",
          2460 => x"81",
          2461 => x"89",
          2462 => x"06",
          2463 => x"73",
          2464 => x"55",
          2465 => x"55",
          2466 => x"81",
          2467 => x"81",
          2468 => x"74",
          2469 => x"75",
          2470 => x"52",
          2471 => x"13",
          2472 => x"08",
          2473 => x"33",
          2474 => x"9c",
          2475 => x"11",
          2476 => x"8a",
          2477 => x"a4",
          2478 => x"96",
          2479 => x"e7",
          2480 => x"a4",
          2481 => x"23",
          2482 => x"e7",
          2483 => x"cb",
          2484 => x"17",
          2485 => x"0d",
          2486 => x"0d",
          2487 => x"5e",
          2488 => x"70",
          2489 => x"55",
          2490 => x"83",
          2491 => x"73",
          2492 => x"91",
          2493 => x"2e",
          2494 => x"1d",
          2495 => x"0c",
          2496 => x"15",
          2497 => x"70",
          2498 => x"56",
          2499 => x"09",
          2500 => x"38",
          2501 => x"80",
          2502 => x"30",
          2503 => x"78",
          2504 => x"54",
          2505 => x"73",
          2506 => x"60",
          2507 => x"54",
          2508 => x"96",
          2509 => x"0b",
          2510 => x"80",
          2511 => x"f6",
          2512 => x"cb",
          2513 => x"85",
          2514 => x"3d",
          2515 => x"5c",
          2516 => x"53",
          2517 => x"51",
          2518 => x"80",
          2519 => x"88",
          2520 => x"5c",
          2521 => x"09",
          2522 => x"d4",
          2523 => x"70",
          2524 => x"71",
          2525 => x"30",
          2526 => x"73",
          2527 => x"51",
          2528 => x"57",
          2529 => x"38",
          2530 => x"75",
          2531 => x"17",
          2532 => x"75",
          2533 => x"30",
          2534 => x"51",
          2535 => x"80",
          2536 => x"38",
          2537 => x"87",
          2538 => x"26",
          2539 => x"77",
          2540 => x"a4",
          2541 => x"27",
          2542 => x"a0",
          2543 => x"39",
          2544 => x"33",
          2545 => x"57",
          2546 => x"27",
          2547 => x"75",
          2548 => x"30",
          2549 => x"32",
          2550 => x"80",
          2551 => x"25",
          2552 => x"56",
          2553 => x"80",
          2554 => x"84",
          2555 => x"58",
          2556 => x"70",
          2557 => x"55",
          2558 => x"09",
          2559 => x"38",
          2560 => x"80",
          2561 => x"30",
          2562 => x"77",
          2563 => x"54",
          2564 => x"81",
          2565 => x"ae",
          2566 => x"06",
          2567 => x"54",
          2568 => x"74",
          2569 => x"80",
          2570 => x"7b",
          2571 => x"30",
          2572 => x"70",
          2573 => x"25",
          2574 => x"07",
          2575 => x"51",
          2576 => x"a7",
          2577 => x"8b",
          2578 => x"39",
          2579 => x"54",
          2580 => x"8c",
          2581 => x"ff",
          2582 => x"80",
          2583 => x"54",
          2584 => x"e1",
          2585 => x"a4",
          2586 => x"b2",
          2587 => x"70",
          2588 => x"71",
          2589 => x"54",
          2590 => x"81",
          2591 => x"80",
          2592 => x"38",
          2593 => x"76",
          2594 => x"df",
          2595 => x"54",
          2596 => x"81",
          2597 => x"55",
          2598 => x"34",
          2599 => x"52",
          2600 => x"51",
          2601 => x"81",
          2602 => x"bf",
          2603 => x"16",
          2604 => x"26",
          2605 => x"16",
          2606 => x"06",
          2607 => x"17",
          2608 => x"34",
          2609 => x"fd",
          2610 => x"19",
          2611 => x"80",
          2612 => x"79",
          2613 => x"81",
          2614 => x"81",
          2615 => x"85",
          2616 => x"54",
          2617 => x"8f",
          2618 => x"86",
          2619 => x"39",
          2620 => x"f3",
          2621 => x"73",
          2622 => x"80",
          2623 => x"52",
          2624 => x"ce",
          2625 => x"a4",
          2626 => x"cb",
          2627 => x"d7",
          2628 => x"08",
          2629 => x"e6",
          2630 => x"cb",
          2631 => x"81",
          2632 => x"80",
          2633 => x"1b",
          2634 => x"55",
          2635 => x"2e",
          2636 => x"8b",
          2637 => x"06",
          2638 => x"1c",
          2639 => x"33",
          2640 => x"70",
          2641 => x"55",
          2642 => x"38",
          2643 => x"52",
          2644 => x"9f",
          2645 => x"a4",
          2646 => x"8b",
          2647 => x"7a",
          2648 => x"3f",
          2649 => x"75",
          2650 => x"57",
          2651 => x"2e",
          2652 => x"84",
          2653 => x"06",
          2654 => x"75",
          2655 => x"81",
          2656 => x"2a",
          2657 => x"73",
          2658 => x"38",
          2659 => x"54",
          2660 => x"fb",
          2661 => x"80",
          2662 => x"34",
          2663 => x"c1",
          2664 => x"06",
          2665 => x"38",
          2666 => x"39",
          2667 => x"70",
          2668 => x"54",
          2669 => x"86",
          2670 => x"84",
          2671 => x"06",
          2672 => x"73",
          2673 => x"38",
          2674 => x"83",
          2675 => x"b4",
          2676 => x"51",
          2677 => x"81",
          2678 => x"88",
          2679 => x"ea",
          2680 => x"cb",
          2681 => x"3d",
          2682 => x"3d",
          2683 => x"ff",
          2684 => x"71",
          2685 => x"5c",
          2686 => x"80",
          2687 => x"38",
          2688 => x"05",
          2689 => x"a0",
          2690 => x"71",
          2691 => x"38",
          2692 => x"71",
          2693 => x"81",
          2694 => x"38",
          2695 => x"11",
          2696 => x"06",
          2697 => x"70",
          2698 => x"38",
          2699 => x"81",
          2700 => x"05",
          2701 => x"76",
          2702 => x"38",
          2703 => x"ba",
          2704 => x"77",
          2705 => x"57",
          2706 => x"05",
          2707 => x"70",
          2708 => x"33",
          2709 => x"53",
          2710 => x"99",
          2711 => x"e0",
          2712 => x"ff",
          2713 => x"ff",
          2714 => x"70",
          2715 => x"38",
          2716 => x"81",
          2717 => x"51",
          2718 => x"9f",
          2719 => x"72",
          2720 => x"81",
          2721 => x"70",
          2722 => x"72",
          2723 => x"32",
          2724 => x"72",
          2725 => x"73",
          2726 => x"53",
          2727 => x"70",
          2728 => x"38",
          2729 => x"19",
          2730 => x"75",
          2731 => x"38",
          2732 => x"83",
          2733 => x"74",
          2734 => x"59",
          2735 => x"39",
          2736 => x"33",
          2737 => x"cb",
          2738 => x"3d",
          2739 => x"3d",
          2740 => x"80",
          2741 => x"34",
          2742 => x"17",
          2743 => x"75",
          2744 => x"3f",
          2745 => x"cb",
          2746 => x"80",
          2747 => x"16",
          2748 => x"3f",
          2749 => x"08",
          2750 => x"06",
          2751 => x"73",
          2752 => x"2e",
          2753 => x"80",
          2754 => x"0b",
          2755 => x"56",
          2756 => x"e9",
          2757 => x"06",
          2758 => x"57",
          2759 => x"32",
          2760 => x"80",
          2761 => x"51",
          2762 => x"8a",
          2763 => x"e8",
          2764 => x"06",
          2765 => x"53",
          2766 => x"52",
          2767 => x"51",
          2768 => x"81",
          2769 => x"55",
          2770 => x"08",
          2771 => x"38",
          2772 => x"ba",
          2773 => x"86",
          2774 => x"97",
          2775 => x"a4",
          2776 => x"cb",
          2777 => x"2e",
          2778 => x"55",
          2779 => x"a4",
          2780 => x"0d",
          2781 => x"0d",
          2782 => x"05",
          2783 => x"33",
          2784 => x"75",
          2785 => x"fc",
          2786 => x"cb",
          2787 => x"8b",
          2788 => x"81",
          2789 => x"24",
          2790 => x"81",
          2791 => x"84",
          2792 => x"c0",
          2793 => x"55",
          2794 => x"73",
          2795 => x"e6",
          2796 => x"0c",
          2797 => x"06",
          2798 => x"57",
          2799 => x"ae",
          2800 => x"33",
          2801 => x"3f",
          2802 => x"08",
          2803 => x"70",
          2804 => x"55",
          2805 => x"76",
          2806 => x"b8",
          2807 => x"2a",
          2808 => x"51",
          2809 => x"72",
          2810 => x"86",
          2811 => x"74",
          2812 => x"15",
          2813 => x"81",
          2814 => x"d7",
          2815 => x"cb",
          2816 => x"ff",
          2817 => x"06",
          2818 => x"56",
          2819 => x"38",
          2820 => x"8f",
          2821 => x"2a",
          2822 => x"51",
          2823 => x"72",
          2824 => x"80",
          2825 => x"52",
          2826 => x"3f",
          2827 => x"08",
          2828 => x"57",
          2829 => x"09",
          2830 => x"e2",
          2831 => x"74",
          2832 => x"56",
          2833 => x"33",
          2834 => x"72",
          2835 => x"38",
          2836 => x"51",
          2837 => x"81",
          2838 => x"57",
          2839 => x"84",
          2840 => x"ff",
          2841 => x"56",
          2842 => x"25",
          2843 => x"0b",
          2844 => x"56",
          2845 => x"05",
          2846 => x"83",
          2847 => x"2e",
          2848 => x"52",
          2849 => x"c6",
          2850 => x"a4",
          2851 => x"06",
          2852 => x"27",
          2853 => x"16",
          2854 => x"27",
          2855 => x"56",
          2856 => x"84",
          2857 => x"56",
          2858 => x"84",
          2859 => x"14",
          2860 => x"3f",
          2861 => x"08",
          2862 => x"06",
          2863 => x"80",
          2864 => x"06",
          2865 => x"80",
          2866 => x"db",
          2867 => x"cb",
          2868 => x"ff",
          2869 => x"77",
          2870 => x"d8",
          2871 => x"de",
          2872 => x"a4",
          2873 => x"9c",
          2874 => x"c4",
          2875 => x"15",
          2876 => x"14",
          2877 => x"70",
          2878 => x"51",
          2879 => x"56",
          2880 => x"84",
          2881 => x"81",
          2882 => x"71",
          2883 => x"16",
          2884 => x"53",
          2885 => x"23",
          2886 => x"8b",
          2887 => x"73",
          2888 => x"80",
          2889 => x"8d",
          2890 => x"39",
          2891 => x"51",
          2892 => x"81",
          2893 => x"53",
          2894 => x"08",
          2895 => x"72",
          2896 => x"8d",
          2897 => x"ce",
          2898 => x"14",
          2899 => x"3f",
          2900 => x"08",
          2901 => x"06",
          2902 => x"38",
          2903 => x"51",
          2904 => x"81",
          2905 => x"55",
          2906 => x"51",
          2907 => x"81",
          2908 => x"83",
          2909 => x"53",
          2910 => x"80",
          2911 => x"38",
          2912 => x"78",
          2913 => x"2a",
          2914 => x"78",
          2915 => x"86",
          2916 => x"22",
          2917 => x"31",
          2918 => x"83",
          2919 => x"a4",
          2920 => x"cb",
          2921 => x"2e",
          2922 => x"81",
          2923 => x"80",
          2924 => x"f5",
          2925 => x"83",
          2926 => x"ff",
          2927 => x"38",
          2928 => x"9f",
          2929 => x"38",
          2930 => x"39",
          2931 => x"80",
          2932 => x"38",
          2933 => x"98",
          2934 => x"a0",
          2935 => x"1c",
          2936 => x"0c",
          2937 => x"17",
          2938 => x"76",
          2939 => x"81",
          2940 => x"80",
          2941 => x"d9",
          2942 => x"cb",
          2943 => x"ff",
          2944 => x"8d",
          2945 => x"8e",
          2946 => x"8a",
          2947 => x"14",
          2948 => x"3f",
          2949 => x"08",
          2950 => x"74",
          2951 => x"a2",
          2952 => x"79",
          2953 => x"ee",
          2954 => x"a8",
          2955 => x"15",
          2956 => x"2e",
          2957 => x"10",
          2958 => x"2a",
          2959 => x"05",
          2960 => x"ff",
          2961 => x"53",
          2962 => x"9c",
          2963 => x"81",
          2964 => x"0b",
          2965 => x"ff",
          2966 => x"0c",
          2967 => x"84",
          2968 => x"83",
          2969 => x"06",
          2970 => x"80",
          2971 => x"d8",
          2972 => x"cb",
          2973 => x"ff",
          2974 => x"72",
          2975 => x"81",
          2976 => x"38",
          2977 => x"73",
          2978 => x"3f",
          2979 => x"08",
          2980 => x"81",
          2981 => x"84",
          2982 => x"b2",
          2983 => x"87",
          2984 => x"a4",
          2985 => x"ff",
          2986 => x"82",
          2987 => x"09",
          2988 => x"c8",
          2989 => x"51",
          2990 => x"81",
          2991 => x"84",
          2992 => x"d2",
          2993 => x"06",
          2994 => x"98",
          2995 => x"ee",
          2996 => x"a4",
          2997 => x"85",
          2998 => x"09",
          2999 => x"38",
          3000 => x"51",
          3001 => x"81",
          3002 => x"90",
          3003 => x"a0",
          3004 => x"ca",
          3005 => x"a4",
          3006 => x"0c",
          3007 => x"81",
          3008 => x"81",
          3009 => x"81",
          3010 => x"72",
          3011 => x"80",
          3012 => x"0c",
          3013 => x"81",
          3014 => x"90",
          3015 => x"fb",
          3016 => x"54",
          3017 => x"80",
          3018 => x"73",
          3019 => x"80",
          3020 => x"72",
          3021 => x"80",
          3022 => x"86",
          3023 => x"15",
          3024 => x"71",
          3025 => x"81",
          3026 => x"81",
          3027 => x"d0",
          3028 => x"cb",
          3029 => x"06",
          3030 => x"38",
          3031 => x"54",
          3032 => x"80",
          3033 => x"71",
          3034 => x"81",
          3035 => x"87",
          3036 => x"fa",
          3037 => x"ab",
          3038 => x"58",
          3039 => x"05",
          3040 => x"e6",
          3041 => x"80",
          3042 => x"a4",
          3043 => x"38",
          3044 => x"08",
          3045 => x"cb",
          3046 => x"08",
          3047 => x"80",
          3048 => x"80",
          3049 => x"54",
          3050 => x"84",
          3051 => x"34",
          3052 => x"75",
          3053 => x"2e",
          3054 => x"53",
          3055 => x"53",
          3056 => x"f7",
          3057 => x"cb",
          3058 => x"73",
          3059 => x"0c",
          3060 => x"04",
          3061 => x"67",
          3062 => x"80",
          3063 => x"59",
          3064 => x"78",
          3065 => x"c8",
          3066 => x"06",
          3067 => x"3d",
          3068 => x"99",
          3069 => x"52",
          3070 => x"3f",
          3071 => x"08",
          3072 => x"a4",
          3073 => x"38",
          3074 => x"52",
          3075 => x"52",
          3076 => x"3f",
          3077 => x"08",
          3078 => x"a4",
          3079 => x"02",
          3080 => x"33",
          3081 => x"55",
          3082 => x"25",
          3083 => x"55",
          3084 => x"54",
          3085 => x"81",
          3086 => x"80",
          3087 => x"74",
          3088 => x"81",
          3089 => x"75",
          3090 => x"3f",
          3091 => x"08",
          3092 => x"02",
          3093 => x"91",
          3094 => x"81",
          3095 => x"82",
          3096 => x"06",
          3097 => x"80",
          3098 => x"88",
          3099 => x"39",
          3100 => x"58",
          3101 => x"38",
          3102 => x"70",
          3103 => x"54",
          3104 => x"81",
          3105 => x"52",
          3106 => x"a5",
          3107 => x"a4",
          3108 => x"88",
          3109 => x"62",
          3110 => x"d4",
          3111 => x"54",
          3112 => x"15",
          3113 => x"62",
          3114 => x"e8",
          3115 => x"52",
          3116 => x"51",
          3117 => x"7a",
          3118 => x"83",
          3119 => x"80",
          3120 => x"38",
          3121 => x"08",
          3122 => x"53",
          3123 => x"3d",
          3124 => x"dd",
          3125 => x"cb",
          3126 => x"81",
          3127 => x"82",
          3128 => x"39",
          3129 => x"38",
          3130 => x"33",
          3131 => x"70",
          3132 => x"55",
          3133 => x"2e",
          3134 => x"55",
          3135 => x"77",
          3136 => x"81",
          3137 => x"73",
          3138 => x"38",
          3139 => x"54",
          3140 => x"a0",
          3141 => x"82",
          3142 => x"52",
          3143 => x"a3",
          3144 => x"a4",
          3145 => x"18",
          3146 => x"55",
          3147 => x"a4",
          3148 => x"38",
          3149 => x"70",
          3150 => x"54",
          3151 => x"86",
          3152 => x"c0",
          3153 => x"b0",
          3154 => x"1b",
          3155 => x"1b",
          3156 => x"70",
          3157 => x"d9",
          3158 => x"a4",
          3159 => x"a4",
          3160 => x"0c",
          3161 => x"52",
          3162 => x"3f",
          3163 => x"08",
          3164 => x"08",
          3165 => x"77",
          3166 => x"86",
          3167 => x"1a",
          3168 => x"1a",
          3169 => x"91",
          3170 => x"0b",
          3171 => x"80",
          3172 => x"0c",
          3173 => x"70",
          3174 => x"54",
          3175 => x"81",
          3176 => x"cb",
          3177 => x"2e",
          3178 => x"81",
          3179 => x"94",
          3180 => x"17",
          3181 => x"2b",
          3182 => x"57",
          3183 => x"52",
          3184 => x"9f",
          3185 => x"a4",
          3186 => x"cb",
          3187 => x"26",
          3188 => x"55",
          3189 => x"08",
          3190 => x"81",
          3191 => x"79",
          3192 => x"31",
          3193 => x"70",
          3194 => x"25",
          3195 => x"76",
          3196 => x"81",
          3197 => x"55",
          3198 => x"38",
          3199 => x"0c",
          3200 => x"75",
          3201 => x"54",
          3202 => x"a2",
          3203 => x"7a",
          3204 => x"3f",
          3205 => x"08",
          3206 => x"55",
          3207 => x"89",
          3208 => x"a4",
          3209 => x"1a",
          3210 => x"80",
          3211 => x"54",
          3212 => x"a4",
          3213 => x"0d",
          3214 => x"0d",
          3215 => x"64",
          3216 => x"59",
          3217 => x"90",
          3218 => x"52",
          3219 => x"cf",
          3220 => x"a4",
          3221 => x"cb",
          3222 => x"38",
          3223 => x"55",
          3224 => x"86",
          3225 => x"82",
          3226 => x"19",
          3227 => x"55",
          3228 => x"80",
          3229 => x"38",
          3230 => x"0b",
          3231 => x"82",
          3232 => x"39",
          3233 => x"1a",
          3234 => x"82",
          3235 => x"19",
          3236 => x"08",
          3237 => x"7c",
          3238 => x"74",
          3239 => x"2e",
          3240 => x"94",
          3241 => x"83",
          3242 => x"56",
          3243 => x"38",
          3244 => x"22",
          3245 => x"89",
          3246 => x"55",
          3247 => x"75",
          3248 => x"19",
          3249 => x"39",
          3250 => x"52",
          3251 => x"93",
          3252 => x"a4",
          3253 => x"75",
          3254 => x"38",
          3255 => x"ff",
          3256 => x"98",
          3257 => x"19",
          3258 => x"51",
          3259 => x"81",
          3260 => x"80",
          3261 => x"38",
          3262 => x"08",
          3263 => x"2a",
          3264 => x"80",
          3265 => x"38",
          3266 => x"8a",
          3267 => x"5c",
          3268 => x"27",
          3269 => x"7a",
          3270 => x"54",
          3271 => x"52",
          3272 => x"51",
          3273 => x"81",
          3274 => x"fe",
          3275 => x"83",
          3276 => x"56",
          3277 => x"9f",
          3278 => x"08",
          3279 => x"74",
          3280 => x"38",
          3281 => x"b4",
          3282 => x"16",
          3283 => x"89",
          3284 => x"51",
          3285 => x"77",
          3286 => x"b9",
          3287 => x"1a",
          3288 => x"08",
          3289 => x"84",
          3290 => x"57",
          3291 => x"27",
          3292 => x"56",
          3293 => x"52",
          3294 => x"c7",
          3295 => x"a4",
          3296 => x"38",
          3297 => x"19",
          3298 => x"06",
          3299 => x"52",
          3300 => x"a2",
          3301 => x"31",
          3302 => x"7f",
          3303 => x"94",
          3304 => x"94",
          3305 => x"5c",
          3306 => x"80",
          3307 => x"cb",
          3308 => x"3d",
          3309 => x"3d",
          3310 => x"65",
          3311 => x"5d",
          3312 => x"0c",
          3313 => x"05",
          3314 => x"f6",
          3315 => x"cb",
          3316 => x"81",
          3317 => x"8a",
          3318 => x"33",
          3319 => x"2e",
          3320 => x"56",
          3321 => x"90",
          3322 => x"81",
          3323 => x"06",
          3324 => x"87",
          3325 => x"2e",
          3326 => x"95",
          3327 => x"91",
          3328 => x"56",
          3329 => x"81",
          3330 => x"34",
          3331 => x"8e",
          3332 => x"08",
          3333 => x"56",
          3334 => x"84",
          3335 => x"5c",
          3336 => x"82",
          3337 => x"18",
          3338 => x"ff",
          3339 => x"74",
          3340 => x"7e",
          3341 => x"ff",
          3342 => x"2a",
          3343 => x"7a",
          3344 => x"8c",
          3345 => x"08",
          3346 => x"38",
          3347 => x"39",
          3348 => x"52",
          3349 => x"e7",
          3350 => x"a4",
          3351 => x"cb",
          3352 => x"2e",
          3353 => x"74",
          3354 => x"91",
          3355 => x"2e",
          3356 => x"74",
          3357 => x"88",
          3358 => x"38",
          3359 => x"0c",
          3360 => x"15",
          3361 => x"08",
          3362 => x"06",
          3363 => x"51",
          3364 => x"81",
          3365 => x"fe",
          3366 => x"18",
          3367 => x"51",
          3368 => x"81",
          3369 => x"80",
          3370 => x"38",
          3371 => x"08",
          3372 => x"2a",
          3373 => x"80",
          3374 => x"38",
          3375 => x"8a",
          3376 => x"5b",
          3377 => x"27",
          3378 => x"7b",
          3379 => x"54",
          3380 => x"52",
          3381 => x"51",
          3382 => x"81",
          3383 => x"fe",
          3384 => x"b0",
          3385 => x"31",
          3386 => x"79",
          3387 => x"84",
          3388 => x"16",
          3389 => x"89",
          3390 => x"52",
          3391 => x"cc",
          3392 => x"55",
          3393 => x"16",
          3394 => x"2b",
          3395 => x"39",
          3396 => x"94",
          3397 => x"93",
          3398 => x"cd",
          3399 => x"cb",
          3400 => x"e3",
          3401 => x"b0",
          3402 => x"76",
          3403 => x"94",
          3404 => x"ff",
          3405 => x"71",
          3406 => x"7b",
          3407 => x"38",
          3408 => x"18",
          3409 => x"51",
          3410 => x"81",
          3411 => x"fd",
          3412 => x"53",
          3413 => x"18",
          3414 => x"06",
          3415 => x"51",
          3416 => x"7e",
          3417 => x"83",
          3418 => x"76",
          3419 => x"17",
          3420 => x"1e",
          3421 => x"18",
          3422 => x"0c",
          3423 => x"58",
          3424 => x"74",
          3425 => x"38",
          3426 => x"8c",
          3427 => x"90",
          3428 => x"33",
          3429 => x"55",
          3430 => x"34",
          3431 => x"81",
          3432 => x"90",
          3433 => x"f8",
          3434 => x"8b",
          3435 => x"53",
          3436 => x"f2",
          3437 => x"cb",
          3438 => x"81",
          3439 => x"80",
          3440 => x"16",
          3441 => x"2a",
          3442 => x"51",
          3443 => x"80",
          3444 => x"38",
          3445 => x"52",
          3446 => x"e7",
          3447 => x"a4",
          3448 => x"cb",
          3449 => x"d4",
          3450 => x"08",
          3451 => x"a0",
          3452 => x"73",
          3453 => x"88",
          3454 => x"74",
          3455 => x"51",
          3456 => x"8c",
          3457 => x"9c",
          3458 => x"fb",
          3459 => x"b2",
          3460 => x"15",
          3461 => x"3f",
          3462 => x"15",
          3463 => x"3f",
          3464 => x"0b",
          3465 => x"78",
          3466 => x"3f",
          3467 => x"08",
          3468 => x"81",
          3469 => x"57",
          3470 => x"34",
          3471 => x"a4",
          3472 => x"0d",
          3473 => x"0d",
          3474 => x"54",
          3475 => x"81",
          3476 => x"53",
          3477 => x"08",
          3478 => x"3d",
          3479 => x"73",
          3480 => x"3f",
          3481 => x"08",
          3482 => x"a4",
          3483 => x"81",
          3484 => x"74",
          3485 => x"cb",
          3486 => x"3d",
          3487 => x"3d",
          3488 => x"51",
          3489 => x"8b",
          3490 => x"81",
          3491 => x"24",
          3492 => x"cb",
          3493 => x"cb",
          3494 => x"52",
          3495 => x"a4",
          3496 => x"0d",
          3497 => x"0d",
          3498 => x"3d",
          3499 => x"94",
          3500 => x"c1",
          3501 => x"a4",
          3502 => x"cb",
          3503 => x"e0",
          3504 => x"63",
          3505 => x"d4",
          3506 => x"8d",
          3507 => x"a4",
          3508 => x"cb",
          3509 => x"38",
          3510 => x"05",
          3511 => x"2b",
          3512 => x"80",
          3513 => x"76",
          3514 => x"0c",
          3515 => x"02",
          3516 => x"70",
          3517 => x"81",
          3518 => x"56",
          3519 => x"9e",
          3520 => x"53",
          3521 => x"db",
          3522 => x"cb",
          3523 => x"15",
          3524 => x"81",
          3525 => x"84",
          3526 => x"06",
          3527 => x"55",
          3528 => x"a4",
          3529 => x"0d",
          3530 => x"0d",
          3531 => x"5b",
          3532 => x"80",
          3533 => x"ff",
          3534 => x"9f",
          3535 => x"b5",
          3536 => x"a4",
          3537 => x"cb",
          3538 => x"fc",
          3539 => x"7a",
          3540 => x"08",
          3541 => x"64",
          3542 => x"2e",
          3543 => x"a0",
          3544 => x"70",
          3545 => x"ea",
          3546 => x"a4",
          3547 => x"cb",
          3548 => x"d4",
          3549 => x"7b",
          3550 => x"3f",
          3551 => x"08",
          3552 => x"a4",
          3553 => x"38",
          3554 => x"51",
          3555 => x"81",
          3556 => x"45",
          3557 => x"51",
          3558 => x"81",
          3559 => x"57",
          3560 => x"08",
          3561 => x"80",
          3562 => x"da",
          3563 => x"cb",
          3564 => x"81",
          3565 => x"a4",
          3566 => x"7b",
          3567 => x"3f",
          3568 => x"a4",
          3569 => x"38",
          3570 => x"51",
          3571 => x"81",
          3572 => x"57",
          3573 => x"08",
          3574 => x"38",
          3575 => x"09",
          3576 => x"38",
          3577 => x"e0",
          3578 => x"dc",
          3579 => x"ff",
          3580 => x"74",
          3581 => x"3f",
          3582 => x"78",
          3583 => x"33",
          3584 => x"56",
          3585 => x"91",
          3586 => x"05",
          3587 => x"81",
          3588 => x"56",
          3589 => x"f5",
          3590 => x"54",
          3591 => x"81",
          3592 => x"80",
          3593 => x"78",
          3594 => x"55",
          3595 => x"11",
          3596 => x"18",
          3597 => x"58",
          3598 => x"34",
          3599 => x"ff",
          3600 => x"55",
          3601 => x"34",
          3602 => x"77",
          3603 => x"81",
          3604 => x"ff",
          3605 => x"55",
          3606 => x"34",
          3607 => x"cb",
          3608 => x"84",
          3609 => x"f0",
          3610 => x"70",
          3611 => x"56",
          3612 => x"76",
          3613 => x"81",
          3614 => x"70",
          3615 => x"56",
          3616 => x"82",
          3617 => x"78",
          3618 => x"80",
          3619 => x"27",
          3620 => x"19",
          3621 => x"7a",
          3622 => x"5c",
          3623 => x"55",
          3624 => x"7a",
          3625 => x"5c",
          3626 => x"2e",
          3627 => x"85",
          3628 => x"94",
          3629 => x"81",
          3630 => x"73",
          3631 => x"81",
          3632 => x"7a",
          3633 => x"38",
          3634 => x"76",
          3635 => x"0c",
          3636 => x"04",
          3637 => x"7b",
          3638 => x"fc",
          3639 => x"53",
          3640 => x"bb",
          3641 => x"a4",
          3642 => x"cb",
          3643 => x"fa",
          3644 => x"33",
          3645 => x"f2",
          3646 => x"08",
          3647 => x"27",
          3648 => x"15",
          3649 => x"2a",
          3650 => x"51",
          3651 => x"83",
          3652 => x"94",
          3653 => x"80",
          3654 => x"0c",
          3655 => x"2e",
          3656 => x"79",
          3657 => x"70",
          3658 => x"51",
          3659 => x"2e",
          3660 => x"52",
          3661 => x"ff",
          3662 => x"81",
          3663 => x"ff",
          3664 => x"70",
          3665 => x"ff",
          3666 => x"81",
          3667 => x"73",
          3668 => x"76",
          3669 => x"06",
          3670 => x"0c",
          3671 => x"98",
          3672 => x"58",
          3673 => x"39",
          3674 => x"54",
          3675 => x"73",
          3676 => x"cd",
          3677 => x"cb",
          3678 => x"81",
          3679 => x"81",
          3680 => x"38",
          3681 => x"08",
          3682 => x"9b",
          3683 => x"a4",
          3684 => x"0c",
          3685 => x"0c",
          3686 => x"81",
          3687 => x"76",
          3688 => x"38",
          3689 => x"94",
          3690 => x"94",
          3691 => x"16",
          3692 => x"2a",
          3693 => x"51",
          3694 => x"72",
          3695 => x"38",
          3696 => x"51",
          3697 => x"81",
          3698 => x"54",
          3699 => x"08",
          3700 => x"cb",
          3701 => x"a7",
          3702 => x"74",
          3703 => x"3f",
          3704 => x"08",
          3705 => x"2e",
          3706 => x"74",
          3707 => x"79",
          3708 => x"14",
          3709 => x"38",
          3710 => x"0c",
          3711 => x"94",
          3712 => x"94",
          3713 => x"83",
          3714 => x"72",
          3715 => x"38",
          3716 => x"51",
          3717 => x"81",
          3718 => x"94",
          3719 => x"91",
          3720 => x"53",
          3721 => x"81",
          3722 => x"34",
          3723 => x"39",
          3724 => x"81",
          3725 => x"05",
          3726 => x"08",
          3727 => x"08",
          3728 => x"38",
          3729 => x"0c",
          3730 => x"80",
          3731 => x"72",
          3732 => x"73",
          3733 => x"53",
          3734 => x"8c",
          3735 => x"16",
          3736 => x"38",
          3737 => x"0c",
          3738 => x"81",
          3739 => x"8b",
          3740 => x"f9",
          3741 => x"56",
          3742 => x"80",
          3743 => x"38",
          3744 => x"3d",
          3745 => x"8a",
          3746 => x"51",
          3747 => x"81",
          3748 => x"55",
          3749 => x"08",
          3750 => x"77",
          3751 => x"52",
          3752 => x"b5",
          3753 => x"a4",
          3754 => x"cb",
          3755 => x"c3",
          3756 => x"33",
          3757 => x"55",
          3758 => x"24",
          3759 => x"16",
          3760 => x"2a",
          3761 => x"51",
          3762 => x"80",
          3763 => x"9c",
          3764 => x"77",
          3765 => x"3f",
          3766 => x"08",
          3767 => x"77",
          3768 => x"22",
          3769 => x"74",
          3770 => x"ce",
          3771 => x"cb",
          3772 => x"74",
          3773 => x"81",
          3774 => x"85",
          3775 => x"74",
          3776 => x"38",
          3777 => x"74",
          3778 => x"cb",
          3779 => x"3d",
          3780 => x"3d",
          3781 => x"3d",
          3782 => x"70",
          3783 => x"ff",
          3784 => x"a4",
          3785 => x"81",
          3786 => x"73",
          3787 => x"0d",
          3788 => x"0d",
          3789 => x"3d",
          3790 => x"71",
          3791 => x"e7",
          3792 => x"cb",
          3793 => x"81",
          3794 => x"80",
          3795 => x"93",
          3796 => x"a4",
          3797 => x"51",
          3798 => x"81",
          3799 => x"53",
          3800 => x"81",
          3801 => x"52",
          3802 => x"ac",
          3803 => x"a4",
          3804 => x"cb",
          3805 => x"2e",
          3806 => x"85",
          3807 => x"87",
          3808 => x"a4",
          3809 => x"74",
          3810 => x"d5",
          3811 => x"52",
          3812 => x"89",
          3813 => x"a4",
          3814 => x"70",
          3815 => x"07",
          3816 => x"81",
          3817 => x"06",
          3818 => x"54",
          3819 => x"a4",
          3820 => x"0d",
          3821 => x"0d",
          3822 => x"53",
          3823 => x"53",
          3824 => x"56",
          3825 => x"81",
          3826 => x"55",
          3827 => x"08",
          3828 => x"52",
          3829 => x"81",
          3830 => x"a4",
          3831 => x"cb",
          3832 => x"38",
          3833 => x"05",
          3834 => x"2b",
          3835 => x"80",
          3836 => x"86",
          3837 => x"76",
          3838 => x"38",
          3839 => x"51",
          3840 => x"74",
          3841 => x"0c",
          3842 => x"04",
          3843 => x"63",
          3844 => x"80",
          3845 => x"ec",
          3846 => x"3d",
          3847 => x"3f",
          3848 => x"08",
          3849 => x"a4",
          3850 => x"38",
          3851 => x"73",
          3852 => x"08",
          3853 => x"13",
          3854 => x"58",
          3855 => x"26",
          3856 => x"7c",
          3857 => x"39",
          3858 => x"cc",
          3859 => x"81",
          3860 => x"cb",
          3861 => x"33",
          3862 => x"81",
          3863 => x"06",
          3864 => x"75",
          3865 => x"52",
          3866 => x"05",
          3867 => x"3f",
          3868 => x"08",
          3869 => x"38",
          3870 => x"08",
          3871 => x"38",
          3872 => x"08",
          3873 => x"cb",
          3874 => x"80",
          3875 => x"81",
          3876 => x"59",
          3877 => x"14",
          3878 => x"ca",
          3879 => x"39",
          3880 => x"81",
          3881 => x"57",
          3882 => x"38",
          3883 => x"18",
          3884 => x"ff",
          3885 => x"81",
          3886 => x"5b",
          3887 => x"08",
          3888 => x"7c",
          3889 => x"12",
          3890 => x"52",
          3891 => x"82",
          3892 => x"06",
          3893 => x"14",
          3894 => x"cb",
          3895 => x"a4",
          3896 => x"ff",
          3897 => x"70",
          3898 => x"82",
          3899 => x"51",
          3900 => x"b4",
          3901 => x"bb",
          3902 => x"cb",
          3903 => x"0a",
          3904 => x"70",
          3905 => x"84",
          3906 => x"51",
          3907 => x"ff",
          3908 => x"56",
          3909 => x"38",
          3910 => x"7c",
          3911 => x"0c",
          3912 => x"81",
          3913 => x"74",
          3914 => x"7a",
          3915 => x"0c",
          3916 => x"04",
          3917 => x"79",
          3918 => x"05",
          3919 => x"57",
          3920 => x"81",
          3921 => x"56",
          3922 => x"08",
          3923 => x"91",
          3924 => x"75",
          3925 => x"90",
          3926 => x"81",
          3927 => x"06",
          3928 => x"87",
          3929 => x"2e",
          3930 => x"94",
          3931 => x"73",
          3932 => x"27",
          3933 => x"73",
          3934 => x"cb",
          3935 => x"88",
          3936 => x"76",
          3937 => x"3f",
          3938 => x"08",
          3939 => x"0c",
          3940 => x"39",
          3941 => x"52",
          3942 => x"bf",
          3943 => x"cb",
          3944 => x"2e",
          3945 => x"83",
          3946 => x"81",
          3947 => x"81",
          3948 => x"06",
          3949 => x"56",
          3950 => x"a0",
          3951 => x"81",
          3952 => x"98",
          3953 => x"94",
          3954 => x"08",
          3955 => x"a4",
          3956 => x"51",
          3957 => x"81",
          3958 => x"56",
          3959 => x"8c",
          3960 => x"17",
          3961 => x"07",
          3962 => x"18",
          3963 => x"2e",
          3964 => x"91",
          3965 => x"55",
          3966 => x"a4",
          3967 => x"0d",
          3968 => x"0d",
          3969 => x"3d",
          3970 => x"52",
          3971 => x"da",
          3972 => x"cb",
          3973 => x"81",
          3974 => x"81",
          3975 => x"45",
          3976 => x"52",
          3977 => x"52",
          3978 => x"3f",
          3979 => x"08",
          3980 => x"a4",
          3981 => x"38",
          3982 => x"05",
          3983 => x"2a",
          3984 => x"51",
          3985 => x"55",
          3986 => x"38",
          3987 => x"54",
          3988 => x"81",
          3989 => x"80",
          3990 => x"70",
          3991 => x"54",
          3992 => x"81",
          3993 => x"52",
          3994 => x"c5",
          3995 => x"a4",
          3996 => x"2a",
          3997 => x"51",
          3998 => x"80",
          3999 => x"38",
          4000 => x"cb",
          4001 => x"15",
          4002 => x"86",
          4003 => x"81",
          4004 => x"5c",
          4005 => x"3d",
          4006 => x"c7",
          4007 => x"cb",
          4008 => x"81",
          4009 => x"80",
          4010 => x"cb",
          4011 => x"73",
          4012 => x"3f",
          4013 => x"08",
          4014 => x"a4",
          4015 => x"87",
          4016 => x"39",
          4017 => x"08",
          4018 => x"38",
          4019 => x"08",
          4020 => x"77",
          4021 => x"3f",
          4022 => x"08",
          4023 => x"08",
          4024 => x"cb",
          4025 => x"80",
          4026 => x"55",
          4027 => x"94",
          4028 => x"2e",
          4029 => x"53",
          4030 => x"51",
          4031 => x"81",
          4032 => x"55",
          4033 => x"78",
          4034 => x"fe",
          4035 => x"a4",
          4036 => x"81",
          4037 => x"a0",
          4038 => x"e9",
          4039 => x"53",
          4040 => x"05",
          4041 => x"51",
          4042 => x"81",
          4043 => x"54",
          4044 => x"08",
          4045 => x"78",
          4046 => x"8e",
          4047 => x"58",
          4048 => x"81",
          4049 => x"54",
          4050 => x"08",
          4051 => x"54",
          4052 => x"81",
          4053 => x"84",
          4054 => x"06",
          4055 => x"02",
          4056 => x"33",
          4057 => x"81",
          4058 => x"86",
          4059 => x"f6",
          4060 => x"74",
          4061 => x"70",
          4062 => x"c3",
          4063 => x"a4",
          4064 => x"56",
          4065 => x"08",
          4066 => x"54",
          4067 => x"08",
          4068 => x"81",
          4069 => x"82",
          4070 => x"a4",
          4071 => x"09",
          4072 => x"38",
          4073 => x"b4",
          4074 => x"b0",
          4075 => x"a4",
          4076 => x"51",
          4077 => x"81",
          4078 => x"54",
          4079 => x"08",
          4080 => x"8b",
          4081 => x"b4",
          4082 => x"b7",
          4083 => x"54",
          4084 => x"15",
          4085 => x"90",
          4086 => x"34",
          4087 => x"0a",
          4088 => x"19",
          4089 => x"9f",
          4090 => x"78",
          4091 => x"51",
          4092 => x"a0",
          4093 => x"11",
          4094 => x"05",
          4095 => x"b6",
          4096 => x"ae",
          4097 => x"15",
          4098 => x"78",
          4099 => x"53",
          4100 => x"3f",
          4101 => x"0b",
          4102 => x"77",
          4103 => x"3f",
          4104 => x"08",
          4105 => x"a4",
          4106 => x"82",
          4107 => x"52",
          4108 => x"51",
          4109 => x"3f",
          4110 => x"52",
          4111 => x"aa",
          4112 => x"90",
          4113 => x"34",
          4114 => x"0b",
          4115 => x"78",
          4116 => x"b6",
          4117 => x"a4",
          4118 => x"39",
          4119 => x"52",
          4120 => x"be",
          4121 => x"81",
          4122 => x"99",
          4123 => x"da",
          4124 => x"3d",
          4125 => x"d2",
          4126 => x"53",
          4127 => x"84",
          4128 => x"3d",
          4129 => x"3f",
          4130 => x"08",
          4131 => x"a4",
          4132 => x"38",
          4133 => x"3d",
          4134 => x"3d",
          4135 => x"cc",
          4136 => x"cb",
          4137 => x"81",
          4138 => x"82",
          4139 => x"81",
          4140 => x"81",
          4141 => x"86",
          4142 => x"aa",
          4143 => x"a4",
          4144 => x"a8",
          4145 => x"05",
          4146 => x"ea",
          4147 => x"77",
          4148 => x"70",
          4149 => x"b4",
          4150 => x"3d",
          4151 => x"51",
          4152 => x"81",
          4153 => x"55",
          4154 => x"08",
          4155 => x"6f",
          4156 => x"06",
          4157 => x"a2",
          4158 => x"92",
          4159 => x"81",
          4160 => x"cb",
          4161 => x"2e",
          4162 => x"81",
          4163 => x"51",
          4164 => x"81",
          4165 => x"55",
          4166 => x"08",
          4167 => x"68",
          4168 => x"a8",
          4169 => x"05",
          4170 => x"51",
          4171 => x"3f",
          4172 => x"33",
          4173 => x"8b",
          4174 => x"84",
          4175 => x"06",
          4176 => x"73",
          4177 => x"a0",
          4178 => x"8b",
          4179 => x"54",
          4180 => x"15",
          4181 => x"33",
          4182 => x"70",
          4183 => x"55",
          4184 => x"2e",
          4185 => x"6e",
          4186 => x"df",
          4187 => x"78",
          4188 => x"3f",
          4189 => x"08",
          4190 => x"ff",
          4191 => x"82",
          4192 => x"a4",
          4193 => x"80",
          4194 => x"cb",
          4195 => x"78",
          4196 => x"af",
          4197 => x"a4",
          4198 => x"d4",
          4199 => x"55",
          4200 => x"08",
          4201 => x"81",
          4202 => x"73",
          4203 => x"81",
          4204 => x"63",
          4205 => x"76",
          4206 => x"3f",
          4207 => x"0b",
          4208 => x"87",
          4209 => x"a4",
          4210 => x"77",
          4211 => x"3f",
          4212 => x"08",
          4213 => x"a4",
          4214 => x"78",
          4215 => x"aa",
          4216 => x"a4",
          4217 => x"81",
          4218 => x"a8",
          4219 => x"ed",
          4220 => x"80",
          4221 => x"02",
          4222 => x"df",
          4223 => x"57",
          4224 => x"3d",
          4225 => x"96",
          4226 => x"e9",
          4227 => x"a4",
          4228 => x"cb",
          4229 => x"cf",
          4230 => x"65",
          4231 => x"d4",
          4232 => x"b5",
          4233 => x"a4",
          4234 => x"cb",
          4235 => x"38",
          4236 => x"05",
          4237 => x"06",
          4238 => x"73",
          4239 => x"a7",
          4240 => x"09",
          4241 => x"71",
          4242 => x"06",
          4243 => x"55",
          4244 => x"15",
          4245 => x"81",
          4246 => x"34",
          4247 => x"b4",
          4248 => x"cb",
          4249 => x"74",
          4250 => x"0c",
          4251 => x"04",
          4252 => x"64",
          4253 => x"93",
          4254 => x"52",
          4255 => x"d1",
          4256 => x"cb",
          4257 => x"81",
          4258 => x"80",
          4259 => x"58",
          4260 => x"3d",
          4261 => x"c8",
          4262 => x"cb",
          4263 => x"81",
          4264 => x"b4",
          4265 => x"c7",
          4266 => x"a0",
          4267 => x"55",
          4268 => x"84",
          4269 => x"17",
          4270 => x"2b",
          4271 => x"96",
          4272 => x"b0",
          4273 => x"54",
          4274 => x"15",
          4275 => x"ff",
          4276 => x"81",
          4277 => x"55",
          4278 => x"a4",
          4279 => x"0d",
          4280 => x"0d",
          4281 => x"5a",
          4282 => x"3d",
          4283 => x"99",
          4284 => x"81",
          4285 => x"a4",
          4286 => x"a4",
          4287 => x"81",
          4288 => x"07",
          4289 => x"55",
          4290 => x"2e",
          4291 => x"81",
          4292 => x"55",
          4293 => x"2e",
          4294 => x"7b",
          4295 => x"80",
          4296 => x"70",
          4297 => x"be",
          4298 => x"cb",
          4299 => x"81",
          4300 => x"80",
          4301 => x"52",
          4302 => x"dc",
          4303 => x"a4",
          4304 => x"cb",
          4305 => x"38",
          4306 => x"08",
          4307 => x"08",
          4308 => x"56",
          4309 => x"19",
          4310 => x"59",
          4311 => x"74",
          4312 => x"56",
          4313 => x"ec",
          4314 => x"75",
          4315 => x"74",
          4316 => x"2e",
          4317 => x"16",
          4318 => x"33",
          4319 => x"73",
          4320 => x"38",
          4321 => x"84",
          4322 => x"06",
          4323 => x"7a",
          4324 => x"76",
          4325 => x"07",
          4326 => x"54",
          4327 => x"80",
          4328 => x"80",
          4329 => x"7b",
          4330 => x"53",
          4331 => x"93",
          4332 => x"a4",
          4333 => x"cb",
          4334 => x"38",
          4335 => x"55",
          4336 => x"56",
          4337 => x"8b",
          4338 => x"56",
          4339 => x"83",
          4340 => x"75",
          4341 => x"51",
          4342 => x"3f",
          4343 => x"08",
          4344 => x"81",
          4345 => x"98",
          4346 => x"e6",
          4347 => x"53",
          4348 => x"b8",
          4349 => x"3d",
          4350 => x"3f",
          4351 => x"08",
          4352 => x"08",
          4353 => x"cb",
          4354 => x"98",
          4355 => x"a0",
          4356 => x"70",
          4357 => x"ae",
          4358 => x"6d",
          4359 => x"81",
          4360 => x"57",
          4361 => x"74",
          4362 => x"38",
          4363 => x"81",
          4364 => x"81",
          4365 => x"52",
          4366 => x"89",
          4367 => x"a4",
          4368 => x"a5",
          4369 => x"33",
          4370 => x"54",
          4371 => x"3f",
          4372 => x"08",
          4373 => x"38",
          4374 => x"76",
          4375 => x"05",
          4376 => x"39",
          4377 => x"08",
          4378 => x"15",
          4379 => x"ff",
          4380 => x"73",
          4381 => x"38",
          4382 => x"83",
          4383 => x"56",
          4384 => x"75",
          4385 => x"81",
          4386 => x"33",
          4387 => x"2e",
          4388 => x"52",
          4389 => x"51",
          4390 => x"3f",
          4391 => x"08",
          4392 => x"ff",
          4393 => x"38",
          4394 => x"88",
          4395 => x"8a",
          4396 => x"38",
          4397 => x"ec",
          4398 => x"75",
          4399 => x"74",
          4400 => x"73",
          4401 => x"05",
          4402 => x"17",
          4403 => x"70",
          4404 => x"34",
          4405 => x"70",
          4406 => x"ff",
          4407 => x"55",
          4408 => x"26",
          4409 => x"8b",
          4410 => x"86",
          4411 => x"e5",
          4412 => x"38",
          4413 => x"99",
          4414 => x"05",
          4415 => x"70",
          4416 => x"73",
          4417 => x"81",
          4418 => x"ff",
          4419 => x"ed",
          4420 => x"80",
          4421 => x"91",
          4422 => x"55",
          4423 => x"3f",
          4424 => x"08",
          4425 => x"a4",
          4426 => x"38",
          4427 => x"51",
          4428 => x"3f",
          4429 => x"08",
          4430 => x"a4",
          4431 => x"76",
          4432 => x"67",
          4433 => x"34",
          4434 => x"81",
          4435 => x"84",
          4436 => x"06",
          4437 => x"80",
          4438 => x"2e",
          4439 => x"81",
          4440 => x"ff",
          4441 => x"81",
          4442 => x"54",
          4443 => x"08",
          4444 => x"53",
          4445 => x"08",
          4446 => x"ff",
          4447 => x"67",
          4448 => x"8b",
          4449 => x"53",
          4450 => x"51",
          4451 => x"3f",
          4452 => x"0b",
          4453 => x"79",
          4454 => x"ee",
          4455 => x"a4",
          4456 => x"55",
          4457 => x"a4",
          4458 => x"0d",
          4459 => x"0d",
          4460 => x"88",
          4461 => x"05",
          4462 => x"fc",
          4463 => x"54",
          4464 => x"d2",
          4465 => x"cb",
          4466 => x"81",
          4467 => x"82",
          4468 => x"1a",
          4469 => x"82",
          4470 => x"80",
          4471 => x"8c",
          4472 => x"78",
          4473 => x"1a",
          4474 => x"2a",
          4475 => x"51",
          4476 => x"90",
          4477 => x"82",
          4478 => x"58",
          4479 => x"81",
          4480 => x"39",
          4481 => x"22",
          4482 => x"70",
          4483 => x"56",
          4484 => x"82",
          4485 => x"14",
          4486 => x"30",
          4487 => x"9f",
          4488 => x"a4",
          4489 => x"19",
          4490 => x"5a",
          4491 => x"81",
          4492 => x"38",
          4493 => x"77",
          4494 => x"82",
          4495 => x"56",
          4496 => x"74",
          4497 => x"ff",
          4498 => x"81",
          4499 => x"55",
          4500 => x"75",
          4501 => x"82",
          4502 => x"a4",
          4503 => x"ff",
          4504 => x"cb",
          4505 => x"2e",
          4506 => x"81",
          4507 => x"8e",
          4508 => x"56",
          4509 => x"09",
          4510 => x"38",
          4511 => x"59",
          4512 => x"77",
          4513 => x"06",
          4514 => x"87",
          4515 => x"39",
          4516 => x"ba",
          4517 => x"55",
          4518 => x"2e",
          4519 => x"15",
          4520 => x"2e",
          4521 => x"83",
          4522 => x"75",
          4523 => x"7e",
          4524 => x"a8",
          4525 => x"a4",
          4526 => x"cb",
          4527 => x"ce",
          4528 => x"16",
          4529 => x"56",
          4530 => x"38",
          4531 => x"19",
          4532 => x"8c",
          4533 => x"7d",
          4534 => x"38",
          4535 => x"0c",
          4536 => x"0c",
          4537 => x"80",
          4538 => x"73",
          4539 => x"98",
          4540 => x"05",
          4541 => x"57",
          4542 => x"26",
          4543 => x"7b",
          4544 => x"0c",
          4545 => x"81",
          4546 => x"84",
          4547 => x"54",
          4548 => x"a4",
          4549 => x"0d",
          4550 => x"0d",
          4551 => x"88",
          4552 => x"05",
          4553 => x"54",
          4554 => x"c5",
          4555 => x"56",
          4556 => x"cb",
          4557 => x"8b",
          4558 => x"cb",
          4559 => x"29",
          4560 => x"05",
          4561 => x"55",
          4562 => x"84",
          4563 => x"34",
          4564 => x"08",
          4565 => x"5f",
          4566 => x"51",
          4567 => x"3f",
          4568 => x"08",
          4569 => x"70",
          4570 => x"57",
          4571 => x"8b",
          4572 => x"82",
          4573 => x"06",
          4574 => x"56",
          4575 => x"38",
          4576 => x"05",
          4577 => x"7e",
          4578 => x"f0",
          4579 => x"a4",
          4580 => x"67",
          4581 => x"2e",
          4582 => x"82",
          4583 => x"8b",
          4584 => x"75",
          4585 => x"80",
          4586 => x"81",
          4587 => x"2e",
          4588 => x"80",
          4589 => x"38",
          4590 => x"0a",
          4591 => x"ff",
          4592 => x"55",
          4593 => x"86",
          4594 => x"8a",
          4595 => x"89",
          4596 => x"2a",
          4597 => x"77",
          4598 => x"59",
          4599 => x"81",
          4600 => x"70",
          4601 => x"07",
          4602 => x"56",
          4603 => x"38",
          4604 => x"05",
          4605 => x"7e",
          4606 => x"80",
          4607 => x"81",
          4608 => x"8a",
          4609 => x"83",
          4610 => x"06",
          4611 => x"08",
          4612 => x"74",
          4613 => x"41",
          4614 => x"56",
          4615 => x"8a",
          4616 => x"61",
          4617 => x"55",
          4618 => x"27",
          4619 => x"93",
          4620 => x"80",
          4621 => x"38",
          4622 => x"70",
          4623 => x"43",
          4624 => x"95",
          4625 => x"06",
          4626 => x"2e",
          4627 => x"77",
          4628 => x"74",
          4629 => x"83",
          4630 => x"06",
          4631 => x"82",
          4632 => x"2e",
          4633 => x"78",
          4634 => x"2e",
          4635 => x"80",
          4636 => x"ae",
          4637 => x"2a",
          4638 => x"81",
          4639 => x"56",
          4640 => x"2e",
          4641 => x"77",
          4642 => x"81",
          4643 => x"79",
          4644 => x"70",
          4645 => x"5a",
          4646 => x"86",
          4647 => x"27",
          4648 => x"52",
          4649 => x"fc",
          4650 => x"cb",
          4651 => x"29",
          4652 => x"70",
          4653 => x"55",
          4654 => x"0b",
          4655 => x"08",
          4656 => x"05",
          4657 => x"ff",
          4658 => x"27",
          4659 => x"88",
          4660 => x"ae",
          4661 => x"2a",
          4662 => x"81",
          4663 => x"56",
          4664 => x"2e",
          4665 => x"77",
          4666 => x"81",
          4667 => x"79",
          4668 => x"70",
          4669 => x"5a",
          4670 => x"86",
          4671 => x"27",
          4672 => x"52",
          4673 => x"fc",
          4674 => x"cb",
          4675 => x"84",
          4676 => x"cb",
          4677 => x"f5",
          4678 => x"81",
          4679 => x"a4",
          4680 => x"cb",
          4681 => x"71",
          4682 => x"83",
          4683 => x"5e",
          4684 => x"89",
          4685 => x"5c",
          4686 => x"1c",
          4687 => x"05",
          4688 => x"ff",
          4689 => x"70",
          4690 => x"31",
          4691 => x"57",
          4692 => x"83",
          4693 => x"06",
          4694 => x"1c",
          4695 => x"5c",
          4696 => x"1d",
          4697 => x"29",
          4698 => x"31",
          4699 => x"55",
          4700 => x"87",
          4701 => x"7c",
          4702 => x"7a",
          4703 => x"31",
          4704 => x"fb",
          4705 => x"cb",
          4706 => x"7d",
          4707 => x"81",
          4708 => x"81",
          4709 => x"83",
          4710 => x"80",
          4711 => x"87",
          4712 => x"81",
          4713 => x"fd",
          4714 => x"f8",
          4715 => x"2e",
          4716 => x"80",
          4717 => x"ff",
          4718 => x"cb",
          4719 => x"a0",
          4720 => x"38",
          4721 => x"74",
          4722 => x"86",
          4723 => x"fd",
          4724 => x"81",
          4725 => x"80",
          4726 => x"83",
          4727 => x"39",
          4728 => x"08",
          4729 => x"92",
          4730 => x"b8",
          4731 => x"59",
          4732 => x"27",
          4733 => x"86",
          4734 => x"55",
          4735 => x"09",
          4736 => x"38",
          4737 => x"f5",
          4738 => x"38",
          4739 => x"55",
          4740 => x"86",
          4741 => x"80",
          4742 => x"7a",
          4743 => x"b9",
          4744 => x"81",
          4745 => x"7a",
          4746 => x"8a",
          4747 => x"52",
          4748 => x"ff",
          4749 => x"79",
          4750 => x"7b",
          4751 => x"06",
          4752 => x"51",
          4753 => x"3f",
          4754 => x"1c",
          4755 => x"32",
          4756 => x"96",
          4757 => x"06",
          4758 => x"91",
          4759 => x"a1",
          4760 => x"55",
          4761 => x"ff",
          4762 => x"74",
          4763 => x"06",
          4764 => x"51",
          4765 => x"3f",
          4766 => x"52",
          4767 => x"ff",
          4768 => x"f8",
          4769 => x"34",
          4770 => x"1b",
          4771 => x"d9",
          4772 => x"52",
          4773 => x"ff",
          4774 => x"60",
          4775 => x"51",
          4776 => x"3f",
          4777 => x"09",
          4778 => x"cb",
          4779 => x"b2",
          4780 => x"c3",
          4781 => x"a0",
          4782 => x"52",
          4783 => x"ff",
          4784 => x"82",
          4785 => x"51",
          4786 => x"3f",
          4787 => x"1b",
          4788 => x"95",
          4789 => x"b2",
          4790 => x"a0",
          4791 => x"80",
          4792 => x"1c",
          4793 => x"80",
          4794 => x"93",
          4795 => x"c8",
          4796 => x"1b",
          4797 => x"82",
          4798 => x"52",
          4799 => x"ff",
          4800 => x"7c",
          4801 => x"06",
          4802 => x"51",
          4803 => x"3f",
          4804 => x"a4",
          4805 => x"0b",
          4806 => x"93",
          4807 => x"dc",
          4808 => x"51",
          4809 => x"3f",
          4810 => x"52",
          4811 => x"70",
          4812 => x"9f",
          4813 => x"54",
          4814 => x"52",
          4815 => x"9b",
          4816 => x"56",
          4817 => x"08",
          4818 => x"7d",
          4819 => x"81",
          4820 => x"38",
          4821 => x"86",
          4822 => x"52",
          4823 => x"9b",
          4824 => x"80",
          4825 => x"7a",
          4826 => x"ed",
          4827 => x"85",
          4828 => x"7a",
          4829 => x"8f",
          4830 => x"85",
          4831 => x"83",
          4832 => x"ff",
          4833 => x"ff",
          4834 => x"e8",
          4835 => x"9e",
          4836 => x"52",
          4837 => x"51",
          4838 => x"3f",
          4839 => x"52",
          4840 => x"9e",
          4841 => x"54",
          4842 => x"53",
          4843 => x"51",
          4844 => x"3f",
          4845 => x"16",
          4846 => x"7e",
          4847 => x"d8",
          4848 => x"80",
          4849 => x"ff",
          4850 => x"7f",
          4851 => x"7d",
          4852 => x"81",
          4853 => x"f8",
          4854 => x"ff",
          4855 => x"ff",
          4856 => x"51",
          4857 => x"3f",
          4858 => x"88",
          4859 => x"39",
          4860 => x"f8",
          4861 => x"2e",
          4862 => x"55",
          4863 => x"51",
          4864 => x"3f",
          4865 => x"57",
          4866 => x"83",
          4867 => x"76",
          4868 => x"7a",
          4869 => x"ff",
          4870 => x"81",
          4871 => x"82",
          4872 => x"80",
          4873 => x"a4",
          4874 => x"51",
          4875 => x"3f",
          4876 => x"78",
          4877 => x"74",
          4878 => x"18",
          4879 => x"2e",
          4880 => x"79",
          4881 => x"2e",
          4882 => x"55",
          4883 => x"62",
          4884 => x"74",
          4885 => x"75",
          4886 => x"7e",
          4887 => x"b8",
          4888 => x"a4",
          4889 => x"38",
          4890 => x"78",
          4891 => x"74",
          4892 => x"56",
          4893 => x"93",
          4894 => x"66",
          4895 => x"26",
          4896 => x"56",
          4897 => x"83",
          4898 => x"64",
          4899 => x"77",
          4900 => x"84",
          4901 => x"52",
          4902 => x"9d",
          4903 => x"d4",
          4904 => x"51",
          4905 => x"3f",
          4906 => x"55",
          4907 => x"81",
          4908 => x"34",
          4909 => x"16",
          4910 => x"16",
          4911 => x"16",
          4912 => x"05",
          4913 => x"c1",
          4914 => x"fe",
          4915 => x"fe",
          4916 => x"34",
          4917 => x"08",
          4918 => x"07",
          4919 => x"16",
          4920 => x"a4",
          4921 => x"34",
          4922 => x"c6",
          4923 => x"9c",
          4924 => x"52",
          4925 => x"51",
          4926 => x"3f",
          4927 => x"53",
          4928 => x"51",
          4929 => x"3f",
          4930 => x"cb",
          4931 => x"38",
          4932 => x"52",
          4933 => x"99",
          4934 => x"56",
          4935 => x"08",
          4936 => x"39",
          4937 => x"39",
          4938 => x"39",
          4939 => x"08",
          4940 => x"cb",
          4941 => x"3d",
          4942 => x"3d",
          4943 => x"71",
          4944 => x"8e",
          4945 => x"29",
          4946 => x"05",
          4947 => x"04",
          4948 => x"51",
          4949 => x"81",
          4950 => x"80",
          4951 => x"bd",
          4952 => x"f2",
          4953 => x"f0",
          4954 => x"39",
          4955 => x"51",
          4956 => x"81",
          4957 => x"80",
          4958 => x"be",
          4959 => x"d6",
          4960 => x"b4",
          4961 => x"39",
          4962 => x"51",
          4963 => x"81",
          4964 => x"80",
          4965 => x"be",
          4966 => x"39",
          4967 => x"51",
          4968 => x"bf",
          4969 => x"39",
          4970 => x"51",
          4971 => x"bf",
          4972 => x"39",
          4973 => x"51",
          4974 => x"c0",
          4975 => x"39",
          4976 => x"51",
          4977 => x"c0",
          4978 => x"39",
          4979 => x"51",
          4980 => x"c0",
          4981 => x"87",
          4982 => x"3d",
          4983 => x"3d",
          4984 => x"56",
          4985 => x"e7",
          4986 => x"74",
          4987 => x"e8",
          4988 => x"39",
          4989 => x"74",
          4990 => x"a3",
          4991 => x"a4",
          4992 => x"51",
          4993 => x"3f",
          4994 => x"08",
          4995 => x"75",
          4996 => x"84",
          4997 => x"a0",
          4998 => x"0d",
          4999 => x"0d",
          5000 => x"02",
          5001 => x"c7",
          5002 => x"73",
          5003 => x"5d",
          5004 => x"5c",
          5005 => x"81",
          5006 => x"ff",
          5007 => x"81",
          5008 => x"ff",
          5009 => x"80",
          5010 => x"27",
          5011 => x"79",
          5012 => x"38",
          5013 => x"a7",
          5014 => x"39",
          5015 => x"72",
          5016 => x"38",
          5017 => x"81",
          5018 => x"ff",
          5019 => x"89",
          5020 => x"c0",
          5021 => x"dc",
          5022 => x"55",
          5023 => x"74",
          5024 => x"78",
          5025 => x"72",
          5026 => x"c1",
          5027 => x"8c",
          5028 => x"39",
          5029 => x"51",
          5030 => x"3f",
          5031 => x"a1",
          5032 => x"53",
          5033 => x"8e",
          5034 => x"52",
          5035 => x"51",
          5036 => x"3f",
          5037 => x"c1",
          5038 => x"86",
          5039 => x"15",
          5040 => x"fe",
          5041 => x"ff",
          5042 => x"c1",
          5043 => x"86",
          5044 => x"55",
          5045 => x"aa",
          5046 => x"70",
          5047 => x"26",
          5048 => x"9f",
          5049 => x"38",
          5050 => x"8b",
          5051 => x"fe",
          5052 => x"73",
          5053 => x"a0",
          5054 => x"d7",
          5055 => x"55",
          5056 => x"c1",
          5057 => x"85",
          5058 => x"16",
          5059 => x"56",
          5060 => x"3f",
          5061 => x"08",
          5062 => x"98",
          5063 => x"74",
          5064 => x"81",
          5065 => x"fe",
          5066 => x"81",
          5067 => x"98",
          5068 => x"2c",
          5069 => x"70",
          5070 => x"07",
          5071 => x"56",
          5072 => x"74",
          5073 => x"38",
          5074 => x"74",
          5075 => x"81",
          5076 => x"80",
          5077 => x"7a",
          5078 => x"76",
          5079 => x"38",
          5080 => x"81",
          5081 => x"8d",
          5082 => x"ec",
          5083 => x"02",
          5084 => x"e3",
          5085 => x"72",
          5086 => x"07",
          5087 => x"87",
          5088 => x"07",
          5089 => x"5a",
          5090 => x"57",
          5091 => x"38",
          5092 => x"52",
          5093 => x"52",
          5094 => x"3f",
          5095 => x"08",
          5096 => x"a4",
          5097 => x"81",
          5098 => x"87",
          5099 => x"0c",
          5100 => x"08",
          5101 => x"d4",
          5102 => x"80",
          5103 => x"76",
          5104 => x"3f",
          5105 => x"08",
          5106 => x"a4",
          5107 => x"7a",
          5108 => x"2e",
          5109 => x"19",
          5110 => x"59",
          5111 => x"3d",
          5112 => x"cc",
          5113 => x"30",
          5114 => x"80",
          5115 => x"79",
          5116 => x"38",
          5117 => x"90",
          5118 => x"dc",
          5119 => x"98",
          5120 => x"78",
          5121 => x"3f",
          5122 => x"81",
          5123 => x"96",
          5124 => x"f9",
          5125 => x"02",
          5126 => x"05",
          5127 => x"ff",
          5128 => x"7a",
          5129 => x"fe",
          5130 => x"cb",
          5131 => x"38",
          5132 => x"88",
          5133 => x"2e",
          5134 => x"39",
          5135 => x"54",
          5136 => x"53",
          5137 => x"51",
          5138 => x"cb",
          5139 => x"83",
          5140 => x"76",
          5141 => x"0c",
          5142 => x"04",
          5143 => x"02",
          5144 => x"81",
          5145 => x"81",
          5146 => x"55",
          5147 => x"3f",
          5148 => x"22",
          5149 => x"e2",
          5150 => x"f8",
          5151 => x"84",
          5152 => x"b5",
          5153 => x"c2",
          5154 => x"88",
          5155 => x"80",
          5156 => x"fe",
          5157 => x"86",
          5158 => x"fe",
          5159 => x"c0",
          5160 => x"53",
          5161 => x"3f",
          5162 => x"f6",
          5163 => x"c2",
          5164 => x"f8",
          5165 => x"51",
          5166 => x"3f",
          5167 => x"70",
          5168 => x"52",
          5169 => x"95",
          5170 => x"fe",
          5171 => x"81",
          5172 => x"fe",
          5173 => x"80",
          5174 => x"dd",
          5175 => x"2a",
          5176 => x"51",
          5177 => x"2e",
          5178 => x"51",
          5179 => x"3f",
          5180 => x"51",
          5181 => x"3f",
          5182 => x"f5",
          5183 => x"83",
          5184 => x"06",
          5185 => x"80",
          5186 => x"81",
          5187 => x"a9",
          5188 => x"e8",
          5189 => x"a1",
          5190 => x"fe",
          5191 => x"72",
          5192 => x"81",
          5193 => x"71",
          5194 => x"38",
          5195 => x"f5",
          5196 => x"c2",
          5197 => x"f7",
          5198 => x"51",
          5199 => x"3f",
          5200 => x"70",
          5201 => x"52",
          5202 => x"95",
          5203 => x"fe",
          5204 => x"81",
          5205 => x"fe",
          5206 => x"80",
          5207 => x"d9",
          5208 => x"2a",
          5209 => x"51",
          5210 => x"2e",
          5211 => x"51",
          5212 => x"3f",
          5213 => x"51",
          5214 => x"3f",
          5215 => x"f4",
          5216 => x"87",
          5217 => x"06",
          5218 => x"80",
          5219 => x"81",
          5220 => x"a5",
          5221 => x"b8",
          5222 => x"9d",
          5223 => x"fe",
          5224 => x"72",
          5225 => x"81",
          5226 => x"71",
          5227 => x"38",
          5228 => x"f4",
          5229 => x"c3",
          5230 => x"f5",
          5231 => x"51",
          5232 => x"3f",
          5233 => x"3f",
          5234 => x"04",
          5235 => x"78",
          5236 => x"55",
          5237 => x"80",
          5238 => x"38",
          5239 => x"77",
          5240 => x"33",
          5241 => x"39",
          5242 => x"80",
          5243 => x"81",
          5244 => x"57",
          5245 => x"2e",
          5246 => x"53",
          5247 => x"84",
          5248 => x"38",
          5249 => x"06",
          5250 => x"2e",
          5251 => x"88",
          5252 => x"70",
          5253 => x"34",
          5254 => x"90",
          5255 => x"d4",
          5256 => x"53",
          5257 => x"55",
          5258 => x"3f",
          5259 => x"08",
          5260 => x"15",
          5261 => x"81",
          5262 => x"38",
          5263 => x"81",
          5264 => x"53",
          5265 => x"d2",
          5266 => x"72",
          5267 => x"0c",
          5268 => x"04",
          5269 => x"80",
          5270 => x"e2",
          5271 => x"5c",
          5272 => x"51",
          5273 => x"3f",
          5274 => x"08",
          5275 => x"59",
          5276 => x"09",
          5277 => x"38",
          5278 => x"52",
          5279 => x"52",
          5280 => x"ca",
          5281 => x"78",
          5282 => x"d4",
          5283 => x"e3",
          5284 => x"a4",
          5285 => x"88",
          5286 => x"90",
          5287 => x"39",
          5288 => x"5c",
          5289 => x"51",
          5290 => x"3f",
          5291 => x"46",
          5292 => x"53",
          5293 => x"51",
          5294 => x"3f",
          5295 => x"64",
          5296 => x"ce",
          5297 => x"fe",
          5298 => x"fd",
          5299 => x"cb",
          5300 => x"2b",
          5301 => x"51",
          5302 => x"c3",
          5303 => x"38",
          5304 => x"24",
          5305 => x"78",
          5306 => x"bc",
          5307 => x"24",
          5308 => x"82",
          5309 => x"38",
          5310 => x"8a",
          5311 => x"2e",
          5312 => x"8d",
          5313 => x"84",
          5314 => x"38",
          5315 => x"82",
          5316 => x"f9",
          5317 => x"c0",
          5318 => x"38",
          5319 => x"24",
          5320 => x"b0",
          5321 => x"38",
          5322 => x"84",
          5323 => x"dd",
          5324 => x"c1",
          5325 => x"38",
          5326 => x"2e",
          5327 => x"8c",
          5328 => x"80",
          5329 => x"ba",
          5330 => x"f8",
          5331 => x"78",
          5332 => x"8a",
          5333 => x"80",
          5334 => x"38",
          5335 => x"2e",
          5336 => x"8c",
          5337 => x"80",
          5338 => x"dc",
          5339 => x"d5",
          5340 => x"38",
          5341 => x"78",
          5342 => x"8b",
          5343 => x"81",
          5344 => x"38",
          5345 => x"2e",
          5346 => x"78",
          5347 => x"8b",
          5348 => x"f9",
          5349 => x"85",
          5350 => x"38",
          5351 => x"2e",
          5352 => x"8b",
          5353 => x"3d",
          5354 => x"53",
          5355 => x"51",
          5356 => x"3f",
          5357 => x"08",
          5358 => x"c4",
          5359 => x"c7",
          5360 => x"fe",
          5361 => x"fe",
          5362 => x"ff",
          5363 => x"81",
          5364 => x"80",
          5365 => x"81",
          5366 => x"38",
          5367 => x"80",
          5368 => x"52",
          5369 => x"05",
          5370 => x"87",
          5371 => x"cb",
          5372 => x"ff",
          5373 => x"8e",
          5374 => x"dc",
          5375 => x"d4",
          5376 => x"fd",
          5377 => x"c4",
          5378 => x"d2",
          5379 => x"fe",
          5380 => x"fe",
          5381 => x"ff",
          5382 => x"81",
          5383 => x"80",
          5384 => x"38",
          5385 => x"52",
          5386 => x"05",
          5387 => x"8b",
          5388 => x"cb",
          5389 => x"81",
          5390 => x"8a",
          5391 => x"3d",
          5392 => x"53",
          5393 => x"51",
          5394 => x"3f",
          5395 => x"08",
          5396 => x"38",
          5397 => x"fc",
          5398 => x"3d",
          5399 => x"53",
          5400 => x"51",
          5401 => x"3f",
          5402 => x"08",
          5403 => x"cb",
          5404 => x"63",
          5405 => x"8c",
          5406 => x"ff",
          5407 => x"02",
          5408 => x"33",
          5409 => x"63",
          5410 => x"81",
          5411 => x"51",
          5412 => x"3f",
          5413 => x"08",
          5414 => x"81",
          5415 => x"fe",
          5416 => x"81",
          5417 => x"39",
          5418 => x"f8",
          5419 => x"ea",
          5420 => x"cb",
          5421 => x"3d",
          5422 => x"52",
          5423 => x"8c",
          5424 => x"81",
          5425 => x"52",
          5426 => x"9f",
          5427 => x"39",
          5428 => x"f8",
          5429 => x"ea",
          5430 => x"cb",
          5431 => x"3d",
          5432 => x"52",
          5433 => x"e4",
          5434 => x"a4",
          5435 => x"fe",
          5436 => x"5a",
          5437 => x"3f",
          5438 => x"08",
          5439 => x"f8",
          5440 => x"fe",
          5441 => x"81",
          5442 => x"81",
          5443 => x"80",
          5444 => x"81",
          5445 => x"81",
          5446 => x"78",
          5447 => x"7a",
          5448 => x"3f",
          5449 => x"08",
          5450 => x"f8",
          5451 => x"a4",
          5452 => x"86",
          5453 => x"39",
          5454 => x"f4",
          5455 => x"f8",
          5456 => x"80",
          5457 => x"cb",
          5458 => x"2e",
          5459 => x"b7",
          5460 => x"11",
          5461 => x"05",
          5462 => x"d1",
          5463 => x"a4",
          5464 => x"fa",
          5465 => x"3d",
          5466 => x"53",
          5467 => x"51",
          5468 => x"3f",
          5469 => x"08",
          5470 => x"cb",
          5471 => x"81",
          5472 => x"fe",
          5473 => x"63",
          5474 => x"79",
          5475 => x"38",
          5476 => x"7a",
          5477 => x"5c",
          5478 => x"26",
          5479 => x"c4",
          5480 => x"ba",
          5481 => x"fe",
          5482 => x"fe",
          5483 => x"fe",
          5484 => x"81",
          5485 => x"80",
          5486 => x"c8",
          5487 => x"78",
          5488 => x"38",
          5489 => x"08",
          5490 => x"81",
          5491 => x"59",
          5492 => x"88",
          5493 => x"98",
          5494 => x"39",
          5495 => x"33",
          5496 => x"38",
          5497 => x"33",
          5498 => x"2e",
          5499 => x"c8",
          5500 => x"89",
          5501 => x"b0",
          5502 => x"05",
          5503 => x"fe",
          5504 => x"fe",
          5505 => x"fe",
          5506 => x"81",
          5507 => x"80",
          5508 => x"c8",
          5509 => x"78",
          5510 => x"38",
          5511 => x"08",
          5512 => x"81",
          5513 => x"59",
          5514 => x"88",
          5515 => x"9c",
          5516 => x"39",
          5517 => x"33",
          5518 => x"38",
          5519 => x"33",
          5520 => x"2e",
          5521 => x"c8",
          5522 => x"88",
          5523 => x"b0",
          5524 => x"43",
          5525 => x"ec",
          5526 => x"f8",
          5527 => x"fe",
          5528 => x"cb",
          5529 => x"2e",
          5530 => x"62",
          5531 => x"88",
          5532 => x"81",
          5533 => x"2e",
          5534 => x"80",
          5535 => x"79",
          5536 => x"38",
          5537 => x"c5",
          5538 => x"f6",
          5539 => x"55",
          5540 => x"53",
          5541 => x"51",
          5542 => x"81",
          5543 => x"84",
          5544 => x"3d",
          5545 => x"53",
          5546 => x"51",
          5547 => x"3f",
          5548 => x"08",
          5549 => x"ec",
          5550 => x"fe",
          5551 => x"fe",
          5552 => x"fe",
          5553 => x"81",
          5554 => x"80",
          5555 => x"63",
          5556 => x"cb",
          5557 => x"34",
          5558 => x"44",
          5559 => x"f0",
          5560 => x"f8",
          5561 => x"fd",
          5562 => x"cb",
          5563 => x"38",
          5564 => x"63",
          5565 => x"52",
          5566 => x"51",
          5567 => x"3f",
          5568 => x"79",
          5569 => x"8a",
          5570 => x"79",
          5571 => x"ae",
          5572 => x"38",
          5573 => x"a0",
          5574 => x"fe",
          5575 => x"fe",
          5576 => x"fe",
          5577 => x"81",
          5578 => x"80",
          5579 => x"63",
          5580 => x"cb",
          5581 => x"34",
          5582 => x"44",
          5583 => x"81",
          5584 => x"fe",
          5585 => x"ff",
          5586 => x"3d",
          5587 => x"53",
          5588 => x"51",
          5589 => x"3f",
          5590 => x"08",
          5591 => x"c4",
          5592 => x"fe",
          5593 => x"fe",
          5594 => x"fe",
          5595 => x"81",
          5596 => x"80",
          5597 => x"60",
          5598 => x"05",
          5599 => x"82",
          5600 => x"78",
          5601 => x"fe",
          5602 => x"fe",
          5603 => x"fe",
          5604 => x"81",
          5605 => x"df",
          5606 => x"39",
          5607 => x"54",
          5608 => x"cc",
          5609 => x"90",
          5610 => x"52",
          5611 => x"fa",
          5612 => x"45",
          5613 => x"78",
          5614 => x"e8",
          5615 => x"26",
          5616 => x"84",
          5617 => x"39",
          5618 => x"e4",
          5619 => x"f8",
          5620 => x"fd",
          5621 => x"cb",
          5622 => x"2e",
          5623 => x"59",
          5624 => x"22",
          5625 => x"05",
          5626 => x"41",
          5627 => x"81",
          5628 => x"fe",
          5629 => x"ff",
          5630 => x"3d",
          5631 => x"53",
          5632 => x"51",
          5633 => x"3f",
          5634 => x"08",
          5635 => x"94",
          5636 => x"fe",
          5637 => x"fe",
          5638 => x"fe",
          5639 => x"81",
          5640 => x"80",
          5641 => x"60",
          5642 => x"59",
          5643 => x"41",
          5644 => x"e4",
          5645 => x"f8",
          5646 => x"fc",
          5647 => x"cb",
          5648 => x"38",
          5649 => x"60",
          5650 => x"52",
          5651 => x"51",
          5652 => x"3f",
          5653 => x"79",
          5654 => x"b6",
          5655 => x"79",
          5656 => x"ae",
          5657 => x"38",
          5658 => x"a8",
          5659 => x"fe",
          5660 => x"fe",
          5661 => x"fe",
          5662 => x"81",
          5663 => x"80",
          5664 => x"7f",
          5665 => x"81",
          5666 => x"fe",
          5667 => x"60",
          5668 => x"59",
          5669 => x"41",
          5670 => x"81",
          5671 => x"fe",
          5672 => x"ff",
          5673 => x"c5",
          5674 => x"f2",
          5675 => x"51",
          5676 => x"3f",
          5677 => x"81",
          5678 => x"fe",
          5679 => x"a2",
          5680 => x"e8",
          5681 => x"39",
          5682 => x"0b",
          5683 => x"84",
          5684 => x"81",
          5685 => x"94",
          5686 => x"c6",
          5687 => x"f1",
          5688 => x"c0",
          5689 => x"a8",
          5690 => x"e8",
          5691 => x"83",
          5692 => x"94",
          5693 => x"80",
          5694 => x"c0",
          5695 => x"f3",
          5696 => x"3d",
          5697 => x"53",
          5698 => x"51",
          5699 => x"3f",
          5700 => x"08",
          5701 => x"8c",
          5702 => x"81",
          5703 => x"fe",
          5704 => x"63",
          5705 => x"b7",
          5706 => x"11",
          5707 => x"05",
          5708 => x"f9",
          5709 => x"a4",
          5710 => x"f2",
          5711 => x"52",
          5712 => x"51",
          5713 => x"3f",
          5714 => x"2d",
          5715 => x"08",
          5716 => x"a4",
          5717 => x"f2",
          5718 => x"cb",
          5719 => x"81",
          5720 => x"fe",
          5721 => x"f2",
          5722 => x"c7",
          5723 => x"f0",
          5724 => x"cd",
          5725 => x"ac",
          5726 => x"ac",
          5727 => x"d4",
          5728 => x"ff",
          5729 => x"ec",
          5730 => x"98",
          5731 => x"33",
          5732 => x"80",
          5733 => x"38",
          5734 => x"80",
          5735 => x"80",
          5736 => x"38",
          5737 => x"f8",
          5738 => x"e0",
          5739 => x"c7",
          5740 => x"cb",
          5741 => x"81",
          5742 => x"80",
          5743 => x"c8",
          5744 => x"70",
          5745 => x"f6",
          5746 => x"c8",
          5747 => x"cb",
          5748 => x"56",
          5749 => x"46",
          5750 => x"80",
          5751 => x"80",
          5752 => x"80",
          5753 => x"ec",
          5754 => x"cb",
          5755 => x"7c",
          5756 => x"81",
          5757 => x"78",
          5758 => x"ff",
          5759 => x"06",
          5760 => x"81",
          5761 => x"fe",
          5762 => x"f1",
          5763 => x"3d",
          5764 => x"81",
          5765 => x"b6",
          5766 => x"0b",
          5767 => x"8c",
          5768 => x"8d",
          5769 => x"c0",
          5770 => x"8c",
          5771 => x"87",
          5772 => x"0c",
          5773 => x"0b",
          5774 => x"94",
          5775 => x"0b",
          5776 => x"0c",
          5777 => x"81",
          5778 => x"fe",
          5779 => x"fe",
          5780 => x"81",
          5781 => x"fe",
          5782 => x"81",
          5783 => x"fe",
          5784 => x"81",
          5785 => x"fe",
          5786 => x"81",
          5787 => x"3f",
          5788 => x"80",
          5789 => x"00",
          5790 => x"00",
          5791 => x"00",
          5792 => x"00",
          5793 => x"00",
          5794 => x"00",
          5795 => x"00",
          5796 => x"00",
          5797 => x"00",
          5798 => x"00",
          5799 => x"00",
          5800 => x"00",
          5801 => x"00",
          5802 => x"00",
          5803 => x"00",
          5804 => x"00",
          5805 => x"00",
          5806 => x"00",
          5807 => x"00",
          5808 => x"00",
          5809 => x"00",
          5810 => x"00",
          5811 => x"00",
          5812 => x"00",
          5813 => x"00",
          5814 => x"64",
          5815 => x"2f",
          5816 => x"25",
          5817 => x"64",
          5818 => x"2e",
          5819 => x"64",
          5820 => x"6f",
          5821 => x"6f",
          5822 => x"67",
          5823 => x"74",
          5824 => x"00",
          5825 => x"28",
          5826 => x"6d",
          5827 => x"43",
          5828 => x"6e",
          5829 => x"29",
          5830 => x"0a",
          5831 => x"69",
          5832 => x"20",
          5833 => x"6c",
          5834 => x"6e",
          5835 => x"3a",
          5836 => x"20",
          5837 => x"4e",
          5838 => x"42",
          5839 => x"20",
          5840 => x"61",
          5841 => x"25",
          5842 => x"2c",
          5843 => x"7a",
          5844 => x"30",
          5845 => x"2e",
          5846 => x"20",
          5847 => x"52",
          5848 => x"28",
          5849 => x"72",
          5850 => x"30",
          5851 => x"20",
          5852 => x"65",
          5853 => x"38",
          5854 => x"0a",
          5855 => x"20",
          5856 => x"41",
          5857 => x"53",
          5858 => x"74",
          5859 => x"38",
          5860 => x"53",
          5861 => x"3d",
          5862 => x"58",
          5863 => x"00",
          5864 => x"20",
          5865 => x"4f",
          5866 => x"0a",
          5867 => x"20",
          5868 => x"53",
          5869 => x"00",
          5870 => x"20",
          5871 => x"50",
          5872 => x"00",
          5873 => x"20",
          5874 => x"44",
          5875 => x"72",
          5876 => x"44",
          5877 => x"63",
          5878 => x"25",
          5879 => x"29",
          5880 => x"00",
          5881 => x"20",
          5882 => x"4e",
          5883 => x"52",
          5884 => x"20",
          5885 => x"54",
          5886 => x"4c",
          5887 => x"00",
          5888 => x"20",
          5889 => x"49",
          5890 => x"31",
          5891 => x"69",
          5892 => x"73",
          5893 => x"31",
          5894 => x"0a",
          5895 => x"64",
          5896 => x"73",
          5897 => x"3a",
          5898 => x"20",
          5899 => x"50",
          5900 => x"65",
          5901 => x"20",
          5902 => x"74",
          5903 => x"41",
          5904 => x"65",
          5905 => x"3d",
          5906 => x"38",
          5907 => x"00",
          5908 => x"20",
          5909 => x"50",
          5910 => x"65",
          5911 => x"79",
          5912 => x"61",
          5913 => x"41",
          5914 => x"65",
          5915 => x"3d",
          5916 => x"38",
          5917 => x"00",
          5918 => x"20",
          5919 => x"74",
          5920 => x"20",
          5921 => x"72",
          5922 => x"64",
          5923 => x"73",
          5924 => x"20",
          5925 => x"3d",
          5926 => x"38",
          5927 => x"00",
          5928 => x"20",
          5929 => x"50",
          5930 => x"64",
          5931 => x"20",
          5932 => x"20",
          5933 => x"20",
          5934 => x"20",
          5935 => x"3d",
          5936 => x"38",
          5937 => x"00",
          5938 => x"20",
          5939 => x"79",
          5940 => x"6d",
          5941 => x"6f",
          5942 => x"46",
          5943 => x"20",
          5944 => x"20",
          5945 => x"3d",
          5946 => x"38",
          5947 => x"00",
          5948 => x"6d",
          5949 => x"00",
          5950 => x"65",
          5951 => x"6d",
          5952 => x"6c",
          5953 => x"00",
          5954 => x"56",
          5955 => x"56",
          5956 => x"6e",
          5957 => x"6e",
          5958 => x"77",
          5959 => x"44",
          5960 => x"2a",
          5961 => x"3b",
          5962 => x"3f",
          5963 => x"7f",
          5964 => x"41",
          5965 => x"41",
          5966 => x"00",
          5967 => x"fe",
          5968 => x"44",
          5969 => x"2e",
          5970 => x"4f",
          5971 => x"4d",
          5972 => x"20",
          5973 => x"54",
          5974 => x"20",
          5975 => x"4f",
          5976 => x"4d",
          5977 => x"20",
          5978 => x"54",
          5979 => x"20",
          5980 => x"00",
          5981 => x"00",
          5982 => x"00",
          5983 => x"00",
          5984 => x"9a",
          5985 => x"41",
          5986 => x"45",
          5987 => x"49",
          5988 => x"92",
          5989 => x"4f",
          5990 => x"99",
          5991 => x"9d",
          5992 => x"49",
          5993 => x"a5",
          5994 => x"a9",
          5995 => x"ad",
          5996 => x"b1",
          5997 => x"b5",
          5998 => x"b9",
          5999 => x"bd",
          6000 => x"c1",
          6001 => x"c5",
          6002 => x"c9",
          6003 => x"cd",
          6004 => x"d1",
          6005 => x"d5",
          6006 => x"d9",
          6007 => x"dd",
          6008 => x"e1",
          6009 => x"e5",
          6010 => x"e9",
          6011 => x"ed",
          6012 => x"f1",
          6013 => x"f5",
          6014 => x"f9",
          6015 => x"fd",
          6016 => x"2e",
          6017 => x"5b",
          6018 => x"22",
          6019 => x"3e",
          6020 => x"00",
          6021 => x"01",
          6022 => x"10",
          6023 => x"00",
          6024 => x"00",
          6025 => x"01",
          6026 => x"04",
          6027 => x"10",
          6028 => x"00",
          6029 => x"69",
          6030 => x"00",
          6031 => x"69",
          6032 => x"6c",
          6033 => x"69",
          6034 => x"00",
          6035 => x"6c",
          6036 => x"00",
          6037 => x"65",
          6038 => x"00",
          6039 => x"63",
          6040 => x"72",
          6041 => x"64",
          6042 => x"00",
          6043 => x"74",
          6044 => x"00",
          6045 => x"65",
          6046 => x"65",
          6047 => x"65",
          6048 => x"69",
          6049 => x"69",
          6050 => x"66",
          6051 => x"66",
          6052 => x"61",
          6053 => x"00",
          6054 => x"6d",
          6055 => x"65",
          6056 => x"72",
          6057 => x"65",
          6058 => x"00",
          6059 => x"6e",
          6060 => x"00",
          6061 => x"65",
          6062 => x"00",
          6063 => x"69",
          6064 => x"45",
          6065 => x"72",
          6066 => x"6e",
          6067 => x"6e",
          6068 => x"65",
          6069 => x"72",
          6070 => x"00",
          6071 => x"69",
          6072 => x"6e",
          6073 => x"72",
          6074 => x"79",
          6075 => x"00",
          6076 => x"6f",
          6077 => x"6c",
          6078 => x"6f",
          6079 => x"2e",
          6080 => x"6f",
          6081 => x"74",
          6082 => x"6f",
          6083 => x"2e",
          6084 => x"6e",
          6085 => x"69",
          6086 => x"69",
          6087 => x"61",
          6088 => x"0a",
          6089 => x"63",
          6090 => x"73",
          6091 => x"6e",
          6092 => x"2e",
          6093 => x"69",
          6094 => x"61",
          6095 => x"61",
          6096 => x"65",
          6097 => x"74",
          6098 => x"00",
          6099 => x"69",
          6100 => x"68",
          6101 => x"6c",
          6102 => x"6e",
          6103 => x"69",
          6104 => x"00",
          6105 => x"44",
          6106 => x"20",
          6107 => x"74",
          6108 => x"72",
          6109 => x"63",
          6110 => x"2e",
          6111 => x"72",
          6112 => x"20",
          6113 => x"62",
          6114 => x"69",
          6115 => x"6e",
          6116 => x"69",
          6117 => x"00",
          6118 => x"69",
          6119 => x"6e",
          6120 => x"65",
          6121 => x"6c",
          6122 => x"0a",
          6123 => x"6f",
          6124 => x"6d",
          6125 => x"69",
          6126 => x"20",
          6127 => x"65",
          6128 => x"74",
          6129 => x"66",
          6130 => x"64",
          6131 => x"20",
          6132 => x"6b",
          6133 => x"00",
          6134 => x"6f",
          6135 => x"74",
          6136 => x"6f",
          6137 => x"64",
          6138 => x"00",
          6139 => x"69",
          6140 => x"75",
          6141 => x"6f",
          6142 => x"61",
          6143 => x"6e",
          6144 => x"6e",
          6145 => x"6c",
          6146 => x"0a",
          6147 => x"69",
          6148 => x"69",
          6149 => x"6f",
          6150 => x"64",
          6151 => x"00",
          6152 => x"6e",
          6153 => x"66",
          6154 => x"65",
          6155 => x"6d",
          6156 => x"72",
          6157 => x"00",
          6158 => x"6f",
          6159 => x"61",
          6160 => x"6f",
          6161 => x"20",
          6162 => x"65",
          6163 => x"00",
          6164 => x"61",
          6165 => x"65",
          6166 => x"73",
          6167 => x"63",
          6168 => x"65",
          6169 => x"0a",
          6170 => x"75",
          6171 => x"73",
          6172 => x"00",
          6173 => x"6e",
          6174 => x"77",
          6175 => x"72",
          6176 => x"2e",
          6177 => x"25",
          6178 => x"62",
          6179 => x"73",
          6180 => x"20",
          6181 => x"25",
          6182 => x"62",
          6183 => x"73",
          6184 => x"63",
          6185 => x"00",
          6186 => x"30",
          6187 => x"00",
          6188 => x"20",
          6189 => x"30",
          6190 => x"00",
          6191 => x"20",
          6192 => x"20",
          6193 => x"00",
          6194 => x"30",
          6195 => x"00",
          6196 => x"20",
          6197 => x"7c",
          6198 => x"0d",
          6199 => x"65",
          6200 => x"00",
          6201 => x"50",
          6202 => x"00",
          6203 => x"2a",
          6204 => x"73",
          6205 => x"00",
          6206 => x"38",
          6207 => x"2f",
          6208 => x"39",
          6209 => x"31",
          6210 => x"00",
          6211 => x"5a",
          6212 => x"20",
          6213 => x"20",
          6214 => x"78",
          6215 => x"73",
          6216 => x"20",
          6217 => x"0a",
          6218 => x"50",
          6219 => x"20",
          6220 => x"65",
          6221 => x"70",
          6222 => x"61",
          6223 => x"65",
          6224 => x"00",
          6225 => x"69",
          6226 => x"20",
          6227 => x"65",
          6228 => x"70",
          6229 => x"00",
          6230 => x"53",
          6231 => x"6e",
          6232 => x"72",
          6233 => x"0a",
          6234 => x"4f",
          6235 => x"20",
          6236 => x"69",
          6237 => x"72",
          6238 => x"74",
          6239 => x"4f",
          6240 => x"20",
          6241 => x"69",
          6242 => x"72",
          6243 => x"74",
          6244 => x"41",
          6245 => x"20",
          6246 => x"69",
          6247 => x"72",
          6248 => x"74",
          6249 => x"41",
          6250 => x"20",
          6251 => x"69",
          6252 => x"72",
          6253 => x"74",
          6254 => x"41",
          6255 => x"20",
          6256 => x"69",
          6257 => x"72",
          6258 => x"74",
          6259 => x"41",
          6260 => x"20",
          6261 => x"69",
          6262 => x"72",
          6263 => x"74",
          6264 => x"65",
          6265 => x"6e",
          6266 => x"70",
          6267 => x"6d",
          6268 => x"2e",
          6269 => x"00",
          6270 => x"6e",
          6271 => x"69",
          6272 => x"74",
          6273 => x"72",
          6274 => x"0a",
          6275 => x"3a",
          6276 => x"61",
          6277 => x"64",
          6278 => x"20",
          6279 => x"74",
          6280 => x"69",
          6281 => x"73",
          6282 => x"61",
          6283 => x"30",
          6284 => x"6c",
          6285 => x"65",
          6286 => x"69",
          6287 => x"61",
          6288 => x"6c",
          6289 => x"0a",
          6290 => x"20",
          6291 => x"61",
          6292 => x"69",
          6293 => x"69",
          6294 => x"00",
          6295 => x"6e",
          6296 => x"61",
          6297 => x"65",
          6298 => x"00",
          6299 => x"61",
          6300 => x"64",
          6301 => x"20",
          6302 => x"74",
          6303 => x"69",
          6304 => x"0a",
          6305 => x"63",
          6306 => x"0a",
          6307 => x"75",
          6308 => x"6c",
          6309 => x"69",
          6310 => x"2e",
          6311 => x"75",
          6312 => x"4d",
          6313 => x"72",
          6314 => x"00",
          6315 => x"43",
          6316 => x"6c",
          6317 => x"2e",
          6318 => x"30",
          6319 => x"25",
          6320 => x"2d",
          6321 => x"3f",
          6322 => x"00",
          6323 => x"30",
          6324 => x"25",
          6325 => x"2d",
          6326 => x"30",
          6327 => x"25",
          6328 => x"2d",
          6329 => x"69",
          6330 => x"6c",
          6331 => x"20",
          6332 => x"65",
          6333 => x"70",
          6334 => x"00",
          6335 => x"6e",
          6336 => x"69",
          6337 => x"69",
          6338 => x"72",
          6339 => x"74",
          6340 => x"00",
          6341 => x"69",
          6342 => x"6c",
          6343 => x"75",
          6344 => x"20",
          6345 => x"6f",
          6346 => x"6e",
          6347 => x"69",
          6348 => x"75",
          6349 => x"20",
          6350 => x"6f",
          6351 => x"78",
          6352 => x"74",
          6353 => x"20",
          6354 => x"65",
          6355 => x"25",
          6356 => x"20",
          6357 => x"0a",
          6358 => x"61",
          6359 => x"6e",
          6360 => x"6f",
          6361 => x"40",
          6362 => x"38",
          6363 => x"2e",
          6364 => x"00",
          6365 => x"61",
          6366 => x"72",
          6367 => x"72",
          6368 => x"20",
          6369 => x"65",
          6370 => x"64",
          6371 => x"00",
          6372 => x"65",
          6373 => x"72",
          6374 => x"67",
          6375 => x"70",
          6376 => x"61",
          6377 => x"6e",
          6378 => x"0a",
          6379 => x"6f",
          6380 => x"72",
          6381 => x"6f",
          6382 => x"67",
          6383 => x"0a",
          6384 => x"50",
          6385 => x"69",
          6386 => x"64",
          6387 => x"73",
          6388 => x"2e",
          6389 => x"00",
          6390 => x"61",
          6391 => x"6f",
          6392 => x"6e",
          6393 => x"00",
          6394 => x"75",
          6395 => x"6e",
          6396 => x"2e",
          6397 => x"6e",
          6398 => x"69",
          6399 => x"69",
          6400 => x"72",
          6401 => x"74",
          6402 => x"2e",
          6403 => x"00",
          6404 => x"00",
          6405 => x"00",
          6406 => x"00",
          6407 => x"00",
          6408 => x"01",
          6409 => x"00",
          6410 => x"00",
          6411 => x"00",
          6412 => x"00",
          6413 => x"00",
          6414 => x"f5",
          6415 => x"01",
          6416 => x"01",
          6417 => x"01",
          6418 => x"00",
          6419 => x"00",
          6420 => x"00",
          6421 => x"00",
          6422 => x"02",
          6423 => x"00",
          6424 => x"00",
          6425 => x"00",
          6426 => x"04",
          6427 => x"00",
          6428 => x"00",
          6429 => x"00",
          6430 => x"14",
          6431 => x"00",
          6432 => x"00",
          6433 => x"00",
          6434 => x"2b",
          6435 => x"00",
          6436 => x"00",
          6437 => x"00",
          6438 => x"30",
          6439 => x"00",
          6440 => x"00",
          6441 => x"00",
          6442 => x"3c",
          6443 => x"00",
          6444 => x"00",
          6445 => x"00",
          6446 => x"40",
          6447 => x"00",
          6448 => x"00",
          6449 => x"00",
          6450 => x"44",
          6451 => x"00",
          6452 => x"00",
          6453 => x"00",
          6454 => x"41",
          6455 => x"00",
          6456 => x"00",
          6457 => x"00",
          6458 => x"42",
          6459 => x"00",
          6460 => x"00",
          6461 => x"00",
          6462 => x"43",
          6463 => x"00",
          6464 => x"00",
          6465 => x"00",
          6466 => x"50",
          6467 => x"00",
          6468 => x"00",
          6469 => x"00",
          6470 => x"51",
          6471 => x"00",
          6472 => x"00",
          6473 => x"00",
          6474 => x"54",
          6475 => x"00",
          6476 => x"00",
          6477 => x"00",
          6478 => x"55",
          6479 => x"00",
          6480 => x"00",
          6481 => x"00",
          6482 => x"79",
          6483 => x"00",
          6484 => x"00",
          6485 => x"00",
          6486 => x"78",
          6487 => x"00",
          6488 => x"00",
          6489 => x"00",
          6490 => x"82",
          6491 => x"00",
          6492 => x"00",
          6493 => x"00",
          6494 => x"83",
          6495 => x"00",
          6496 => x"00",
          6497 => x"00",
          6498 => x"85",
          6499 => x"00",
          6500 => x"00",
          6501 => x"00",
          6502 => x"87",
          6503 => x"00",
          6504 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"80",
             2 => x"0b",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"80",
            10 => x"0b",
            11 => x"0b",
            12 => x"93",
            13 => x"0b",
            14 => x"0b",
            15 => x"b1",
            16 => x"0b",
            17 => x"0b",
            18 => x"cf",
            19 => x"0b",
            20 => x"0b",
            21 => x"ed",
            22 => x"0b",
            23 => x"0b",
            24 => x"8b",
            25 => x"0b",
            26 => x"0b",
            27 => x"a9",
            28 => x"0b",
            29 => x"0b",
            30 => x"c7",
            31 => x"0b",
            32 => x"0b",
            33 => x"e5",
            34 => x"0b",
            35 => x"0b",
            36 => x"83",
            37 => x"0b",
            38 => x"0b",
            39 => x"a3",
            40 => x"0b",
            41 => x"0b",
            42 => x"c3",
            43 => x"0b",
            44 => x"0b",
            45 => x"e3",
            46 => x"0b",
            47 => x"0b",
            48 => x"83",
            49 => x"0b",
            50 => x"0b",
            51 => x"a3",
            52 => x"0b",
            53 => x"0b",
            54 => x"c3",
            55 => x"0b",
            56 => x"0b",
            57 => x"e3",
            58 => x"0b",
            59 => x"0b",
            60 => x"83",
            61 => x"0b",
            62 => x"0b",
            63 => x"a3",
            64 => x"0b",
            65 => x"0b",
            66 => x"c3",
            67 => x"0b",
            68 => x"0b",
            69 => x"e3",
            70 => x"0b",
            71 => x"0b",
            72 => x"83",
            73 => x"0b",
            74 => x"0b",
            75 => x"a2",
            76 => x"0b",
            77 => x"0b",
            78 => x"c0",
            79 => x"0b",
            80 => x"0b",
            81 => x"de",
            82 => x"0b",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"00",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"00",
           137 => x"00",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"00",
           145 => x"00",
           146 => x"00",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"00",
           153 => x"00",
           154 => x"00",
           155 => x"00",
           156 => x"00",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"00",
           161 => x"00",
           162 => x"00",
           163 => x"00",
           164 => x"00",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"00",
           169 => x"00",
           170 => x"00",
           171 => x"00",
           172 => x"00",
           173 => x"00",
           174 => x"00",
           175 => x"00",
           176 => x"00",
           177 => x"00",
           178 => x"00",
           179 => x"00",
           180 => x"00",
           181 => x"00",
           182 => x"00",
           183 => x"00",
           184 => x"00",
           185 => x"00",
           186 => x"00",
           187 => x"00",
           188 => x"00",
           189 => x"00",
           190 => x"00",
           191 => x"00",
           192 => x"00",
           193 => x"00",
           194 => x"00",
           195 => x"00",
           196 => x"00",
           197 => x"00",
           198 => x"00",
           199 => x"00",
           200 => x"00",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"00",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"00",
           233 => x"00",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"00",
           249 => x"00",
           250 => x"00",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"81",
           258 => x"98",
           259 => x"cb",
           260 => x"e4",
           261 => x"cb",
           262 => x"f5",
           263 => x"b0",
           264 => x"90",
           265 => x"b0",
           266 => x"2d",
           267 => x"08",
           268 => x"04",
           269 => x"0c",
           270 => x"81",
           271 => x"81",
           272 => x"81",
           273 => x"aa",
           274 => x"cb",
           275 => x"e4",
           276 => x"cb",
           277 => x"8e",
           278 => x"b0",
           279 => x"90",
           280 => x"b0",
           281 => x"2d",
           282 => x"08",
           283 => x"04",
           284 => x"0c",
           285 => x"81",
           286 => x"81",
           287 => x"81",
           288 => x"ad",
           289 => x"cb",
           290 => x"e4",
           291 => x"cb",
           292 => x"b6",
           293 => x"b0",
           294 => x"90",
           295 => x"b0",
           296 => x"2d",
           297 => x"08",
           298 => x"04",
           299 => x"0c",
           300 => x"81",
           301 => x"81",
           302 => x"81",
           303 => x"9a",
           304 => x"cb",
           305 => x"e4",
           306 => x"cb",
           307 => x"a3",
           308 => x"b0",
           309 => x"90",
           310 => x"b0",
           311 => x"2d",
           312 => x"08",
           313 => x"04",
           314 => x"0c",
           315 => x"81",
           316 => x"81",
           317 => x"81",
           318 => x"96",
           319 => x"cb",
           320 => x"e4",
           321 => x"cb",
           322 => x"df",
           323 => x"cb",
           324 => x"e4",
           325 => x"cb",
           326 => x"ec",
           327 => x"cb",
           328 => x"e4",
           329 => x"cb",
           330 => x"e4",
           331 => x"cb",
           332 => x"e4",
           333 => x"cb",
           334 => x"e7",
           335 => x"cb",
           336 => x"e4",
           337 => x"cb",
           338 => x"f1",
           339 => x"cb",
           340 => x"e4",
           341 => x"cb",
           342 => x"fa",
           343 => x"cb",
           344 => x"e4",
           345 => x"cb",
           346 => x"eb",
           347 => x"cb",
           348 => x"e4",
           349 => x"cb",
           350 => x"f4",
           351 => x"cb",
           352 => x"e4",
           353 => x"cb",
           354 => x"f6",
           355 => x"cb",
           356 => x"e4",
           357 => x"cb",
           358 => x"f6",
           359 => x"cb",
           360 => x"e4",
           361 => x"cb",
           362 => x"fe",
           363 => x"cb",
           364 => x"e4",
           365 => x"cb",
           366 => x"fb",
           367 => x"cb",
           368 => x"e4",
           369 => x"cb",
           370 => x"80",
           371 => x"cb",
           372 => x"e4",
           373 => x"cb",
           374 => x"f7",
           375 => x"cb",
           376 => x"e4",
           377 => x"cb",
           378 => x"83",
           379 => x"cb",
           380 => x"e4",
           381 => x"cb",
           382 => x"84",
           383 => x"cb",
           384 => x"e4",
           385 => x"cb",
           386 => x"ed",
           387 => x"cb",
           388 => x"e4",
           389 => x"cb",
           390 => x"ec",
           391 => x"cb",
           392 => x"e4",
           393 => x"cb",
           394 => x"ee",
           395 => x"cb",
           396 => x"e4",
           397 => x"cb",
           398 => x"f8",
           399 => x"cb",
           400 => x"e4",
           401 => x"cb",
           402 => x"85",
           403 => x"cb",
           404 => x"e4",
           405 => x"cb",
           406 => x"87",
           407 => x"cb",
           408 => x"e4",
           409 => x"cb",
           410 => x"8b",
           411 => x"cb",
           412 => x"e4",
           413 => x"cb",
           414 => x"de",
           415 => x"cb",
           416 => x"e4",
           417 => x"cb",
           418 => x"8e",
           419 => x"cb",
           420 => x"e4",
           421 => x"cb",
           422 => x"ac",
           423 => x"b0",
           424 => x"90",
           425 => x"b0",
           426 => x"2d",
           427 => x"08",
           428 => x"04",
           429 => x"0c",
           430 => x"81",
           431 => x"81",
           432 => x"81",
           433 => x"93",
           434 => x"cb",
           435 => x"e4",
           436 => x"cb",
           437 => x"ca",
           438 => x"b0",
           439 => x"90",
           440 => x"b0",
           441 => x"2d",
           442 => x"08",
           443 => x"04",
           444 => x"0c",
           445 => x"2d",
           446 => x"08",
           447 => x"04",
           448 => x"70",
           449 => x"27",
           450 => x"71",
           451 => x"53",
           452 => x"0b",
           453 => x"88",
           454 => x"b4",
           455 => x"04",
           456 => x"08",
           457 => x"b0",
           458 => x"0d",
           459 => x"cb",
           460 => x"05",
           461 => x"cb",
           462 => x"05",
           463 => x"c5",
           464 => x"a4",
           465 => x"cb",
           466 => x"85",
           467 => x"cb",
           468 => x"81",
           469 => x"02",
           470 => x"0c",
           471 => x"81",
           472 => x"b0",
           473 => x"08",
           474 => x"b0",
           475 => x"08",
           476 => x"81",
           477 => x"70",
           478 => x"0c",
           479 => x"0d",
           480 => x"0c",
           481 => x"b0",
           482 => x"cb",
           483 => x"3d",
           484 => x"81",
           485 => x"fc",
           486 => x"0b",
           487 => x"08",
           488 => x"81",
           489 => x"8c",
           490 => x"cb",
           491 => x"05",
           492 => x"38",
           493 => x"08",
           494 => x"80",
           495 => x"80",
           496 => x"b0",
           497 => x"08",
           498 => x"81",
           499 => x"8c",
           500 => x"81",
           501 => x"8c",
           502 => x"cb",
           503 => x"05",
           504 => x"cb",
           505 => x"05",
           506 => x"39",
           507 => x"08",
           508 => x"80",
           509 => x"38",
           510 => x"08",
           511 => x"81",
           512 => x"88",
           513 => x"ad",
           514 => x"b0",
           515 => x"08",
           516 => x"08",
           517 => x"31",
           518 => x"08",
           519 => x"81",
           520 => x"f8",
           521 => x"cb",
           522 => x"05",
           523 => x"cb",
           524 => x"05",
           525 => x"b0",
           526 => x"08",
           527 => x"cb",
           528 => x"05",
           529 => x"b0",
           530 => x"08",
           531 => x"cb",
           532 => x"05",
           533 => x"39",
           534 => x"08",
           535 => x"80",
           536 => x"81",
           537 => x"88",
           538 => x"81",
           539 => x"f4",
           540 => x"91",
           541 => x"b0",
           542 => x"08",
           543 => x"b0",
           544 => x"0c",
           545 => x"b0",
           546 => x"08",
           547 => x"0c",
           548 => x"81",
           549 => x"04",
           550 => x"76",
           551 => x"8c",
           552 => x"33",
           553 => x"55",
           554 => x"8a",
           555 => x"06",
           556 => x"2e",
           557 => x"12",
           558 => x"2e",
           559 => x"73",
           560 => x"55",
           561 => x"52",
           562 => x"09",
           563 => x"38",
           564 => x"a4",
           565 => x"0d",
           566 => x"88",
           567 => x"70",
           568 => x"07",
           569 => x"8f",
           570 => x"38",
           571 => x"84",
           572 => x"72",
           573 => x"05",
           574 => x"71",
           575 => x"53",
           576 => x"70",
           577 => x"0c",
           578 => x"71",
           579 => x"38",
           580 => x"90",
           581 => x"70",
           582 => x"0c",
           583 => x"71",
           584 => x"38",
           585 => x"8e",
           586 => x"0d",
           587 => x"72",
           588 => x"53",
           589 => x"93",
           590 => x"73",
           591 => x"54",
           592 => x"2e",
           593 => x"73",
           594 => x"71",
           595 => x"ff",
           596 => x"70",
           597 => x"38",
           598 => x"70",
           599 => x"81",
           600 => x"81",
           601 => x"71",
           602 => x"ff",
           603 => x"54",
           604 => x"38",
           605 => x"73",
           606 => x"75",
           607 => x"71",
           608 => x"cb",
           609 => x"52",
           610 => x"04",
           611 => x"f7",
           612 => x"14",
           613 => x"84",
           614 => x"06",
           615 => x"70",
           616 => x"14",
           617 => x"08",
           618 => x"71",
           619 => x"dc",
           620 => x"54",
           621 => x"39",
           622 => x"cb",
           623 => x"3d",
           624 => x"3d",
           625 => x"83",
           626 => x"2b",
           627 => x"3f",
           628 => x"08",
           629 => x"72",
           630 => x"54",
           631 => x"25",
           632 => x"81",
           633 => x"84",
           634 => x"fb",
           635 => x"70",
           636 => x"53",
           637 => x"2e",
           638 => x"71",
           639 => x"a0",
           640 => x"06",
           641 => x"12",
           642 => x"71",
           643 => x"81",
           644 => x"73",
           645 => x"ff",
           646 => x"55",
           647 => x"83",
           648 => x"70",
           649 => x"38",
           650 => x"73",
           651 => x"51",
           652 => x"09",
           653 => x"38",
           654 => x"81",
           655 => x"72",
           656 => x"51",
           657 => x"a4",
           658 => x"0d",
           659 => x"0d",
           660 => x"08",
           661 => x"38",
           662 => x"05",
           663 => x"98",
           664 => x"cb",
           665 => x"38",
           666 => x"39",
           667 => x"81",
           668 => x"86",
           669 => x"fc",
           670 => x"82",
           671 => x"05",
           672 => x"52",
           673 => x"81",
           674 => x"13",
           675 => x"51",
           676 => x"9e",
           677 => x"38",
           678 => x"51",
           679 => x"97",
           680 => x"38",
           681 => x"51",
           682 => x"bb",
           683 => x"38",
           684 => x"51",
           685 => x"bb",
           686 => x"38",
           687 => x"55",
           688 => x"87",
           689 => x"d9",
           690 => x"22",
           691 => x"73",
           692 => x"80",
           693 => x"0b",
           694 => x"9c",
           695 => x"87",
           696 => x"0c",
           697 => x"87",
           698 => x"0c",
           699 => x"87",
           700 => x"0c",
           701 => x"87",
           702 => x"0c",
           703 => x"87",
           704 => x"0c",
           705 => x"87",
           706 => x"0c",
           707 => x"98",
           708 => x"87",
           709 => x"0c",
           710 => x"c0",
           711 => x"80",
           712 => x"cb",
           713 => x"3d",
           714 => x"3d",
           715 => x"87",
           716 => x"5d",
           717 => x"87",
           718 => x"08",
           719 => x"23",
           720 => x"b8",
           721 => x"82",
           722 => x"c0",
           723 => x"5a",
           724 => x"34",
           725 => x"b0",
           726 => x"84",
           727 => x"c0",
           728 => x"5a",
           729 => x"34",
           730 => x"a8",
           731 => x"86",
           732 => x"c0",
           733 => x"5c",
           734 => x"23",
           735 => x"a0",
           736 => x"8a",
           737 => x"7d",
           738 => x"ff",
           739 => x"7b",
           740 => x"06",
           741 => x"33",
           742 => x"33",
           743 => x"33",
           744 => x"33",
           745 => x"33",
           746 => x"ff",
           747 => x"81",
           748 => x"92",
           749 => x"3d",
           750 => x"3d",
           751 => x"05",
           752 => x"70",
           753 => x"52",
           754 => x"0b",
           755 => x"34",
           756 => x"04",
           757 => x"77",
           758 => x"c8",
           759 => x"81",
           760 => x"55",
           761 => x"94",
           762 => x"80",
           763 => x"87",
           764 => x"51",
           765 => x"96",
           766 => x"06",
           767 => x"70",
           768 => x"38",
           769 => x"70",
           770 => x"51",
           771 => x"72",
           772 => x"81",
           773 => x"70",
           774 => x"38",
           775 => x"70",
           776 => x"51",
           777 => x"38",
           778 => x"06",
           779 => x"94",
           780 => x"80",
           781 => x"87",
           782 => x"52",
           783 => x"75",
           784 => x"0c",
           785 => x"04",
           786 => x"02",
           787 => x"0b",
           788 => x"8c",
           789 => x"ff",
           790 => x"56",
           791 => x"84",
           792 => x"2e",
           793 => x"c0",
           794 => x"70",
           795 => x"2a",
           796 => x"53",
           797 => x"80",
           798 => x"71",
           799 => x"81",
           800 => x"70",
           801 => x"81",
           802 => x"06",
           803 => x"80",
           804 => x"71",
           805 => x"81",
           806 => x"70",
           807 => x"73",
           808 => x"51",
           809 => x"80",
           810 => x"2e",
           811 => x"c0",
           812 => x"75",
           813 => x"3d",
           814 => x"3d",
           815 => x"80",
           816 => x"81",
           817 => x"53",
           818 => x"2e",
           819 => x"71",
           820 => x"81",
           821 => x"81",
           822 => x"70",
           823 => x"59",
           824 => x"87",
           825 => x"51",
           826 => x"86",
           827 => x"94",
           828 => x"08",
           829 => x"70",
           830 => x"54",
           831 => x"2e",
           832 => x"91",
           833 => x"06",
           834 => x"d7",
           835 => x"32",
           836 => x"51",
           837 => x"2e",
           838 => x"93",
           839 => x"06",
           840 => x"ff",
           841 => x"81",
           842 => x"87",
           843 => x"52",
           844 => x"86",
           845 => x"94",
           846 => x"72",
           847 => x"74",
           848 => x"ff",
           849 => x"57",
           850 => x"38",
           851 => x"a4",
           852 => x"0d",
           853 => x"0d",
           854 => x"c8",
           855 => x"81",
           856 => x"52",
           857 => x"84",
           858 => x"2e",
           859 => x"c0",
           860 => x"70",
           861 => x"2a",
           862 => x"51",
           863 => x"80",
           864 => x"71",
           865 => x"51",
           866 => x"80",
           867 => x"2e",
           868 => x"c0",
           869 => x"71",
           870 => x"ff",
           871 => x"a4",
           872 => x"3d",
           873 => x"3d",
           874 => x"81",
           875 => x"70",
           876 => x"52",
           877 => x"94",
           878 => x"80",
           879 => x"87",
           880 => x"52",
           881 => x"82",
           882 => x"06",
           883 => x"ff",
           884 => x"2e",
           885 => x"81",
           886 => x"87",
           887 => x"52",
           888 => x"86",
           889 => x"94",
           890 => x"08",
           891 => x"70",
           892 => x"53",
           893 => x"cb",
           894 => x"3d",
           895 => x"3d",
           896 => x"9e",
           897 => x"9c",
           898 => x"51",
           899 => x"2e",
           900 => x"87",
           901 => x"08",
           902 => x"0c",
           903 => x"a0",
           904 => x"94",
           905 => x"9e",
           906 => x"c8",
           907 => x"c0",
           908 => x"81",
           909 => x"87",
           910 => x"08",
           911 => x"0c",
           912 => x"98",
           913 => x"a4",
           914 => x"9e",
           915 => x"c8",
           916 => x"c0",
           917 => x"81",
           918 => x"87",
           919 => x"08",
           920 => x"0c",
           921 => x"80",
           922 => x"81",
           923 => x"87",
           924 => x"08",
           925 => x"0c",
           926 => x"c8",
           927 => x"0b",
           928 => x"88",
           929 => x"80",
           930 => x"52",
           931 => x"83",
           932 => x"71",
           933 => x"34",
           934 => x"c0",
           935 => x"70",
           936 => x"06",
           937 => x"70",
           938 => x"38",
           939 => x"81",
           940 => x"80",
           941 => x"9e",
           942 => x"80",
           943 => x"51",
           944 => x"80",
           945 => x"81",
           946 => x"c8",
           947 => x"0b",
           948 => x"88",
           949 => x"80",
           950 => x"52",
           951 => x"83",
           952 => x"71",
           953 => x"34",
           954 => x"c0",
           955 => x"70",
           956 => x"51",
           957 => x"80",
           958 => x"81",
           959 => x"c8",
           960 => x"0b",
           961 => x"88",
           962 => x"80",
           963 => x"52",
           964 => x"83",
           965 => x"71",
           966 => x"34",
           967 => x"c0",
           968 => x"70",
           969 => x"51",
           970 => x"80",
           971 => x"81",
           972 => x"c8",
           973 => x"0b",
           974 => x"88",
           975 => x"80",
           976 => x"52",
           977 => x"83",
           978 => x"71",
           979 => x"34",
           980 => x"88",
           981 => x"e0",
           982 => x"2c",
           983 => x"70",
           984 => x"34",
           985 => x"c0",
           986 => x"70",
           987 => x"52",
           988 => x"2e",
           989 => x"52",
           990 => x"c6",
           991 => x"87",
           992 => x"08",
           993 => x"51",
           994 => x"80",
           995 => x"81",
           996 => x"c8",
           997 => x"c0",
           998 => x"70",
           999 => x"51",
          1000 => x"c8",
          1001 => x"0d",
          1002 => x"0d",
          1003 => x"51",
          1004 => x"81",
          1005 => x"54",
          1006 => x"88",
          1007 => x"84",
          1008 => x"3f",
          1009 => x"51",
          1010 => x"81",
          1011 => x"54",
          1012 => x"92",
          1013 => x"94",
          1014 => x"c8",
          1015 => x"81",
          1016 => x"89",
          1017 => x"c8",
          1018 => x"73",
          1019 => x"38",
          1020 => x"08",
          1021 => x"98",
          1022 => x"b6",
          1023 => x"b9",
          1024 => x"bf",
          1025 => x"8b",
          1026 => x"c0",
          1027 => x"80",
          1028 => x"81",
          1029 => x"53",
          1030 => x"08",
          1031 => x"fc",
          1032 => x"3f",
          1033 => x"33",
          1034 => x"2e",
          1035 => x"b7",
          1036 => x"a1",
          1037 => x"c2",
          1038 => x"80",
          1039 => x"81",
          1040 => x"83",
          1041 => x"c8",
          1042 => x"73",
          1043 => x"38",
          1044 => x"51",
          1045 => x"81",
          1046 => x"54",
          1047 => x"8d",
          1048 => x"c5",
          1049 => x"b7",
          1050 => x"cd",
          1051 => x"c6",
          1052 => x"80",
          1053 => x"81",
          1054 => x"82",
          1055 => x"c8",
          1056 => x"73",
          1057 => x"38",
          1058 => x"33",
          1059 => x"80",
          1060 => x"3f",
          1061 => x"51",
          1062 => x"81",
          1063 => x"52",
          1064 => x"51",
          1065 => x"81",
          1066 => x"52",
          1067 => x"51",
          1068 => x"81",
          1069 => x"52",
          1070 => x"51",
          1071 => x"81",
          1072 => x"52",
          1073 => x"51",
          1074 => x"81",
          1075 => x"52",
          1076 => x"51",
          1077 => x"85",
          1078 => x"fe",
          1079 => x"92",
          1080 => x"05",
          1081 => x"26",
          1082 => x"84",
          1083 => x"81",
          1084 => x"52",
          1085 => x"81",
          1086 => x"9d",
          1087 => x"f8",
          1088 => x"81",
          1089 => x"91",
          1090 => x"88",
          1091 => x"81",
          1092 => x"85",
          1093 => x"94",
          1094 => x"3f",
          1095 => x"04",
          1096 => x"0c",
          1097 => x"87",
          1098 => x"0c",
          1099 => x"0d",
          1100 => x"84",
          1101 => x"52",
          1102 => x"70",
          1103 => x"81",
          1104 => x"72",
          1105 => x"0d",
          1106 => x"0d",
          1107 => x"84",
          1108 => x"c8",
          1109 => x"80",
          1110 => x"09",
          1111 => x"cc",
          1112 => x"81",
          1113 => x"73",
          1114 => x"3d",
          1115 => x"c8",
          1116 => x"c0",
          1117 => x"04",
          1118 => x"02",
          1119 => x"53",
          1120 => x"09",
          1121 => x"38",
          1122 => x"3f",
          1123 => x"08",
          1124 => x"2e",
          1125 => x"72",
          1126 => x"bc",
          1127 => x"81",
          1128 => x"8f",
          1129 => x"b4",
          1130 => x"80",
          1131 => x"72",
          1132 => x"84",
          1133 => x"fe",
          1134 => x"97",
          1135 => x"cb",
          1136 => x"81",
          1137 => x"54",
          1138 => x"3f",
          1139 => x"b4",
          1140 => x"0d",
          1141 => x"0d",
          1142 => x"33",
          1143 => x"06",
          1144 => x"80",
          1145 => x"72",
          1146 => x"51",
          1147 => x"ff",
          1148 => x"39",
          1149 => x"04",
          1150 => x"77",
          1151 => x"08",
          1152 => x"b4",
          1153 => x"73",
          1154 => x"ff",
          1155 => x"71",
          1156 => x"38",
          1157 => x"06",
          1158 => x"54",
          1159 => x"e7",
          1160 => x"cb",
          1161 => x"3d",
          1162 => x"3d",
          1163 => x"59",
          1164 => x"81",
          1165 => x"56",
          1166 => x"84",
          1167 => x"a5",
          1168 => x"06",
          1169 => x"80",
          1170 => x"81",
          1171 => x"58",
          1172 => x"b0",
          1173 => x"06",
          1174 => x"5a",
          1175 => x"ad",
          1176 => x"06",
          1177 => x"5a",
          1178 => x"05",
          1179 => x"75",
          1180 => x"81",
          1181 => x"77",
          1182 => x"08",
          1183 => x"05",
          1184 => x"5d",
          1185 => x"39",
          1186 => x"72",
          1187 => x"38",
          1188 => x"7b",
          1189 => x"05",
          1190 => x"70",
          1191 => x"33",
          1192 => x"39",
          1193 => x"32",
          1194 => x"72",
          1195 => x"78",
          1196 => x"70",
          1197 => x"07",
          1198 => x"07",
          1199 => x"51",
          1200 => x"80",
          1201 => x"79",
          1202 => x"70",
          1203 => x"33",
          1204 => x"80",
          1205 => x"38",
          1206 => x"e0",
          1207 => x"38",
          1208 => x"81",
          1209 => x"53",
          1210 => x"2e",
          1211 => x"73",
          1212 => x"a2",
          1213 => x"c3",
          1214 => x"38",
          1215 => x"24",
          1216 => x"80",
          1217 => x"8c",
          1218 => x"39",
          1219 => x"2e",
          1220 => x"81",
          1221 => x"80",
          1222 => x"80",
          1223 => x"d5",
          1224 => x"73",
          1225 => x"8e",
          1226 => x"39",
          1227 => x"2e",
          1228 => x"80",
          1229 => x"84",
          1230 => x"56",
          1231 => x"74",
          1232 => x"72",
          1233 => x"38",
          1234 => x"15",
          1235 => x"54",
          1236 => x"38",
          1237 => x"56",
          1238 => x"81",
          1239 => x"72",
          1240 => x"38",
          1241 => x"90",
          1242 => x"06",
          1243 => x"2e",
          1244 => x"51",
          1245 => x"74",
          1246 => x"53",
          1247 => x"fd",
          1248 => x"51",
          1249 => x"ef",
          1250 => x"19",
          1251 => x"53",
          1252 => x"39",
          1253 => x"39",
          1254 => x"39",
          1255 => x"39",
          1256 => x"39",
          1257 => x"d0",
          1258 => x"39",
          1259 => x"70",
          1260 => x"53",
          1261 => x"88",
          1262 => x"19",
          1263 => x"39",
          1264 => x"54",
          1265 => x"74",
          1266 => x"70",
          1267 => x"07",
          1268 => x"55",
          1269 => x"80",
          1270 => x"72",
          1271 => x"38",
          1272 => x"90",
          1273 => x"80",
          1274 => x"5e",
          1275 => x"74",
          1276 => x"3f",
          1277 => x"08",
          1278 => x"7c",
          1279 => x"54",
          1280 => x"81",
          1281 => x"55",
          1282 => x"92",
          1283 => x"53",
          1284 => x"2e",
          1285 => x"14",
          1286 => x"ff",
          1287 => x"14",
          1288 => x"70",
          1289 => x"34",
          1290 => x"30",
          1291 => x"9f",
          1292 => x"57",
          1293 => x"85",
          1294 => x"b1",
          1295 => x"2a",
          1296 => x"51",
          1297 => x"2e",
          1298 => x"3d",
          1299 => x"05",
          1300 => x"34",
          1301 => x"76",
          1302 => x"54",
          1303 => x"72",
          1304 => x"54",
          1305 => x"70",
          1306 => x"56",
          1307 => x"81",
          1308 => x"7b",
          1309 => x"73",
          1310 => x"3f",
          1311 => x"53",
          1312 => x"74",
          1313 => x"53",
          1314 => x"eb",
          1315 => x"77",
          1316 => x"53",
          1317 => x"14",
          1318 => x"54",
          1319 => x"3f",
          1320 => x"74",
          1321 => x"53",
          1322 => x"fb",
          1323 => x"51",
          1324 => x"ef",
          1325 => x"0d",
          1326 => x"0d",
          1327 => x"70",
          1328 => x"08",
          1329 => x"51",
          1330 => x"85",
          1331 => x"fe",
          1332 => x"81",
          1333 => x"85",
          1334 => x"52",
          1335 => x"ca",
          1336 => x"bc",
          1337 => x"73",
          1338 => x"81",
          1339 => x"84",
          1340 => x"fd",
          1341 => x"cb",
          1342 => x"81",
          1343 => x"87",
          1344 => x"53",
          1345 => x"fa",
          1346 => x"81",
          1347 => x"85",
          1348 => x"fb",
          1349 => x"79",
          1350 => x"08",
          1351 => x"57",
          1352 => x"71",
          1353 => x"e0",
          1354 => x"b8",
          1355 => x"2d",
          1356 => x"08",
          1357 => x"53",
          1358 => x"80",
          1359 => x"8d",
          1360 => x"72",
          1361 => x"30",
          1362 => x"51",
          1363 => x"80",
          1364 => x"71",
          1365 => x"38",
          1366 => x"97",
          1367 => x"25",
          1368 => x"16",
          1369 => x"25",
          1370 => x"14",
          1371 => x"34",
          1372 => x"72",
          1373 => x"3f",
          1374 => x"73",
          1375 => x"72",
          1376 => x"f7",
          1377 => x"53",
          1378 => x"a4",
          1379 => x"0d",
          1380 => x"0d",
          1381 => x"08",
          1382 => x"b8",
          1383 => x"76",
          1384 => x"ef",
          1385 => x"cb",
          1386 => x"3d",
          1387 => x"3d",
          1388 => x"5a",
          1389 => x"7a",
          1390 => x"08",
          1391 => x"53",
          1392 => x"09",
          1393 => x"38",
          1394 => x"0c",
          1395 => x"ad",
          1396 => x"06",
          1397 => x"76",
          1398 => x"0c",
          1399 => x"33",
          1400 => x"73",
          1401 => x"81",
          1402 => x"38",
          1403 => x"05",
          1404 => x"08",
          1405 => x"53",
          1406 => x"2e",
          1407 => x"57",
          1408 => x"2e",
          1409 => x"39",
          1410 => x"13",
          1411 => x"08",
          1412 => x"53",
          1413 => x"55",
          1414 => x"80",
          1415 => x"14",
          1416 => x"88",
          1417 => x"27",
          1418 => x"eb",
          1419 => x"53",
          1420 => x"89",
          1421 => x"38",
          1422 => x"55",
          1423 => x"8a",
          1424 => x"a0",
          1425 => x"c2",
          1426 => x"74",
          1427 => x"e0",
          1428 => x"ff",
          1429 => x"d0",
          1430 => x"ff",
          1431 => x"90",
          1432 => x"38",
          1433 => x"81",
          1434 => x"53",
          1435 => x"ca",
          1436 => x"27",
          1437 => x"77",
          1438 => x"08",
          1439 => x"0c",
          1440 => x"33",
          1441 => x"ff",
          1442 => x"80",
          1443 => x"74",
          1444 => x"79",
          1445 => x"74",
          1446 => x"0c",
          1447 => x"04",
          1448 => x"7a",
          1449 => x"80",
          1450 => x"58",
          1451 => x"33",
          1452 => x"a0",
          1453 => x"06",
          1454 => x"13",
          1455 => x"39",
          1456 => x"09",
          1457 => x"38",
          1458 => x"11",
          1459 => x"08",
          1460 => x"54",
          1461 => x"2e",
          1462 => x"80",
          1463 => x"08",
          1464 => x"0c",
          1465 => x"33",
          1466 => x"80",
          1467 => x"38",
          1468 => x"80",
          1469 => x"38",
          1470 => x"57",
          1471 => x"0c",
          1472 => x"33",
          1473 => x"39",
          1474 => x"74",
          1475 => x"38",
          1476 => x"80",
          1477 => x"89",
          1478 => x"38",
          1479 => x"d0",
          1480 => x"55",
          1481 => x"80",
          1482 => x"39",
          1483 => x"d9",
          1484 => x"80",
          1485 => x"27",
          1486 => x"80",
          1487 => x"89",
          1488 => x"70",
          1489 => x"55",
          1490 => x"70",
          1491 => x"55",
          1492 => x"27",
          1493 => x"14",
          1494 => x"06",
          1495 => x"74",
          1496 => x"73",
          1497 => x"38",
          1498 => x"14",
          1499 => x"05",
          1500 => x"08",
          1501 => x"54",
          1502 => x"39",
          1503 => x"84",
          1504 => x"55",
          1505 => x"81",
          1506 => x"cb",
          1507 => x"3d",
          1508 => x"3d",
          1509 => x"05",
          1510 => x"52",
          1511 => x"87",
          1512 => x"d0",
          1513 => x"71",
          1514 => x"0c",
          1515 => x"04",
          1516 => x"02",
          1517 => x"02",
          1518 => x"05",
          1519 => x"83",
          1520 => x"26",
          1521 => x"72",
          1522 => x"c0",
          1523 => x"53",
          1524 => x"74",
          1525 => x"38",
          1526 => x"73",
          1527 => x"c0",
          1528 => x"51",
          1529 => x"85",
          1530 => x"98",
          1531 => x"52",
          1532 => x"82",
          1533 => x"70",
          1534 => x"38",
          1535 => x"8c",
          1536 => x"ec",
          1537 => x"fc",
          1538 => x"52",
          1539 => x"87",
          1540 => x"08",
          1541 => x"2e",
          1542 => x"81",
          1543 => x"34",
          1544 => x"13",
          1545 => x"81",
          1546 => x"86",
          1547 => x"f3",
          1548 => x"62",
          1549 => x"05",
          1550 => x"57",
          1551 => x"83",
          1552 => x"fe",
          1553 => x"cb",
          1554 => x"06",
          1555 => x"71",
          1556 => x"71",
          1557 => x"2b",
          1558 => x"80",
          1559 => x"92",
          1560 => x"c0",
          1561 => x"41",
          1562 => x"5a",
          1563 => x"87",
          1564 => x"0c",
          1565 => x"84",
          1566 => x"08",
          1567 => x"70",
          1568 => x"53",
          1569 => x"2e",
          1570 => x"08",
          1571 => x"70",
          1572 => x"34",
          1573 => x"80",
          1574 => x"53",
          1575 => x"2e",
          1576 => x"53",
          1577 => x"26",
          1578 => x"80",
          1579 => x"87",
          1580 => x"08",
          1581 => x"38",
          1582 => x"8c",
          1583 => x"80",
          1584 => x"78",
          1585 => x"99",
          1586 => x"0c",
          1587 => x"8c",
          1588 => x"08",
          1589 => x"51",
          1590 => x"38",
          1591 => x"8d",
          1592 => x"17",
          1593 => x"81",
          1594 => x"53",
          1595 => x"2e",
          1596 => x"fc",
          1597 => x"52",
          1598 => x"7d",
          1599 => x"ed",
          1600 => x"80",
          1601 => x"71",
          1602 => x"38",
          1603 => x"53",
          1604 => x"a4",
          1605 => x"0d",
          1606 => x"0d",
          1607 => x"02",
          1608 => x"05",
          1609 => x"58",
          1610 => x"80",
          1611 => x"fc",
          1612 => x"cb",
          1613 => x"06",
          1614 => x"71",
          1615 => x"81",
          1616 => x"38",
          1617 => x"2b",
          1618 => x"80",
          1619 => x"92",
          1620 => x"c0",
          1621 => x"40",
          1622 => x"5a",
          1623 => x"c0",
          1624 => x"76",
          1625 => x"76",
          1626 => x"75",
          1627 => x"2a",
          1628 => x"51",
          1629 => x"80",
          1630 => x"7a",
          1631 => x"5c",
          1632 => x"81",
          1633 => x"81",
          1634 => x"06",
          1635 => x"80",
          1636 => x"87",
          1637 => x"08",
          1638 => x"38",
          1639 => x"8c",
          1640 => x"80",
          1641 => x"77",
          1642 => x"99",
          1643 => x"0c",
          1644 => x"8c",
          1645 => x"08",
          1646 => x"51",
          1647 => x"38",
          1648 => x"8d",
          1649 => x"70",
          1650 => x"84",
          1651 => x"5b",
          1652 => x"2e",
          1653 => x"fc",
          1654 => x"52",
          1655 => x"7d",
          1656 => x"f8",
          1657 => x"80",
          1658 => x"71",
          1659 => x"38",
          1660 => x"53",
          1661 => x"a4",
          1662 => x"0d",
          1663 => x"0d",
          1664 => x"05",
          1665 => x"02",
          1666 => x"05",
          1667 => x"54",
          1668 => x"fe",
          1669 => x"a4",
          1670 => x"53",
          1671 => x"80",
          1672 => x"0b",
          1673 => x"8c",
          1674 => x"71",
          1675 => x"dc",
          1676 => x"24",
          1677 => x"84",
          1678 => x"92",
          1679 => x"54",
          1680 => x"8d",
          1681 => x"39",
          1682 => x"80",
          1683 => x"cb",
          1684 => x"70",
          1685 => x"81",
          1686 => x"52",
          1687 => x"8a",
          1688 => x"98",
          1689 => x"71",
          1690 => x"c0",
          1691 => x"52",
          1692 => x"81",
          1693 => x"c0",
          1694 => x"53",
          1695 => x"82",
          1696 => x"71",
          1697 => x"39",
          1698 => x"39",
          1699 => x"77",
          1700 => x"81",
          1701 => x"72",
          1702 => x"84",
          1703 => x"73",
          1704 => x"0c",
          1705 => x"04",
          1706 => x"74",
          1707 => x"71",
          1708 => x"2b",
          1709 => x"a4",
          1710 => x"84",
          1711 => x"fd",
          1712 => x"83",
          1713 => x"12",
          1714 => x"2b",
          1715 => x"07",
          1716 => x"70",
          1717 => x"2b",
          1718 => x"07",
          1719 => x"0c",
          1720 => x"56",
          1721 => x"3d",
          1722 => x"3d",
          1723 => x"84",
          1724 => x"22",
          1725 => x"72",
          1726 => x"54",
          1727 => x"2a",
          1728 => x"34",
          1729 => x"04",
          1730 => x"73",
          1731 => x"70",
          1732 => x"05",
          1733 => x"88",
          1734 => x"72",
          1735 => x"54",
          1736 => x"2a",
          1737 => x"70",
          1738 => x"34",
          1739 => x"51",
          1740 => x"83",
          1741 => x"fe",
          1742 => x"75",
          1743 => x"51",
          1744 => x"92",
          1745 => x"81",
          1746 => x"73",
          1747 => x"55",
          1748 => x"51",
          1749 => x"3d",
          1750 => x"3d",
          1751 => x"76",
          1752 => x"72",
          1753 => x"05",
          1754 => x"11",
          1755 => x"38",
          1756 => x"04",
          1757 => x"78",
          1758 => x"56",
          1759 => x"81",
          1760 => x"74",
          1761 => x"56",
          1762 => x"31",
          1763 => x"52",
          1764 => x"80",
          1765 => x"71",
          1766 => x"38",
          1767 => x"a4",
          1768 => x"0d",
          1769 => x"0d",
          1770 => x"51",
          1771 => x"73",
          1772 => x"81",
          1773 => x"33",
          1774 => x"38",
          1775 => x"cb",
          1776 => x"3d",
          1777 => x"0b",
          1778 => x"0c",
          1779 => x"81",
          1780 => x"04",
          1781 => x"7b",
          1782 => x"83",
          1783 => x"5a",
          1784 => x"80",
          1785 => x"54",
          1786 => x"53",
          1787 => x"53",
          1788 => x"52",
          1789 => x"3f",
          1790 => x"08",
          1791 => x"81",
          1792 => x"81",
          1793 => x"83",
          1794 => x"16",
          1795 => x"18",
          1796 => x"18",
          1797 => x"58",
          1798 => x"9f",
          1799 => x"33",
          1800 => x"2e",
          1801 => x"93",
          1802 => x"76",
          1803 => x"52",
          1804 => x"51",
          1805 => x"83",
          1806 => x"79",
          1807 => x"0c",
          1808 => x"04",
          1809 => x"78",
          1810 => x"80",
          1811 => x"17",
          1812 => x"38",
          1813 => x"fc",
          1814 => x"a4",
          1815 => x"cb",
          1816 => x"38",
          1817 => x"53",
          1818 => x"81",
          1819 => x"f7",
          1820 => x"cb",
          1821 => x"2e",
          1822 => x"55",
          1823 => x"b0",
          1824 => x"81",
          1825 => x"88",
          1826 => x"f8",
          1827 => x"70",
          1828 => x"c0",
          1829 => x"a4",
          1830 => x"cb",
          1831 => x"91",
          1832 => x"55",
          1833 => x"09",
          1834 => x"f0",
          1835 => x"33",
          1836 => x"2e",
          1837 => x"80",
          1838 => x"80",
          1839 => x"a4",
          1840 => x"17",
          1841 => x"fd",
          1842 => x"d4",
          1843 => x"b2",
          1844 => x"96",
          1845 => x"85",
          1846 => x"75",
          1847 => x"3f",
          1848 => x"e4",
          1849 => x"98",
          1850 => x"9c",
          1851 => x"08",
          1852 => x"17",
          1853 => x"3f",
          1854 => x"52",
          1855 => x"51",
          1856 => x"a0",
          1857 => x"05",
          1858 => x"0c",
          1859 => x"75",
          1860 => x"33",
          1861 => x"3f",
          1862 => x"34",
          1863 => x"52",
          1864 => x"51",
          1865 => x"81",
          1866 => x"80",
          1867 => x"81",
          1868 => x"cb",
          1869 => x"3d",
          1870 => x"3d",
          1871 => x"1a",
          1872 => x"fe",
          1873 => x"54",
          1874 => x"73",
          1875 => x"8a",
          1876 => x"71",
          1877 => x"08",
          1878 => x"75",
          1879 => x"0c",
          1880 => x"04",
          1881 => x"7a",
          1882 => x"56",
          1883 => x"77",
          1884 => x"38",
          1885 => x"08",
          1886 => x"38",
          1887 => x"54",
          1888 => x"2e",
          1889 => x"72",
          1890 => x"38",
          1891 => x"8d",
          1892 => x"39",
          1893 => x"81",
          1894 => x"b6",
          1895 => x"2a",
          1896 => x"2a",
          1897 => x"05",
          1898 => x"55",
          1899 => x"81",
          1900 => x"81",
          1901 => x"83",
          1902 => x"b4",
          1903 => x"17",
          1904 => x"a4",
          1905 => x"55",
          1906 => x"57",
          1907 => x"3f",
          1908 => x"08",
          1909 => x"74",
          1910 => x"14",
          1911 => x"70",
          1912 => x"07",
          1913 => x"71",
          1914 => x"52",
          1915 => x"72",
          1916 => x"75",
          1917 => x"58",
          1918 => x"76",
          1919 => x"15",
          1920 => x"73",
          1921 => x"3f",
          1922 => x"08",
          1923 => x"76",
          1924 => x"06",
          1925 => x"05",
          1926 => x"3f",
          1927 => x"08",
          1928 => x"06",
          1929 => x"76",
          1930 => x"15",
          1931 => x"73",
          1932 => x"3f",
          1933 => x"08",
          1934 => x"82",
          1935 => x"06",
          1936 => x"05",
          1937 => x"3f",
          1938 => x"08",
          1939 => x"58",
          1940 => x"58",
          1941 => x"a4",
          1942 => x"0d",
          1943 => x"0d",
          1944 => x"5a",
          1945 => x"59",
          1946 => x"82",
          1947 => x"98",
          1948 => x"82",
          1949 => x"33",
          1950 => x"2e",
          1951 => x"72",
          1952 => x"38",
          1953 => x"8d",
          1954 => x"39",
          1955 => x"81",
          1956 => x"f7",
          1957 => x"2a",
          1958 => x"2a",
          1959 => x"05",
          1960 => x"55",
          1961 => x"81",
          1962 => x"59",
          1963 => x"08",
          1964 => x"74",
          1965 => x"16",
          1966 => x"16",
          1967 => x"59",
          1968 => x"53",
          1969 => x"8f",
          1970 => x"2b",
          1971 => x"74",
          1972 => x"71",
          1973 => x"72",
          1974 => x"0b",
          1975 => x"74",
          1976 => x"17",
          1977 => x"75",
          1978 => x"3f",
          1979 => x"08",
          1980 => x"a4",
          1981 => x"38",
          1982 => x"06",
          1983 => x"78",
          1984 => x"54",
          1985 => x"77",
          1986 => x"33",
          1987 => x"71",
          1988 => x"51",
          1989 => x"34",
          1990 => x"76",
          1991 => x"17",
          1992 => x"75",
          1993 => x"3f",
          1994 => x"08",
          1995 => x"a4",
          1996 => x"38",
          1997 => x"ff",
          1998 => x"10",
          1999 => x"76",
          2000 => x"51",
          2001 => x"be",
          2002 => x"2a",
          2003 => x"05",
          2004 => x"f9",
          2005 => x"cb",
          2006 => x"81",
          2007 => x"ab",
          2008 => x"0a",
          2009 => x"2b",
          2010 => x"70",
          2011 => x"70",
          2012 => x"54",
          2013 => x"81",
          2014 => x"8f",
          2015 => x"07",
          2016 => x"f7",
          2017 => x"0b",
          2018 => x"78",
          2019 => x"0c",
          2020 => x"04",
          2021 => x"7a",
          2022 => x"08",
          2023 => x"59",
          2024 => x"a4",
          2025 => x"17",
          2026 => x"38",
          2027 => x"aa",
          2028 => x"73",
          2029 => x"fd",
          2030 => x"cb",
          2031 => x"81",
          2032 => x"80",
          2033 => x"39",
          2034 => x"eb",
          2035 => x"80",
          2036 => x"cb",
          2037 => x"80",
          2038 => x"52",
          2039 => x"84",
          2040 => x"a4",
          2041 => x"cb",
          2042 => x"2e",
          2043 => x"81",
          2044 => x"81",
          2045 => x"81",
          2046 => x"ff",
          2047 => x"80",
          2048 => x"75",
          2049 => x"3f",
          2050 => x"08",
          2051 => x"16",
          2052 => x"90",
          2053 => x"55",
          2054 => x"27",
          2055 => x"15",
          2056 => x"84",
          2057 => x"07",
          2058 => x"17",
          2059 => x"76",
          2060 => x"a6",
          2061 => x"73",
          2062 => x"0c",
          2063 => x"04",
          2064 => x"7c",
          2065 => x"59",
          2066 => x"95",
          2067 => x"08",
          2068 => x"2e",
          2069 => x"17",
          2070 => x"b2",
          2071 => x"ae",
          2072 => x"7a",
          2073 => x"3f",
          2074 => x"81",
          2075 => x"27",
          2076 => x"81",
          2077 => x"55",
          2078 => x"08",
          2079 => x"d2",
          2080 => x"08",
          2081 => x"08",
          2082 => x"38",
          2083 => x"17",
          2084 => x"54",
          2085 => x"82",
          2086 => x"7a",
          2087 => x"06",
          2088 => x"81",
          2089 => x"17",
          2090 => x"83",
          2091 => x"75",
          2092 => x"f9",
          2093 => x"59",
          2094 => x"08",
          2095 => x"81",
          2096 => x"81",
          2097 => x"59",
          2098 => x"08",
          2099 => x"70",
          2100 => x"25",
          2101 => x"81",
          2102 => x"54",
          2103 => x"55",
          2104 => x"38",
          2105 => x"08",
          2106 => x"38",
          2107 => x"54",
          2108 => x"90",
          2109 => x"18",
          2110 => x"38",
          2111 => x"39",
          2112 => x"38",
          2113 => x"16",
          2114 => x"08",
          2115 => x"38",
          2116 => x"78",
          2117 => x"38",
          2118 => x"51",
          2119 => x"81",
          2120 => x"80",
          2121 => x"80",
          2122 => x"a4",
          2123 => x"09",
          2124 => x"38",
          2125 => x"08",
          2126 => x"a4",
          2127 => x"30",
          2128 => x"80",
          2129 => x"07",
          2130 => x"55",
          2131 => x"38",
          2132 => x"09",
          2133 => x"ae",
          2134 => x"80",
          2135 => x"53",
          2136 => x"51",
          2137 => x"81",
          2138 => x"81",
          2139 => x"30",
          2140 => x"a4",
          2141 => x"25",
          2142 => x"79",
          2143 => x"38",
          2144 => x"8f",
          2145 => x"79",
          2146 => x"f9",
          2147 => x"cb",
          2148 => x"74",
          2149 => x"8c",
          2150 => x"17",
          2151 => x"90",
          2152 => x"54",
          2153 => x"86",
          2154 => x"90",
          2155 => x"17",
          2156 => x"54",
          2157 => x"34",
          2158 => x"56",
          2159 => x"90",
          2160 => x"80",
          2161 => x"81",
          2162 => x"55",
          2163 => x"56",
          2164 => x"81",
          2165 => x"8c",
          2166 => x"f8",
          2167 => x"70",
          2168 => x"f0",
          2169 => x"a4",
          2170 => x"56",
          2171 => x"08",
          2172 => x"7b",
          2173 => x"f6",
          2174 => x"cb",
          2175 => x"cb",
          2176 => x"17",
          2177 => x"80",
          2178 => x"b4",
          2179 => x"57",
          2180 => x"77",
          2181 => x"81",
          2182 => x"15",
          2183 => x"78",
          2184 => x"81",
          2185 => x"53",
          2186 => x"15",
          2187 => x"e9",
          2188 => x"a4",
          2189 => x"df",
          2190 => x"22",
          2191 => x"30",
          2192 => x"70",
          2193 => x"51",
          2194 => x"81",
          2195 => x"8a",
          2196 => x"f8",
          2197 => x"7c",
          2198 => x"56",
          2199 => x"80",
          2200 => x"f1",
          2201 => x"06",
          2202 => x"e9",
          2203 => x"18",
          2204 => x"08",
          2205 => x"38",
          2206 => x"82",
          2207 => x"38",
          2208 => x"54",
          2209 => x"74",
          2210 => x"82",
          2211 => x"22",
          2212 => x"79",
          2213 => x"38",
          2214 => x"98",
          2215 => x"cd",
          2216 => x"22",
          2217 => x"54",
          2218 => x"26",
          2219 => x"52",
          2220 => x"b0",
          2221 => x"a4",
          2222 => x"cb",
          2223 => x"2e",
          2224 => x"0b",
          2225 => x"08",
          2226 => x"98",
          2227 => x"cb",
          2228 => x"85",
          2229 => x"bd",
          2230 => x"31",
          2231 => x"73",
          2232 => x"f4",
          2233 => x"cb",
          2234 => x"18",
          2235 => x"18",
          2236 => x"08",
          2237 => x"72",
          2238 => x"38",
          2239 => x"58",
          2240 => x"89",
          2241 => x"18",
          2242 => x"ff",
          2243 => x"05",
          2244 => x"80",
          2245 => x"cb",
          2246 => x"3d",
          2247 => x"3d",
          2248 => x"08",
          2249 => x"a0",
          2250 => x"54",
          2251 => x"77",
          2252 => x"80",
          2253 => x"0c",
          2254 => x"53",
          2255 => x"80",
          2256 => x"38",
          2257 => x"06",
          2258 => x"b5",
          2259 => x"98",
          2260 => x"14",
          2261 => x"92",
          2262 => x"2a",
          2263 => x"56",
          2264 => x"26",
          2265 => x"80",
          2266 => x"16",
          2267 => x"77",
          2268 => x"53",
          2269 => x"38",
          2270 => x"51",
          2271 => x"81",
          2272 => x"53",
          2273 => x"0b",
          2274 => x"08",
          2275 => x"38",
          2276 => x"cb",
          2277 => x"2e",
          2278 => x"98",
          2279 => x"cb",
          2280 => x"80",
          2281 => x"8a",
          2282 => x"15",
          2283 => x"80",
          2284 => x"14",
          2285 => x"51",
          2286 => x"81",
          2287 => x"53",
          2288 => x"cb",
          2289 => x"2e",
          2290 => x"82",
          2291 => x"a4",
          2292 => x"ba",
          2293 => x"81",
          2294 => x"ff",
          2295 => x"81",
          2296 => x"52",
          2297 => x"f3",
          2298 => x"a4",
          2299 => x"72",
          2300 => x"72",
          2301 => x"f2",
          2302 => x"cb",
          2303 => x"15",
          2304 => x"15",
          2305 => x"b4",
          2306 => x"0c",
          2307 => x"81",
          2308 => x"8a",
          2309 => x"f7",
          2310 => x"7d",
          2311 => x"5b",
          2312 => x"76",
          2313 => x"3f",
          2314 => x"08",
          2315 => x"a4",
          2316 => x"38",
          2317 => x"08",
          2318 => x"08",
          2319 => x"f0",
          2320 => x"cb",
          2321 => x"81",
          2322 => x"80",
          2323 => x"cb",
          2324 => x"18",
          2325 => x"51",
          2326 => x"81",
          2327 => x"81",
          2328 => x"81",
          2329 => x"a4",
          2330 => x"83",
          2331 => x"77",
          2332 => x"72",
          2333 => x"38",
          2334 => x"75",
          2335 => x"81",
          2336 => x"a5",
          2337 => x"a4",
          2338 => x"52",
          2339 => x"8e",
          2340 => x"a4",
          2341 => x"cb",
          2342 => x"2e",
          2343 => x"73",
          2344 => x"81",
          2345 => x"87",
          2346 => x"cb",
          2347 => x"3d",
          2348 => x"3d",
          2349 => x"11",
          2350 => x"ec",
          2351 => x"a4",
          2352 => x"ff",
          2353 => x"33",
          2354 => x"71",
          2355 => x"81",
          2356 => x"94",
          2357 => x"d0",
          2358 => x"a4",
          2359 => x"73",
          2360 => x"81",
          2361 => x"85",
          2362 => x"fc",
          2363 => x"79",
          2364 => x"ff",
          2365 => x"12",
          2366 => x"eb",
          2367 => x"70",
          2368 => x"72",
          2369 => x"81",
          2370 => x"73",
          2371 => x"94",
          2372 => x"d6",
          2373 => x"0d",
          2374 => x"0d",
          2375 => x"55",
          2376 => x"5a",
          2377 => x"08",
          2378 => x"8a",
          2379 => x"08",
          2380 => x"ee",
          2381 => x"cb",
          2382 => x"81",
          2383 => x"80",
          2384 => x"15",
          2385 => x"55",
          2386 => x"38",
          2387 => x"e6",
          2388 => x"33",
          2389 => x"70",
          2390 => x"58",
          2391 => x"86",
          2392 => x"cb",
          2393 => x"73",
          2394 => x"83",
          2395 => x"73",
          2396 => x"38",
          2397 => x"06",
          2398 => x"80",
          2399 => x"75",
          2400 => x"38",
          2401 => x"08",
          2402 => x"54",
          2403 => x"2e",
          2404 => x"83",
          2405 => x"73",
          2406 => x"38",
          2407 => x"51",
          2408 => x"81",
          2409 => x"58",
          2410 => x"08",
          2411 => x"15",
          2412 => x"38",
          2413 => x"0b",
          2414 => x"77",
          2415 => x"0c",
          2416 => x"04",
          2417 => x"77",
          2418 => x"54",
          2419 => x"51",
          2420 => x"81",
          2421 => x"55",
          2422 => x"08",
          2423 => x"14",
          2424 => x"51",
          2425 => x"81",
          2426 => x"55",
          2427 => x"08",
          2428 => x"53",
          2429 => x"08",
          2430 => x"08",
          2431 => x"3f",
          2432 => x"14",
          2433 => x"08",
          2434 => x"3f",
          2435 => x"17",
          2436 => x"cb",
          2437 => x"3d",
          2438 => x"3d",
          2439 => x"08",
          2440 => x"54",
          2441 => x"53",
          2442 => x"81",
          2443 => x"8d",
          2444 => x"08",
          2445 => x"34",
          2446 => x"15",
          2447 => x"0d",
          2448 => x"0d",
          2449 => x"57",
          2450 => x"17",
          2451 => x"08",
          2452 => x"82",
          2453 => x"89",
          2454 => x"55",
          2455 => x"14",
          2456 => x"16",
          2457 => x"71",
          2458 => x"38",
          2459 => x"09",
          2460 => x"38",
          2461 => x"73",
          2462 => x"81",
          2463 => x"ae",
          2464 => x"05",
          2465 => x"15",
          2466 => x"70",
          2467 => x"34",
          2468 => x"8a",
          2469 => x"38",
          2470 => x"05",
          2471 => x"81",
          2472 => x"17",
          2473 => x"12",
          2474 => x"34",
          2475 => x"9c",
          2476 => x"e8",
          2477 => x"cb",
          2478 => x"0c",
          2479 => x"e7",
          2480 => x"cb",
          2481 => x"17",
          2482 => x"51",
          2483 => x"81",
          2484 => x"84",
          2485 => x"3d",
          2486 => x"3d",
          2487 => x"08",
          2488 => x"61",
          2489 => x"55",
          2490 => x"2e",
          2491 => x"55",
          2492 => x"2e",
          2493 => x"80",
          2494 => x"94",
          2495 => x"1c",
          2496 => x"81",
          2497 => x"61",
          2498 => x"56",
          2499 => x"2e",
          2500 => x"83",
          2501 => x"73",
          2502 => x"70",
          2503 => x"25",
          2504 => x"51",
          2505 => x"38",
          2506 => x"0c",
          2507 => x"51",
          2508 => x"26",
          2509 => x"80",
          2510 => x"34",
          2511 => x"51",
          2512 => x"81",
          2513 => x"55",
          2514 => x"91",
          2515 => x"1d",
          2516 => x"8b",
          2517 => x"79",
          2518 => x"3f",
          2519 => x"57",
          2520 => x"55",
          2521 => x"2e",
          2522 => x"80",
          2523 => x"18",
          2524 => x"1a",
          2525 => x"70",
          2526 => x"2a",
          2527 => x"07",
          2528 => x"5a",
          2529 => x"8c",
          2530 => x"54",
          2531 => x"81",
          2532 => x"39",
          2533 => x"70",
          2534 => x"2a",
          2535 => x"75",
          2536 => x"8c",
          2537 => x"2e",
          2538 => x"a0",
          2539 => x"38",
          2540 => x"0c",
          2541 => x"76",
          2542 => x"38",
          2543 => x"b8",
          2544 => x"70",
          2545 => x"5a",
          2546 => x"76",
          2547 => x"38",
          2548 => x"70",
          2549 => x"dc",
          2550 => x"72",
          2551 => x"80",
          2552 => x"51",
          2553 => x"73",
          2554 => x"38",
          2555 => x"18",
          2556 => x"1a",
          2557 => x"55",
          2558 => x"2e",
          2559 => x"83",
          2560 => x"73",
          2561 => x"70",
          2562 => x"25",
          2563 => x"51",
          2564 => x"38",
          2565 => x"75",
          2566 => x"81",
          2567 => x"81",
          2568 => x"27",
          2569 => x"73",
          2570 => x"38",
          2571 => x"70",
          2572 => x"32",
          2573 => x"80",
          2574 => x"2a",
          2575 => x"56",
          2576 => x"81",
          2577 => x"57",
          2578 => x"f5",
          2579 => x"2b",
          2580 => x"25",
          2581 => x"80",
          2582 => x"bb",
          2583 => x"57",
          2584 => x"e6",
          2585 => x"cb",
          2586 => x"2e",
          2587 => x"18",
          2588 => x"1a",
          2589 => x"56",
          2590 => x"3f",
          2591 => x"08",
          2592 => x"e8",
          2593 => x"54",
          2594 => x"80",
          2595 => x"17",
          2596 => x"34",
          2597 => x"11",
          2598 => x"74",
          2599 => x"75",
          2600 => x"a0",
          2601 => x"3f",
          2602 => x"08",
          2603 => x"9f",
          2604 => x"99",
          2605 => x"e0",
          2606 => x"ff",
          2607 => x"79",
          2608 => x"74",
          2609 => x"57",
          2610 => x"77",
          2611 => x"76",
          2612 => x"38",
          2613 => x"73",
          2614 => x"09",
          2615 => x"38",
          2616 => x"84",
          2617 => x"27",
          2618 => x"39",
          2619 => x"f2",
          2620 => x"80",
          2621 => x"54",
          2622 => x"34",
          2623 => x"58",
          2624 => x"f2",
          2625 => x"cb",
          2626 => x"81",
          2627 => x"80",
          2628 => x"1b",
          2629 => x"51",
          2630 => x"81",
          2631 => x"56",
          2632 => x"08",
          2633 => x"9c",
          2634 => x"33",
          2635 => x"80",
          2636 => x"38",
          2637 => x"bf",
          2638 => x"86",
          2639 => x"15",
          2640 => x"2a",
          2641 => x"51",
          2642 => x"92",
          2643 => x"79",
          2644 => x"e4",
          2645 => x"cb",
          2646 => x"2e",
          2647 => x"52",
          2648 => x"ba",
          2649 => x"39",
          2650 => x"33",
          2651 => x"80",
          2652 => x"74",
          2653 => x"81",
          2654 => x"38",
          2655 => x"70",
          2656 => x"82",
          2657 => x"54",
          2658 => x"96",
          2659 => x"06",
          2660 => x"2e",
          2661 => x"ff",
          2662 => x"1c",
          2663 => x"80",
          2664 => x"81",
          2665 => x"ba",
          2666 => x"b6",
          2667 => x"2a",
          2668 => x"51",
          2669 => x"38",
          2670 => x"70",
          2671 => x"81",
          2672 => x"55",
          2673 => x"e1",
          2674 => x"08",
          2675 => x"1d",
          2676 => x"7c",
          2677 => x"3f",
          2678 => x"08",
          2679 => x"fa",
          2680 => x"81",
          2681 => x"8f",
          2682 => x"f6",
          2683 => x"5b",
          2684 => x"70",
          2685 => x"59",
          2686 => x"73",
          2687 => x"c6",
          2688 => x"81",
          2689 => x"70",
          2690 => x"52",
          2691 => x"8d",
          2692 => x"38",
          2693 => x"09",
          2694 => x"a5",
          2695 => x"d0",
          2696 => x"ff",
          2697 => x"53",
          2698 => x"91",
          2699 => x"73",
          2700 => x"d0",
          2701 => x"71",
          2702 => x"f7",
          2703 => x"81",
          2704 => x"55",
          2705 => x"55",
          2706 => x"81",
          2707 => x"74",
          2708 => x"56",
          2709 => x"12",
          2710 => x"70",
          2711 => x"38",
          2712 => x"81",
          2713 => x"51",
          2714 => x"51",
          2715 => x"89",
          2716 => x"70",
          2717 => x"53",
          2718 => x"70",
          2719 => x"51",
          2720 => x"09",
          2721 => x"38",
          2722 => x"38",
          2723 => x"77",
          2724 => x"70",
          2725 => x"2a",
          2726 => x"07",
          2727 => x"51",
          2728 => x"8f",
          2729 => x"84",
          2730 => x"83",
          2731 => x"94",
          2732 => x"74",
          2733 => x"38",
          2734 => x"0c",
          2735 => x"86",
          2736 => x"d4",
          2737 => x"81",
          2738 => x"8c",
          2739 => x"fa",
          2740 => x"56",
          2741 => x"17",
          2742 => x"b0",
          2743 => x"52",
          2744 => x"e0",
          2745 => x"81",
          2746 => x"81",
          2747 => x"b2",
          2748 => x"b4",
          2749 => x"a4",
          2750 => x"ff",
          2751 => x"55",
          2752 => x"d5",
          2753 => x"06",
          2754 => x"80",
          2755 => x"33",
          2756 => x"81",
          2757 => x"81",
          2758 => x"81",
          2759 => x"eb",
          2760 => x"70",
          2761 => x"07",
          2762 => x"73",
          2763 => x"81",
          2764 => x"81",
          2765 => x"83",
          2766 => x"b0",
          2767 => x"16",
          2768 => x"3f",
          2769 => x"08",
          2770 => x"a4",
          2771 => x"9d",
          2772 => x"81",
          2773 => x"81",
          2774 => x"e0",
          2775 => x"cb",
          2776 => x"81",
          2777 => x"80",
          2778 => x"82",
          2779 => x"cb",
          2780 => x"3d",
          2781 => x"3d",
          2782 => x"84",
          2783 => x"05",
          2784 => x"80",
          2785 => x"51",
          2786 => x"81",
          2787 => x"58",
          2788 => x"0b",
          2789 => x"08",
          2790 => x"38",
          2791 => x"08",
          2792 => x"cb",
          2793 => x"08",
          2794 => x"56",
          2795 => x"86",
          2796 => x"75",
          2797 => x"fe",
          2798 => x"54",
          2799 => x"2e",
          2800 => x"14",
          2801 => x"ca",
          2802 => x"a4",
          2803 => x"06",
          2804 => x"54",
          2805 => x"38",
          2806 => x"86",
          2807 => x"82",
          2808 => x"06",
          2809 => x"56",
          2810 => x"38",
          2811 => x"80",
          2812 => x"81",
          2813 => x"52",
          2814 => x"51",
          2815 => x"81",
          2816 => x"81",
          2817 => x"81",
          2818 => x"83",
          2819 => x"87",
          2820 => x"2e",
          2821 => x"82",
          2822 => x"06",
          2823 => x"56",
          2824 => x"38",
          2825 => x"74",
          2826 => x"a3",
          2827 => x"a4",
          2828 => x"06",
          2829 => x"2e",
          2830 => x"80",
          2831 => x"3d",
          2832 => x"83",
          2833 => x"15",
          2834 => x"53",
          2835 => x"8d",
          2836 => x"15",
          2837 => x"3f",
          2838 => x"08",
          2839 => x"70",
          2840 => x"0c",
          2841 => x"16",
          2842 => x"80",
          2843 => x"80",
          2844 => x"54",
          2845 => x"84",
          2846 => x"5b",
          2847 => x"80",
          2848 => x"7a",
          2849 => x"fc",
          2850 => x"cb",
          2851 => x"ff",
          2852 => x"77",
          2853 => x"81",
          2854 => x"76",
          2855 => x"81",
          2856 => x"2e",
          2857 => x"8d",
          2858 => x"26",
          2859 => x"bf",
          2860 => x"f4",
          2861 => x"a4",
          2862 => x"ff",
          2863 => x"84",
          2864 => x"81",
          2865 => x"38",
          2866 => x"51",
          2867 => x"81",
          2868 => x"83",
          2869 => x"58",
          2870 => x"80",
          2871 => x"db",
          2872 => x"cb",
          2873 => x"77",
          2874 => x"80",
          2875 => x"82",
          2876 => x"c4",
          2877 => x"11",
          2878 => x"06",
          2879 => x"8d",
          2880 => x"26",
          2881 => x"74",
          2882 => x"78",
          2883 => x"c1",
          2884 => x"59",
          2885 => x"15",
          2886 => x"2e",
          2887 => x"13",
          2888 => x"72",
          2889 => x"38",
          2890 => x"eb",
          2891 => x"14",
          2892 => x"3f",
          2893 => x"08",
          2894 => x"a4",
          2895 => x"23",
          2896 => x"57",
          2897 => x"83",
          2898 => x"c7",
          2899 => x"d8",
          2900 => x"a4",
          2901 => x"ff",
          2902 => x"8d",
          2903 => x"14",
          2904 => x"3f",
          2905 => x"08",
          2906 => x"14",
          2907 => x"3f",
          2908 => x"08",
          2909 => x"06",
          2910 => x"72",
          2911 => x"97",
          2912 => x"22",
          2913 => x"84",
          2914 => x"5a",
          2915 => x"83",
          2916 => x"14",
          2917 => x"79",
          2918 => x"b3",
          2919 => x"cb",
          2920 => x"81",
          2921 => x"80",
          2922 => x"38",
          2923 => x"08",
          2924 => x"ff",
          2925 => x"38",
          2926 => x"83",
          2927 => x"83",
          2928 => x"74",
          2929 => x"85",
          2930 => x"89",
          2931 => x"76",
          2932 => x"c3",
          2933 => x"70",
          2934 => x"7b",
          2935 => x"73",
          2936 => x"17",
          2937 => x"ac",
          2938 => x"55",
          2939 => x"09",
          2940 => x"38",
          2941 => x"51",
          2942 => x"81",
          2943 => x"83",
          2944 => x"53",
          2945 => x"82",
          2946 => x"82",
          2947 => x"e0",
          2948 => x"ab",
          2949 => x"a4",
          2950 => x"0c",
          2951 => x"53",
          2952 => x"56",
          2953 => x"81",
          2954 => x"13",
          2955 => x"74",
          2956 => x"82",
          2957 => x"74",
          2958 => x"81",
          2959 => x"06",
          2960 => x"83",
          2961 => x"2a",
          2962 => x"72",
          2963 => x"26",
          2964 => x"ff",
          2965 => x"0c",
          2966 => x"15",
          2967 => x"0b",
          2968 => x"76",
          2969 => x"81",
          2970 => x"38",
          2971 => x"51",
          2972 => x"81",
          2973 => x"83",
          2974 => x"53",
          2975 => x"09",
          2976 => x"f9",
          2977 => x"52",
          2978 => x"b8",
          2979 => x"a4",
          2980 => x"38",
          2981 => x"08",
          2982 => x"84",
          2983 => x"d8",
          2984 => x"cb",
          2985 => x"ff",
          2986 => x"72",
          2987 => x"2e",
          2988 => x"80",
          2989 => x"14",
          2990 => x"3f",
          2991 => x"08",
          2992 => x"a4",
          2993 => x"81",
          2994 => x"84",
          2995 => x"d7",
          2996 => x"cb",
          2997 => x"8a",
          2998 => x"2e",
          2999 => x"9d",
          3000 => x"14",
          3001 => x"3f",
          3002 => x"08",
          3003 => x"84",
          3004 => x"d7",
          3005 => x"cb",
          3006 => x"15",
          3007 => x"34",
          3008 => x"22",
          3009 => x"72",
          3010 => x"23",
          3011 => x"23",
          3012 => x"15",
          3013 => x"75",
          3014 => x"0c",
          3015 => x"04",
          3016 => x"77",
          3017 => x"73",
          3018 => x"38",
          3019 => x"72",
          3020 => x"38",
          3021 => x"71",
          3022 => x"38",
          3023 => x"84",
          3024 => x"52",
          3025 => x"09",
          3026 => x"38",
          3027 => x"51",
          3028 => x"81",
          3029 => x"81",
          3030 => x"88",
          3031 => x"08",
          3032 => x"39",
          3033 => x"73",
          3034 => x"74",
          3035 => x"0c",
          3036 => x"04",
          3037 => x"02",
          3038 => x"7a",
          3039 => x"fc",
          3040 => x"f4",
          3041 => x"54",
          3042 => x"cb",
          3043 => x"bc",
          3044 => x"a4",
          3045 => x"81",
          3046 => x"70",
          3047 => x"73",
          3048 => x"38",
          3049 => x"78",
          3050 => x"2e",
          3051 => x"74",
          3052 => x"0c",
          3053 => x"80",
          3054 => x"80",
          3055 => x"70",
          3056 => x"51",
          3057 => x"81",
          3058 => x"54",
          3059 => x"a4",
          3060 => x"0d",
          3061 => x"0d",
          3062 => x"05",
          3063 => x"33",
          3064 => x"54",
          3065 => x"84",
          3066 => x"bf",
          3067 => x"98",
          3068 => x"53",
          3069 => x"05",
          3070 => x"fa",
          3071 => x"a4",
          3072 => x"cb",
          3073 => x"a4",
          3074 => x"68",
          3075 => x"70",
          3076 => x"c6",
          3077 => x"a4",
          3078 => x"cb",
          3079 => x"38",
          3080 => x"05",
          3081 => x"2b",
          3082 => x"80",
          3083 => x"86",
          3084 => x"06",
          3085 => x"2e",
          3086 => x"74",
          3087 => x"38",
          3088 => x"09",
          3089 => x"38",
          3090 => x"f8",
          3091 => x"a4",
          3092 => x"39",
          3093 => x"33",
          3094 => x"73",
          3095 => x"77",
          3096 => x"81",
          3097 => x"73",
          3098 => x"38",
          3099 => x"bc",
          3100 => x"07",
          3101 => x"b4",
          3102 => x"2a",
          3103 => x"51",
          3104 => x"2e",
          3105 => x"62",
          3106 => x"e8",
          3107 => x"cb",
          3108 => x"82",
          3109 => x"52",
          3110 => x"51",
          3111 => x"62",
          3112 => x"8b",
          3113 => x"53",
          3114 => x"51",
          3115 => x"80",
          3116 => x"05",
          3117 => x"3f",
          3118 => x"0b",
          3119 => x"75",
          3120 => x"f1",
          3121 => x"11",
          3122 => x"80",
          3123 => x"97",
          3124 => x"51",
          3125 => x"81",
          3126 => x"55",
          3127 => x"08",
          3128 => x"b7",
          3129 => x"c4",
          3130 => x"05",
          3131 => x"2a",
          3132 => x"51",
          3133 => x"80",
          3134 => x"84",
          3135 => x"39",
          3136 => x"70",
          3137 => x"54",
          3138 => x"a9",
          3139 => x"06",
          3140 => x"2e",
          3141 => x"55",
          3142 => x"73",
          3143 => x"d6",
          3144 => x"cb",
          3145 => x"ff",
          3146 => x"0c",
          3147 => x"cb",
          3148 => x"f8",
          3149 => x"2a",
          3150 => x"51",
          3151 => x"2e",
          3152 => x"80",
          3153 => x"7a",
          3154 => x"a0",
          3155 => x"a4",
          3156 => x"53",
          3157 => x"e6",
          3158 => x"cb",
          3159 => x"cb",
          3160 => x"1b",
          3161 => x"05",
          3162 => x"d3",
          3163 => x"a4",
          3164 => x"a4",
          3165 => x"0c",
          3166 => x"56",
          3167 => x"84",
          3168 => x"90",
          3169 => x"0b",
          3170 => x"80",
          3171 => x"0c",
          3172 => x"1a",
          3173 => x"2a",
          3174 => x"51",
          3175 => x"2e",
          3176 => x"81",
          3177 => x"80",
          3178 => x"38",
          3179 => x"08",
          3180 => x"8a",
          3181 => x"89",
          3182 => x"59",
          3183 => x"76",
          3184 => x"d7",
          3185 => x"cb",
          3186 => x"81",
          3187 => x"81",
          3188 => x"82",
          3189 => x"a4",
          3190 => x"09",
          3191 => x"38",
          3192 => x"78",
          3193 => x"30",
          3194 => x"80",
          3195 => x"77",
          3196 => x"38",
          3197 => x"06",
          3198 => x"c3",
          3199 => x"1a",
          3200 => x"38",
          3201 => x"06",
          3202 => x"2e",
          3203 => x"52",
          3204 => x"a6",
          3205 => x"a4",
          3206 => x"82",
          3207 => x"75",
          3208 => x"cb",
          3209 => x"9c",
          3210 => x"39",
          3211 => x"74",
          3212 => x"cb",
          3213 => x"3d",
          3214 => x"3d",
          3215 => x"65",
          3216 => x"5d",
          3217 => x"0c",
          3218 => x"05",
          3219 => x"f9",
          3220 => x"cb",
          3221 => x"81",
          3222 => x"8a",
          3223 => x"33",
          3224 => x"2e",
          3225 => x"56",
          3226 => x"90",
          3227 => x"06",
          3228 => x"74",
          3229 => x"b6",
          3230 => x"82",
          3231 => x"34",
          3232 => x"aa",
          3233 => x"91",
          3234 => x"56",
          3235 => x"8c",
          3236 => x"1a",
          3237 => x"74",
          3238 => x"38",
          3239 => x"80",
          3240 => x"38",
          3241 => x"70",
          3242 => x"56",
          3243 => x"b2",
          3244 => x"11",
          3245 => x"77",
          3246 => x"5b",
          3247 => x"38",
          3248 => x"88",
          3249 => x"8f",
          3250 => x"08",
          3251 => x"d5",
          3252 => x"cb",
          3253 => x"81",
          3254 => x"9f",
          3255 => x"2e",
          3256 => x"74",
          3257 => x"98",
          3258 => x"7e",
          3259 => x"3f",
          3260 => x"08",
          3261 => x"83",
          3262 => x"a4",
          3263 => x"89",
          3264 => x"77",
          3265 => x"d6",
          3266 => x"7f",
          3267 => x"58",
          3268 => x"75",
          3269 => x"75",
          3270 => x"77",
          3271 => x"7c",
          3272 => x"33",
          3273 => x"3f",
          3274 => x"08",
          3275 => x"7e",
          3276 => x"56",
          3277 => x"2e",
          3278 => x"16",
          3279 => x"55",
          3280 => x"94",
          3281 => x"53",
          3282 => x"b0",
          3283 => x"31",
          3284 => x"05",
          3285 => x"3f",
          3286 => x"56",
          3287 => x"9c",
          3288 => x"19",
          3289 => x"06",
          3290 => x"31",
          3291 => x"76",
          3292 => x"7b",
          3293 => x"08",
          3294 => x"d1",
          3295 => x"cb",
          3296 => x"81",
          3297 => x"94",
          3298 => x"ff",
          3299 => x"05",
          3300 => x"cf",
          3301 => x"76",
          3302 => x"17",
          3303 => x"1e",
          3304 => x"18",
          3305 => x"5e",
          3306 => x"39",
          3307 => x"81",
          3308 => x"90",
          3309 => x"f2",
          3310 => x"63",
          3311 => x"40",
          3312 => x"7e",
          3313 => x"fc",
          3314 => x"51",
          3315 => x"81",
          3316 => x"55",
          3317 => x"08",
          3318 => x"18",
          3319 => x"80",
          3320 => x"74",
          3321 => x"39",
          3322 => x"70",
          3323 => x"81",
          3324 => x"56",
          3325 => x"80",
          3326 => x"38",
          3327 => x"0b",
          3328 => x"82",
          3329 => x"39",
          3330 => x"19",
          3331 => x"83",
          3332 => x"18",
          3333 => x"56",
          3334 => x"27",
          3335 => x"09",
          3336 => x"2e",
          3337 => x"94",
          3338 => x"83",
          3339 => x"56",
          3340 => x"38",
          3341 => x"22",
          3342 => x"89",
          3343 => x"55",
          3344 => x"75",
          3345 => x"18",
          3346 => x"9c",
          3347 => x"85",
          3348 => x"08",
          3349 => x"d7",
          3350 => x"cb",
          3351 => x"81",
          3352 => x"80",
          3353 => x"38",
          3354 => x"ff",
          3355 => x"ff",
          3356 => x"38",
          3357 => x"0c",
          3358 => x"85",
          3359 => x"19",
          3360 => x"b0",
          3361 => x"19",
          3362 => x"81",
          3363 => x"74",
          3364 => x"3f",
          3365 => x"08",
          3366 => x"98",
          3367 => x"7e",
          3368 => x"3f",
          3369 => x"08",
          3370 => x"d2",
          3371 => x"a4",
          3372 => x"89",
          3373 => x"78",
          3374 => x"d5",
          3375 => x"7f",
          3376 => x"58",
          3377 => x"75",
          3378 => x"75",
          3379 => x"78",
          3380 => x"7c",
          3381 => x"33",
          3382 => x"3f",
          3383 => x"08",
          3384 => x"7e",
          3385 => x"78",
          3386 => x"74",
          3387 => x"38",
          3388 => x"b0",
          3389 => x"31",
          3390 => x"05",
          3391 => x"51",
          3392 => x"7e",
          3393 => x"83",
          3394 => x"89",
          3395 => x"db",
          3396 => x"08",
          3397 => x"26",
          3398 => x"51",
          3399 => x"81",
          3400 => x"fd",
          3401 => x"77",
          3402 => x"55",
          3403 => x"0c",
          3404 => x"83",
          3405 => x"80",
          3406 => x"55",
          3407 => x"83",
          3408 => x"9c",
          3409 => x"7e",
          3410 => x"3f",
          3411 => x"08",
          3412 => x"75",
          3413 => x"94",
          3414 => x"ff",
          3415 => x"05",
          3416 => x"3f",
          3417 => x"0b",
          3418 => x"7b",
          3419 => x"08",
          3420 => x"76",
          3421 => x"08",
          3422 => x"1c",
          3423 => x"08",
          3424 => x"5c",
          3425 => x"83",
          3426 => x"74",
          3427 => x"fd",
          3428 => x"18",
          3429 => x"07",
          3430 => x"19",
          3431 => x"75",
          3432 => x"0c",
          3433 => x"04",
          3434 => x"7a",
          3435 => x"05",
          3436 => x"56",
          3437 => x"81",
          3438 => x"57",
          3439 => x"08",
          3440 => x"90",
          3441 => x"86",
          3442 => x"06",
          3443 => x"73",
          3444 => x"e9",
          3445 => x"08",
          3446 => x"cc",
          3447 => x"cb",
          3448 => x"81",
          3449 => x"80",
          3450 => x"16",
          3451 => x"33",
          3452 => x"55",
          3453 => x"34",
          3454 => x"53",
          3455 => x"08",
          3456 => x"3f",
          3457 => x"52",
          3458 => x"c9",
          3459 => x"88",
          3460 => x"96",
          3461 => x"f0",
          3462 => x"92",
          3463 => x"ca",
          3464 => x"81",
          3465 => x"34",
          3466 => x"df",
          3467 => x"a4",
          3468 => x"33",
          3469 => x"55",
          3470 => x"17",
          3471 => x"cb",
          3472 => x"3d",
          3473 => x"3d",
          3474 => x"52",
          3475 => x"3f",
          3476 => x"08",
          3477 => x"a4",
          3478 => x"86",
          3479 => x"52",
          3480 => x"bc",
          3481 => x"a4",
          3482 => x"cb",
          3483 => x"38",
          3484 => x"08",
          3485 => x"81",
          3486 => x"86",
          3487 => x"ff",
          3488 => x"3d",
          3489 => x"3f",
          3490 => x"0b",
          3491 => x"08",
          3492 => x"81",
          3493 => x"81",
          3494 => x"80",
          3495 => x"cb",
          3496 => x"3d",
          3497 => x"3d",
          3498 => x"93",
          3499 => x"52",
          3500 => x"e9",
          3501 => x"cb",
          3502 => x"81",
          3503 => x"80",
          3504 => x"58",
          3505 => x"3d",
          3506 => x"e0",
          3507 => x"cb",
          3508 => x"81",
          3509 => x"bc",
          3510 => x"c7",
          3511 => x"98",
          3512 => x"73",
          3513 => x"38",
          3514 => x"12",
          3515 => x"39",
          3516 => x"33",
          3517 => x"70",
          3518 => x"55",
          3519 => x"2e",
          3520 => x"7f",
          3521 => x"54",
          3522 => x"81",
          3523 => x"94",
          3524 => x"39",
          3525 => x"08",
          3526 => x"81",
          3527 => x"85",
          3528 => x"cb",
          3529 => x"3d",
          3530 => x"3d",
          3531 => x"5b",
          3532 => x"34",
          3533 => x"3d",
          3534 => x"52",
          3535 => x"e8",
          3536 => x"cb",
          3537 => x"81",
          3538 => x"82",
          3539 => x"43",
          3540 => x"11",
          3541 => x"58",
          3542 => x"80",
          3543 => x"38",
          3544 => x"3d",
          3545 => x"d5",
          3546 => x"cb",
          3547 => x"81",
          3548 => x"82",
          3549 => x"52",
          3550 => x"c8",
          3551 => x"a4",
          3552 => x"cb",
          3553 => x"c1",
          3554 => x"7b",
          3555 => x"3f",
          3556 => x"08",
          3557 => x"74",
          3558 => x"3f",
          3559 => x"08",
          3560 => x"a4",
          3561 => x"38",
          3562 => x"51",
          3563 => x"81",
          3564 => x"57",
          3565 => x"08",
          3566 => x"52",
          3567 => x"f2",
          3568 => x"cb",
          3569 => x"a6",
          3570 => x"74",
          3571 => x"3f",
          3572 => x"08",
          3573 => x"a4",
          3574 => x"cc",
          3575 => x"2e",
          3576 => x"86",
          3577 => x"81",
          3578 => x"81",
          3579 => x"3d",
          3580 => x"52",
          3581 => x"c9",
          3582 => x"3d",
          3583 => x"11",
          3584 => x"5a",
          3585 => x"2e",
          3586 => x"b9",
          3587 => x"16",
          3588 => x"33",
          3589 => x"73",
          3590 => x"16",
          3591 => x"26",
          3592 => x"75",
          3593 => x"38",
          3594 => x"05",
          3595 => x"6f",
          3596 => x"ff",
          3597 => x"55",
          3598 => x"74",
          3599 => x"38",
          3600 => x"11",
          3601 => x"74",
          3602 => x"39",
          3603 => x"09",
          3604 => x"38",
          3605 => x"11",
          3606 => x"74",
          3607 => x"81",
          3608 => x"70",
          3609 => x"ba",
          3610 => x"08",
          3611 => x"5c",
          3612 => x"73",
          3613 => x"38",
          3614 => x"1a",
          3615 => x"55",
          3616 => x"38",
          3617 => x"73",
          3618 => x"38",
          3619 => x"76",
          3620 => x"74",
          3621 => x"33",
          3622 => x"05",
          3623 => x"15",
          3624 => x"ba",
          3625 => x"05",
          3626 => x"ff",
          3627 => x"06",
          3628 => x"57",
          3629 => x"18",
          3630 => x"54",
          3631 => x"70",
          3632 => x"34",
          3633 => x"ee",
          3634 => x"34",
          3635 => x"a4",
          3636 => x"0d",
          3637 => x"0d",
          3638 => x"3d",
          3639 => x"71",
          3640 => x"ec",
          3641 => x"cb",
          3642 => x"81",
          3643 => x"82",
          3644 => x"15",
          3645 => x"82",
          3646 => x"15",
          3647 => x"76",
          3648 => x"90",
          3649 => x"81",
          3650 => x"06",
          3651 => x"72",
          3652 => x"56",
          3653 => x"54",
          3654 => x"17",
          3655 => x"78",
          3656 => x"38",
          3657 => x"22",
          3658 => x"59",
          3659 => x"78",
          3660 => x"76",
          3661 => x"51",
          3662 => x"3f",
          3663 => x"08",
          3664 => x"54",
          3665 => x"53",
          3666 => x"3f",
          3667 => x"08",
          3668 => x"38",
          3669 => x"75",
          3670 => x"18",
          3671 => x"31",
          3672 => x"57",
          3673 => x"b1",
          3674 => x"08",
          3675 => x"38",
          3676 => x"51",
          3677 => x"81",
          3678 => x"54",
          3679 => x"08",
          3680 => x"9a",
          3681 => x"a4",
          3682 => x"81",
          3683 => x"cb",
          3684 => x"16",
          3685 => x"16",
          3686 => x"2e",
          3687 => x"76",
          3688 => x"dc",
          3689 => x"31",
          3690 => x"18",
          3691 => x"90",
          3692 => x"81",
          3693 => x"06",
          3694 => x"56",
          3695 => x"9a",
          3696 => x"74",
          3697 => x"3f",
          3698 => x"08",
          3699 => x"a4",
          3700 => x"81",
          3701 => x"56",
          3702 => x"52",
          3703 => x"84",
          3704 => x"a4",
          3705 => x"ff",
          3706 => x"81",
          3707 => x"38",
          3708 => x"98",
          3709 => x"a6",
          3710 => x"16",
          3711 => x"39",
          3712 => x"16",
          3713 => x"75",
          3714 => x"53",
          3715 => x"aa",
          3716 => x"79",
          3717 => x"3f",
          3718 => x"08",
          3719 => x"0b",
          3720 => x"82",
          3721 => x"39",
          3722 => x"16",
          3723 => x"bb",
          3724 => x"2a",
          3725 => x"08",
          3726 => x"15",
          3727 => x"15",
          3728 => x"90",
          3729 => x"16",
          3730 => x"33",
          3731 => x"53",
          3732 => x"34",
          3733 => x"06",
          3734 => x"2e",
          3735 => x"9c",
          3736 => x"85",
          3737 => x"16",
          3738 => x"72",
          3739 => x"0c",
          3740 => x"04",
          3741 => x"79",
          3742 => x"75",
          3743 => x"8a",
          3744 => x"89",
          3745 => x"52",
          3746 => x"05",
          3747 => x"3f",
          3748 => x"08",
          3749 => x"a4",
          3750 => x"38",
          3751 => x"7a",
          3752 => x"d8",
          3753 => x"cb",
          3754 => x"81",
          3755 => x"80",
          3756 => x"16",
          3757 => x"2b",
          3758 => x"74",
          3759 => x"86",
          3760 => x"84",
          3761 => x"06",
          3762 => x"73",
          3763 => x"38",
          3764 => x"52",
          3765 => x"da",
          3766 => x"a4",
          3767 => x"0c",
          3768 => x"14",
          3769 => x"23",
          3770 => x"51",
          3771 => x"81",
          3772 => x"55",
          3773 => x"09",
          3774 => x"38",
          3775 => x"39",
          3776 => x"84",
          3777 => x"0c",
          3778 => x"81",
          3779 => x"89",
          3780 => x"fc",
          3781 => x"87",
          3782 => x"53",
          3783 => x"e7",
          3784 => x"cb",
          3785 => x"38",
          3786 => x"08",
          3787 => x"3d",
          3788 => x"3d",
          3789 => x"89",
          3790 => x"54",
          3791 => x"54",
          3792 => x"81",
          3793 => x"53",
          3794 => x"08",
          3795 => x"74",
          3796 => x"cb",
          3797 => x"73",
          3798 => x"3f",
          3799 => x"08",
          3800 => x"39",
          3801 => x"08",
          3802 => x"d3",
          3803 => x"cb",
          3804 => x"81",
          3805 => x"84",
          3806 => x"06",
          3807 => x"53",
          3808 => x"cb",
          3809 => x"38",
          3810 => x"51",
          3811 => x"72",
          3812 => x"cf",
          3813 => x"cb",
          3814 => x"32",
          3815 => x"72",
          3816 => x"70",
          3817 => x"08",
          3818 => x"54",
          3819 => x"cb",
          3820 => x"3d",
          3821 => x"3d",
          3822 => x"80",
          3823 => x"70",
          3824 => x"52",
          3825 => x"3f",
          3826 => x"08",
          3827 => x"a4",
          3828 => x"64",
          3829 => x"d6",
          3830 => x"cb",
          3831 => x"81",
          3832 => x"a0",
          3833 => x"cb",
          3834 => x"98",
          3835 => x"73",
          3836 => x"38",
          3837 => x"39",
          3838 => x"88",
          3839 => x"75",
          3840 => x"3f",
          3841 => x"a4",
          3842 => x"0d",
          3843 => x"0d",
          3844 => x"5c",
          3845 => x"3d",
          3846 => x"93",
          3847 => x"d6",
          3848 => x"a4",
          3849 => x"cb",
          3850 => x"80",
          3851 => x"0c",
          3852 => x"11",
          3853 => x"90",
          3854 => x"56",
          3855 => x"74",
          3856 => x"75",
          3857 => x"e4",
          3858 => x"81",
          3859 => x"5b",
          3860 => x"81",
          3861 => x"75",
          3862 => x"73",
          3863 => x"81",
          3864 => x"82",
          3865 => x"76",
          3866 => x"f0",
          3867 => x"f4",
          3868 => x"a4",
          3869 => x"d1",
          3870 => x"a4",
          3871 => x"ce",
          3872 => x"a4",
          3873 => x"81",
          3874 => x"07",
          3875 => x"05",
          3876 => x"53",
          3877 => x"98",
          3878 => x"26",
          3879 => x"f9",
          3880 => x"08",
          3881 => x"08",
          3882 => x"98",
          3883 => x"81",
          3884 => x"58",
          3885 => x"3f",
          3886 => x"08",
          3887 => x"a4",
          3888 => x"38",
          3889 => x"77",
          3890 => x"5d",
          3891 => x"74",
          3892 => x"81",
          3893 => x"b4",
          3894 => x"bb",
          3895 => x"cb",
          3896 => x"ff",
          3897 => x"30",
          3898 => x"1b",
          3899 => x"5b",
          3900 => x"39",
          3901 => x"ff",
          3902 => x"81",
          3903 => x"f0",
          3904 => x"30",
          3905 => x"1b",
          3906 => x"5b",
          3907 => x"83",
          3908 => x"58",
          3909 => x"92",
          3910 => x"0c",
          3911 => x"12",
          3912 => x"33",
          3913 => x"54",
          3914 => x"34",
          3915 => x"a4",
          3916 => x"0d",
          3917 => x"0d",
          3918 => x"fc",
          3919 => x"52",
          3920 => x"3f",
          3921 => x"08",
          3922 => x"a4",
          3923 => x"38",
          3924 => x"56",
          3925 => x"38",
          3926 => x"70",
          3927 => x"81",
          3928 => x"55",
          3929 => x"80",
          3930 => x"38",
          3931 => x"54",
          3932 => x"08",
          3933 => x"38",
          3934 => x"81",
          3935 => x"53",
          3936 => x"52",
          3937 => x"8c",
          3938 => x"a4",
          3939 => x"19",
          3940 => x"c9",
          3941 => x"08",
          3942 => x"ff",
          3943 => x"81",
          3944 => x"ff",
          3945 => x"06",
          3946 => x"56",
          3947 => x"08",
          3948 => x"81",
          3949 => x"82",
          3950 => x"75",
          3951 => x"54",
          3952 => x"08",
          3953 => x"27",
          3954 => x"17",
          3955 => x"cb",
          3956 => x"76",
          3957 => x"3f",
          3958 => x"08",
          3959 => x"08",
          3960 => x"90",
          3961 => x"c0",
          3962 => x"90",
          3963 => x"80",
          3964 => x"75",
          3965 => x"75",
          3966 => x"cb",
          3967 => x"3d",
          3968 => x"3d",
          3969 => x"a0",
          3970 => x"05",
          3971 => x"51",
          3972 => x"81",
          3973 => x"55",
          3974 => x"08",
          3975 => x"78",
          3976 => x"08",
          3977 => x"70",
          3978 => x"ae",
          3979 => x"a4",
          3980 => x"cb",
          3981 => x"db",
          3982 => x"fb",
          3983 => x"85",
          3984 => x"06",
          3985 => x"86",
          3986 => x"c7",
          3987 => x"2b",
          3988 => x"24",
          3989 => x"02",
          3990 => x"33",
          3991 => x"58",
          3992 => x"76",
          3993 => x"6b",
          3994 => x"cc",
          3995 => x"cb",
          3996 => x"84",
          3997 => x"06",
          3998 => x"73",
          3999 => x"d4",
          4000 => x"81",
          4001 => x"94",
          4002 => x"81",
          4003 => x"5a",
          4004 => x"08",
          4005 => x"8a",
          4006 => x"54",
          4007 => x"81",
          4008 => x"55",
          4009 => x"08",
          4010 => x"81",
          4011 => x"52",
          4012 => x"e5",
          4013 => x"a4",
          4014 => x"cb",
          4015 => x"38",
          4016 => x"cf",
          4017 => x"a4",
          4018 => x"88",
          4019 => x"a4",
          4020 => x"38",
          4021 => x"c2",
          4022 => x"a4",
          4023 => x"a4",
          4024 => x"81",
          4025 => x"07",
          4026 => x"55",
          4027 => x"2e",
          4028 => x"80",
          4029 => x"80",
          4030 => x"77",
          4031 => x"3f",
          4032 => x"08",
          4033 => x"38",
          4034 => x"ba",
          4035 => x"cb",
          4036 => x"74",
          4037 => x"0c",
          4038 => x"04",
          4039 => x"82",
          4040 => x"c0",
          4041 => x"3d",
          4042 => x"3f",
          4043 => x"08",
          4044 => x"a4",
          4045 => x"38",
          4046 => x"52",
          4047 => x"52",
          4048 => x"3f",
          4049 => x"08",
          4050 => x"a4",
          4051 => x"88",
          4052 => x"39",
          4053 => x"08",
          4054 => x"81",
          4055 => x"38",
          4056 => x"05",
          4057 => x"2a",
          4058 => x"55",
          4059 => x"81",
          4060 => x"5a",
          4061 => x"3d",
          4062 => x"c1",
          4063 => x"cb",
          4064 => x"55",
          4065 => x"a4",
          4066 => x"87",
          4067 => x"a4",
          4068 => x"09",
          4069 => x"38",
          4070 => x"cb",
          4071 => x"2e",
          4072 => x"86",
          4073 => x"81",
          4074 => x"81",
          4075 => x"cb",
          4076 => x"78",
          4077 => x"3f",
          4078 => x"08",
          4079 => x"a4",
          4080 => x"38",
          4081 => x"52",
          4082 => x"ff",
          4083 => x"78",
          4084 => x"b4",
          4085 => x"54",
          4086 => x"15",
          4087 => x"b2",
          4088 => x"ca",
          4089 => x"b6",
          4090 => x"53",
          4091 => x"53",
          4092 => x"3f",
          4093 => x"b4",
          4094 => x"d4",
          4095 => x"b6",
          4096 => x"54",
          4097 => x"d5",
          4098 => x"53",
          4099 => x"11",
          4100 => x"d7",
          4101 => x"81",
          4102 => x"34",
          4103 => x"a4",
          4104 => x"a4",
          4105 => x"cb",
          4106 => x"38",
          4107 => x"0a",
          4108 => x"05",
          4109 => x"d0",
          4110 => x"64",
          4111 => x"c9",
          4112 => x"54",
          4113 => x"15",
          4114 => x"81",
          4115 => x"34",
          4116 => x"b8",
          4117 => x"cb",
          4118 => x"8b",
          4119 => x"75",
          4120 => x"ff",
          4121 => x"73",
          4122 => x"0c",
          4123 => x"04",
          4124 => x"a9",
          4125 => x"51",
          4126 => x"82",
          4127 => x"ff",
          4128 => x"a9",
          4129 => x"ee",
          4130 => x"a4",
          4131 => x"cb",
          4132 => x"d3",
          4133 => x"a9",
          4134 => x"9d",
          4135 => x"58",
          4136 => x"81",
          4137 => x"55",
          4138 => x"08",
          4139 => x"02",
          4140 => x"33",
          4141 => x"54",
          4142 => x"82",
          4143 => x"53",
          4144 => x"52",
          4145 => x"88",
          4146 => x"b4",
          4147 => x"53",
          4148 => x"3d",
          4149 => x"ff",
          4150 => x"aa",
          4151 => x"73",
          4152 => x"3f",
          4153 => x"08",
          4154 => x"a4",
          4155 => x"63",
          4156 => x"81",
          4157 => x"65",
          4158 => x"2e",
          4159 => x"55",
          4160 => x"81",
          4161 => x"84",
          4162 => x"06",
          4163 => x"73",
          4164 => x"3f",
          4165 => x"08",
          4166 => x"a4",
          4167 => x"38",
          4168 => x"53",
          4169 => x"95",
          4170 => x"16",
          4171 => x"87",
          4172 => x"05",
          4173 => x"34",
          4174 => x"70",
          4175 => x"81",
          4176 => x"55",
          4177 => x"74",
          4178 => x"73",
          4179 => x"78",
          4180 => x"83",
          4181 => x"16",
          4182 => x"2a",
          4183 => x"51",
          4184 => x"80",
          4185 => x"38",
          4186 => x"80",
          4187 => x"52",
          4188 => x"be",
          4189 => x"a4",
          4190 => x"51",
          4191 => x"3f",
          4192 => x"cb",
          4193 => x"2e",
          4194 => x"81",
          4195 => x"52",
          4196 => x"b5",
          4197 => x"cb",
          4198 => x"80",
          4199 => x"58",
          4200 => x"a4",
          4201 => x"38",
          4202 => x"54",
          4203 => x"09",
          4204 => x"38",
          4205 => x"52",
          4206 => x"af",
          4207 => x"81",
          4208 => x"34",
          4209 => x"cb",
          4210 => x"38",
          4211 => x"ca",
          4212 => x"a4",
          4213 => x"cb",
          4214 => x"38",
          4215 => x"b5",
          4216 => x"cb",
          4217 => x"74",
          4218 => x"0c",
          4219 => x"04",
          4220 => x"02",
          4221 => x"33",
          4222 => x"80",
          4223 => x"57",
          4224 => x"95",
          4225 => x"52",
          4226 => x"d2",
          4227 => x"cb",
          4228 => x"81",
          4229 => x"80",
          4230 => x"5a",
          4231 => x"3d",
          4232 => x"c9",
          4233 => x"cb",
          4234 => x"81",
          4235 => x"b8",
          4236 => x"cf",
          4237 => x"a0",
          4238 => x"55",
          4239 => x"75",
          4240 => x"71",
          4241 => x"33",
          4242 => x"74",
          4243 => x"57",
          4244 => x"8b",
          4245 => x"54",
          4246 => x"15",
          4247 => x"ff",
          4248 => x"81",
          4249 => x"55",
          4250 => x"a4",
          4251 => x"0d",
          4252 => x"0d",
          4253 => x"53",
          4254 => x"05",
          4255 => x"51",
          4256 => x"81",
          4257 => x"55",
          4258 => x"08",
          4259 => x"76",
          4260 => x"93",
          4261 => x"51",
          4262 => x"81",
          4263 => x"55",
          4264 => x"08",
          4265 => x"80",
          4266 => x"81",
          4267 => x"86",
          4268 => x"38",
          4269 => x"86",
          4270 => x"90",
          4271 => x"54",
          4272 => x"ff",
          4273 => x"76",
          4274 => x"83",
          4275 => x"51",
          4276 => x"3f",
          4277 => x"08",
          4278 => x"cb",
          4279 => x"3d",
          4280 => x"3d",
          4281 => x"5c",
          4282 => x"98",
          4283 => x"52",
          4284 => x"d1",
          4285 => x"cb",
          4286 => x"cb",
          4287 => x"70",
          4288 => x"08",
          4289 => x"51",
          4290 => x"80",
          4291 => x"38",
          4292 => x"06",
          4293 => x"80",
          4294 => x"38",
          4295 => x"5f",
          4296 => x"3d",
          4297 => x"ff",
          4298 => x"81",
          4299 => x"57",
          4300 => x"08",
          4301 => x"74",
          4302 => x"c3",
          4303 => x"cb",
          4304 => x"81",
          4305 => x"bf",
          4306 => x"a4",
          4307 => x"a4",
          4308 => x"59",
          4309 => x"81",
          4310 => x"56",
          4311 => x"33",
          4312 => x"16",
          4313 => x"27",
          4314 => x"56",
          4315 => x"80",
          4316 => x"80",
          4317 => x"ff",
          4318 => x"70",
          4319 => x"56",
          4320 => x"e8",
          4321 => x"76",
          4322 => x"81",
          4323 => x"80",
          4324 => x"57",
          4325 => x"78",
          4326 => x"51",
          4327 => x"2e",
          4328 => x"73",
          4329 => x"38",
          4330 => x"08",
          4331 => x"b1",
          4332 => x"cb",
          4333 => x"81",
          4334 => x"a7",
          4335 => x"33",
          4336 => x"c3",
          4337 => x"2e",
          4338 => x"e4",
          4339 => x"2e",
          4340 => x"56",
          4341 => x"05",
          4342 => x"e3",
          4343 => x"a4",
          4344 => x"76",
          4345 => x"0c",
          4346 => x"04",
          4347 => x"82",
          4348 => x"ff",
          4349 => x"9d",
          4350 => x"fa",
          4351 => x"a4",
          4352 => x"a4",
          4353 => x"81",
          4354 => x"83",
          4355 => x"53",
          4356 => x"3d",
          4357 => x"ff",
          4358 => x"73",
          4359 => x"70",
          4360 => x"52",
          4361 => x"9f",
          4362 => x"bc",
          4363 => x"74",
          4364 => x"6d",
          4365 => x"70",
          4366 => x"af",
          4367 => x"cb",
          4368 => x"2e",
          4369 => x"70",
          4370 => x"57",
          4371 => x"fd",
          4372 => x"a4",
          4373 => x"8d",
          4374 => x"2b",
          4375 => x"81",
          4376 => x"86",
          4377 => x"a4",
          4378 => x"9f",
          4379 => x"ff",
          4380 => x"54",
          4381 => x"8a",
          4382 => x"70",
          4383 => x"06",
          4384 => x"ff",
          4385 => x"38",
          4386 => x"15",
          4387 => x"80",
          4388 => x"74",
          4389 => x"80",
          4390 => x"89",
          4391 => x"a4",
          4392 => x"81",
          4393 => x"88",
          4394 => x"26",
          4395 => x"39",
          4396 => x"86",
          4397 => x"81",
          4398 => x"ff",
          4399 => x"38",
          4400 => x"54",
          4401 => x"81",
          4402 => x"81",
          4403 => x"78",
          4404 => x"5a",
          4405 => x"6d",
          4406 => x"81",
          4407 => x"57",
          4408 => x"9f",
          4409 => x"38",
          4410 => x"54",
          4411 => x"81",
          4412 => x"b1",
          4413 => x"2e",
          4414 => x"a7",
          4415 => x"15",
          4416 => x"54",
          4417 => x"09",
          4418 => x"38",
          4419 => x"76",
          4420 => x"41",
          4421 => x"52",
          4422 => x"52",
          4423 => x"b3",
          4424 => x"a4",
          4425 => x"cb",
          4426 => x"f7",
          4427 => x"74",
          4428 => x"e5",
          4429 => x"a4",
          4430 => x"cb",
          4431 => x"38",
          4432 => x"38",
          4433 => x"74",
          4434 => x"39",
          4435 => x"08",
          4436 => x"81",
          4437 => x"38",
          4438 => x"74",
          4439 => x"38",
          4440 => x"51",
          4441 => x"3f",
          4442 => x"08",
          4443 => x"a4",
          4444 => x"a0",
          4445 => x"a4",
          4446 => x"51",
          4447 => x"3f",
          4448 => x"0b",
          4449 => x"8b",
          4450 => x"67",
          4451 => x"a7",
          4452 => x"81",
          4453 => x"34",
          4454 => x"ad",
          4455 => x"cb",
          4456 => x"73",
          4457 => x"cb",
          4458 => x"3d",
          4459 => x"3d",
          4460 => x"02",
          4461 => x"cb",
          4462 => x"3d",
          4463 => x"72",
          4464 => x"5a",
          4465 => x"81",
          4466 => x"58",
          4467 => x"08",
          4468 => x"91",
          4469 => x"77",
          4470 => x"7c",
          4471 => x"38",
          4472 => x"59",
          4473 => x"90",
          4474 => x"81",
          4475 => x"06",
          4476 => x"73",
          4477 => x"54",
          4478 => x"82",
          4479 => x"39",
          4480 => x"8b",
          4481 => x"11",
          4482 => x"2b",
          4483 => x"54",
          4484 => x"ff",
          4485 => x"ff",
          4486 => x"70",
          4487 => x"07",
          4488 => x"cb",
          4489 => x"8c",
          4490 => x"40",
          4491 => x"55",
          4492 => x"88",
          4493 => x"08",
          4494 => x"38",
          4495 => x"77",
          4496 => x"56",
          4497 => x"51",
          4498 => x"3f",
          4499 => x"55",
          4500 => x"08",
          4501 => x"38",
          4502 => x"cb",
          4503 => x"2e",
          4504 => x"81",
          4505 => x"ff",
          4506 => x"38",
          4507 => x"08",
          4508 => x"16",
          4509 => x"2e",
          4510 => x"87",
          4511 => x"74",
          4512 => x"74",
          4513 => x"81",
          4514 => x"38",
          4515 => x"ff",
          4516 => x"2e",
          4517 => x"7b",
          4518 => x"80",
          4519 => x"81",
          4520 => x"81",
          4521 => x"06",
          4522 => x"56",
          4523 => x"52",
          4524 => x"af",
          4525 => x"cb",
          4526 => x"81",
          4527 => x"80",
          4528 => x"81",
          4529 => x"56",
          4530 => x"d3",
          4531 => x"ff",
          4532 => x"7c",
          4533 => x"55",
          4534 => x"b3",
          4535 => x"1b",
          4536 => x"1b",
          4537 => x"33",
          4538 => x"54",
          4539 => x"34",
          4540 => x"fe",
          4541 => x"08",
          4542 => x"74",
          4543 => x"75",
          4544 => x"16",
          4545 => x"33",
          4546 => x"73",
          4547 => x"77",
          4548 => x"cb",
          4549 => x"3d",
          4550 => x"3d",
          4551 => x"02",
          4552 => x"eb",
          4553 => x"3d",
          4554 => x"59",
          4555 => x"8b",
          4556 => x"81",
          4557 => x"24",
          4558 => x"81",
          4559 => x"84",
          4560 => x"c0",
          4561 => x"51",
          4562 => x"2e",
          4563 => x"75",
          4564 => x"a4",
          4565 => x"06",
          4566 => x"7e",
          4567 => x"d0",
          4568 => x"a4",
          4569 => x"06",
          4570 => x"56",
          4571 => x"74",
          4572 => x"76",
          4573 => x"81",
          4574 => x"8a",
          4575 => x"b2",
          4576 => x"fc",
          4577 => x"52",
          4578 => x"a4",
          4579 => x"cb",
          4580 => x"38",
          4581 => x"80",
          4582 => x"74",
          4583 => x"26",
          4584 => x"15",
          4585 => x"74",
          4586 => x"38",
          4587 => x"80",
          4588 => x"84",
          4589 => x"92",
          4590 => x"80",
          4591 => x"38",
          4592 => x"06",
          4593 => x"2e",
          4594 => x"56",
          4595 => x"78",
          4596 => x"89",
          4597 => x"2b",
          4598 => x"43",
          4599 => x"38",
          4600 => x"30",
          4601 => x"77",
          4602 => x"91",
          4603 => x"c2",
          4604 => x"f8",
          4605 => x"52",
          4606 => x"a4",
          4607 => x"56",
          4608 => x"08",
          4609 => x"77",
          4610 => x"77",
          4611 => x"a4",
          4612 => x"45",
          4613 => x"bf",
          4614 => x"8e",
          4615 => x"26",
          4616 => x"74",
          4617 => x"48",
          4618 => x"75",
          4619 => x"38",
          4620 => x"81",
          4621 => x"fa",
          4622 => x"2a",
          4623 => x"56",
          4624 => x"2e",
          4625 => x"87",
          4626 => x"82",
          4627 => x"38",
          4628 => x"55",
          4629 => x"83",
          4630 => x"81",
          4631 => x"56",
          4632 => x"80",
          4633 => x"38",
          4634 => x"83",
          4635 => x"06",
          4636 => x"78",
          4637 => x"91",
          4638 => x"0b",
          4639 => x"22",
          4640 => x"80",
          4641 => x"74",
          4642 => x"38",
          4643 => x"56",
          4644 => x"17",
          4645 => x"57",
          4646 => x"2e",
          4647 => x"75",
          4648 => x"79",
          4649 => x"fe",
          4650 => x"81",
          4651 => x"84",
          4652 => x"05",
          4653 => x"5e",
          4654 => x"80",
          4655 => x"a4",
          4656 => x"8a",
          4657 => x"fd",
          4658 => x"75",
          4659 => x"38",
          4660 => x"78",
          4661 => x"8c",
          4662 => x"0b",
          4663 => x"22",
          4664 => x"80",
          4665 => x"74",
          4666 => x"38",
          4667 => x"56",
          4668 => x"17",
          4669 => x"57",
          4670 => x"2e",
          4671 => x"75",
          4672 => x"79",
          4673 => x"fe",
          4674 => x"81",
          4675 => x"10",
          4676 => x"81",
          4677 => x"9f",
          4678 => x"38",
          4679 => x"cb",
          4680 => x"81",
          4681 => x"05",
          4682 => x"2a",
          4683 => x"56",
          4684 => x"17",
          4685 => x"81",
          4686 => x"60",
          4687 => x"65",
          4688 => x"12",
          4689 => x"30",
          4690 => x"74",
          4691 => x"59",
          4692 => x"7d",
          4693 => x"81",
          4694 => x"76",
          4695 => x"41",
          4696 => x"76",
          4697 => x"90",
          4698 => x"62",
          4699 => x"51",
          4700 => x"26",
          4701 => x"75",
          4702 => x"31",
          4703 => x"65",
          4704 => x"fe",
          4705 => x"81",
          4706 => x"58",
          4707 => x"09",
          4708 => x"38",
          4709 => x"08",
          4710 => x"26",
          4711 => x"78",
          4712 => x"79",
          4713 => x"78",
          4714 => x"86",
          4715 => x"82",
          4716 => x"06",
          4717 => x"83",
          4718 => x"81",
          4719 => x"27",
          4720 => x"8f",
          4721 => x"55",
          4722 => x"26",
          4723 => x"59",
          4724 => x"62",
          4725 => x"74",
          4726 => x"38",
          4727 => x"88",
          4728 => x"a4",
          4729 => x"26",
          4730 => x"86",
          4731 => x"1a",
          4732 => x"79",
          4733 => x"38",
          4734 => x"80",
          4735 => x"2e",
          4736 => x"83",
          4737 => x"9f",
          4738 => x"8b",
          4739 => x"06",
          4740 => x"74",
          4741 => x"84",
          4742 => x"52",
          4743 => x"a2",
          4744 => x"53",
          4745 => x"52",
          4746 => x"a2",
          4747 => x"80",
          4748 => x"51",
          4749 => x"3f",
          4750 => x"34",
          4751 => x"ff",
          4752 => x"1b",
          4753 => x"a2",
          4754 => x"90",
          4755 => x"83",
          4756 => x"70",
          4757 => x"80",
          4758 => x"55",
          4759 => x"ff",
          4760 => x"66",
          4761 => x"ff",
          4762 => x"38",
          4763 => x"ff",
          4764 => x"1b",
          4765 => x"f2",
          4766 => x"74",
          4767 => x"51",
          4768 => x"3f",
          4769 => x"1c",
          4770 => x"98",
          4771 => x"a0",
          4772 => x"ff",
          4773 => x"51",
          4774 => x"3f",
          4775 => x"1b",
          4776 => x"e4",
          4777 => x"2e",
          4778 => x"80",
          4779 => x"88",
          4780 => x"80",
          4781 => x"ff",
          4782 => x"7c",
          4783 => x"51",
          4784 => x"3f",
          4785 => x"1b",
          4786 => x"bc",
          4787 => x"b0",
          4788 => x"a0",
          4789 => x"52",
          4790 => x"ff",
          4791 => x"ff",
          4792 => x"c0",
          4793 => x"0b",
          4794 => x"34",
          4795 => x"ba",
          4796 => x"c7",
          4797 => x"39",
          4798 => x"0a",
          4799 => x"51",
          4800 => x"3f",
          4801 => x"ff",
          4802 => x"1b",
          4803 => x"da",
          4804 => x"0b",
          4805 => x"a9",
          4806 => x"34",
          4807 => x"ba",
          4808 => x"1b",
          4809 => x"8f",
          4810 => x"d5",
          4811 => x"1b",
          4812 => x"ff",
          4813 => x"81",
          4814 => x"7a",
          4815 => x"ff",
          4816 => x"81",
          4817 => x"a4",
          4818 => x"38",
          4819 => x"09",
          4820 => x"ee",
          4821 => x"60",
          4822 => x"7a",
          4823 => x"ff",
          4824 => x"84",
          4825 => x"52",
          4826 => x"9f",
          4827 => x"8b",
          4828 => x"52",
          4829 => x"9f",
          4830 => x"8a",
          4831 => x"52",
          4832 => x"51",
          4833 => x"3f",
          4834 => x"83",
          4835 => x"ff",
          4836 => x"82",
          4837 => x"1b",
          4838 => x"ec",
          4839 => x"d5",
          4840 => x"ff",
          4841 => x"75",
          4842 => x"05",
          4843 => x"7e",
          4844 => x"e5",
          4845 => x"60",
          4846 => x"52",
          4847 => x"9a",
          4848 => x"53",
          4849 => x"51",
          4850 => x"3f",
          4851 => x"58",
          4852 => x"09",
          4853 => x"38",
          4854 => x"51",
          4855 => x"3f",
          4856 => x"1b",
          4857 => x"a0",
          4858 => x"52",
          4859 => x"91",
          4860 => x"ff",
          4861 => x"81",
          4862 => x"f8",
          4863 => x"7a",
          4864 => x"84",
          4865 => x"61",
          4866 => x"26",
          4867 => x"57",
          4868 => x"53",
          4869 => x"51",
          4870 => x"3f",
          4871 => x"08",
          4872 => x"84",
          4873 => x"cb",
          4874 => x"7a",
          4875 => x"aa",
          4876 => x"75",
          4877 => x"56",
          4878 => x"81",
          4879 => x"80",
          4880 => x"38",
          4881 => x"83",
          4882 => x"63",
          4883 => x"74",
          4884 => x"38",
          4885 => x"54",
          4886 => x"52",
          4887 => x"99",
          4888 => x"cb",
          4889 => x"c1",
          4890 => x"75",
          4891 => x"56",
          4892 => x"8c",
          4893 => x"2e",
          4894 => x"56",
          4895 => x"ff",
          4896 => x"84",
          4897 => x"2e",
          4898 => x"56",
          4899 => x"58",
          4900 => x"38",
          4901 => x"77",
          4902 => x"ff",
          4903 => x"82",
          4904 => x"78",
          4905 => x"c2",
          4906 => x"1b",
          4907 => x"34",
          4908 => x"16",
          4909 => x"82",
          4910 => x"83",
          4911 => x"84",
          4912 => x"67",
          4913 => x"fd",
          4914 => x"51",
          4915 => x"3f",
          4916 => x"16",
          4917 => x"a4",
          4918 => x"bf",
          4919 => x"86",
          4920 => x"cb",
          4921 => x"16",
          4922 => x"83",
          4923 => x"ff",
          4924 => x"66",
          4925 => x"1b",
          4926 => x"8c",
          4927 => x"77",
          4928 => x"7e",
          4929 => x"91",
          4930 => x"81",
          4931 => x"a2",
          4932 => x"80",
          4933 => x"ff",
          4934 => x"81",
          4935 => x"a4",
          4936 => x"89",
          4937 => x"8a",
          4938 => x"86",
          4939 => x"a4",
          4940 => x"81",
          4941 => x"99",
          4942 => x"ff",
          4943 => x"52",
          4944 => x"81",
          4945 => x"84",
          4946 => x"88",
          4947 => x"08",
          4948 => x"bc",
          4949 => x"39",
          4950 => x"51",
          4951 => x"81",
          4952 => x"80",
          4953 => x"bd",
          4954 => x"eb",
          4955 => x"80",
          4956 => x"39",
          4957 => x"51",
          4958 => x"81",
          4959 => x"80",
          4960 => x"be",
          4961 => x"cf",
          4962 => x"cc",
          4963 => x"39",
          4964 => x"51",
          4965 => x"81",
          4966 => x"bb",
          4967 => x"98",
          4968 => x"81",
          4969 => x"af",
          4970 => x"d8",
          4971 => x"81",
          4972 => x"a3",
          4973 => x"8c",
          4974 => x"81",
          4975 => x"97",
          4976 => x"b8",
          4977 => x"81",
          4978 => x"8b",
          4979 => x"e8",
          4980 => x"81",
          4981 => x"ff",
          4982 => x"83",
          4983 => x"fb",
          4984 => x"79",
          4985 => x"87",
          4986 => x"38",
          4987 => x"87",
          4988 => x"91",
          4989 => x"52",
          4990 => x"f2",
          4991 => x"cb",
          4992 => x"75",
          4993 => x"98",
          4994 => x"a4",
          4995 => x"53",
          4996 => x"c1",
          4997 => x"8d",
          4998 => x"3d",
          4999 => x"3d",
          5000 => x"61",
          5001 => x"80",
          5002 => x"73",
          5003 => x"5f",
          5004 => x"5c",
          5005 => x"52",
          5006 => x"51",
          5007 => x"3f",
          5008 => x"51",
          5009 => x"3f",
          5010 => x"77",
          5011 => x"38",
          5012 => x"89",
          5013 => x"2e",
          5014 => x"c6",
          5015 => x"53",
          5016 => x"8e",
          5017 => x"52",
          5018 => x"51",
          5019 => x"3f",
          5020 => x"c1",
          5021 => x"86",
          5022 => x"15",
          5023 => x"39",
          5024 => x"72",
          5025 => x"38",
          5026 => x"81",
          5027 => x"ff",
          5028 => x"89",
          5029 => x"bc",
          5030 => x"b9",
          5031 => x"55",
          5032 => x"16",
          5033 => x"27",
          5034 => x"33",
          5035 => x"c8",
          5036 => x"85",
          5037 => x"81",
          5038 => x"ff",
          5039 => x"81",
          5040 => x"51",
          5041 => x"3f",
          5042 => x"81",
          5043 => x"ff",
          5044 => x"80",
          5045 => x"27",
          5046 => x"16",
          5047 => x"72",
          5048 => x"53",
          5049 => x"90",
          5050 => x"2e",
          5051 => x"80",
          5052 => x"38",
          5053 => x"39",
          5054 => x"f9",
          5055 => x"15",
          5056 => x"81",
          5057 => x"ff",
          5058 => x"76",
          5059 => x"5a",
          5060 => x"92",
          5061 => x"a4",
          5062 => x"70",
          5063 => x"55",
          5064 => x"09",
          5065 => x"38",
          5066 => x"3f",
          5067 => x"08",
          5068 => x"98",
          5069 => x"32",
          5070 => x"72",
          5071 => x"51",
          5072 => x"55",
          5073 => x"8c",
          5074 => x"38",
          5075 => x"09",
          5076 => x"38",
          5077 => x"39",
          5078 => x"72",
          5079 => x"d6",
          5080 => x"72",
          5081 => x"0c",
          5082 => x"04",
          5083 => x"66",
          5084 => x"80",
          5085 => x"69",
          5086 => x"74",
          5087 => x"70",
          5088 => x"27",
          5089 => x"58",
          5090 => x"93",
          5091 => x"fb",
          5092 => x"75",
          5093 => x"70",
          5094 => x"b9",
          5095 => x"a4",
          5096 => x"cb",
          5097 => x"38",
          5098 => x"08",
          5099 => x"88",
          5100 => x"a4",
          5101 => x"3d",
          5102 => x"84",
          5103 => x"52",
          5104 => x"f6",
          5105 => x"a4",
          5106 => x"cb",
          5107 => x"38",
          5108 => x"80",
          5109 => x"74",
          5110 => x"59",
          5111 => x"96",
          5112 => x"51",
          5113 => x"75",
          5114 => x"07",
          5115 => x"55",
          5116 => x"95",
          5117 => x"2e",
          5118 => x"c1",
          5119 => x"c0",
          5120 => x"52",
          5121 => x"d7",
          5122 => x"76",
          5123 => x"0c",
          5124 => x"04",
          5125 => x"7b",
          5126 => x"b3",
          5127 => x"58",
          5128 => x"53",
          5129 => x"51",
          5130 => x"81",
          5131 => x"a4",
          5132 => x"2e",
          5133 => x"81",
          5134 => x"98",
          5135 => x"7f",
          5136 => x"a4",
          5137 => x"7d",
          5138 => x"81",
          5139 => x"57",
          5140 => x"04",
          5141 => x"a4",
          5142 => x"0d",
          5143 => x"0d",
          5144 => x"33",
          5145 => x"53",
          5146 => x"52",
          5147 => x"c9",
          5148 => x"b4",
          5149 => x"80",
          5150 => x"c1",
          5151 => x"c2",
          5152 => x"c8",
          5153 => x"81",
          5154 => x"ff",
          5155 => x"74",
          5156 => x"38",
          5157 => x"3f",
          5158 => x"04",
          5159 => x"87",
          5160 => x"08",
          5161 => x"fd",
          5162 => x"fe",
          5163 => x"81",
          5164 => x"fe",
          5165 => x"80",
          5166 => x"fe",
          5167 => x"2a",
          5168 => x"51",
          5169 => x"2e",
          5170 => x"51",
          5171 => x"3f",
          5172 => x"51",
          5173 => x"3f",
          5174 => x"f5",
          5175 => x"82",
          5176 => x"06",
          5177 => x"80",
          5178 => x"81",
          5179 => x"ca",
          5180 => x"d8",
          5181 => x"c2",
          5182 => x"fe",
          5183 => x"72",
          5184 => x"81",
          5185 => x"71",
          5186 => x"38",
          5187 => x"f5",
          5188 => x"c2",
          5189 => x"f7",
          5190 => x"51",
          5191 => x"3f",
          5192 => x"70",
          5193 => x"52",
          5194 => x"95",
          5195 => x"fe",
          5196 => x"81",
          5197 => x"fe",
          5198 => x"80",
          5199 => x"fa",
          5200 => x"2a",
          5201 => x"51",
          5202 => x"2e",
          5203 => x"51",
          5204 => x"3f",
          5205 => x"51",
          5206 => x"3f",
          5207 => x"f4",
          5208 => x"86",
          5209 => x"06",
          5210 => x"80",
          5211 => x"81",
          5212 => x"c6",
          5213 => x"a4",
          5214 => x"be",
          5215 => x"fe",
          5216 => x"72",
          5217 => x"81",
          5218 => x"71",
          5219 => x"38",
          5220 => x"f4",
          5221 => x"c3",
          5222 => x"f6",
          5223 => x"51",
          5224 => x"3f",
          5225 => x"70",
          5226 => x"52",
          5227 => x"95",
          5228 => x"fe",
          5229 => x"81",
          5230 => x"fe",
          5231 => x"80",
          5232 => x"f6",
          5233 => x"a6",
          5234 => x"0d",
          5235 => x"0d",
          5236 => x"70",
          5237 => x"73",
          5238 => x"f0",
          5239 => x"73",
          5240 => x"15",
          5241 => x"e4",
          5242 => x"54",
          5243 => x"70",
          5244 => x"57",
          5245 => x"a0",
          5246 => x"81",
          5247 => x"2e",
          5248 => x"e5",
          5249 => x"ff",
          5250 => x"a0",
          5251 => x"06",
          5252 => x"74",
          5253 => x"56",
          5254 => x"75",
          5255 => x"c8",
          5256 => x"08",
          5257 => x"52",
          5258 => x"fd",
          5259 => x"a4",
          5260 => x"84",
          5261 => x"72",
          5262 => x"a3",
          5263 => x"70",
          5264 => x"57",
          5265 => x"27",
          5266 => x"53",
          5267 => x"a4",
          5268 => x"0d",
          5269 => x"0d",
          5270 => x"81",
          5271 => x"5e",
          5272 => x"7b",
          5273 => x"c8",
          5274 => x"a4",
          5275 => x"06",
          5276 => x"2e",
          5277 => x"a2",
          5278 => x"8c",
          5279 => x"70",
          5280 => x"84",
          5281 => x"53",
          5282 => x"cc",
          5283 => x"b9",
          5284 => x"cb",
          5285 => x"2e",
          5286 => x"c4",
          5287 => x"e8",
          5288 => x"5e",
          5289 => x"c8",
          5290 => x"a9",
          5291 => x"70",
          5292 => x"f8",
          5293 => x"79",
          5294 => x"dc",
          5295 => x"52",
          5296 => x"84",
          5297 => x"3d",
          5298 => x"51",
          5299 => x"81",
          5300 => x"90",
          5301 => x"2c",
          5302 => x"80",
          5303 => x"9b",
          5304 => x"c3",
          5305 => x"38",
          5306 => x"83",
          5307 => x"ab",
          5308 => x"78",
          5309 => x"af",
          5310 => x"24",
          5311 => x"80",
          5312 => x"38",
          5313 => x"78",
          5314 => x"82",
          5315 => x"2e",
          5316 => x"8c",
          5317 => x"80",
          5318 => x"8a",
          5319 => x"c0",
          5320 => x"78",
          5321 => x"a9",
          5322 => x"2e",
          5323 => x"8c",
          5324 => x"80",
          5325 => x"eb",
          5326 => x"c2",
          5327 => x"38",
          5328 => x"78",
          5329 => x"8b",
          5330 => x"80",
          5331 => x"38",
          5332 => x"2e",
          5333 => x"78",
          5334 => x"8b",
          5335 => x"d0",
          5336 => x"38",
          5337 => x"78",
          5338 => x"8a",
          5339 => x"80",
          5340 => x"f2",
          5341 => x"39",
          5342 => x"2e",
          5343 => x"78",
          5344 => x"92",
          5345 => x"f9",
          5346 => x"38",
          5347 => x"2e",
          5348 => x"8b",
          5349 => x"81",
          5350 => x"eb",
          5351 => x"87",
          5352 => x"38",
          5353 => x"b7",
          5354 => x"11",
          5355 => x"05",
          5356 => x"fa",
          5357 => x"a4",
          5358 => x"81",
          5359 => x"8c",
          5360 => x"3d",
          5361 => x"53",
          5362 => x"51",
          5363 => x"3f",
          5364 => x"08",
          5365 => x"38",
          5366 => x"83",
          5367 => x"02",
          5368 => x"33",
          5369 => x"cf",
          5370 => x"ff",
          5371 => x"81",
          5372 => x"81",
          5373 => x"78",
          5374 => x"c4",
          5375 => x"fb",
          5376 => x"5d",
          5377 => x"81",
          5378 => x"89",
          5379 => x"3d",
          5380 => x"53",
          5381 => x"51",
          5382 => x"3f",
          5383 => x"08",
          5384 => x"81",
          5385 => x"80",
          5386 => x"cf",
          5387 => x"ff",
          5388 => x"81",
          5389 => x"52",
          5390 => x"51",
          5391 => x"b7",
          5392 => x"11",
          5393 => x"05",
          5394 => x"e2",
          5395 => x"a4",
          5396 => x"87",
          5397 => x"26",
          5398 => x"b7",
          5399 => x"11",
          5400 => x"05",
          5401 => x"c6",
          5402 => x"a4",
          5403 => x"81",
          5404 => x"43",
          5405 => x"c5",
          5406 => x"51",
          5407 => x"3f",
          5408 => x"05",
          5409 => x"52",
          5410 => x"29",
          5411 => x"05",
          5412 => x"e0",
          5413 => x"a4",
          5414 => x"38",
          5415 => x"51",
          5416 => x"3f",
          5417 => x"fd",
          5418 => x"fe",
          5419 => x"fe",
          5420 => x"81",
          5421 => x"b8",
          5422 => x"05",
          5423 => x"eb",
          5424 => x"53",
          5425 => x"08",
          5426 => x"f5",
          5427 => x"d5",
          5428 => x"fe",
          5429 => x"fe",
          5430 => x"81",
          5431 => x"b8",
          5432 => x"05",
          5433 => x"ea",
          5434 => x"cb",
          5435 => x"3d",
          5436 => x"52",
          5437 => x"d5",
          5438 => x"a4",
          5439 => x"fe",
          5440 => x"59",
          5441 => x"3f",
          5442 => x"58",
          5443 => x"57",
          5444 => x"55",
          5445 => x"08",
          5446 => x"54",
          5447 => x"52",
          5448 => x"f0",
          5449 => x"a4",
          5450 => x"fa",
          5451 => x"cb",
          5452 => x"f0",
          5453 => x"ed",
          5454 => x"fe",
          5455 => x"fe",
          5456 => x"ff",
          5457 => x"81",
          5458 => x"80",
          5459 => x"38",
          5460 => x"f0",
          5461 => x"f8",
          5462 => x"80",
          5463 => x"cb",
          5464 => x"2e",
          5465 => x"b7",
          5466 => x"11",
          5467 => x"05",
          5468 => x"ba",
          5469 => x"a4",
          5470 => x"81",
          5471 => x"42",
          5472 => x"51",
          5473 => x"3f",
          5474 => x"5a",
          5475 => x"8f",
          5476 => x"78",
          5477 => x"05",
          5478 => x"7a",
          5479 => x"81",
          5480 => x"86",
          5481 => x"3d",
          5482 => x"53",
          5483 => x"51",
          5484 => x"3f",
          5485 => x"08",
          5486 => x"81",
          5487 => x"59",
          5488 => x"88",
          5489 => x"90",
          5490 => x"39",
          5491 => x"33",
          5492 => x"2e",
          5493 => x"c8",
          5494 => x"a2",
          5495 => x"bf",
          5496 => x"8b",
          5497 => x"c0",
          5498 => x"80",
          5499 => x"81",
          5500 => x"44",
          5501 => x"c8",
          5502 => x"80",
          5503 => x"3d",
          5504 => x"53",
          5505 => x"51",
          5506 => x"3f",
          5507 => x"08",
          5508 => x"81",
          5509 => x"59",
          5510 => x"88",
          5511 => x"94",
          5512 => x"39",
          5513 => x"33",
          5514 => x"2e",
          5515 => x"c8",
          5516 => x"a1",
          5517 => x"bf",
          5518 => x"8b",
          5519 => x"c0",
          5520 => x"80",
          5521 => x"81",
          5522 => x"43",
          5523 => x"c8",
          5524 => x"05",
          5525 => x"fe",
          5526 => x"fe",
          5527 => x"fe",
          5528 => x"81",
          5529 => x"80",
          5530 => x"80",
          5531 => x"79",
          5532 => x"38",
          5533 => x"90",
          5534 => x"78",
          5535 => x"38",
          5536 => x"83",
          5537 => x"81",
          5538 => x"fe",
          5539 => x"a0",
          5540 => x"61",
          5541 => x"63",
          5542 => x"3f",
          5543 => x"51",
          5544 => x"b7",
          5545 => x"11",
          5546 => x"05",
          5547 => x"fe",
          5548 => x"a4",
          5549 => x"f7",
          5550 => x"3d",
          5551 => x"53",
          5552 => x"51",
          5553 => x"3f",
          5554 => x"08",
          5555 => x"38",
          5556 => x"80",
          5557 => x"79",
          5558 => x"05",
          5559 => x"fe",
          5560 => x"fe",
          5561 => x"fe",
          5562 => x"81",
          5563 => x"e0",
          5564 => x"39",
          5565 => x"54",
          5566 => x"b8",
          5567 => x"b9",
          5568 => x"52",
          5569 => x"fc",
          5570 => x"45",
          5571 => x"78",
          5572 => x"91",
          5573 => x"27",
          5574 => x"3d",
          5575 => x"53",
          5576 => x"51",
          5577 => x"3f",
          5578 => x"08",
          5579 => x"38",
          5580 => x"80",
          5581 => x"79",
          5582 => x"05",
          5583 => x"39",
          5584 => x"51",
          5585 => x"3f",
          5586 => x"b7",
          5587 => x"11",
          5588 => x"05",
          5589 => x"c8",
          5590 => x"a4",
          5591 => x"f6",
          5592 => x"3d",
          5593 => x"53",
          5594 => x"51",
          5595 => x"3f",
          5596 => x"08",
          5597 => x"38",
          5598 => x"be",
          5599 => x"70",
          5600 => x"23",
          5601 => x"3d",
          5602 => x"53",
          5603 => x"51",
          5604 => x"3f",
          5605 => x"08",
          5606 => x"89",
          5607 => x"22",
          5608 => x"c5",
          5609 => x"fa",
          5610 => x"f8",
          5611 => x"fe",
          5612 => x"79",
          5613 => x"59",
          5614 => x"f5",
          5615 => x"9f",
          5616 => x"60",
          5617 => x"d5",
          5618 => x"fe",
          5619 => x"fe",
          5620 => x"fe",
          5621 => x"81",
          5622 => x"80",
          5623 => x"60",
          5624 => x"05",
          5625 => x"82",
          5626 => x"78",
          5627 => x"39",
          5628 => x"51",
          5629 => x"3f",
          5630 => x"b7",
          5631 => x"11",
          5632 => x"05",
          5633 => x"98",
          5634 => x"a4",
          5635 => x"f5",
          5636 => x"3d",
          5637 => x"53",
          5638 => x"51",
          5639 => x"3f",
          5640 => x"08",
          5641 => x"38",
          5642 => x"0c",
          5643 => x"05",
          5644 => x"fe",
          5645 => x"fe",
          5646 => x"fe",
          5647 => x"81",
          5648 => x"e4",
          5649 => x"39",
          5650 => x"54",
          5651 => x"d8",
          5652 => x"e5",
          5653 => x"52",
          5654 => x"f9",
          5655 => x"45",
          5656 => x"78",
          5657 => x"bd",
          5658 => x"27",
          5659 => x"3d",
          5660 => x"53",
          5661 => x"51",
          5662 => x"3f",
          5663 => x"08",
          5664 => x"38",
          5665 => x"52",
          5666 => x"51",
          5667 => x"3f",
          5668 => x"0c",
          5669 => x"05",
          5670 => x"39",
          5671 => x"51",
          5672 => x"3f",
          5673 => x"81",
          5674 => x"fe",
          5675 => x"82",
          5676 => x"95",
          5677 => x"39",
          5678 => x"51",
          5679 => x"3f",
          5680 => x"f0",
          5681 => x"dd",
          5682 => x"81",
          5683 => x"94",
          5684 => x"80",
          5685 => x"c0",
          5686 => x"81",
          5687 => x"fe",
          5688 => x"f3",
          5689 => x"c6",
          5690 => x"f1",
          5691 => x"80",
          5692 => x"c0",
          5693 => x"8c",
          5694 => x"87",
          5695 => x"0c",
          5696 => x"b7",
          5697 => x"11",
          5698 => x"05",
          5699 => x"9e",
          5700 => x"a4",
          5701 => x"f3",
          5702 => x"52",
          5703 => x"51",
          5704 => x"3f",
          5705 => x"04",
          5706 => x"f4",
          5707 => x"f8",
          5708 => x"f8",
          5709 => x"cb",
          5710 => x"2e",
          5711 => x"63",
          5712 => x"d8",
          5713 => x"f1",
          5714 => x"78",
          5715 => x"a4",
          5716 => x"cb",
          5717 => x"2e",
          5718 => x"81",
          5719 => x"52",
          5720 => x"51",
          5721 => x"3f",
          5722 => x"81",
          5723 => x"fe",
          5724 => x"fe",
          5725 => x"f2",
          5726 => x"c7",
          5727 => x"f0",
          5728 => x"59",
          5729 => x"fe",
          5730 => x"f2",
          5731 => x"70",
          5732 => x"78",
          5733 => x"8d",
          5734 => x"2e",
          5735 => x"7c",
          5736 => x"cc",
          5737 => x"fe",
          5738 => x"fe",
          5739 => x"81",
          5740 => x"81",
          5741 => x"55",
          5742 => x"54",
          5743 => x"c7",
          5744 => x"3d",
          5745 => x"fe",
          5746 => x"81",
          5747 => x"81",
          5748 => x"80",
          5749 => x"11",
          5750 => x"55",
          5751 => x"e4",
          5752 => x"e4",
          5753 => x"51",
          5754 => x"81",
          5755 => x"5e",
          5756 => x"7c",
          5757 => x"59",
          5758 => x"7d",
          5759 => x"81",
          5760 => x"38",
          5761 => x"51",
          5762 => x"3f",
          5763 => x"80",
          5764 => x"0b",
          5765 => x"34",
          5766 => x"c8",
          5767 => x"94",
          5768 => x"a0",
          5769 => x"87",
          5770 => x"0c",
          5771 => x"0b",
          5772 => x"84",
          5773 => x"83",
          5774 => x"94",
          5775 => x"d1",
          5776 => x"b4",
          5777 => x"0b",
          5778 => x"0c",
          5779 => x"3f",
          5780 => x"3f",
          5781 => x"51",
          5782 => x"3f",
          5783 => x"51",
          5784 => x"3f",
          5785 => x"51",
          5786 => x"3f",
          5787 => x"ed",
          5788 => x"3f",
          5789 => x"00",
          5790 => x"00",
          5791 => x"00",
          5792 => x"00",
          5793 => x"00",
          5794 => x"00",
          5795 => x"00",
          5796 => x"00",
          5797 => x"00",
          5798 => x"00",
          5799 => x"00",
          5800 => x"00",
          5801 => x"00",
          5802 => x"00",
          5803 => x"00",
          5804 => x"00",
          5805 => x"00",
          5806 => x"00",
          5807 => x"00",
          5808 => x"00",
          5809 => x"00",
          5810 => x"00",
          5811 => x"00",
          5812 => x"00",
          5813 => x"00",
          5814 => x"25",
          5815 => x"64",
          5816 => x"20",
          5817 => x"25",
          5818 => x"64",
          5819 => x"25",
          5820 => x"53",
          5821 => x"43",
          5822 => x"69",
          5823 => x"61",
          5824 => x"6e",
          5825 => x"20",
          5826 => x"6f",
          5827 => x"6f",
          5828 => x"6f",
          5829 => x"67",
          5830 => x"3a",
          5831 => x"76",
          5832 => x"73",
          5833 => x"70",
          5834 => x"65",
          5835 => x"64",
          5836 => x"20",
          5837 => x"49",
          5838 => x"20",
          5839 => x"4d",
          5840 => x"74",
          5841 => x"3d",
          5842 => x"58",
          5843 => x"69",
          5844 => x"25",
          5845 => x"29",
          5846 => x"20",
          5847 => x"42",
          5848 => x"20",
          5849 => x"61",
          5850 => x"25",
          5851 => x"2c",
          5852 => x"7a",
          5853 => x"30",
          5854 => x"2e",
          5855 => x"20",
          5856 => x"52",
          5857 => x"28",
          5858 => x"72",
          5859 => x"30",
          5860 => x"20",
          5861 => x"65",
          5862 => x"38",
          5863 => x"0a",
          5864 => x"20",
          5865 => x"49",
          5866 => x"4c",
          5867 => x"20",
          5868 => x"50",
          5869 => x"00",
          5870 => x"20",
          5871 => x"53",
          5872 => x"00",
          5873 => x"20",
          5874 => x"53",
          5875 => x"61",
          5876 => x"28",
          5877 => x"69",
          5878 => x"3d",
          5879 => x"58",
          5880 => x"00",
          5881 => x"20",
          5882 => x"49",
          5883 => x"52",
          5884 => x"54",
          5885 => x"4e",
          5886 => x"4c",
          5887 => x"0a",
          5888 => x"20",
          5889 => x"54",
          5890 => x"52",
          5891 => x"54",
          5892 => x"72",
          5893 => x"30",
          5894 => x"2e",
          5895 => x"41",
          5896 => x"65",
          5897 => x"73",
          5898 => x"20",
          5899 => x"43",
          5900 => x"52",
          5901 => x"74",
          5902 => x"63",
          5903 => x"20",
          5904 => x"72",
          5905 => x"20",
          5906 => x"30",
          5907 => x"00",
          5908 => x"20",
          5909 => x"43",
          5910 => x"4d",
          5911 => x"72",
          5912 => x"74",
          5913 => x"20",
          5914 => x"72",
          5915 => x"20",
          5916 => x"30",
          5917 => x"00",
          5918 => x"20",
          5919 => x"53",
          5920 => x"6b",
          5921 => x"61",
          5922 => x"41",
          5923 => x"65",
          5924 => x"20",
          5925 => x"20",
          5926 => x"30",
          5927 => x"00",
          5928 => x"20",
          5929 => x"5a",
          5930 => x"49",
          5931 => x"20",
          5932 => x"20",
          5933 => x"20",
          5934 => x"20",
          5935 => x"20",
          5936 => x"30",
          5937 => x"00",
          5938 => x"20",
          5939 => x"53",
          5940 => x"65",
          5941 => x"6c",
          5942 => x"20",
          5943 => x"71",
          5944 => x"20",
          5945 => x"20",
          5946 => x"30",
          5947 => x"00",
          5948 => x"53",
          5949 => x"6c",
          5950 => x"4d",
          5951 => x"75",
          5952 => x"46",
          5953 => x"00",
          5954 => x"45",
          5955 => x"45",
          5956 => x"69",
          5957 => x"55",
          5958 => x"6f",
          5959 => x"53",
          5960 => x"22",
          5961 => x"3a",
          5962 => x"3e",
          5963 => x"7c",
          5964 => x"46",
          5965 => x"46",
          5966 => x"32",
          5967 => x"eb",
          5968 => x"53",
          5969 => x"35",
          5970 => x"4e",
          5971 => x"41",
          5972 => x"20",
          5973 => x"41",
          5974 => x"20",
          5975 => x"4e",
          5976 => x"41",
          5977 => x"20",
          5978 => x"41",
          5979 => x"20",
          5980 => x"00",
          5981 => x"00",
          5982 => x"00",
          5983 => x"00",
          5984 => x"80",
          5985 => x"8e",
          5986 => x"45",
          5987 => x"49",
          5988 => x"90",
          5989 => x"99",
          5990 => x"59",
          5991 => x"9c",
          5992 => x"41",
          5993 => x"a5",
          5994 => x"a8",
          5995 => x"ac",
          5996 => x"b0",
          5997 => x"b4",
          5998 => x"b8",
          5999 => x"bc",
          6000 => x"c0",
          6001 => x"c4",
          6002 => x"c8",
          6003 => x"cc",
          6004 => x"d0",
          6005 => x"d4",
          6006 => x"d8",
          6007 => x"dc",
          6008 => x"e0",
          6009 => x"e4",
          6010 => x"e8",
          6011 => x"ec",
          6012 => x"f0",
          6013 => x"f4",
          6014 => x"f8",
          6015 => x"fc",
          6016 => x"2b",
          6017 => x"3d",
          6018 => x"5c",
          6019 => x"3c",
          6020 => x"7f",
          6021 => x"00",
          6022 => x"00",
          6023 => x"01",
          6024 => x"00",
          6025 => x"00",
          6026 => x"00",
          6027 => x"00",
          6028 => x"00",
          6029 => x"64",
          6030 => x"74",
          6031 => x"64",
          6032 => x"74",
          6033 => x"66",
          6034 => x"74",
          6035 => x"66",
          6036 => x"64",
          6037 => x"66",
          6038 => x"63",
          6039 => x"6d",
          6040 => x"61",
          6041 => x"6d",
          6042 => x"70",
          6043 => x"6d",
          6044 => x"74",
          6045 => x"6d",
          6046 => x"6d",
          6047 => x"6d",
          6048 => x"68",
          6049 => x"68",
          6050 => x"68",
          6051 => x"68",
          6052 => x"63",
          6053 => x"00",
          6054 => x"6a",
          6055 => x"72",
          6056 => x"61",
          6057 => x"72",
          6058 => x"74",
          6059 => x"69",
          6060 => x"00",
          6061 => x"74",
          6062 => x"00",
          6063 => x"44",
          6064 => x"20",
          6065 => x"6f",
          6066 => x"49",
          6067 => x"72",
          6068 => x"20",
          6069 => x"6f",
          6070 => x"00",
          6071 => x"44",
          6072 => x"20",
          6073 => x"20",
          6074 => x"64",
          6075 => x"00",
          6076 => x"4e",
          6077 => x"69",
          6078 => x"66",
          6079 => x"64",
          6080 => x"4e",
          6081 => x"61",
          6082 => x"66",
          6083 => x"64",
          6084 => x"49",
          6085 => x"6c",
          6086 => x"66",
          6087 => x"6e",
          6088 => x"2e",
          6089 => x"41",
          6090 => x"73",
          6091 => x"65",
          6092 => x"64",
          6093 => x"46",
          6094 => x"20",
          6095 => x"65",
          6096 => x"20",
          6097 => x"73",
          6098 => x"0a",
          6099 => x"46",
          6100 => x"20",
          6101 => x"64",
          6102 => x"69",
          6103 => x"6c",
          6104 => x"0a",
          6105 => x"53",
          6106 => x"73",
          6107 => x"69",
          6108 => x"70",
          6109 => x"65",
          6110 => x"64",
          6111 => x"44",
          6112 => x"65",
          6113 => x"6d",
          6114 => x"20",
          6115 => x"69",
          6116 => x"6c",
          6117 => x"0a",
          6118 => x"44",
          6119 => x"20",
          6120 => x"20",
          6121 => x"62",
          6122 => x"2e",
          6123 => x"4e",
          6124 => x"6f",
          6125 => x"74",
          6126 => x"65",
          6127 => x"6c",
          6128 => x"73",
          6129 => x"20",
          6130 => x"6e",
          6131 => x"6e",
          6132 => x"73",
          6133 => x"00",
          6134 => x"46",
          6135 => x"61",
          6136 => x"62",
          6137 => x"65",
          6138 => x"00",
          6139 => x"54",
          6140 => x"6f",
          6141 => x"20",
          6142 => x"72",
          6143 => x"6f",
          6144 => x"61",
          6145 => x"6c",
          6146 => x"2e",
          6147 => x"46",
          6148 => x"20",
          6149 => x"6c",
          6150 => x"65",
          6151 => x"00",
          6152 => x"49",
          6153 => x"66",
          6154 => x"69",
          6155 => x"20",
          6156 => x"6f",
          6157 => x"0a",
          6158 => x"54",
          6159 => x"6d",
          6160 => x"20",
          6161 => x"6e",
          6162 => x"6c",
          6163 => x"0a",
          6164 => x"50",
          6165 => x"6d",
          6166 => x"72",
          6167 => x"6e",
          6168 => x"72",
          6169 => x"2e",
          6170 => x"53",
          6171 => x"65",
          6172 => x"0a",
          6173 => x"55",
          6174 => x"6f",
          6175 => x"65",
          6176 => x"72",
          6177 => x"0a",
          6178 => x"20",
          6179 => x"65",
          6180 => x"73",
          6181 => x"20",
          6182 => x"20",
          6183 => x"65",
          6184 => x"65",
          6185 => x"00",
          6186 => x"25",
          6187 => x"00",
          6188 => x"3a",
          6189 => x"25",
          6190 => x"00",
          6191 => x"20",
          6192 => x"20",
          6193 => x"00",
          6194 => x"25",
          6195 => x"00",
          6196 => x"20",
          6197 => x"20",
          6198 => x"7c",
          6199 => x"72",
          6200 => x"00",
          6201 => x"5a",
          6202 => x"41",
          6203 => x"0a",
          6204 => x"25",
          6205 => x"00",
          6206 => x"31",
          6207 => x"37",
          6208 => x"31",
          6209 => x"76",
          6210 => x"00",
          6211 => x"20",
          6212 => x"2c",
          6213 => x"76",
          6214 => x"32",
          6215 => x"25",
          6216 => x"73",
          6217 => x"0a",
          6218 => x"5a",
          6219 => x"41",
          6220 => x"74",
          6221 => x"75",
          6222 => x"48",
          6223 => x"6c",
          6224 => x"00",
          6225 => x"54",
          6226 => x"72",
          6227 => x"74",
          6228 => x"75",
          6229 => x"00",
          6230 => x"50",
          6231 => x"69",
          6232 => x"72",
          6233 => x"74",
          6234 => x"49",
          6235 => x"4c",
          6236 => x"20",
          6237 => x"65",
          6238 => x"70",
          6239 => x"49",
          6240 => x"4c",
          6241 => x"20",
          6242 => x"65",
          6243 => x"70",
          6244 => x"55",
          6245 => x"30",
          6246 => x"20",
          6247 => x"65",
          6248 => x"70",
          6249 => x"55",
          6250 => x"30",
          6251 => x"20",
          6252 => x"65",
          6253 => x"70",
          6254 => x"55",
          6255 => x"31",
          6256 => x"20",
          6257 => x"65",
          6258 => x"70",
          6259 => x"55",
          6260 => x"31",
          6261 => x"20",
          6262 => x"65",
          6263 => x"70",
          6264 => x"53",
          6265 => x"69",
          6266 => x"75",
          6267 => x"69",
          6268 => x"2e",
          6269 => x"00",
          6270 => x"45",
          6271 => x"6c",
          6272 => x"20",
          6273 => x"65",
          6274 => x"2e",
          6275 => x"30",
          6276 => x"46",
          6277 => x"65",
          6278 => x"6f",
          6279 => x"69",
          6280 => x"6c",
          6281 => x"20",
          6282 => x"63",
          6283 => x"20",
          6284 => x"70",
          6285 => x"73",
          6286 => x"6e",
          6287 => x"6d",
          6288 => x"61",
          6289 => x"2e",
          6290 => x"2a",
          6291 => x"42",
          6292 => x"64",
          6293 => x"20",
          6294 => x"0a",
          6295 => x"49",
          6296 => x"69",
          6297 => x"73",
          6298 => x"0a",
          6299 => x"46",
          6300 => x"65",
          6301 => x"6f",
          6302 => x"69",
          6303 => x"6c",
          6304 => x"2e",
          6305 => x"72",
          6306 => x"64",
          6307 => x"25",
          6308 => x"43",
          6309 => x"72",
          6310 => x"2e",
          6311 => x"44",
          6312 => x"20",
          6313 => x"6f",
          6314 => x"00",
          6315 => x"0a",
          6316 => x"70",
          6317 => x"65",
          6318 => x"25",
          6319 => x"20",
          6320 => x"58",
          6321 => x"3f",
          6322 => x"00",
          6323 => x"25",
          6324 => x"20",
          6325 => x"58",
          6326 => x"25",
          6327 => x"20",
          6328 => x"58",
          6329 => x"44",
          6330 => x"62",
          6331 => x"67",
          6332 => x"74",
          6333 => x"75",
          6334 => x"0a",
          6335 => x"45",
          6336 => x"6c",
          6337 => x"20",
          6338 => x"65",
          6339 => x"70",
          6340 => x"00",
          6341 => x"44",
          6342 => x"62",
          6343 => x"20",
          6344 => x"74",
          6345 => x"66",
          6346 => x"45",
          6347 => x"6c",
          6348 => x"20",
          6349 => x"74",
          6350 => x"66",
          6351 => x"45",
          6352 => x"75",
          6353 => x"67",
          6354 => x"64",
          6355 => x"20",
          6356 => x"78",
          6357 => x"2e",
          6358 => x"43",
          6359 => x"69",
          6360 => x"63",
          6361 => x"20",
          6362 => x"30",
          6363 => x"2e",
          6364 => x"00",
          6365 => x"43",
          6366 => x"20",
          6367 => x"75",
          6368 => x"64",
          6369 => x"64",
          6370 => x"25",
          6371 => x"0a",
          6372 => x"52",
          6373 => x"61",
          6374 => x"6e",
          6375 => x"70",
          6376 => x"63",
          6377 => x"6f",
          6378 => x"2e",
          6379 => x"43",
          6380 => x"20",
          6381 => x"6f",
          6382 => x"6e",
          6383 => x"2e",
          6384 => x"5a",
          6385 => x"62",
          6386 => x"25",
          6387 => x"25",
          6388 => x"73",
          6389 => x"00",
          6390 => x"42",
          6391 => x"63",
          6392 => x"61",
          6393 => x"0a",
          6394 => x"52",
          6395 => x"69",
          6396 => x"2e",
          6397 => x"45",
          6398 => x"6c",
          6399 => x"20",
          6400 => x"65",
          6401 => x"70",
          6402 => x"2e",
          6403 => x"00",
          6404 => x"00",
          6405 => x"00",
          6406 => x"00",
          6407 => x"00",
          6408 => x"00",
          6409 => x"00",
          6410 => x"00",
          6411 => x"00",
          6412 => x"00",
          6413 => x"00",
          6414 => x"05",
          6415 => x"00",
          6416 => x"01",
          6417 => x"80",
          6418 => x"01",
          6419 => x"00",
          6420 => x"01",
          6421 => x"00",
          6422 => x"01",
          6423 => x"00",
          6424 => x"00",
          6425 => x"00",
          6426 => x"01",
          6427 => x"00",
          6428 => x"00",
          6429 => x"00",
          6430 => x"01",
          6431 => x"00",
          6432 => x"00",
          6433 => x"00",
          6434 => x"01",
          6435 => x"00",
          6436 => x"00",
          6437 => x"00",
          6438 => x"01",
          6439 => x"00",
          6440 => x"00",
          6441 => x"00",
          6442 => x"01",
          6443 => x"00",
          6444 => x"00",
          6445 => x"00",
          6446 => x"01",
          6447 => x"00",
          6448 => x"00",
          6449 => x"00",
          6450 => x"01",
          6451 => x"00",
          6452 => x"00",
          6453 => x"00",
          6454 => x"01",
          6455 => x"00",
          6456 => x"00",
          6457 => x"00",
          6458 => x"01",
          6459 => x"00",
          6460 => x"00",
          6461 => x"00",
          6462 => x"01",
          6463 => x"00",
          6464 => x"00",
          6465 => x"00",
          6466 => x"01",
          6467 => x"00",
          6468 => x"00",
          6469 => x"00",
          6470 => x"01",
          6471 => x"00",
          6472 => x"00",
          6473 => x"00",
          6474 => x"01",
          6475 => x"00",
          6476 => x"00",
          6477 => x"00",
          6478 => x"01",
          6479 => x"00",
          6480 => x"00",
          6481 => x"00",
          6482 => x"01",
          6483 => x"00",
          6484 => x"00",
          6485 => x"00",
          6486 => x"01",
          6487 => x"00",
          6488 => x"00",
          6489 => x"00",
          6490 => x"01",
          6491 => x"00",
          6492 => x"00",
          6493 => x"00",
          6494 => x"01",
          6495 => x"00",
          6496 => x"00",
          6497 => x"00",
          6498 => x"01",
          6499 => x"00",
          6500 => x"00",
          6501 => x"00",
          6502 => x"01",
          6503 => x"00",
          6504 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
