-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.softZPU_pkg.all;

entity DualPortBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBRAM;

architecture arch of DualPortBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"ff",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"80",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"ac",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"c5",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"c7",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"84",
           386 => x"97",
           387 => x"84",
           388 => x"90",
           389 => x"84",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"82",
           395 => x"84",
           396 => x"82",
           397 => x"af",
           398 => x"d5",
           399 => x"80",
           400 => x"d5",
           401 => x"ad",
           402 => x"84",
           403 => x"90",
           404 => x"84",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"82",
           418 => x"84",
           419 => x"82",
           420 => x"96",
           421 => x"d5",
           422 => x"80",
           423 => x"d5",
           424 => x"cd",
           425 => x"84",
           426 => x"90",
           427 => x"84",
           428 => x"c1",
           429 => x"84",
           430 => x"90",
           431 => x"84",
           432 => x"9f",
           433 => x"84",
           434 => x"90",
           435 => x"84",
           436 => x"dc",
           437 => x"84",
           438 => x"90",
           439 => x"84",
           440 => x"d3",
           441 => x"84",
           442 => x"90",
           443 => x"84",
           444 => x"86",
           445 => x"84",
           446 => x"90",
           447 => x"84",
           448 => x"eb",
           449 => x"84",
           450 => x"90",
           451 => x"84",
           452 => x"ea",
           453 => x"84",
           454 => x"90",
           455 => x"84",
           456 => x"d0",
           457 => x"84",
           458 => x"90",
           459 => x"84",
           460 => x"d0",
           461 => x"84",
           462 => x"90",
           463 => x"84",
           464 => x"a8",
           465 => x"84",
           466 => x"90",
           467 => x"84",
           468 => x"91",
           469 => x"84",
           470 => x"90",
           471 => x"84",
           472 => x"c7",
           473 => x"84",
           474 => x"90",
           475 => x"84",
           476 => x"cb",
           477 => x"84",
           478 => x"90",
           479 => x"84",
           480 => x"eb",
           481 => x"84",
           482 => x"90",
           483 => x"84",
           484 => x"8a",
           485 => x"84",
           486 => x"90",
           487 => x"84",
           488 => x"fe",
           489 => x"84",
           490 => x"90",
           491 => x"84",
           492 => x"e0",
           493 => x"84",
           494 => x"90",
           495 => x"84",
           496 => x"da",
           497 => x"84",
           498 => x"90",
           499 => x"84",
           500 => x"90",
           501 => x"84",
           502 => x"90",
           503 => x"84",
           504 => x"df",
           505 => x"84",
           506 => x"90",
           507 => x"84",
           508 => x"e0",
           509 => x"84",
           510 => x"90",
           511 => x"84",
           512 => x"ca",
           513 => x"84",
           514 => x"90",
           515 => x"84",
           516 => x"a3",
           517 => x"84",
           518 => x"90",
           519 => x"84",
           520 => x"ce",
           521 => x"84",
           522 => x"90",
           523 => x"84",
           524 => x"e7",
           525 => x"84",
           526 => x"90",
           527 => x"84",
           528 => x"d1",
           529 => x"84",
           530 => x"90",
           531 => x"84",
           532 => x"dc",
           533 => x"84",
           534 => x"90",
           535 => x"84",
           536 => x"e3",
           537 => x"84",
           538 => x"90",
           539 => x"84",
           540 => x"8a",
           541 => x"84",
           542 => x"90",
           543 => x"84",
           544 => x"cf",
           545 => x"84",
           546 => x"90",
           547 => x"84",
           548 => x"84",
           549 => x"84",
           550 => x"90",
           551 => x"84",
           552 => x"f0",
           553 => x"84",
           554 => x"90",
           555 => x"84",
           556 => x"92",
           557 => x"84",
           558 => x"90",
           559 => x"84",
           560 => x"fc",
           561 => x"84",
           562 => x"90",
           563 => x"84",
           564 => x"e0",
           565 => x"84",
           566 => x"90",
           567 => x"84",
           568 => x"85",
           569 => x"84",
           570 => x"90",
           571 => x"84",
           572 => x"a9",
           573 => x"84",
           574 => x"90",
           575 => x"84",
           576 => x"8c",
           577 => x"84",
           578 => x"90",
           579 => x"84",
           580 => x"bf",
           581 => x"84",
           582 => x"90",
           583 => x"84",
           584 => x"a6",
           585 => x"84",
           586 => x"90",
           587 => x"84",
           588 => x"ce",
           589 => x"84",
           590 => x"90",
           591 => x"84",
           592 => x"c6",
           593 => x"84",
           594 => x"90",
           595 => x"84",
           596 => x"90",
           597 => x"84",
           598 => x"90",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"00",
           609 => x"ff",
           610 => x"06",
           611 => x"83",
           612 => x"10",
           613 => x"fc",
           614 => x"51",
           615 => x"80",
           616 => x"ff",
           617 => x"06",
           618 => x"52",
           619 => x"0a",
           620 => x"38",
           621 => x"51",
           622 => x"f8",
           623 => x"e4",
           624 => x"80",
           625 => x"05",
           626 => x"0b",
           627 => x"04",
           628 => x"80",
           629 => x"00",
           630 => x"08",
           631 => x"84",
           632 => x"0d",
           633 => x"08",
           634 => x"82",
           635 => x"fc",
           636 => x"d5",
           637 => x"05",
           638 => x"d5",
           639 => x"05",
           640 => x"f0",
           641 => x"54",
           642 => x"82",
           643 => x"70",
           644 => x"08",
           645 => x"82",
           646 => x"f8",
           647 => x"82",
           648 => x"51",
           649 => x"0d",
           650 => x"0c",
           651 => x"84",
           652 => x"d5",
           653 => x"3d",
           654 => x"84",
           655 => x"08",
           656 => x"70",
           657 => x"81",
           658 => x"51",
           659 => x"38",
           660 => x"d5",
           661 => x"05",
           662 => x"38",
           663 => x"0b",
           664 => x"08",
           665 => x"81",
           666 => x"d5",
           667 => x"05",
           668 => x"82",
           669 => x"8c",
           670 => x"0b",
           671 => x"08",
           672 => x"82",
           673 => x"88",
           674 => x"d5",
           675 => x"05",
           676 => x"84",
           677 => x"08",
           678 => x"f6",
           679 => x"82",
           680 => x"8c",
           681 => x"80",
           682 => x"d5",
           683 => x"05",
           684 => x"90",
           685 => x"f8",
           686 => x"d5",
           687 => x"05",
           688 => x"d5",
           689 => x"05",
           690 => x"09",
           691 => x"38",
           692 => x"d5",
           693 => x"05",
           694 => x"39",
           695 => x"08",
           696 => x"82",
           697 => x"f8",
           698 => x"53",
           699 => x"82",
           700 => x"8c",
           701 => x"05",
           702 => x"08",
           703 => x"82",
           704 => x"fc",
           705 => x"05",
           706 => x"08",
           707 => x"ff",
           708 => x"d5",
           709 => x"05",
           710 => x"72",
           711 => x"84",
           712 => x"08",
           713 => x"84",
           714 => x"0c",
           715 => x"84",
           716 => x"08",
           717 => x"0c",
           718 => x"82",
           719 => x"04",
           720 => x"08",
           721 => x"84",
           722 => x"0d",
           723 => x"d5",
           724 => x"05",
           725 => x"84",
           726 => x"08",
           727 => x"08",
           728 => x"fe",
           729 => x"d5",
           730 => x"05",
           731 => x"84",
           732 => x"70",
           733 => x"08",
           734 => x"82",
           735 => x"fc",
           736 => x"82",
           737 => x"8c",
           738 => x"82",
           739 => x"e0",
           740 => x"51",
           741 => x"3f",
           742 => x"08",
           743 => x"84",
           744 => x"0c",
           745 => x"08",
           746 => x"82",
           747 => x"88",
           748 => x"51",
           749 => x"34",
           750 => x"08",
           751 => x"70",
           752 => x"0c",
           753 => x"0d",
           754 => x"0c",
           755 => x"84",
           756 => x"d5",
           757 => x"3d",
           758 => x"84",
           759 => x"70",
           760 => x"08",
           761 => x"82",
           762 => x"fc",
           763 => x"82",
           764 => x"8c",
           765 => x"82",
           766 => x"88",
           767 => x"54",
           768 => x"d4",
           769 => x"82",
           770 => x"f8",
           771 => x"d5",
           772 => x"05",
           773 => x"d4",
           774 => x"54",
           775 => x"82",
           776 => x"04",
           777 => x"08",
           778 => x"84",
           779 => x"0d",
           780 => x"d5",
           781 => x"05",
           782 => x"84",
           783 => x"08",
           784 => x"8c",
           785 => x"d5",
           786 => x"05",
           787 => x"33",
           788 => x"70",
           789 => x"81",
           790 => x"51",
           791 => x"80",
           792 => x"ff",
           793 => x"84",
           794 => x"0c",
           795 => x"82",
           796 => x"8c",
           797 => x"72",
           798 => x"82",
           799 => x"f8",
           800 => x"81",
           801 => x"72",
           802 => x"fa",
           803 => x"84",
           804 => x"08",
           805 => x"d5",
           806 => x"05",
           807 => x"84",
           808 => x"22",
           809 => x"51",
           810 => x"2e",
           811 => x"82",
           812 => x"f8",
           813 => x"af",
           814 => x"fc",
           815 => x"84",
           816 => x"33",
           817 => x"26",
           818 => x"82",
           819 => x"f8",
           820 => x"72",
           821 => x"81",
           822 => x"38",
           823 => x"08",
           824 => x"70",
           825 => x"98",
           826 => x"53",
           827 => x"82",
           828 => x"e4",
           829 => x"83",
           830 => x"32",
           831 => x"51",
           832 => x"72",
           833 => x"38",
           834 => x"08",
           835 => x"70",
           836 => x"51",
           837 => x"d5",
           838 => x"05",
           839 => x"39",
           840 => x"08",
           841 => x"70",
           842 => x"98",
           843 => x"83",
           844 => x"73",
           845 => x"51",
           846 => x"53",
           847 => x"84",
           848 => x"34",
           849 => x"08",
           850 => x"54",
           851 => x"08",
           852 => x"70",
           853 => x"51",
           854 => x"82",
           855 => x"e8",
           856 => x"d5",
           857 => x"05",
           858 => x"2b",
           859 => x"51",
           860 => x"80",
           861 => x"80",
           862 => x"d5",
           863 => x"05",
           864 => x"84",
           865 => x"22",
           866 => x"70",
           867 => x"51",
           868 => x"db",
           869 => x"84",
           870 => x"33",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"d5",
           876 => x"05",
           877 => x"39",
           878 => x"08",
           879 => x"70",
           880 => x"81",
           881 => x"53",
           882 => x"9d",
           883 => x"84",
           884 => x"33",
           885 => x"70",
           886 => x"51",
           887 => x"38",
           888 => x"d5",
           889 => x"05",
           890 => x"84",
           891 => x"33",
           892 => x"d5",
           893 => x"05",
           894 => x"d5",
           895 => x"05",
           896 => x"26",
           897 => x"82",
           898 => x"c4",
           899 => x"82",
           900 => x"f8",
           901 => x"51",
           902 => x"72",
           903 => x"84",
           904 => x"22",
           905 => x"51",
           906 => x"d5",
           907 => x"05",
           908 => x"84",
           909 => x"22",
           910 => x"51",
           911 => x"d5",
           912 => x"05",
           913 => x"39",
           914 => x"08",
           915 => x"70",
           916 => x"51",
           917 => x"d5",
           918 => x"05",
           919 => x"39",
           920 => x"08",
           921 => x"70",
           922 => x"51",
           923 => x"d5",
           924 => x"05",
           925 => x"39",
           926 => x"08",
           927 => x"70",
           928 => x"53",
           929 => x"84",
           930 => x"23",
           931 => x"d5",
           932 => x"05",
           933 => x"39",
           934 => x"08",
           935 => x"70",
           936 => x"53",
           937 => x"84",
           938 => x"23",
           939 => x"bf",
           940 => x"84",
           941 => x"34",
           942 => x"08",
           943 => x"ff",
           944 => x"72",
           945 => x"08",
           946 => x"80",
           947 => x"d5",
           948 => x"05",
           949 => x"39",
           950 => x"08",
           951 => x"82",
           952 => x"90",
           953 => x"05",
           954 => x"08",
           955 => x"70",
           956 => x"72",
           957 => x"08",
           958 => x"82",
           959 => x"ec",
           960 => x"11",
           961 => x"82",
           962 => x"ec",
           963 => x"ef",
           964 => x"84",
           965 => x"08",
           966 => x"08",
           967 => x"84",
           968 => x"84",
           969 => x"0c",
           970 => x"d5",
           971 => x"05",
           972 => x"84",
           973 => x"22",
           974 => x"70",
           975 => x"51",
           976 => x"80",
           977 => x"82",
           978 => x"e8",
           979 => x"98",
           980 => x"98",
           981 => x"d5",
           982 => x"05",
           983 => x"a4",
           984 => x"d4",
           985 => x"72",
           986 => x"08",
           987 => x"99",
           988 => x"84",
           989 => x"08",
           990 => x"3f",
           991 => x"08",
           992 => x"d5",
           993 => x"05",
           994 => x"84",
           995 => x"22",
           996 => x"84",
           997 => x"22",
           998 => x"54",
           999 => x"d5",
          1000 => x"05",
          1001 => x"39",
          1002 => x"08",
          1003 => x"82",
          1004 => x"90",
          1005 => x"05",
          1006 => x"08",
          1007 => x"70",
          1008 => x"84",
          1009 => x"0c",
          1010 => x"08",
          1011 => x"70",
          1012 => x"81",
          1013 => x"51",
          1014 => x"2e",
          1015 => x"d5",
          1016 => x"05",
          1017 => x"2b",
          1018 => x"2c",
          1019 => x"84",
          1020 => x"08",
          1021 => x"ec",
          1022 => x"f8",
          1023 => x"82",
          1024 => x"f4",
          1025 => x"39",
          1026 => x"08",
          1027 => x"51",
          1028 => x"82",
          1029 => x"53",
          1030 => x"84",
          1031 => x"23",
          1032 => x"08",
          1033 => x"53",
          1034 => x"08",
          1035 => x"73",
          1036 => x"54",
          1037 => x"84",
          1038 => x"23",
          1039 => x"82",
          1040 => x"e4",
          1041 => x"82",
          1042 => x"06",
          1043 => x"72",
          1044 => x"38",
          1045 => x"08",
          1046 => x"82",
          1047 => x"90",
          1048 => x"05",
          1049 => x"08",
          1050 => x"70",
          1051 => x"84",
          1052 => x"0c",
          1053 => x"82",
          1054 => x"90",
          1055 => x"d5",
          1056 => x"05",
          1057 => x"82",
          1058 => x"90",
          1059 => x"08",
          1060 => x"08",
          1061 => x"53",
          1062 => x"08",
          1063 => x"82",
          1064 => x"fc",
          1065 => x"d5",
          1066 => x"05",
          1067 => x"a4",
          1068 => x"84",
          1069 => x"22",
          1070 => x"51",
          1071 => x"d5",
          1072 => x"05",
          1073 => x"84",
          1074 => x"08",
          1075 => x"84",
          1076 => x"0c",
          1077 => x"08",
          1078 => x"70",
          1079 => x"51",
          1080 => x"d5",
          1081 => x"05",
          1082 => x"39",
          1083 => x"d5",
          1084 => x"05",
          1085 => x"82",
          1086 => x"e4",
          1087 => x"80",
          1088 => x"53",
          1089 => x"84",
          1090 => x"23",
          1091 => x"82",
          1092 => x"f8",
          1093 => x"0b",
          1094 => x"08",
          1095 => x"82",
          1096 => x"e4",
          1097 => x"82",
          1098 => x"06",
          1099 => x"72",
          1100 => x"38",
          1101 => x"08",
          1102 => x"82",
          1103 => x"90",
          1104 => x"05",
          1105 => x"08",
          1106 => x"70",
          1107 => x"84",
          1108 => x"0c",
          1109 => x"82",
          1110 => x"90",
          1111 => x"d5",
          1112 => x"05",
          1113 => x"82",
          1114 => x"90",
          1115 => x"08",
          1116 => x"08",
          1117 => x"53",
          1118 => x"08",
          1119 => x"82",
          1120 => x"fc",
          1121 => x"d5",
          1122 => x"05",
          1123 => x"06",
          1124 => x"82",
          1125 => x"e4",
          1126 => x"d5",
          1127 => x"d5",
          1128 => x"05",
          1129 => x"84",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"fc",
          1134 => x"55",
          1135 => x"54",
          1136 => x"3f",
          1137 => x"08",
          1138 => x"34",
          1139 => x"08",
          1140 => x"82",
          1141 => x"d4",
          1142 => x"d5",
          1143 => x"05",
          1144 => x"51",
          1145 => x"27",
          1146 => x"d5",
          1147 => x"05",
          1148 => x"33",
          1149 => x"84",
          1150 => x"33",
          1151 => x"11",
          1152 => x"72",
          1153 => x"08",
          1154 => x"97",
          1155 => x"84",
          1156 => x"08",
          1157 => x"b0",
          1158 => x"72",
          1159 => x"08",
          1160 => x"82",
          1161 => x"d4",
          1162 => x"82",
          1163 => x"d0",
          1164 => x"34",
          1165 => x"08",
          1166 => x"81",
          1167 => x"84",
          1168 => x"0c",
          1169 => x"08",
          1170 => x"70",
          1171 => x"84",
          1172 => x"08",
          1173 => x"d6",
          1174 => x"f8",
          1175 => x"d5",
          1176 => x"05",
          1177 => x"d5",
          1178 => x"05",
          1179 => x"84",
          1180 => x"39",
          1181 => x"08",
          1182 => x"82",
          1183 => x"55",
          1184 => x"70",
          1185 => x"53",
          1186 => x"84",
          1187 => x"34",
          1188 => x"08",
          1189 => x"70",
          1190 => x"53",
          1191 => x"94",
          1192 => x"84",
          1193 => x"22",
          1194 => x"53",
          1195 => x"84",
          1196 => x"23",
          1197 => x"08",
          1198 => x"70",
          1199 => x"81",
          1200 => x"53",
          1201 => x"80",
          1202 => x"d5",
          1203 => x"05",
          1204 => x"2b",
          1205 => x"08",
          1206 => x"82",
          1207 => x"cc",
          1208 => x"2c",
          1209 => x"08",
          1210 => x"82",
          1211 => x"f4",
          1212 => x"53",
          1213 => x"09",
          1214 => x"38",
          1215 => x"08",
          1216 => x"fe",
          1217 => x"82",
          1218 => x"c8",
          1219 => x"39",
          1220 => x"08",
          1221 => x"ff",
          1222 => x"82",
          1223 => x"c8",
          1224 => x"d5",
          1225 => x"05",
          1226 => x"84",
          1227 => x"23",
          1228 => x"08",
          1229 => x"70",
          1230 => x"81",
          1231 => x"53",
          1232 => x"80",
          1233 => x"d5",
          1234 => x"05",
          1235 => x"2b",
          1236 => x"82",
          1237 => x"fc",
          1238 => x"51",
          1239 => x"74",
          1240 => x"82",
          1241 => x"e4",
          1242 => x"f7",
          1243 => x"72",
          1244 => x"08",
          1245 => x"9d",
          1246 => x"84",
          1247 => x"33",
          1248 => x"84",
          1249 => x"33",
          1250 => x"54",
          1251 => x"d5",
          1252 => x"05",
          1253 => x"84",
          1254 => x"22",
          1255 => x"70",
          1256 => x"51",
          1257 => x"2e",
          1258 => x"d5",
          1259 => x"05",
          1260 => x"2b",
          1261 => x"70",
          1262 => x"88",
          1263 => x"51",
          1264 => x"54",
          1265 => x"08",
          1266 => x"70",
          1267 => x"53",
          1268 => x"84",
          1269 => x"23",
          1270 => x"d5",
          1271 => x"05",
          1272 => x"2b",
          1273 => x"70",
          1274 => x"88",
          1275 => x"51",
          1276 => x"54",
          1277 => x"08",
          1278 => x"70",
          1279 => x"53",
          1280 => x"84",
          1281 => x"23",
          1282 => x"08",
          1283 => x"70",
          1284 => x"51",
          1285 => x"38",
          1286 => x"08",
          1287 => x"ff",
          1288 => x"72",
          1289 => x"08",
          1290 => x"73",
          1291 => x"90",
          1292 => x"80",
          1293 => x"38",
          1294 => x"08",
          1295 => x"52",
          1296 => x"ee",
          1297 => x"82",
          1298 => x"e4",
          1299 => x"81",
          1300 => x"06",
          1301 => x"72",
          1302 => x"38",
          1303 => x"08",
          1304 => x"52",
          1305 => x"ca",
          1306 => x"39",
          1307 => x"08",
          1308 => x"70",
          1309 => x"81",
          1310 => x"53",
          1311 => x"90",
          1312 => x"84",
          1313 => x"08",
          1314 => x"8a",
          1315 => x"39",
          1316 => x"08",
          1317 => x"70",
          1318 => x"81",
          1319 => x"53",
          1320 => x"8e",
          1321 => x"84",
          1322 => x"08",
          1323 => x"8a",
          1324 => x"d5",
          1325 => x"05",
          1326 => x"2a",
          1327 => x"51",
          1328 => x"80",
          1329 => x"82",
          1330 => x"88",
          1331 => x"b0",
          1332 => x"3f",
          1333 => x"08",
          1334 => x"53",
          1335 => x"09",
          1336 => x"38",
          1337 => x"08",
          1338 => x"52",
          1339 => x"08",
          1340 => x"51",
          1341 => x"82",
          1342 => x"e4",
          1343 => x"88",
          1344 => x"06",
          1345 => x"72",
          1346 => x"38",
          1347 => x"08",
          1348 => x"ff",
          1349 => x"72",
          1350 => x"08",
          1351 => x"73",
          1352 => x"90",
          1353 => x"80",
          1354 => x"38",
          1355 => x"08",
          1356 => x"52",
          1357 => x"fa",
          1358 => x"82",
          1359 => x"e4",
          1360 => x"83",
          1361 => x"06",
          1362 => x"72",
          1363 => x"38",
          1364 => x"08",
          1365 => x"ff",
          1366 => x"72",
          1367 => x"08",
          1368 => x"73",
          1369 => x"98",
          1370 => x"80",
          1371 => x"38",
          1372 => x"08",
          1373 => x"52",
          1374 => x"b6",
          1375 => x"82",
          1376 => x"e4",
          1377 => x"87",
          1378 => x"06",
          1379 => x"72",
          1380 => x"d5",
          1381 => x"05",
          1382 => x"54",
          1383 => x"d5",
          1384 => x"05",
          1385 => x"2b",
          1386 => x"51",
          1387 => x"25",
          1388 => x"d5",
          1389 => x"05",
          1390 => x"51",
          1391 => x"d2",
          1392 => x"84",
          1393 => x"33",
          1394 => x"e3",
          1395 => x"06",
          1396 => x"d5",
          1397 => x"05",
          1398 => x"d5",
          1399 => x"05",
          1400 => x"ce",
          1401 => x"39",
          1402 => x"08",
          1403 => x"53",
          1404 => x"2e",
          1405 => x"80",
          1406 => x"d5",
          1407 => x"05",
          1408 => x"51",
          1409 => x"d5",
          1410 => x"05",
          1411 => x"ff",
          1412 => x"72",
          1413 => x"2e",
          1414 => x"82",
          1415 => x"88",
          1416 => x"82",
          1417 => x"fc",
          1418 => x"33",
          1419 => x"84",
          1420 => x"08",
          1421 => x"d5",
          1422 => x"05",
          1423 => x"f2",
          1424 => x"39",
          1425 => x"08",
          1426 => x"53",
          1427 => x"2e",
          1428 => x"80",
          1429 => x"d5",
          1430 => x"05",
          1431 => x"51",
          1432 => x"d5",
          1433 => x"05",
          1434 => x"ff",
          1435 => x"72",
          1436 => x"2e",
          1437 => x"82",
          1438 => x"88",
          1439 => x"82",
          1440 => x"fc",
          1441 => x"33",
          1442 => x"a6",
          1443 => x"84",
          1444 => x"08",
          1445 => x"d5",
          1446 => x"05",
          1447 => x"39",
          1448 => x"08",
          1449 => x"82",
          1450 => x"a9",
          1451 => x"84",
          1452 => x"08",
          1453 => x"84",
          1454 => x"08",
          1455 => x"d5",
          1456 => x"05",
          1457 => x"84",
          1458 => x"08",
          1459 => x"53",
          1460 => x"cc",
          1461 => x"84",
          1462 => x"22",
          1463 => x"70",
          1464 => x"51",
          1465 => x"2e",
          1466 => x"82",
          1467 => x"ec",
          1468 => x"11",
          1469 => x"82",
          1470 => x"ec",
          1471 => x"90",
          1472 => x"2c",
          1473 => x"73",
          1474 => x"82",
          1475 => x"88",
          1476 => x"a0",
          1477 => x"3f",
          1478 => x"d5",
          1479 => x"05",
          1480 => x"d5",
          1481 => x"05",
          1482 => x"86",
          1483 => x"82",
          1484 => x"e4",
          1485 => x"b7",
          1486 => x"84",
          1487 => x"33",
          1488 => x"2e",
          1489 => x"a8",
          1490 => x"82",
          1491 => x"e4",
          1492 => x"0b",
          1493 => x"08",
          1494 => x"80",
          1495 => x"84",
          1496 => x"34",
          1497 => x"d5",
          1498 => x"05",
          1499 => x"39",
          1500 => x"08",
          1501 => x"52",
          1502 => x"08",
          1503 => x"51",
          1504 => x"e9",
          1505 => x"d5",
          1506 => x"05",
          1507 => x"08",
          1508 => x"84",
          1509 => x"0c",
          1510 => x"d5",
          1511 => x"05",
          1512 => x"f8",
          1513 => x"0d",
          1514 => x"0c",
          1515 => x"84",
          1516 => x"d5",
          1517 => x"3d",
          1518 => x"d8",
          1519 => x"d5",
          1520 => x"05",
          1521 => x"d5",
          1522 => x"05",
          1523 => x"dd",
          1524 => x"f8",
          1525 => x"d4",
          1526 => x"85",
          1527 => x"d5",
          1528 => x"82",
          1529 => x"02",
          1530 => x"0c",
          1531 => x"80",
          1532 => x"84",
          1533 => x"0c",
          1534 => x"08",
          1535 => x"70",
          1536 => x"81",
          1537 => x"06",
          1538 => x"51",
          1539 => x"2e",
          1540 => x"0b",
          1541 => x"08",
          1542 => x"81",
          1543 => x"d5",
          1544 => x"05",
          1545 => x"33",
          1546 => x"08",
          1547 => x"81",
          1548 => x"84",
          1549 => x"0c",
          1550 => x"d5",
          1551 => x"05",
          1552 => x"ff",
          1553 => x"80",
          1554 => x"82",
          1555 => x"82",
          1556 => x"53",
          1557 => x"08",
          1558 => x"52",
          1559 => x"51",
          1560 => x"82",
          1561 => x"53",
          1562 => x"ff",
          1563 => x"0b",
          1564 => x"08",
          1565 => x"ff",
          1566 => x"f0",
          1567 => x"f0",
          1568 => x"53",
          1569 => x"13",
          1570 => x"2d",
          1571 => x"08",
          1572 => x"2e",
          1573 => x"0b",
          1574 => x"08",
          1575 => x"82",
          1576 => x"f8",
          1577 => x"82",
          1578 => x"f4",
          1579 => x"82",
          1580 => x"f4",
          1581 => x"d4",
          1582 => x"3d",
          1583 => x"84",
          1584 => x"d5",
          1585 => x"82",
          1586 => x"fb",
          1587 => x"0b",
          1588 => x"08",
          1589 => x"82",
          1590 => x"8c",
          1591 => x"11",
          1592 => x"2a",
          1593 => x"70",
          1594 => x"51",
          1595 => x"72",
          1596 => x"38",
          1597 => x"d5",
          1598 => x"05",
          1599 => x"39",
          1600 => x"08",
          1601 => x"53",
          1602 => x"d5",
          1603 => x"05",
          1604 => x"82",
          1605 => x"88",
          1606 => x"72",
          1607 => x"08",
          1608 => x"72",
          1609 => x"53",
          1610 => x"b6",
          1611 => x"84",
          1612 => x"08",
          1613 => x"08",
          1614 => x"53",
          1615 => x"08",
          1616 => x"52",
          1617 => x"51",
          1618 => x"82",
          1619 => x"53",
          1620 => x"ff",
          1621 => x"0b",
          1622 => x"08",
          1623 => x"ff",
          1624 => x"d5",
          1625 => x"05",
          1626 => x"d5",
          1627 => x"05",
          1628 => x"d5",
          1629 => x"05",
          1630 => x"f8",
          1631 => x"0d",
          1632 => x"0c",
          1633 => x"84",
          1634 => x"d5",
          1635 => x"3d",
          1636 => x"dc",
          1637 => x"d5",
          1638 => x"05",
          1639 => x"3f",
          1640 => x"08",
          1641 => x"f8",
          1642 => x"3d",
          1643 => x"84",
          1644 => x"d5",
          1645 => x"82",
          1646 => x"fb",
          1647 => x"d5",
          1648 => x"05",
          1649 => x"33",
          1650 => x"70",
          1651 => x"81",
          1652 => x"51",
          1653 => x"80",
          1654 => x"ff",
          1655 => x"84",
          1656 => x"0c",
          1657 => x"82",
          1658 => x"8c",
          1659 => x"11",
          1660 => x"2a",
          1661 => x"51",
          1662 => x"72",
          1663 => x"db",
          1664 => x"84",
          1665 => x"08",
          1666 => x"08",
          1667 => x"54",
          1668 => x"08",
          1669 => x"25",
          1670 => x"d5",
          1671 => x"05",
          1672 => x"70",
          1673 => x"08",
          1674 => x"52",
          1675 => x"72",
          1676 => x"08",
          1677 => x"0c",
          1678 => x"08",
          1679 => x"8c",
          1680 => x"05",
          1681 => x"82",
          1682 => x"88",
          1683 => x"82",
          1684 => x"fc",
          1685 => x"53",
          1686 => x"82",
          1687 => x"8c",
          1688 => x"d5",
          1689 => x"05",
          1690 => x"d5",
          1691 => x"05",
          1692 => x"ff",
          1693 => x"12",
          1694 => x"54",
          1695 => x"d4",
          1696 => x"72",
          1697 => x"d5",
          1698 => x"05",
          1699 => x"08",
          1700 => x"12",
          1701 => x"84",
          1702 => x"08",
          1703 => x"84",
          1704 => x"0c",
          1705 => x"39",
          1706 => x"d5",
          1707 => x"05",
          1708 => x"84",
          1709 => x"08",
          1710 => x"0c",
          1711 => x"82",
          1712 => x"04",
          1713 => x"08",
          1714 => x"84",
          1715 => x"0d",
          1716 => x"08",
          1717 => x"85",
          1718 => x"81",
          1719 => x"06",
          1720 => x"52",
          1721 => x"8d",
          1722 => x"82",
          1723 => x"f8",
          1724 => x"94",
          1725 => x"84",
          1726 => x"08",
          1727 => x"70",
          1728 => x"81",
          1729 => x"51",
          1730 => x"2e",
          1731 => x"82",
          1732 => x"88",
          1733 => x"d5",
          1734 => x"05",
          1735 => x"85",
          1736 => x"ff",
          1737 => x"52",
          1738 => x"34",
          1739 => x"08",
          1740 => x"8c",
          1741 => x"05",
          1742 => x"82",
          1743 => x"88",
          1744 => x"11",
          1745 => x"d5",
          1746 => x"05",
          1747 => x"52",
          1748 => x"82",
          1749 => x"88",
          1750 => x"11",
          1751 => x"2a",
          1752 => x"51",
          1753 => x"71",
          1754 => x"d7",
          1755 => x"84",
          1756 => x"08",
          1757 => x"33",
          1758 => x"08",
          1759 => x"51",
          1760 => x"84",
          1761 => x"08",
          1762 => x"d5",
          1763 => x"05",
          1764 => x"84",
          1765 => x"08",
          1766 => x"12",
          1767 => x"07",
          1768 => x"85",
          1769 => x"0b",
          1770 => x"08",
          1771 => x"81",
          1772 => x"d5",
          1773 => x"05",
          1774 => x"81",
          1775 => x"52",
          1776 => x"82",
          1777 => x"88",
          1778 => x"d5",
          1779 => x"05",
          1780 => x"11",
          1781 => x"71",
          1782 => x"f8",
          1783 => x"d5",
          1784 => x"05",
          1785 => x"d5",
          1786 => x"05",
          1787 => x"80",
          1788 => x"d5",
          1789 => x"05",
          1790 => x"84",
          1791 => x"0c",
          1792 => x"08",
          1793 => x"85",
          1794 => x"d5",
          1795 => x"05",
          1796 => x"d5",
          1797 => x"05",
          1798 => x"09",
          1799 => x"38",
          1800 => x"08",
          1801 => x"90",
          1802 => x"82",
          1803 => x"ec",
          1804 => x"39",
          1805 => x"08",
          1806 => x"a0",
          1807 => x"82",
          1808 => x"ec",
          1809 => x"d5",
          1810 => x"05",
          1811 => x"d5",
          1812 => x"05",
          1813 => x"34",
          1814 => x"d5",
          1815 => x"05",
          1816 => x"82",
          1817 => x"88",
          1818 => x"11",
          1819 => x"8c",
          1820 => x"d5",
          1821 => x"05",
          1822 => x"ff",
          1823 => x"d5",
          1824 => x"05",
          1825 => x"52",
          1826 => x"08",
          1827 => x"82",
          1828 => x"89",
          1829 => x"d5",
          1830 => x"82",
          1831 => x"02",
          1832 => x"0c",
          1833 => x"82",
          1834 => x"88",
          1835 => x"d5",
          1836 => x"05",
          1837 => x"84",
          1838 => x"08",
          1839 => x"08",
          1840 => x"82",
          1841 => x"90",
          1842 => x"2e",
          1843 => x"82",
          1844 => x"f8",
          1845 => x"d5",
          1846 => x"05",
          1847 => x"ac",
          1848 => x"84",
          1849 => x"08",
          1850 => x"08",
          1851 => x"05",
          1852 => x"84",
          1853 => x"08",
          1854 => x"90",
          1855 => x"84",
          1856 => x"08",
          1857 => x"08",
          1858 => x"05",
          1859 => x"08",
          1860 => x"82",
          1861 => x"f8",
          1862 => x"d5",
          1863 => x"05",
          1864 => x"d5",
          1865 => x"05",
          1866 => x"84",
          1867 => x"08",
          1868 => x"d5",
          1869 => x"05",
          1870 => x"84",
          1871 => x"08",
          1872 => x"d5",
          1873 => x"05",
          1874 => x"84",
          1875 => x"08",
          1876 => x"9c",
          1877 => x"84",
          1878 => x"08",
          1879 => x"d5",
          1880 => x"05",
          1881 => x"84",
          1882 => x"08",
          1883 => x"d5",
          1884 => x"05",
          1885 => x"84",
          1886 => x"08",
          1887 => x"08",
          1888 => x"53",
          1889 => x"71",
          1890 => x"39",
          1891 => x"08",
          1892 => x"81",
          1893 => x"84",
          1894 => x"0c",
          1895 => x"08",
          1896 => x"ff",
          1897 => x"84",
          1898 => x"0c",
          1899 => x"08",
          1900 => x"80",
          1901 => x"82",
          1902 => x"f8",
          1903 => x"70",
          1904 => x"84",
          1905 => x"08",
          1906 => x"d5",
          1907 => x"05",
          1908 => x"84",
          1909 => x"08",
          1910 => x"71",
          1911 => x"84",
          1912 => x"08",
          1913 => x"d5",
          1914 => x"05",
          1915 => x"39",
          1916 => x"08",
          1917 => x"70",
          1918 => x"0c",
          1919 => x"0d",
          1920 => x"0c",
          1921 => x"84",
          1922 => x"d5",
          1923 => x"3d",
          1924 => x"84",
          1925 => x"08",
          1926 => x"08",
          1927 => x"82",
          1928 => x"fc",
          1929 => x"71",
          1930 => x"84",
          1931 => x"08",
          1932 => x"d5",
          1933 => x"05",
          1934 => x"ff",
          1935 => x"70",
          1936 => x"38",
          1937 => x"d5",
          1938 => x"05",
          1939 => x"82",
          1940 => x"fc",
          1941 => x"d5",
          1942 => x"05",
          1943 => x"84",
          1944 => x"08",
          1945 => x"d4",
          1946 => x"84",
          1947 => x"d5",
          1948 => x"82",
          1949 => x"02",
          1950 => x"0c",
          1951 => x"82",
          1952 => x"88",
          1953 => x"d5",
          1954 => x"05",
          1955 => x"84",
          1956 => x"08",
          1957 => x"82",
          1958 => x"8c",
          1959 => x"05",
          1960 => x"08",
          1961 => x"82",
          1962 => x"fc",
          1963 => x"51",
          1964 => x"82",
          1965 => x"fc",
          1966 => x"05",
          1967 => x"08",
          1968 => x"70",
          1969 => x"51",
          1970 => x"84",
          1971 => x"39",
          1972 => x"08",
          1973 => x"70",
          1974 => x"0c",
          1975 => x"0d",
          1976 => x"0c",
          1977 => x"84",
          1978 => x"d5",
          1979 => x"3d",
          1980 => x"84",
          1981 => x"08",
          1982 => x"08",
          1983 => x"82",
          1984 => x"8c",
          1985 => x"d5",
          1986 => x"05",
          1987 => x"84",
          1988 => x"08",
          1989 => x"e5",
          1990 => x"84",
          1991 => x"08",
          1992 => x"d5",
          1993 => x"05",
          1994 => x"84",
          1995 => x"08",
          1996 => x"d5",
          1997 => x"05",
          1998 => x"84",
          1999 => x"08",
          2000 => x"38",
          2001 => x"08",
          2002 => x"51",
          2003 => x"d5",
          2004 => x"05",
          2005 => x"82",
          2006 => x"f8",
          2007 => x"d5",
          2008 => x"05",
          2009 => x"71",
          2010 => x"d5",
          2011 => x"05",
          2012 => x"82",
          2013 => x"fc",
          2014 => x"ad",
          2015 => x"84",
          2016 => x"08",
          2017 => x"f8",
          2018 => x"3d",
          2019 => x"84",
          2020 => x"d5",
          2021 => x"82",
          2022 => x"fd",
          2023 => x"d5",
          2024 => x"05",
          2025 => x"81",
          2026 => x"d5",
          2027 => x"05",
          2028 => x"33",
          2029 => x"08",
          2030 => x"81",
          2031 => x"84",
          2032 => x"0c",
          2033 => x"08",
          2034 => x"70",
          2035 => x"ff",
          2036 => x"54",
          2037 => x"2e",
          2038 => x"ce",
          2039 => x"84",
          2040 => x"08",
          2041 => x"82",
          2042 => x"88",
          2043 => x"05",
          2044 => x"08",
          2045 => x"70",
          2046 => x"51",
          2047 => x"38",
          2048 => x"d5",
          2049 => x"05",
          2050 => x"39",
          2051 => x"08",
          2052 => x"ff",
          2053 => x"84",
          2054 => x"0c",
          2055 => x"08",
          2056 => x"80",
          2057 => x"ff",
          2058 => x"d5",
          2059 => x"05",
          2060 => x"80",
          2061 => x"d5",
          2062 => x"05",
          2063 => x"52",
          2064 => x"38",
          2065 => x"d5",
          2066 => x"05",
          2067 => x"39",
          2068 => x"08",
          2069 => x"ff",
          2070 => x"84",
          2071 => x"0c",
          2072 => x"08",
          2073 => x"70",
          2074 => x"70",
          2075 => x"0b",
          2076 => x"08",
          2077 => x"ae",
          2078 => x"84",
          2079 => x"08",
          2080 => x"d5",
          2081 => x"05",
          2082 => x"72",
          2083 => x"82",
          2084 => x"fc",
          2085 => x"55",
          2086 => x"8a",
          2087 => x"82",
          2088 => x"fc",
          2089 => x"d5",
          2090 => x"05",
          2091 => x"f8",
          2092 => x"0d",
          2093 => x"0c",
          2094 => x"84",
          2095 => x"d5",
          2096 => x"3d",
          2097 => x"84",
          2098 => x"08",
          2099 => x"84",
          2100 => x"08",
          2101 => x"3f",
          2102 => x"08",
          2103 => x"84",
          2104 => x"0c",
          2105 => x"08",
          2106 => x"81",
          2107 => x"51",
          2108 => x"b2",
          2109 => x"f8",
          2110 => x"d5",
          2111 => x"05",
          2112 => x"d5",
          2113 => x"05",
          2114 => x"80",
          2115 => x"84",
          2116 => x"0c",
          2117 => x"d5",
          2118 => x"05",
          2119 => x"84",
          2120 => x"08",
          2121 => x"74",
          2122 => x"84",
          2123 => x"08",
          2124 => x"84",
          2125 => x"08",
          2126 => x"84",
          2127 => x"08",
          2128 => x"3f",
          2129 => x"08",
          2130 => x"84",
          2131 => x"0c",
          2132 => x"84",
          2133 => x"08",
          2134 => x"0c",
          2135 => x"82",
          2136 => x"04",
          2137 => x"08",
          2138 => x"84",
          2139 => x"0d",
          2140 => x"08",
          2141 => x"82",
          2142 => x"f8",
          2143 => x"d5",
          2144 => x"05",
          2145 => x"80",
          2146 => x"84",
          2147 => x"0c",
          2148 => x"82",
          2149 => x"f8",
          2150 => x"71",
          2151 => x"84",
          2152 => x"08",
          2153 => x"d5",
          2154 => x"05",
          2155 => x"ff",
          2156 => x"70",
          2157 => x"38",
          2158 => x"08",
          2159 => x"ff",
          2160 => x"84",
          2161 => x"0c",
          2162 => x"08",
          2163 => x"ff",
          2164 => x"ff",
          2165 => x"d5",
          2166 => x"05",
          2167 => x"82",
          2168 => x"f8",
          2169 => x"d5",
          2170 => x"05",
          2171 => x"84",
          2172 => x"08",
          2173 => x"d5",
          2174 => x"05",
          2175 => x"d5",
          2176 => x"05",
          2177 => x"f8",
          2178 => x"0d",
          2179 => x"0c",
          2180 => x"84",
          2181 => x"d5",
          2182 => x"3d",
          2183 => x"84",
          2184 => x"08",
          2185 => x"08",
          2186 => x"82",
          2187 => x"90",
          2188 => x"2e",
          2189 => x"82",
          2190 => x"90",
          2191 => x"05",
          2192 => x"08",
          2193 => x"82",
          2194 => x"90",
          2195 => x"05",
          2196 => x"08",
          2197 => x"82",
          2198 => x"90",
          2199 => x"2e",
          2200 => x"d5",
          2201 => x"05",
          2202 => x"82",
          2203 => x"fc",
          2204 => x"52",
          2205 => x"82",
          2206 => x"fc",
          2207 => x"05",
          2208 => x"08",
          2209 => x"ff",
          2210 => x"d5",
          2211 => x"05",
          2212 => x"d4",
          2213 => x"84",
          2214 => x"d5",
          2215 => x"82",
          2216 => x"02",
          2217 => x"0c",
          2218 => x"80",
          2219 => x"84",
          2220 => x"0c",
          2221 => x"08",
          2222 => x"80",
          2223 => x"82",
          2224 => x"88",
          2225 => x"82",
          2226 => x"88",
          2227 => x"0b",
          2228 => x"08",
          2229 => x"82",
          2230 => x"fc",
          2231 => x"38",
          2232 => x"d5",
          2233 => x"05",
          2234 => x"84",
          2235 => x"08",
          2236 => x"08",
          2237 => x"82",
          2238 => x"8c",
          2239 => x"25",
          2240 => x"d5",
          2241 => x"05",
          2242 => x"d5",
          2243 => x"05",
          2244 => x"82",
          2245 => x"f0",
          2246 => x"d5",
          2247 => x"05",
          2248 => x"81",
          2249 => x"84",
          2250 => x"0c",
          2251 => x"08",
          2252 => x"82",
          2253 => x"fc",
          2254 => x"53",
          2255 => x"08",
          2256 => x"52",
          2257 => x"08",
          2258 => x"51",
          2259 => x"82",
          2260 => x"70",
          2261 => x"08",
          2262 => x"54",
          2263 => x"08",
          2264 => x"80",
          2265 => x"82",
          2266 => x"f8",
          2267 => x"82",
          2268 => x"f8",
          2269 => x"d5",
          2270 => x"05",
          2271 => x"d4",
          2272 => x"89",
          2273 => x"d5",
          2274 => x"82",
          2275 => x"02",
          2276 => x"0c",
          2277 => x"80",
          2278 => x"84",
          2279 => x"0c",
          2280 => x"08",
          2281 => x"80",
          2282 => x"82",
          2283 => x"88",
          2284 => x"82",
          2285 => x"88",
          2286 => x"0b",
          2287 => x"08",
          2288 => x"82",
          2289 => x"8c",
          2290 => x"25",
          2291 => x"d5",
          2292 => x"05",
          2293 => x"d5",
          2294 => x"05",
          2295 => x"82",
          2296 => x"8c",
          2297 => x"82",
          2298 => x"88",
          2299 => x"81",
          2300 => x"d4",
          2301 => x"82",
          2302 => x"f8",
          2303 => x"82",
          2304 => x"fc",
          2305 => x"2e",
          2306 => x"d5",
          2307 => x"05",
          2308 => x"d5",
          2309 => x"05",
          2310 => x"84",
          2311 => x"08",
          2312 => x"f8",
          2313 => x"3d",
          2314 => x"84",
          2315 => x"d5",
          2316 => x"82",
          2317 => x"fd",
          2318 => x"53",
          2319 => x"08",
          2320 => x"52",
          2321 => x"08",
          2322 => x"51",
          2323 => x"82",
          2324 => x"70",
          2325 => x"0c",
          2326 => x"0d",
          2327 => x"0c",
          2328 => x"84",
          2329 => x"d5",
          2330 => x"3d",
          2331 => x"82",
          2332 => x"8c",
          2333 => x"82",
          2334 => x"88",
          2335 => x"93",
          2336 => x"f8",
          2337 => x"d4",
          2338 => x"85",
          2339 => x"d5",
          2340 => x"82",
          2341 => x"02",
          2342 => x"0c",
          2343 => x"81",
          2344 => x"84",
          2345 => x"0c",
          2346 => x"d5",
          2347 => x"05",
          2348 => x"84",
          2349 => x"08",
          2350 => x"08",
          2351 => x"27",
          2352 => x"d5",
          2353 => x"05",
          2354 => x"ae",
          2355 => x"82",
          2356 => x"8c",
          2357 => x"a2",
          2358 => x"84",
          2359 => x"08",
          2360 => x"84",
          2361 => x"0c",
          2362 => x"08",
          2363 => x"10",
          2364 => x"08",
          2365 => x"ff",
          2366 => x"d5",
          2367 => x"05",
          2368 => x"80",
          2369 => x"d5",
          2370 => x"05",
          2371 => x"84",
          2372 => x"08",
          2373 => x"82",
          2374 => x"88",
          2375 => x"d5",
          2376 => x"05",
          2377 => x"d5",
          2378 => x"05",
          2379 => x"84",
          2380 => x"08",
          2381 => x"08",
          2382 => x"07",
          2383 => x"08",
          2384 => x"82",
          2385 => x"fc",
          2386 => x"2a",
          2387 => x"08",
          2388 => x"82",
          2389 => x"8c",
          2390 => x"2a",
          2391 => x"08",
          2392 => x"ff",
          2393 => x"d5",
          2394 => x"05",
          2395 => x"93",
          2396 => x"84",
          2397 => x"08",
          2398 => x"84",
          2399 => x"0c",
          2400 => x"82",
          2401 => x"f8",
          2402 => x"82",
          2403 => x"f4",
          2404 => x"82",
          2405 => x"f4",
          2406 => x"d4",
          2407 => x"3d",
          2408 => x"84",
          2409 => x"d5",
          2410 => x"82",
          2411 => x"f7",
          2412 => x"0b",
          2413 => x"08",
          2414 => x"82",
          2415 => x"8c",
          2416 => x"80",
          2417 => x"d5",
          2418 => x"05",
          2419 => x"51",
          2420 => x"53",
          2421 => x"84",
          2422 => x"34",
          2423 => x"06",
          2424 => x"2e",
          2425 => x"91",
          2426 => x"84",
          2427 => x"08",
          2428 => x"05",
          2429 => x"ce",
          2430 => x"84",
          2431 => x"33",
          2432 => x"2e",
          2433 => x"a4",
          2434 => x"82",
          2435 => x"f0",
          2436 => x"d5",
          2437 => x"05",
          2438 => x"81",
          2439 => x"70",
          2440 => x"72",
          2441 => x"84",
          2442 => x"34",
          2443 => x"08",
          2444 => x"53",
          2445 => x"09",
          2446 => x"dc",
          2447 => x"84",
          2448 => x"08",
          2449 => x"05",
          2450 => x"08",
          2451 => x"33",
          2452 => x"08",
          2453 => x"82",
          2454 => x"f8",
          2455 => x"d5",
          2456 => x"05",
          2457 => x"84",
          2458 => x"08",
          2459 => x"b6",
          2460 => x"84",
          2461 => x"08",
          2462 => x"84",
          2463 => x"39",
          2464 => x"d5",
          2465 => x"05",
          2466 => x"84",
          2467 => x"08",
          2468 => x"05",
          2469 => x"08",
          2470 => x"33",
          2471 => x"08",
          2472 => x"81",
          2473 => x"0b",
          2474 => x"08",
          2475 => x"82",
          2476 => x"88",
          2477 => x"08",
          2478 => x"0c",
          2479 => x"53",
          2480 => x"d5",
          2481 => x"05",
          2482 => x"39",
          2483 => x"08",
          2484 => x"53",
          2485 => x"8d",
          2486 => x"82",
          2487 => x"ec",
          2488 => x"80",
          2489 => x"84",
          2490 => x"33",
          2491 => x"27",
          2492 => x"d5",
          2493 => x"05",
          2494 => x"b9",
          2495 => x"8d",
          2496 => x"82",
          2497 => x"ec",
          2498 => x"d8",
          2499 => x"82",
          2500 => x"f4",
          2501 => x"39",
          2502 => x"08",
          2503 => x"53",
          2504 => x"90",
          2505 => x"84",
          2506 => x"33",
          2507 => x"26",
          2508 => x"39",
          2509 => x"d5",
          2510 => x"05",
          2511 => x"39",
          2512 => x"d5",
          2513 => x"05",
          2514 => x"82",
          2515 => x"fc",
          2516 => x"d5",
          2517 => x"05",
          2518 => x"73",
          2519 => x"38",
          2520 => x"08",
          2521 => x"53",
          2522 => x"27",
          2523 => x"d5",
          2524 => x"05",
          2525 => x"51",
          2526 => x"d5",
          2527 => x"05",
          2528 => x"84",
          2529 => x"33",
          2530 => x"53",
          2531 => x"84",
          2532 => x"34",
          2533 => x"08",
          2534 => x"53",
          2535 => x"ad",
          2536 => x"84",
          2537 => x"33",
          2538 => x"53",
          2539 => x"84",
          2540 => x"34",
          2541 => x"08",
          2542 => x"53",
          2543 => x"8d",
          2544 => x"82",
          2545 => x"ec",
          2546 => x"98",
          2547 => x"84",
          2548 => x"33",
          2549 => x"08",
          2550 => x"54",
          2551 => x"26",
          2552 => x"0b",
          2553 => x"08",
          2554 => x"80",
          2555 => x"d5",
          2556 => x"05",
          2557 => x"d5",
          2558 => x"05",
          2559 => x"d5",
          2560 => x"05",
          2561 => x"82",
          2562 => x"fc",
          2563 => x"d5",
          2564 => x"05",
          2565 => x"81",
          2566 => x"70",
          2567 => x"52",
          2568 => x"33",
          2569 => x"08",
          2570 => x"fe",
          2571 => x"d5",
          2572 => x"05",
          2573 => x"80",
          2574 => x"82",
          2575 => x"fc",
          2576 => x"82",
          2577 => x"fc",
          2578 => x"d5",
          2579 => x"05",
          2580 => x"84",
          2581 => x"08",
          2582 => x"81",
          2583 => x"84",
          2584 => x"0c",
          2585 => x"08",
          2586 => x"82",
          2587 => x"8b",
          2588 => x"d5",
          2589 => x"82",
          2590 => x"02",
          2591 => x"0c",
          2592 => x"80",
          2593 => x"84",
          2594 => x"34",
          2595 => x"08",
          2596 => x"53",
          2597 => x"82",
          2598 => x"88",
          2599 => x"08",
          2600 => x"33",
          2601 => x"d5",
          2602 => x"05",
          2603 => x"ff",
          2604 => x"a0",
          2605 => x"06",
          2606 => x"d5",
          2607 => x"05",
          2608 => x"81",
          2609 => x"53",
          2610 => x"d5",
          2611 => x"05",
          2612 => x"ad",
          2613 => x"06",
          2614 => x"0b",
          2615 => x"08",
          2616 => x"82",
          2617 => x"88",
          2618 => x"08",
          2619 => x"0c",
          2620 => x"53",
          2621 => x"d5",
          2622 => x"05",
          2623 => x"84",
          2624 => x"33",
          2625 => x"2e",
          2626 => x"81",
          2627 => x"d5",
          2628 => x"05",
          2629 => x"81",
          2630 => x"70",
          2631 => x"72",
          2632 => x"84",
          2633 => x"34",
          2634 => x"08",
          2635 => x"82",
          2636 => x"e8",
          2637 => x"d5",
          2638 => x"05",
          2639 => x"2e",
          2640 => x"d5",
          2641 => x"05",
          2642 => x"2e",
          2643 => x"cd",
          2644 => x"82",
          2645 => x"f4",
          2646 => x"d5",
          2647 => x"05",
          2648 => x"81",
          2649 => x"70",
          2650 => x"72",
          2651 => x"84",
          2652 => x"34",
          2653 => x"82",
          2654 => x"84",
          2655 => x"34",
          2656 => x"08",
          2657 => x"70",
          2658 => x"71",
          2659 => x"51",
          2660 => x"82",
          2661 => x"f8",
          2662 => x"fe",
          2663 => x"84",
          2664 => x"33",
          2665 => x"26",
          2666 => x"0b",
          2667 => x"08",
          2668 => x"83",
          2669 => x"d5",
          2670 => x"05",
          2671 => x"73",
          2672 => x"82",
          2673 => x"f8",
          2674 => x"72",
          2675 => x"38",
          2676 => x"0b",
          2677 => x"08",
          2678 => x"82",
          2679 => x"0b",
          2680 => x"08",
          2681 => x"b2",
          2682 => x"84",
          2683 => x"33",
          2684 => x"27",
          2685 => x"d5",
          2686 => x"05",
          2687 => x"b9",
          2688 => x"8d",
          2689 => x"82",
          2690 => x"ec",
          2691 => x"a5",
          2692 => x"82",
          2693 => x"f4",
          2694 => x"0b",
          2695 => x"08",
          2696 => x"82",
          2697 => x"f8",
          2698 => x"a0",
          2699 => x"cf",
          2700 => x"84",
          2701 => x"33",
          2702 => x"73",
          2703 => x"82",
          2704 => x"f8",
          2705 => x"11",
          2706 => x"82",
          2707 => x"f8",
          2708 => x"d5",
          2709 => x"05",
          2710 => x"51",
          2711 => x"d5",
          2712 => x"05",
          2713 => x"84",
          2714 => x"33",
          2715 => x"27",
          2716 => x"d5",
          2717 => x"05",
          2718 => x"51",
          2719 => x"d5",
          2720 => x"05",
          2721 => x"84",
          2722 => x"33",
          2723 => x"26",
          2724 => x"0b",
          2725 => x"08",
          2726 => x"81",
          2727 => x"d5",
          2728 => x"05",
          2729 => x"84",
          2730 => x"33",
          2731 => x"74",
          2732 => x"80",
          2733 => x"84",
          2734 => x"0c",
          2735 => x"82",
          2736 => x"f4",
          2737 => x"82",
          2738 => x"fc",
          2739 => x"82",
          2740 => x"f8",
          2741 => x"12",
          2742 => x"08",
          2743 => x"82",
          2744 => x"88",
          2745 => x"08",
          2746 => x"0c",
          2747 => x"51",
          2748 => x"72",
          2749 => x"84",
          2750 => x"34",
          2751 => x"82",
          2752 => x"f0",
          2753 => x"72",
          2754 => x"38",
          2755 => x"08",
          2756 => x"30",
          2757 => x"08",
          2758 => x"82",
          2759 => x"8c",
          2760 => x"d5",
          2761 => x"05",
          2762 => x"53",
          2763 => x"d5",
          2764 => x"05",
          2765 => x"84",
          2766 => x"08",
          2767 => x"0c",
          2768 => x"82",
          2769 => x"04",
          2770 => x"7a",
          2771 => x"56",
          2772 => x"80",
          2773 => x"38",
          2774 => x"15",
          2775 => x"16",
          2776 => x"d2",
          2777 => x"54",
          2778 => x"09",
          2779 => x"38",
          2780 => x"f1",
          2781 => x"76",
          2782 => x"cf",
          2783 => x"08",
          2784 => x"81",
          2785 => x"f8",
          2786 => x"f8",
          2787 => x"53",
          2788 => x"58",
          2789 => x"82",
          2790 => x"8b",
          2791 => x"33",
          2792 => x"2e",
          2793 => x"81",
          2794 => x"ff",
          2795 => x"99",
          2796 => x"38",
          2797 => x"82",
          2798 => x"8a",
          2799 => x"ff",
          2800 => x"52",
          2801 => x"81",
          2802 => x"84",
          2803 => x"98",
          2804 => x"08",
          2805 => x"88",
          2806 => x"39",
          2807 => x"51",
          2808 => x"82",
          2809 => x"80",
          2810 => x"b2",
          2811 => x"eb",
          2812 => x"c4",
          2813 => x"39",
          2814 => x"51",
          2815 => x"82",
          2816 => x"80",
          2817 => x"b2",
          2818 => x"cf",
          2819 => x"90",
          2820 => x"39",
          2821 => x"51",
          2822 => x"82",
          2823 => x"bb",
          2824 => x"dc",
          2825 => x"82",
          2826 => x"af",
          2827 => x"98",
          2828 => x"82",
          2829 => x"a3",
          2830 => x"c8",
          2831 => x"82",
          2832 => x"97",
          2833 => x"f0",
          2834 => x"82",
          2835 => x"8b",
          2836 => x"a0",
          2837 => x"82",
          2838 => x"d7",
          2839 => x"3d",
          2840 => x"3d",
          2841 => x"56",
          2842 => x"e7",
          2843 => x"74",
          2844 => x"e8",
          2845 => x"39",
          2846 => x"74",
          2847 => x"3f",
          2848 => x"08",
          2849 => x"ef",
          2850 => x"d4",
          2851 => x"79",
          2852 => x"82",
          2853 => x"ff",
          2854 => x"87",
          2855 => x"ec",
          2856 => x"02",
          2857 => x"e3",
          2858 => x"57",
          2859 => x"30",
          2860 => x"73",
          2861 => x"59",
          2862 => x"77",
          2863 => x"83",
          2864 => x"74",
          2865 => x"81",
          2866 => x"55",
          2867 => x"81",
          2868 => x"53",
          2869 => x"3d",
          2870 => x"81",
          2871 => x"82",
          2872 => x"57",
          2873 => x"08",
          2874 => x"d4",
          2875 => x"c0",
          2876 => x"82",
          2877 => x"59",
          2878 => x"05",
          2879 => x"53",
          2880 => x"51",
          2881 => x"3f",
          2882 => x"08",
          2883 => x"f8",
          2884 => x"7a",
          2885 => x"2e",
          2886 => x"19",
          2887 => x"59",
          2888 => x"3d",
          2889 => x"81",
          2890 => x"76",
          2891 => x"07",
          2892 => x"30",
          2893 => x"72",
          2894 => x"51",
          2895 => x"2e",
          2896 => x"b5",
          2897 => x"c0",
          2898 => x"52",
          2899 => x"92",
          2900 => x"75",
          2901 => x"0c",
          2902 => x"04",
          2903 => x"7d",
          2904 => x"bb",
          2905 => x"5a",
          2906 => x"53",
          2907 => x"51",
          2908 => x"82",
          2909 => x"80",
          2910 => x"80",
          2911 => x"77",
          2912 => x"38",
          2913 => x"f0",
          2914 => x"f0",
          2915 => x"f0",
          2916 => x"f0",
          2917 => x"82",
          2918 => x"53",
          2919 => x"08",
          2920 => x"e8",
          2921 => x"b0",
          2922 => x"d8",
          2923 => x"61",
          2924 => x"f8",
          2925 => x"7f",
          2926 => x"82",
          2927 => x"59",
          2928 => x"04",
          2929 => x"f8",
          2930 => x"0d",
          2931 => x"0d",
          2932 => x"02",
          2933 => x"cf",
          2934 => x"73",
          2935 => x"5f",
          2936 => x"5e",
          2937 => x"82",
          2938 => x"ff",
          2939 => x"82",
          2940 => x"ff",
          2941 => x"80",
          2942 => x"27",
          2943 => x"7b",
          2944 => x"38",
          2945 => x"a7",
          2946 => x"39",
          2947 => x"72",
          2948 => x"38",
          2949 => x"82",
          2950 => x"ff",
          2951 => x"89",
          2952 => x"b4",
          2953 => x"b0",
          2954 => x"55",
          2955 => x"74",
          2956 => x"7a",
          2957 => x"72",
          2958 => x"b6",
          2959 => x"b7",
          2960 => x"39",
          2961 => x"51",
          2962 => x"3f",
          2963 => x"a1",
          2964 => x"53",
          2965 => x"8e",
          2966 => x"52",
          2967 => x"51",
          2968 => x"3f",
          2969 => x"b6",
          2970 => x"b6",
          2971 => x"15",
          2972 => x"dc",
          2973 => x"51",
          2974 => x"fe",
          2975 => x"b6",
          2976 => x"b6",
          2977 => x"55",
          2978 => x"80",
          2979 => x"18",
          2980 => x"53",
          2981 => x"7a",
          2982 => x"81",
          2983 => x"9f",
          2984 => x"38",
          2985 => x"73",
          2986 => x"ff",
          2987 => x"72",
          2988 => x"38",
          2989 => x"26",
          2990 => x"f0",
          2991 => x"73",
          2992 => x"82",
          2993 => x"52",
          2994 => x"e6",
          2995 => x"55",
          2996 => x"82",
          2997 => x"d2",
          2998 => x"18",
          2999 => x"58",
          3000 => x"82",
          3001 => x"98",
          3002 => x"2c",
          3003 => x"a0",
          3004 => x"06",
          3005 => x"a7",
          3006 => x"f8",
          3007 => x"70",
          3008 => x"a0",
          3009 => x"72",
          3010 => x"30",
          3011 => x"73",
          3012 => x"51",
          3013 => x"57",
          3014 => x"73",
          3015 => x"76",
          3016 => x"81",
          3017 => x"80",
          3018 => x"7c",
          3019 => x"78",
          3020 => x"38",
          3021 => x"82",
          3022 => x"8f",
          3023 => x"fc",
          3024 => x"9b",
          3025 => x"b6",
          3026 => x"b6",
          3027 => x"ff",
          3028 => x"82",
          3029 => x"51",
          3030 => x"82",
          3031 => x"82",
          3032 => x"82",
          3033 => x"52",
          3034 => x"51",
          3035 => x"3f",
          3036 => x"84",
          3037 => x"3f",
          3038 => x"04",
          3039 => x"87",
          3040 => x"08",
          3041 => x"3f",
          3042 => x"80",
          3043 => x"90",
          3044 => x"3f",
          3045 => x"f4",
          3046 => x"2a",
          3047 => x"51",
          3048 => x"2e",
          3049 => x"51",
          3050 => x"82",
          3051 => x"99",
          3052 => x"51",
          3053 => x"72",
          3054 => x"81",
          3055 => x"71",
          3056 => x"38",
          3057 => x"c4",
          3058 => x"b8",
          3059 => x"3f",
          3060 => x"b8",
          3061 => x"2a",
          3062 => x"51",
          3063 => x"2e",
          3064 => x"51",
          3065 => x"82",
          3066 => x"99",
          3067 => x"51",
          3068 => x"72",
          3069 => x"81",
          3070 => x"71",
          3071 => x"38",
          3072 => x"88",
          3073 => x"dc",
          3074 => x"3f",
          3075 => x"fc",
          3076 => x"2a",
          3077 => x"51",
          3078 => x"2e",
          3079 => x"51",
          3080 => x"82",
          3081 => x"98",
          3082 => x"51",
          3083 => x"72",
          3084 => x"81",
          3085 => x"71",
          3086 => x"38",
          3087 => x"cc",
          3088 => x"84",
          3089 => x"3f",
          3090 => x"c0",
          3091 => x"2a",
          3092 => x"51",
          3093 => x"2e",
          3094 => x"51",
          3095 => x"82",
          3096 => x"98",
          3097 => x"51",
          3098 => x"72",
          3099 => x"81",
          3100 => x"71",
          3101 => x"38",
          3102 => x"90",
          3103 => x"ac",
          3104 => x"3f",
          3105 => x"84",
          3106 => x"3f",
          3107 => x"04",
          3108 => x"77",
          3109 => x"a3",
          3110 => x"55",
          3111 => x"52",
          3112 => x"ed",
          3113 => x"82",
          3114 => x"54",
          3115 => x"81",
          3116 => x"e8",
          3117 => x"88",
          3118 => x"af",
          3119 => x"f8",
          3120 => x"82",
          3121 => x"07",
          3122 => x"71",
          3123 => x"54",
          3124 => x"82",
          3125 => x"0b",
          3126 => x"f4",
          3127 => x"81",
          3128 => x"06",
          3129 => x"ec",
          3130 => x"52",
          3131 => x"c4",
          3132 => x"d4",
          3133 => x"2e",
          3134 => x"d4",
          3135 => x"cd",
          3136 => x"39",
          3137 => x"51",
          3138 => x"3f",
          3139 => x"0b",
          3140 => x"34",
          3141 => x"cf",
          3142 => x"73",
          3143 => x"81",
          3144 => x"82",
          3145 => x"74",
          3146 => x"aa",
          3147 => x"0b",
          3148 => x"0c",
          3149 => x"04",
          3150 => x"80",
          3151 => x"ff",
          3152 => x"84",
          3153 => x"52",
          3154 => x"c7",
          3155 => x"d4",
          3156 => x"ff",
          3157 => x"7e",
          3158 => x"06",
          3159 => x"3d",
          3160 => x"82",
          3161 => x"78",
          3162 => x"3f",
          3163 => x"52",
          3164 => x"51",
          3165 => x"3f",
          3166 => x"08",
          3167 => x"38",
          3168 => x"51",
          3169 => x"81",
          3170 => x"82",
          3171 => x"ff",
          3172 => x"97",
          3173 => x"5a",
          3174 => x"79",
          3175 => x"3f",
          3176 => x"84",
          3177 => x"a0",
          3178 => x"f8",
          3179 => x"70",
          3180 => x"59",
          3181 => x"2e",
          3182 => x"78",
          3183 => x"b2",
          3184 => x"2e",
          3185 => x"78",
          3186 => x"38",
          3187 => x"ff",
          3188 => x"bc",
          3189 => x"38",
          3190 => x"78",
          3191 => x"83",
          3192 => x"80",
          3193 => x"cd",
          3194 => x"2e",
          3195 => x"8a",
          3196 => x"80",
          3197 => x"db",
          3198 => x"f9",
          3199 => x"78",
          3200 => x"88",
          3201 => x"80",
          3202 => x"a3",
          3203 => x"39",
          3204 => x"2e",
          3205 => x"78",
          3206 => x"8b",
          3207 => x"82",
          3208 => x"38",
          3209 => x"78",
          3210 => x"89",
          3211 => x"80",
          3212 => x"ff",
          3213 => x"ff",
          3214 => x"ec",
          3215 => x"d4",
          3216 => x"2e",
          3217 => x"b5",
          3218 => x"11",
          3219 => x"05",
          3220 => x"3f",
          3221 => x"08",
          3222 => x"af",
          3223 => x"fe",
          3224 => x"ff",
          3225 => x"ec",
          3226 => x"d4",
          3227 => x"38",
          3228 => x"08",
          3229 => x"c0",
          3230 => x"dc",
          3231 => x"5c",
          3232 => x"27",
          3233 => x"62",
          3234 => x"70",
          3235 => x"0c",
          3236 => x"f5",
          3237 => x"39",
          3238 => x"80",
          3239 => x"84",
          3240 => x"d3",
          3241 => x"f8",
          3242 => x"fd",
          3243 => x"3d",
          3244 => x"53",
          3245 => x"51",
          3246 => x"82",
          3247 => x"80",
          3248 => x"38",
          3249 => x"f8",
          3250 => x"84",
          3251 => x"a7",
          3252 => x"f8",
          3253 => x"fd",
          3254 => x"b9",
          3255 => x"ad",
          3256 => x"5a",
          3257 => x"81",
          3258 => x"59",
          3259 => x"05",
          3260 => x"34",
          3261 => x"43",
          3262 => x"3d",
          3263 => x"53",
          3264 => x"51",
          3265 => x"82",
          3266 => x"80",
          3267 => x"38",
          3268 => x"fc",
          3269 => x"84",
          3270 => x"db",
          3271 => x"f8",
          3272 => x"fc",
          3273 => x"3d",
          3274 => x"53",
          3275 => x"51",
          3276 => x"82",
          3277 => x"80",
          3278 => x"38",
          3279 => x"51",
          3280 => x"3f",
          3281 => x"64",
          3282 => x"62",
          3283 => x"33",
          3284 => x"78",
          3285 => x"38",
          3286 => x"54",
          3287 => x"79",
          3288 => x"ec",
          3289 => x"f0",
          3290 => x"63",
          3291 => x"5a",
          3292 => x"51",
          3293 => x"fc",
          3294 => x"3d",
          3295 => x"53",
          3296 => x"51",
          3297 => x"82",
          3298 => x"80",
          3299 => x"d3",
          3300 => x"78",
          3301 => x"38",
          3302 => x"08",
          3303 => x"39",
          3304 => x"33",
          3305 => x"2e",
          3306 => x"d3",
          3307 => x"bc",
          3308 => x"e6",
          3309 => x"80",
          3310 => x"82",
          3311 => x"45",
          3312 => x"d3",
          3313 => x"78",
          3314 => x"38",
          3315 => x"08",
          3316 => x"82",
          3317 => x"59",
          3318 => x"88",
          3319 => x"bc",
          3320 => x"39",
          3321 => x"08",
          3322 => x"45",
          3323 => x"fc",
          3324 => x"84",
          3325 => x"ff",
          3326 => x"f8",
          3327 => x"38",
          3328 => x"33",
          3329 => x"2e",
          3330 => x"d3",
          3331 => x"80",
          3332 => x"d3",
          3333 => x"78",
          3334 => x"38",
          3335 => x"08",
          3336 => x"82",
          3337 => x"59",
          3338 => x"88",
          3339 => x"b0",
          3340 => x"39",
          3341 => x"33",
          3342 => x"2e",
          3343 => x"d3",
          3344 => x"99",
          3345 => x"e2",
          3346 => x"80",
          3347 => x"82",
          3348 => x"44",
          3349 => x"d3",
          3350 => x"05",
          3351 => x"fe",
          3352 => x"ff",
          3353 => x"e8",
          3354 => x"d4",
          3355 => x"2e",
          3356 => x"63",
          3357 => x"88",
          3358 => x"81",
          3359 => x"32",
          3360 => x"72",
          3361 => x"70",
          3362 => x"51",
          3363 => x"80",
          3364 => x"7a",
          3365 => x"38",
          3366 => x"ba",
          3367 => x"c3",
          3368 => x"64",
          3369 => x"63",
          3370 => x"f2",
          3371 => x"ba",
          3372 => x"b1",
          3373 => x"ff",
          3374 => x"ff",
          3375 => x"e7",
          3376 => x"d4",
          3377 => x"2e",
          3378 => x"b5",
          3379 => x"11",
          3380 => x"05",
          3381 => x"3f",
          3382 => x"08",
          3383 => x"38",
          3384 => x"80",
          3385 => x"79",
          3386 => x"05",
          3387 => x"fe",
          3388 => x"ff",
          3389 => x"e6",
          3390 => x"d4",
          3391 => x"38",
          3392 => x"64",
          3393 => x"52",
          3394 => x"51",
          3395 => x"3f",
          3396 => x"08",
          3397 => x"52",
          3398 => x"aa",
          3399 => x"46",
          3400 => x"78",
          3401 => x"e3",
          3402 => x"27",
          3403 => x"3d",
          3404 => x"53",
          3405 => x"51",
          3406 => x"82",
          3407 => x"80",
          3408 => x"64",
          3409 => x"cf",
          3410 => x"34",
          3411 => x"45",
          3412 => x"82",
          3413 => x"c5",
          3414 => x"a7",
          3415 => x"fe",
          3416 => x"ff",
          3417 => x"e0",
          3418 => x"d4",
          3419 => x"2e",
          3420 => x"b5",
          3421 => x"11",
          3422 => x"05",
          3423 => x"3f",
          3424 => x"08",
          3425 => x"38",
          3426 => x"80",
          3427 => x"79",
          3428 => x"5b",
          3429 => x"b5",
          3430 => x"11",
          3431 => x"05",
          3432 => x"3f",
          3433 => x"08",
          3434 => x"df",
          3435 => x"22",
          3436 => x"ba",
          3437 => x"a8",
          3438 => x"f0",
          3439 => x"80",
          3440 => x"51",
          3441 => x"3f",
          3442 => x"33",
          3443 => x"2e",
          3444 => x"78",
          3445 => x"38",
          3446 => x"42",
          3447 => x"3d",
          3448 => x"53",
          3449 => x"51",
          3450 => x"82",
          3451 => x"80",
          3452 => x"61",
          3453 => x"c2",
          3454 => x"70",
          3455 => x"23",
          3456 => x"a9",
          3457 => x"ac",
          3458 => x"3f",
          3459 => x"b5",
          3460 => x"11",
          3461 => x"05",
          3462 => x"3f",
          3463 => x"08",
          3464 => x"e7",
          3465 => x"fe",
          3466 => x"ff",
          3467 => x"de",
          3468 => x"d4",
          3469 => x"2e",
          3470 => x"61",
          3471 => x"61",
          3472 => x"b5",
          3473 => x"11",
          3474 => x"05",
          3475 => x"3f",
          3476 => x"08",
          3477 => x"b3",
          3478 => x"08",
          3479 => x"ba",
          3480 => x"a6",
          3481 => x"f0",
          3482 => x"80",
          3483 => x"51",
          3484 => x"3f",
          3485 => x"33",
          3486 => x"2e",
          3487 => x"9f",
          3488 => x"38",
          3489 => x"f0",
          3490 => x"84",
          3491 => x"96",
          3492 => x"f8",
          3493 => x"8d",
          3494 => x"71",
          3495 => x"84",
          3496 => x"b5",
          3497 => x"ac",
          3498 => x"3f",
          3499 => x"b5",
          3500 => x"11",
          3501 => x"05",
          3502 => x"3f",
          3503 => x"08",
          3504 => x"c7",
          3505 => x"82",
          3506 => x"ff",
          3507 => x"64",
          3508 => x"b5",
          3509 => x"11",
          3510 => x"05",
          3511 => x"3f",
          3512 => x"08",
          3513 => x"a3",
          3514 => x"82",
          3515 => x"ff",
          3516 => x"64",
          3517 => x"82",
          3518 => x"80",
          3519 => x"38",
          3520 => x"08",
          3521 => x"84",
          3522 => x"cc",
          3523 => x"39",
          3524 => x"51",
          3525 => x"ff",
          3526 => x"f4",
          3527 => x"bb",
          3528 => x"bf",
          3529 => x"ff",
          3530 => x"95",
          3531 => x"39",
          3532 => x"59",
          3533 => x"f4",
          3534 => x"f8",
          3535 => x"d2",
          3536 => x"d4",
          3537 => x"82",
          3538 => x"80",
          3539 => x"38",
          3540 => x"08",
          3541 => x"ff",
          3542 => x"84",
          3543 => x"d4",
          3544 => x"7f",
          3545 => x"78",
          3546 => x"d2",
          3547 => x"f8",
          3548 => x"91",
          3549 => x"f8",
          3550 => x"81",
          3551 => x"5b",
          3552 => x"b2",
          3553 => x"24",
          3554 => x"81",
          3555 => x"80",
          3556 => x"83",
          3557 => x"80",
          3558 => x"bb",
          3559 => x"55",
          3560 => x"54",
          3561 => x"bb",
          3562 => x"3d",
          3563 => x"51",
          3564 => x"3f",
          3565 => x"52",
          3566 => x"b0",
          3567 => x"b3",
          3568 => x"7b",
          3569 => x"d4",
          3570 => x"82",
          3571 => x"b5",
          3572 => x"05",
          3573 => x"e8",
          3574 => x"7b",
          3575 => x"82",
          3576 => x"b5",
          3577 => x"05",
          3578 => x"d4",
          3579 => x"9c",
          3580 => x"a8",
          3581 => x"65",
          3582 => x"84",
          3583 => x"84",
          3584 => x"b5",
          3585 => x"05",
          3586 => x"3f",
          3587 => x"08",
          3588 => x"08",
          3589 => x"70",
          3590 => x"25",
          3591 => x"5f",
          3592 => x"83",
          3593 => x"81",
          3594 => x"06",
          3595 => x"2e",
          3596 => x"1b",
          3597 => x"06",
          3598 => x"fe",
          3599 => x"81",
          3600 => x"32",
          3601 => x"89",
          3602 => x"2e",
          3603 => x"89",
          3604 => x"fc",
          3605 => x"8b",
          3606 => x"b1",
          3607 => x"ab",
          3608 => x"8c",
          3609 => x"fb",
          3610 => x"39",
          3611 => x"80",
          3612 => x"a8",
          3613 => x"94",
          3614 => x"87",
          3615 => x"72",
          3616 => x"3f",
          3617 => x"08",
          3618 => x"c0",
          3619 => x"55",
          3620 => x"80",
          3621 => x"d7",
          3622 => x"82",
          3623 => x"07",
          3624 => x"8c",
          3625 => x"94",
          3626 => x"87",
          3627 => x"72",
          3628 => x"3f",
          3629 => x"08",
          3630 => x"c0",
          3631 => x"55",
          3632 => x"80",
          3633 => x"d6",
          3634 => x"82",
          3635 => x"07",
          3636 => x"9c",
          3637 => x"83",
          3638 => x"94",
          3639 => x"80",
          3640 => x"c0",
          3641 => x"ae",
          3642 => x"88",
          3643 => x"73",
          3644 => x"55",
          3645 => x"ff",
          3646 => x"ef",
          3647 => x"0a",
          3648 => x"b6",
          3649 => x"70",
          3650 => x"0c",
          3651 => x"fe",
          3652 => x"38",
          3653 => x"59",
          3654 => x"5a",
          3655 => x"05",
          3656 => x"80",
          3657 => x"70",
          3658 => x"0c",
          3659 => x"d8",
          3660 => x"dc",
          3661 => x"3f",
          3662 => x"82",
          3663 => x"ff",
          3664 => x"82",
          3665 => x"ff",
          3666 => x"80",
          3667 => x"92",
          3668 => x"51",
          3669 => x"ef",
          3670 => x"04",
          3671 => x"80",
          3672 => x"71",
          3673 => x"87",
          3674 => x"d4",
          3675 => x"ff",
          3676 => x"ff",
          3677 => x"72",
          3678 => x"38",
          3679 => x"f8",
          3680 => x"0d",
          3681 => x"0d",
          3682 => x"54",
          3683 => x"52",
          3684 => x"2e",
          3685 => x"72",
          3686 => x"a0",
          3687 => x"06",
          3688 => x"13",
          3689 => x"72",
          3690 => x"a2",
          3691 => x"06",
          3692 => x"13",
          3693 => x"72",
          3694 => x"2e",
          3695 => x"9f",
          3696 => x"81",
          3697 => x"72",
          3698 => x"70",
          3699 => x"38",
          3700 => x"80",
          3701 => x"73",
          3702 => x"39",
          3703 => x"80",
          3704 => x"54",
          3705 => x"83",
          3706 => x"70",
          3707 => x"38",
          3708 => x"80",
          3709 => x"54",
          3710 => x"09",
          3711 => x"38",
          3712 => x"a2",
          3713 => x"70",
          3714 => x"07",
          3715 => x"70",
          3716 => x"38",
          3717 => x"81",
          3718 => x"71",
          3719 => x"51",
          3720 => x"f8",
          3721 => x"0d",
          3722 => x"0d",
          3723 => x"08",
          3724 => x"38",
          3725 => x"05",
          3726 => x"d6",
          3727 => x"d4",
          3728 => x"38",
          3729 => x"39",
          3730 => x"82",
          3731 => x"86",
          3732 => x"fc",
          3733 => x"82",
          3734 => x"05",
          3735 => x"52",
          3736 => x"81",
          3737 => x"13",
          3738 => x"51",
          3739 => x"9e",
          3740 => x"38",
          3741 => x"51",
          3742 => x"97",
          3743 => x"38",
          3744 => x"51",
          3745 => x"bb",
          3746 => x"38",
          3747 => x"51",
          3748 => x"bb",
          3749 => x"38",
          3750 => x"55",
          3751 => x"87",
          3752 => x"d9",
          3753 => x"22",
          3754 => x"73",
          3755 => x"80",
          3756 => x"0b",
          3757 => x"9c",
          3758 => x"87",
          3759 => x"0c",
          3760 => x"87",
          3761 => x"0c",
          3762 => x"87",
          3763 => x"0c",
          3764 => x"87",
          3765 => x"0c",
          3766 => x"87",
          3767 => x"0c",
          3768 => x"87",
          3769 => x"0c",
          3770 => x"98",
          3771 => x"87",
          3772 => x"0c",
          3773 => x"c0",
          3774 => x"80",
          3775 => x"d4",
          3776 => x"3d",
          3777 => x"3d",
          3778 => x"87",
          3779 => x"5d",
          3780 => x"87",
          3781 => x"08",
          3782 => x"23",
          3783 => x"b8",
          3784 => x"82",
          3785 => x"c0",
          3786 => x"5a",
          3787 => x"34",
          3788 => x"b0",
          3789 => x"84",
          3790 => x"c0",
          3791 => x"5a",
          3792 => x"34",
          3793 => x"a8",
          3794 => x"86",
          3795 => x"c0",
          3796 => x"5c",
          3797 => x"23",
          3798 => x"a0",
          3799 => x"8a",
          3800 => x"7d",
          3801 => x"ff",
          3802 => x"7b",
          3803 => x"06",
          3804 => x"33",
          3805 => x"33",
          3806 => x"33",
          3807 => x"33",
          3808 => x"33",
          3809 => x"ff",
          3810 => x"82",
          3811 => x"ff",
          3812 => x"8f",
          3813 => x"fb",
          3814 => x"9f",
          3815 => x"d3",
          3816 => x"81",
          3817 => x"55",
          3818 => x"94",
          3819 => x"80",
          3820 => x"87",
          3821 => x"51",
          3822 => x"96",
          3823 => x"06",
          3824 => x"70",
          3825 => x"38",
          3826 => x"70",
          3827 => x"51",
          3828 => x"72",
          3829 => x"81",
          3830 => x"70",
          3831 => x"38",
          3832 => x"70",
          3833 => x"51",
          3834 => x"38",
          3835 => x"06",
          3836 => x"94",
          3837 => x"80",
          3838 => x"87",
          3839 => x"52",
          3840 => x"74",
          3841 => x"0c",
          3842 => x"04",
          3843 => x"02",
          3844 => x"70",
          3845 => x"2a",
          3846 => x"70",
          3847 => x"34",
          3848 => x"04",
          3849 => x"02",
          3850 => x"58",
          3851 => x"09",
          3852 => x"38",
          3853 => x"51",
          3854 => x"d3",
          3855 => x"81",
          3856 => x"56",
          3857 => x"84",
          3858 => x"2e",
          3859 => x"c0",
          3860 => x"72",
          3861 => x"2a",
          3862 => x"55",
          3863 => x"80",
          3864 => x"73",
          3865 => x"81",
          3866 => x"72",
          3867 => x"81",
          3868 => x"06",
          3869 => x"80",
          3870 => x"73",
          3871 => x"81",
          3872 => x"72",
          3873 => x"75",
          3874 => x"53",
          3875 => x"80",
          3876 => x"2e",
          3877 => x"c0",
          3878 => x"77",
          3879 => x"0b",
          3880 => x"0c",
          3881 => x"04",
          3882 => x"79",
          3883 => x"33",
          3884 => x"06",
          3885 => x"70",
          3886 => x"fc",
          3887 => x"ff",
          3888 => x"82",
          3889 => x"70",
          3890 => x"59",
          3891 => x"87",
          3892 => x"51",
          3893 => x"86",
          3894 => x"94",
          3895 => x"08",
          3896 => x"70",
          3897 => x"54",
          3898 => x"2e",
          3899 => x"91",
          3900 => x"06",
          3901 => x"d7",
          3902 => x"32",
          3903 => x"51",
          3904 => x"2e",
          3905 => x"93",
          3906 => x"06",
          3907 => x"ff",
          3908 => x"81",
          3909 => x"87",
          3910 => x"52",
          3911 => x"86",
          3912 => x"94",
          3913 => x"72",
          3914 => x"74",
          3915 => x"ff",
          3916 => x"57",
          3917 => x"38",
          3918 => x"f8",
          3919 => x"0d",
          3920 => x"0d",
          3921 => x"33",
          3922 => x"06",
          3923 => x"c0",
          3924 => x"72",
          3925 => x"38",
          3926 => x"94",
          3927 => x"70",
          3928 => x"81",
          3929 => x"51",
          3930 => x"e2",
          3931 => x"ff",
          3932 => x"c0",
          3933 => x"70",
          3934 => x"38",
          3935 => x"90",
          3936 => x"70",
          3937 => x"82",
          3938 => x"51",
          3939 => x"04",
          3940 => x"82",
          3941 => x"81",
          3942 => x"d4",
          3943 => x"fe",
          3944 => x"d3",
          3945 => x"81",
          3946 => x"53",
          3947 => x"84",
          3948 => x"2e",
          3949 => x"c0",
          3950 => x"71",
          3951 => x"2a",
          3952 => x"51",
          3953 => x"52",
          3954 => x"a0",
          3955 => x"ff",
          3956 => x"c0",
          3957 => x"70",
          3958 => x"38",
          3959 => x"90",
          3960 => x"70",
          3961 => x"98",
          3962 => x"51",
          3963 => x"f8",
          3964 => x"0d",
          3965 => x"0d",
          3966 => x"80",
          3967 => x"2a",
          3968 => x"51",
          3969 => x"84",
          3970 => x"c0",
          3971 => x"82",
          3972 => x"87",
          3973 => x"08",
          3974 => x"0c",
          3975 => x"94",
          3976 => x"a4",
          3977 => x"9e",
          3978 => x"d3",
          3979 => x"c0",
          3980 => x"82",
          3981 => x"87",
          3982 => x"08",
          3983 => x"0c",
          3984 => x"ac",
          3985 => x"b4",
          3986 => x"9e",
          3987 => x"d3",
          3988 => x"c0",
          3989 => x"82",
          3990 => x"87",
          3991 => x"08",
          3992 => x"0c",
          3993 => x"bc",
          3994 => x"c4",
          3995 => x"9e",
          3996 => x"d3",
          3997 => x"c0",
          3998 => x"82",
          3999 => x"87",
          4000 => x"08",
          4001 => x"d3",
          4002 => x"c0",
          4003 => x"82",
          4004 => x"87",
          4005 => x"08",
          4006 => x"0c",
          4007 => x"8c",
          4008 => x"dc",
          4009 => x"82",
          4010 => x"80",
          4011 => x"9e",
          4012 => x"84",
          4013 => x"51",
          4014 => x"80",
          4015 => x"81",
          4016 => x"d3",
          4017 => x"0b",
          4018 => x"90",
          4019 => x"80",
          4020 => x"52",
          4021 => x"2e",
          4022 => x"52",
          4023 => x"e2",
          4024 => x"87",
          4025 => x"08",
          4026 => x"0a",
          4027 => x"52",
          4028 => x"83",
          4029 => x"71",
          4030 => x"34",
          4031 => x"c0",
          4032 => x"70",
          4033 => x"06",
          4034 => x"70",
          4035 => x"38",
          4036 => x"82",
          4037 => x"80",
          4038 => x"9e",
          4039 => x"a0",
          4040 => x"51",
          4041 => x"80",
          4042 => x"81",
          4043 => x"d3",
          4044 => x"0b",
          4045 => x"90",
          4046 => x"80",
          4047 => x"52",
          4048 => x"2e",
          4049 => x"52",
          4050 => x"e6",
          4051 => x"87",
          4052 => x"08",
          4053 => x"80",
          4054 => x"52",
          4055 => x"83",
          4056 => x"71",
          4057 => x"34",
          4058 => x"c0",
          4059 => x"70",
          4060 => x"06",
          4061 => x"70",
          4062 => x"38",
          4063 => x"82",
          4064 => x"80",
          4065 => x"9e",
          4066 => x"81",
          4067 => x"51",
          4068 => x"80",
          4069 => x"81",
          4070 => x"d3",
          4071 => x"0b",
          4072 => x"90",
          4073 => x"c0",
          4074 => x"52",
          4075 => x"2e",
          4076 => x"52",
          4077 => x"ea",
          4078 => x"87",
          4079 => x"08",
          4080 => x"06",
          4081 => x"70",
          4082 => x"38",
          4083 => x"82",
          4084 => x"87",
          4085 => x"08",
          4086 => x"06",
          4087 => x"51",
          4088 => x"82",
          4089 => x"80",
          4090 => x"9e",
          4091 => x"84",
          4092 => x"52",
          4093 => x"2e",
          4094 => x"52",
          4095 => x"ed",
          4096 => x"9e",
          4097 => x"83",
          4098 => x"84",
          4099 => x"51",
          4100 => x"ee",
          4101 => x"87",
          4102 => x"08",
          4103 => x"51",
          4104 => x"80",
          4105 => x"81",
          4106 => x"d3",
          4107 => x"c0",
          4108 => x"70",
          4109 => x"51",
          4110 => x"f0",
          4111 => x"0d",
          4112 => x"0d",
          4113 => x"51",
          4114 => x"3f",
          4115 => x"33",
          4116 => x"2e",
          4117 => x"bd",
          4118 => x"92",
          4119 => x"bd",
          4120 => x"ae",
          4121 => x"d3",
          4122 => x"73",
          4123 => x"38",
          4124 => x"08",
          4125 => x"08",
          4126 => x"82",
          4127 => x"ff",
          4128 => x"82",
          4129 => x"54",
          4130 => x"94",
          4131 => x"b4",
          4132 => x"b8",
          4133 => x"52",
          4134 => x"51",
          4135 => x"3f",
          4136 => x"33",
          4137 => x"2e",
          4138 => x"d3",
          4139 => x"d3",
          4140 => x"54",
          4141 => x"ec",
          4142 => x"9c",
          4143 => x"e5",
          4144 => x"80",
          4145 => x"82",
          4146 => x"82",
          4147 => x"11",
          4148 => x"be",
          4149 => x"91",
          4150 => x"d3",
          4151 => x"73",
          4152 => x"38",
          4153 => x"08",
          4154 => x"08",
          4155 => x"82",
          4156 => x"ff",
          4157 => x"82",
          4158 => x"54",
          4159 => x"8e",
          4160 => x"ec",
          4161 => x"be",
          4162 => x"91",
          4163 => x"d3",
          4164 => x"73",
          4165 => x"38",
          4166 => x"33",
          4167 => x"e0",
          4168 => x"b4",
          4169 => x"ed",
          4170 => x"80",
          4171 => x"82",
          4172 => x"52",
          4173 => x"51",
          4174 => x"3f",
          4175 => x"33",
          4176 => x"2e",
          4177 => x"bf",
          4178 => x"ad",
          4179 => x"d3",
          4180 => x"73",
          4181 => x"38",
          4182 => x"51",
          4183 => x"3f",
          4184 => x"33",
          4185 => x"2e",
          4186 => x"bf",
          4187 => x"ac",
          4188 => x"d3",
          4189 => x"73",
          4190 => x"38",
          4191 => x"51",
          4192 => x"3f",
          4193 => x"33",
          4194 => x"2e",
          4195 => x"bf",
          4196 => x"ac",
          4197 => x"bf",
          4198 => x"ac",
          4199 => x"d3",
          4200 => x"82",
          4201 => x"ff",
          4202 => x"82",
          4203 => x"52",
          4204 => x"51",
          4205 => x"3f",
          4206 => x"08",
          4207 => x"b8",
          4208 => x"94",
          4209 => x"e0",
          4210 => x"97",
          4211 => x"d0",
          4212 => x"c0",
          4213 => x"8f",
          4214 => x"d3",
          4215 => x"bd",
          4216 => x"75",
          4217 => x"3f",
          4218 => x"08",
          4219 => x"29",
          4220 => x"54",
          4221 => x"f8",
          4222 => x"c1",
          4223 => x"8f",
          4224 => x"d3",
          4225 => x"73",
          4226 => x"38",
          4227 => x"08",
          4228 => x"c0",
          4229 => x"c4",
          4230 => x"d4",
          4231 => x"84",
          4232 => x"71",
          4233 => x"82",
          4234 => x"52",
          4235 => x"51",
          4236 => x"3f",
          4237 => x"33",
          4238 => x"2e",
          4239 => x"d3",
          4240 => x"bd",
          4241 => x"75",
          4242 => x"3f",
          4243 => x"08",
          4244 => x"29",
          4245 => x"54",
          4246 => x"f8",
          4247 => x"c1",
          4248 => x"8e",
          4249 => x"51",
          4250 => x"3f",
          4251 => x"04",
          4252 => x"02",
          4253 => x"ff",
          4254 => x"84",
          4255 => x"71",
          4256 => x"ac",
          4257 => x"71",
          4258 => x"c2",
          4259 => x"39",
          4260 => x"51",
          4261 => x"c2",
          4262 => x"39",
          4263 => x"51",
          4264 => x"c2",
          4265 => x"39",
          4266 => x"51",
          4267 => x"3f",
          4268 => x"04",
          4269 => x"0c",
          4270 => x"87",
          4271 => x"0c",
          4272 => x"f4",
          4273 => x"96",
          4274 => x"fd",
          4275 => x"98",
          4276 => x"2c",
          4277 => x"70",
          4278 => x"10",
          4279 => x"2b",
          4280 => x"54",
          4281 => x"0b",
          4282 => x"12",
          4283 => x"71",
          4284 => x"38",
          4285 => x"11",
          4286 => x"84",
          4287 => x"33",
          4288 => x"52",
          4289 => x"2e",
          4290 => x"83",
          4291 => x"72",
          4292 => x"0c",
          4293 => x"04",
          4294 => x"79",
          4295 => x"a3",
          4296 => x"33",
          4297 => x"72",
          4298 => x"38",
          4299 => x"08",
          4300 => x"ff",
          4301 => x"82",
          4302 => x"52",
          4303 => x"ac",
          4304 => x"f0",
          4305 => x"88",
          4306 => x"e6",
          4307 => x"ff",
          4308 => x"74",
          4309 => x"ff",
          4310 => x"39",
          4311 => x"8c",
          4312 => x"74",
          4313 => x"0d",
          4314 => x"0d",
          4315 => x"05",
          4316 => x"02",
          4317 => x"05",
          4318 => x"d0",
          4319 => x"29",
          4320 => x"05",
          4321 => x"59",
          4322 => x"59",
          4323 => x"86",
          4324 => x"9a",
          4325 => x"d4",
          4326 => x"84",
          4327 => x"f8",
          4328 => x"70",
          4329 => x"5a",
          4330 => x"82",
          4331 => x"75",
          4332 => x"d0",
          4333 => x"29",
          4334 => x"05",
          4335 => x"56",
          4336 => x"2e",
          4337 => x"53",
          4338 => x"51",
          4339 => x"3f",
          4340 => x"33",
          4341 => x"74",
          4342 => x"34",
          4343 => x"06",
          4344 => x"27",
          4345 => x"0b",
          4346 => x"34",
          4347 => x"b6",
          4348 => x"cc",
          4349 => x"80",
          4350 => x"82",
          4351 => x"55",
          4352 => x"8c",
          4353 => x"54",
          4354 => x"52",
          4355 => x"eb",
          4356 => x"d4",
          4357 => x"8a",
          4358 => x"e8",
          4359 => x"cc",
          4360 => x"ef",
          4361 => x"3d",
          4362 => x"3d",
          4363 => x"f8",
          4364 => x"72",
          4365 => x"80",
          4366 => x"71",
          4367 => x"3f",
          4368 => x"ff",
          4369 => x"54",
          4370 => x"25",
          4371 => x"0b",
          4372 => x"34",
          4373 => x"08",
          4374 => x"2e",
          4375 => x"51",
          4376 => x"3f",
          4377 => x"08",
          4378 => x"3f",
          4379 => x"d4",
          4380 => x"3d",
          4381 => x"3d",
          4382 => x"80",
          4383 => x"cc",
          4384 => x"f5",
          4385 => x"d4",
          4386 => x"d3",
          4387 => x"cc",
          4388 => x"f8",
          4389 => x"70",
          4390 => x"9d",
          4391 => x"d4",
          4392 => x"2e",
          4393 => x"51",
          4394 => x"3f",
          4395 => x"08",
          4396 => x"82",
          4397 => x"25",
          4398 => x"d4",
          4399 => x"05",
          4400 => x"55",
          4401 => x"75",
          4402 => x"81",
          4403 => x"b4",
          4404 => x"8a",
          4405 => x"ff",
          4406 => x"06",
          4407 => x"a6",
          4408 => x"d9",
          4409 => x"3d",
          4410 => x"08",
          4411 => x"70",
          4412 => x"52",
          4413 => x"08",
          4414 => x"ac",
          4415 => x"f8",
          4416 => x"38",
          4417 => x"d4",
          4418 => x"55",
          4419 => x"8b",
          4420 => x"56",
          4421 => x"3f",
          4422 => x"08",
          4423 => x"38",
          4424 => x"b1",
          4425 => x"d4",
          4426 => x"18",
          4427 => x"0b",
          4428 => x"08",
          4429 => x"82",
          4430 => x"ff",
          4431 => x"55",
          4432 => x"34",
          4433 => x"30",
          4434 => x"9f",
          4435 => x"55",
          4436 => x"85",
          4437 => x"ac",
          4438 => x"cc",
          4439 => x"08",
          4440 => x"f3",
          4441 => x"d4",
          4442 => x"2e",
          4443 => x"c5",
          4444 => x"88",
          4445 => x"77",
          4446 => x"06",
          4447 => x"52",
          4448 => x"b1",
          4449 => x"51",
          4450 => x"3f",
          4451 => x"54",
          4452 => x"08",
          4453 => x"58",
          4454 => x"f8",
          4455 => x"0d",
          4456 => x"0d",
          4457 => x"5c",
          4458 => x"57",
          4459 => x"73",
          4460 => x"81",
          4461 => x"78",
          4462 => x"56",
          4463 => x"98",
          4464 => x"70",
          4465 => x"33",
          4466 => x"73",
          4467 => x"81",
          4468 => x"75",
          4469 => x"38",
          4470 => x"88",
          4471 => x"d4",
          4472 => x"52",
          4473 => x"9d",
          4474 => x"f8",
          4475 => x"52",
          4476 => x"ff",
          4477 => x"82",
          4478 => x"80",
          4479 => x"15",
          4480 => x"81",
          4481 => x"74",
          4482 => x"38",
          4483 => x"e6",
          4484 => x"81",
          4485 => x"3d",
          4486 => x"f8",
          4487 => x"d7",
          4488 => x"f8",
          4489 => x"9a",
          4490 => x"53",
          4491 => x"51",
          4492 => x"82",
          4493 => x"81",
          4494 => x"74",
          4495 => x"54",
          4496 => x"14",
          4497 => x"06",
          4498 => x"74",
          4499 => x"38",
          4500 => x"82",
          4501 => x"8c",
          4502 => x"d3",
          4503 => x"3d",
          4504 => x"08",
          4505 => x"59",
          4506 => x"0b",
          4507 => x"82",
          4508 => x"82",
          4509 => x"55",
          4510 => x"cb",
          4511 => x"d4",
          4512 => x"55",
          4513 => x"81",
          4514 => x"2e",
          4515 => x"81",
          4516 => x"55",
          4517 => x"2e",
          4518 => x"a8",
          4519 => x"3f",
          4520 => x"08",
          4521 => x"0c",
          4522 => x"08",
          4523 => x"92",
          4524 => x"76",
          4525 => x"f8",
          4526 => x"de",
          4527 => x"d4",
          4528 => x"2e",
          4529 => x"c5",
          4530 => x"a2",
          4531 => x"f7",
          4532 => x"f8",
          4533 => x"d4",
          4534 => x"80",
          4535 => x"3d",
          4536 => x"81",
          4537 => x"82",
          4538 => x"56",
          4539 => x"08",
          4540 => x"81",
          4541 => x"38",
          4542 => x"08",
          4543 => x"85",
          4544 => x"f8",
          4545 => x"0b",
          4546 => x"08",
          4547 => x"82",
          4548 => x"ff",
          4549 => x"55",
          4550 => x"34",
          4551 => x"81",
          4552 => x"75",
          4553 => x"3f",
          4554 => x"81",
          4555 => x"54",
          4556 => x"83",
          4557 => x"74",
          4558 => x"81",
          4559 => x"38",
          4560 => x"82",
          4561 => x"76",
          4562 => x"d4",
          4563 => x"2e",
          4564 => x"d6",
          4565 => x"5d",
          4566 => x"82",
          4567 => x"98",
          4568 => x"2c",
          4569 => x"ff",
          4570 => x"78",
          4571 => x"82",
          4572 => x"70",
          4573 => x"98",
          4574 => x"b0",
          4575 => x"2b",
          4576 => x"71",
          4577 => x"70",
          4578 => x"c2",
          4579 => x"08",
          4580 => x"51",
          4581 => x"59",
          4582 => x"5d",
          4583 => x"73",
          4584 => x"e9",
          4585 => x"27",
          4586 => x"81",
          4587 => x"81",
          4588 => x"70",
          4589 => x"55",
          4590 => x"80",
          4591 => x"53",
          4592 => x"51",
          4593 => x"82",
          4594 => x"81",
          4595 => x"73",
          4596 => x"38",
          4597 => x"b0",
          4598 => x"b1",
          4599 => x"80",
          4600 => x"80",
          4601 => x"98",
          4602 => x"ff",
          4603 => x"55",
          4604 => x"97",
          4605 => x"74",
          4606 => x"f5",
          4607 => x"d4",
          4608 => x"ff",
          4609 => x"cc",
          4610 => x"80",
          4611 => x"2e",
          4612 => x"81",
          4613 => x"82",
          4614 => x"74",
          4615 => x"98",
          4616 => x"b0",
          4617 => x"2b",
          4618 => x"70",
          4619 => x"82",
          4620 => x"c4",
          4621 => x"51",
          4622 => x"58",
          4623 => x"77",
          4624 => x"06",
          4625 => x"82",
          4626 => x"08",
          4627 => x"0b",
          4628 => x"34",
          4629 => x"ec",
          4630 => x"39",
          4631 => x"b4",
          4632 => x"ec",
          4633 => x"af",
          4634 => x"7d",
          4635 => x"73",
          4636 => x"e1",
          4637 => x"29",
          4638 => x"05",
          4639 => x"04",
          4640 => x"33",
          4641 => x"2e",
          4642 => x"82",
          4643 => x"55",
          4644 => x"ab",
          4645 => x"2b",
          4646 => x"51",
          4647 => x"24",
          4648 => x"1a",
          4649 => x"81",
          4650 => x"81",
          4651 => x"81",
          4652 => x"70",
          4653 => x"ec",
          4654 => x"51",
          4655 => x"82",
          4656 => x"81",
          4657 => x"74",
          4658 => x"34",
          4659 => x"ae",
          4660 => x"34",
          4661 => x"33",
          4662 => x"25",
          4663 => x"14",
          4664 => x"ec",
          4665 => x"ec",
          4666 => x"81",
          4667 => x"81",
          4668 => x"70",
          4669 => x"ec",
          4670 => x"51",
          4671 => x"77",
          4672 => x"82",
          4673 => x"52",
          4674 => x"33",
          4675 => x"a1",
          4676 => x"81",
          4677 => x"81",
          4678 => x"70",
          4679 => x"ec",
          4680 => x"51",
          4681 => x"24",
          4682 => x"ec",
          4683 => x"98",
          4684 => x"2c",
          4685 => x"33",
          4686 => x"56",
          4687 => x"fc",
          4688 => x"f0",
          4689 => x"88",
          4690 => x"e6",
          4691 => x"80",
          4692 => x"80",
          4693 => x"98",
          4694 => x"b8",
          4695 => x"55",
          4696 => x"de",
          4697 => x"39",
          4698 => x"80",
          4699 => x"34",
          4700 => x"53",
          4701 => x"b5",
          4702 => x"9c",
          4703 => x"39",
          4704 => x"33",
          4705 => x"06",
          4706 => x"80",
          4707 => x"38",
          4708 => x"33",
          4709 => x"73",
          4710 => x"34",
          4711 => x"73",
          4712 => x"34",
          4713 => x"08",
          4714 => x"ff",
          4715 => x"82",
          4716 => x"70",
          4717 => x"98",
          4718 => x"b8",
          4719 => x"56",
          4720 => x"25",
          4721 => x"1a",
          4722 => x"33",
          4723 => x"f0",
          4724 => x"73",
          4725 => x"9f",
          4726 => x"81",
          4727 => x"81",
          4728 => x"70",
          4729 => x"ec",
          4730 => x"51",
          4731 => x"24",
          4732 => x"f0",
          4733 => x"a0",
          4734 => x"b6",
          4735 => x"bc",
          4736 => x"2b",
          4737 => x"82",
          4738 => x"57",
          4739 => x"74",
          4740 => x"c1",
          4741 => x"dc",
          4742 => x"51",
          4743 => x"3f",
          4744 => x"0a",
          4745 => x"0a",
          4746 => x"2c",
          4747 => x"33",
          4748 => x"75",
          4749 => x"38",
          4750 => x"82",
          4751 => x"7a",
          4752 => x"74",
          4753 => x"dc",
          4754 => x"51",
          4755 => x"3f",
          4756 => x"52",
          4757 => x"c9",
          4758 => x"f8",
          4759 => x"06",
          4760 => x"38",
          4761 => x"33",
          4762 => x"2e",
          4763 => x"53",
          4764 => x"51",
          4765 => x"84",
          4766 => x"34",
          4767 => x"ec",
          4768 => x"0b",
          4769 => x"34",
          4770 => x"f8",
          4771 => x"0d",
          4772 => x"bc",
          4773 => x"80",
          4774 => x"38",
          4775 => x"08",
          4776 => x"ff",
          4777 => x"82",
          4778 => x"ff",
          4779 => x"82",
          4780 => x"73",
          4781 => x"54",
          4782 => x"ec",
          4783 => x"ec",
          4784 => x"55",
          4785 => x"f9",
          4786 => x"14",
          4787 => x"ec",
          4788 => x"98",
          4789 => x"2c",
          4790 => x"06",
          4791 => x"74",
          4792 => x"38",
          4793 => x"81",
          4794 => x"34",
          4795 => x"08",
          4796 => x"51",
          4797 => x"3f",
          4798 => x"0a",
          4799 => x"0a",
          4800 => x"2c",
          4801 => x"33",
          4802 => x"75",
          4803 => x"38",
          4804 => x"08",
          4805 => x"ff",
          4806 => x"82",
          4807 => x"70",
          4808 => x"98",
          4809 => x"b8",
          4810 => x"56",
          4811 => x"24",
          4812 => x"82",
          4813 => x"52",
          4814 => x"9c",
          4815 => x"81",
          4816 => x"81",
          4817 => x"70",
          4818 => x"ec",
          4819 => x"51",
          4820 => x"25",
          4821 => x"fd",
          4822 => x"bc",
          4823 => x"ff",
          4824 => x"b8",
          4825 => x"54",
          4826 => x"f7",
          4827 => x"f0",
          4828 => x"81",
          4829 => x"82",
          4830 => x"74",
          4831 => x"52",
          4832 => x"ae",
          4833 => x"bc",
          4834 => x"ff",
          4835 => x"b8",
          4836 => x"54",
          4837 => x"d6",
          4838 => x"39",
          4839 => x"53",
          4840 => x"b5",
          4841 => x"f0",
          4842 => x"82",
          4843 => x"80",
          4844 => x"b8",
          4845 => x"39",
          4846 => x"82",
          4847 => x"55",
          4848 => x"a6",
          4849 => x"ff",
          4850 => x"82",
          4851 => x"82",
          4852 => x"82",
          4853 => x"81",
          4854 => x"05",
          4855 => x"79",
          4856 => x"81",
          4857 => x"81",
          4858 => x"84",
          4859 => x"f8",
          4860 => x"08",
          4861 => x"80",
          4862 => x"74",
          4863 => x"85",
          4864 => x"f8",
          4865 => x"b8",
          4866 => x"f8",
          4867 => x"06",
          4868 => x"74",
          4869 => x"ff",
          4870 => x"ff",
          4871 => x"fa",
          4872 => x"55",
          4873 => x"f6",
          4874 => x"51",
          4875 => x"3f",
          4876 => x"93",
          4877 => x"06",
          4878 => x"d3",
          4879 => x"74",
          4880 => x"38",
          4881 => x"a3",
          4882 => x"d4",
          4883 => x"ec",
          4884 => x"d4",
          4885 => x"ff",
          4886 => x"53",
          4887 => x"51",
          4888 => x"3f",
          4889 => x"7a",
          4890 => x"d3",
          4891 => x"08",
          4892 => x"80",
          4893 => x"74",
          4894 => x"89",
          4895 => x"f8",
          4896 => x"b8",
          4897 => x"f8",
          4898 => x"06",
          4899 => x"74",
          4900 => x"ff",
          4901 => x"81",
          4902 => x"81",
          4903 => x"89",
          4904 => x"ec",
          4905 => x"7a",
          4906 => x"bc",
          4907 => x"b8",
          4908 => x"51",
          4909 => x"f5",
          4910 => x"ec",
          4911 => x"81",
          4912 => x"ec",
          4913 => x"56",
          4914 => x"27",
          4915 => x"82",
          4916 => x"52",
          4917 => x"73",
          4918 => x"34",
          4919 => x"33",
          4920 => x"99",
          4921 => x"ed",
          4922 => x"bc",
          4923 => x"80",
          4924 => x"38",
          4925 => x"08",
          4926 => x"ff",
          4927 => x"82",
          4928 => x"ff",
          4929 => x"82",
          4930 => x"f4",
          4931 => x"3d",
          4932 => x"f4",
          4933 => x"f0",
          4934 => x"0b",
          4935 => x"23",
          4936 => x"53",
          4937 => x"ff",
          4938 => x"a9",
          4939 => x"d4",
          4940 => x"80",
          4941 => x"34",
          4942 => x"81",
          4943 => x"d4",
          4944 => x"77",
          4945 => x"76",
          4946 => x"82",
          4947 => x"54",
          4948 => x"34",
          4949 => x"34",
          4950 => x"08",
          4951 => x"22",
          4952 => x"80",
          4953 => x"83",
          4954 => x"70",
          4955 => x"51",
          4956 => x"88",
          4957 => x"89",
          4958 => x"d4",
          4959 => x"88",
          4960 => x"f0",
          4961 => x"11",
          4962 => x"77",
          4963 => x"76",
          4964 => x"89",
          4965 => x"ff",
          4966 => x"52",
          4967 => x"72",
          4968 => x"fb",
          4969 => x"82",
          4970 => x"ff",
          4971 => x"51",
          4972 => x"d4",
          4973 => x"3d",
          4974 => x"3d",
          4975 => x"05",
          4976 => x"05",
          4977 => x"71",
          4978 => x"f0",
          4979 => x"2b",
          4980 => x"83",
          4981 => x"70",
          4982 => x"33",
          4983 => x"07",
          4984 => x"ae",
          4985 => x"81",
          4986 => x"07",
          4987 => x"53",
          4988 => x"54",
          4989 => x"53",
          4990 => x"77",
          4991 => x"18",
          4992 => x"f0",
          4993 => x"88",
          4994 => x"70",
          4995 => x"74",
          4996 => x"82",
          4997 => x"70",
          4998 => x"81",
          4999 => x"88",
          5000 => x"83",
          5001 => x"f8",
          5002 => x"56",
          5003 => x"73",
          5004 => x"06",
          5005 => x"54",
          5006 => x"82",
          5007 => x"81",
          5008 => x"72",
          5009 => x"82",
          5010 => x"16",
          5011 => x"34",
          5012 => x"34",
          5013 => x"04",
          5014 => x"82",
          5015 => x"02",
          5016 => x"05",
          5017 => x"2b",
          5018 => x"11",
          5019 => x"33",
          5020 => x"71",
          5021 => x"58",
          5022 => x"55",
          5023 => x"84",
          5024 => x"13",
          5025 => x"2b",
          5026 => x"2a",
          5027 => x"52",
          5028 => x"34",
          5029 => x"34",
          5030 => x"08",
          5031 => x"11",
          5032 => x"33",
          5033 => x"71",
          5034 => x"56",
          5035 => x"72",
          5036 => x"33",
          5037 => x"71",
          5038 => x"70",
          5039 => x"56",
          5040 => x"86",
          5041 => x"87",
          5042 => x"d4",
          5043 => x"70",
          5044 => x"33",
          5045 => x"07",
          5046 => x"ff",
          5047 => x"2a",
          5048 => x"53",
          5049 => x"34",
          5050 => x"34",
          5051 => x"04",
          5052 => x"02",
          5053 => x"82",
          5054 => x"71",
          5055 => x"11",
          5056 => x"12",
          5057 => x"2b",
          5058 => x"29",
          5059 => x"81",
          5060 => x"98",
          5061 => x"2b",
          5062 => x"53",
          5063 => x"56",
          5064 => x"71",
          5065 => x"f6",
          5066 => x"fe",
          5067 => x"d4",
          5068 => x"16",
          5069 => x"12",
          5070 => x"2b",
          5071 => x"07",
          5072 => x"33",
          5073 => x"71",
          5074 => x"70",
          5075 => x"ff",
          5076 => x"52",
          5077 => x"5a",
          5078 => x"05",
          5079 => x"54",
          5080 => x"13",
          5081 => x"13",
          5082 => x"f0",
          5083 => x"70",
          5084 => x"33",
          5085 => x"71",
          5086 => x"56",
          5087 => x"72",
          5088 => x"81",
          5089 => x"88",
          5090 => x"81",
          5091 => x"70",
          5092 => x"51",
          5093 => x"72",
          5094 => x"81",
          5095 => x"3d",
          5096 => x"3d",
          5097 => x"f0",
          5098 => x"05",
          5099 => x"70",
          5100 => x"11",
          5101 => x"83",
          5102 => x"8b",
          5103 => x"2b",
          5104 => x"59",
          5105 => x"73",
          5106 => x"81",
          5107 => x"88",
          5108 => x"8c",
          5109 => x"22",
          5110 => x"88",
          5111 => x"53",
          5112 => x"73",
          5113 => x"14",
          5114 => x"f0",
          5115 => x"70",
          5116 => x"33",
          5117 => x"71",
          5118 => x"56",
          5119 => x"72",
          5120 => x"33",
          5121 => x"71",
          5122 => x"70",
          5123 => x"55",
          5124 => x"82",
          5125 => x"83",
          5126 => x"d4",
          5127 => x"82",
          5128 => x"12",
          5129 => x"2b",
          5130 => x"f8",
          5131 => x"87",
          5132 => x"f7",
          5133 => x"82",
          5134 => x"31",
          5135 => x"83",
          5136 => x"70",
          5137 => x"fd",
          5138 => x"d4",
          5139 => x"83",
          5140 => x"82",
          5141 => x"12",
          5142 => x"2b",
          5143 => x"07",
          5144 => x"33",
          5145 => x"71",
          5146 => x"90",
          5147 => x"42",
          5148 => x"5b",
          5149 => x"54",
          5150 => x"8d",
          5151 => x"80",
          5152 => x"fe",
          5153 => x"84",
          5154 => x"33",
          5155 => x"71",
          5156 => x"83",
          5157 => x"11",
          5158 => x"53",
          5159 => x"55",
          5160 => x"34",
          5161 => x"06",
          5162 => x"14",
          5163 => x"f0",
          5164 => x"84",
          5165 => x"13",
          5166 => x"2b",
          5167 => x"2a",
          5168 => x"56",
          5169 => x"16",
          5170 => x"16",
          5171 => x"f0",
          5172 => x"80",
          5173 => x"34",
          5174 => x"14",
          5175 => x"f0",
          5176 => x"84",
          5177 => x"85",
          5178 => x"d4",
          5179 => x"70",
          5180 => x"33",
          5181 => x"07",
          5182 => x"80",
          5183 => x"2a",
          5184 => x"56",
          5185 => x"34",
          5186 => x"34",
          5187 => x"04",
          5188 => x"73",
          5189 => x"f0",
          5190 => x"f7",
          5191 => x"80",
          5192 => x"71",
          5193 => x"3f",
          5194 => x"04",
          5195 => x"80",
          5196 => x"f8",
          5197 => x"d4",
          5198 => x"ff",
          5199 => x"d4",
          5200 => x"11",
          5201 => x"33",
          5202 => x"07",
          5203 => x"56",
          5204 => x"ff",
          5205 => x"78",
          5206 => x"38",
          5207 => x"17",
          5208 => x"12",
          5209 => x"2b",
          5210 => x"ff",
          5211 => x"31",
          5212 => x"ff",
          5213 => x"27",
          5214 => x"56",
          5215 => x"79",
          5216 => x"73",
          5217 => x"38",
          5218 => x"5b",
          5219 => x"85",
          5220 => x"88",
          5221 => x"54",
          5222 => x"78",
          5223 => x"2e",
          5224 => x"79",
          5225 => x"76",
          5226 => x"d4",
          5227 => x"70",
          5228 => x"33",
          5229 => x"07",
          5230 => x"ff",
          5231 => x"5a",
          5232 => x"73",
          5233 => x"38",
          5234 => x"54",
          5235 => x"81",
          5236 => x"54",
          5237 => x"81",
          5238 => x"7a",
          5239 => x"06",
          5240 => x"51",
          5241 => x"81",
          5242 => x"80",
          5243 => x"52",
          5244 => x"c6",
          5245 => x"f0",
          5246 => x"86",
          5247 => x"12",
          5248 => x"2b",
          5249 => x"07",
          5250 => x"55",
          5251 => x"17",
          5252 => x"ff",
          5253 => x"2a",
          5254 => x"54",
          5255 => x"34",
          5256 => x"06",
          5257 => x"15",
          5258 => x"f0",
          5259 => x"2b",
          5260 => x"1e",
          5261 => x"87",
          5262 => x"88",
          5263 => x"88",
          5264 => x"5e",
          5265 => x"54",
          5266 => x"34",
          5267 => x"34",
          5268 => x"08",
          5269 => x"11",
          5270 => x"33",
          5271 => x"71",
          5272 => x"53",
          5273 => x"74",
          5274 => x"86",
          5275 => x"87",
          5276 => x"d4",
          5277 => x"16",
          5278 => x"11",
          5279 => x"33",
          5280 => x"07",
          5281 => x"53",
          5282 => x"56",
          5283 => x"16",
          5284 => x"16",
          5285 => x"f0",
          5286 => x"05",
          5287 => x"d4",
          5288 => x"3d",
          5289 => x"3d",
          5290 => x"82",
          5291 => x"84",
          5292 => x"3f",
          5293 => x"80",
          5294 => x"71",
          5295 => x"3f",
          5296 => x"08",
          5297 => x"d4",
          5298 => x"3d",
          5299 => x"3d",
          5300 => x"40",
          5301 => x"42",
          5302 => x"f0",
          5303 => x"09",
          5304 => x"38",
          5305 => x"7b",
          5306 => x"51",
          5307 => x"82",
          5308 => x"54",
          5309 => x"7e",
          5310 => x"51",
          5311 => x"7e",
          5312 => x"39",
          5313 => x"8f",
          5314 => x"f8",
          5315 => x"ff",
          5316 => x"f0",
          5317 => x"31",
          5318 => x"83",
          5319 => x"70",
          5320 => x"11",
          5321 => x"12",
          5322 => x"2b",
          5323 => x"31",
          5324 => x"ff",
          5325 => x"29",
          5326 => x"88",
          5327 => x"33",
          5328 => x"71",
          5329 => x"70",
          5330 => x"44",
          5331 => x"41",
          5332 => x"5b",
          5333 => x"5b",
          5334 => x"25",
          5335 => x"81",
          5336 => x"75",
          5337 => x"ff",
          5338 => x"54",
          5339 => x"83",
          5340 => x"88",
          5341 => x"88",
          5342 => x"33",
          5343 => x"71",
          5344 => x"90",
          5345 => x"47",
          5346 => x"54",
          5347 => x"8b",
          5348 => x"31",
          5349 => x"ff",
          5350 => x"77",
          5351 => x"fe",
          5352 => x"54",
          5353 => x"09",
          5354 => x"38",
          5355 => x"c0",
          5356 => x"ff",
          5357 => x"81",
          5358 => x"8e",
          5359 => x"24",
          5360 => x"51",
          5361 => x"81",
          5362 => x"18",
          5363 => x"24",
          5364 => x"79",
          5365 => x"33",
          5366 => x"71",
          5367 => x"53",
          5368 => x"f4",
          5369 => x"78",
          5370 => x"3f",
          5371 => x"08",
          5372 => x"06",
          5373 => x"53",
          5374 => x"82",
          5375 => x"11",
          5376 => x"55",
          5377 => x"93",
          5378 => x"f0",
          5379 => x"05",
          5380 => x"ff",
          5381 => x"81",
          5382 => x"15",
          5383 => x"24",
          5384 => x"78",
          5385 => x"3f",
          5386 => x"08",
          5387 => x"33",
          5388 => x"71",
          5389 => x"53",
          5390 => x"9c",
          5391 => x"78",
          5392 => x"3f",
          5393 => x"08",
          5394 => x"06",
          5395 => x"53",
          5396 => x"82",
          5397 => x"11",
          5398 => x"55",
          5399 => x"bb",
          5400 => x"f0",
          5401 => x"05",
          5402 => x"19",
          5403 => x"83",
          5404 => x"58",
          5405 => x"7f",
          5406 => x"b0",
          5407 => x"f8",
          5408 => x"d4",
          5409 => x"2e",
          5410 => x"53",
          5411 => x"d4",
          5412 => x"ff",
          5413 => x"73",
          5414 => x"3f",
          5415 => x"78",
          5416 => x"80",
          5417 => x"78",
          5418 => x"3f",
          5419 => x"2b",
          5420 => x"08",
          5421 => x"51",
          5422 => x"7b",
          5423 => x"d4",
          5424 => x"3d",
          5425 => x"3d",
          5426 => x"29",
          5427 => x"fb",
          5428 => x"d4",
          5429 => x"82",
          5430 => x"80",
          5431 => x"73",
          5432 => x"82",
          5433 => x"51",
          5434 => x"3f",
          5435 => x"f8",
          5436 => x"0d",
          5437 => x"0d",
          5438 => x"33",
          5439 => x"70",
          5440 => x"38",
          5441 => x"11",
          5442 => x"82",
          5443 => x"83",
          5444 => x"fc",
          5445 => x"9b",
          5446 => x"84",
          5447 => x"33",
          5448 => x"51",
          5449 => x"80",
          5450 => x"84",
          5451 => x"92",
          5452 => x"51",
          5453 => x"80",
          5454 => x"81",
          5455 => x"72",
          5456 => x"92",
          5457 => x"81",
          5458 => x"0b",
          5459 => x"8c",
          5460 => x"71",
          5461 => x"06",
          5462 => x"80",
          5463 => x"87",
          5464 => x"08",
          5465 => x"38",
          5466 => x"80",
          5467 => x"71",
          5468 => x"c0",
          5469 => x"51",
          5470 => x"87",
          5471 => x"d4",
          5472 => x"82",
          5473 => x"33",
          5474 => x"d4",
          5475 => x"3d",
          5476 => x"3d",
          5477 => x"64",
          5478 => x"bf",
          5479 => x"40",
          5480 => x"74",
          5481 => x"cd",
          5482 => x"f8",
          5483 => x"7a",
          5484 => x"81",
          5485 => x"72",
          5486 => x"87",
          5487 => x"11",
          5488 => x"8c",
          5489 => x"92",
          5490 => x"5a",
          5491 => x"58",
          5492 => x"c0",
          5493 => x"76",
          5494 => x"76",
          5495 => x"70",
          5496 => x"81",
          5497 => x"54",
          5498 => x"8e",
          5499 => x"52",
          5500 => x"81",
          5501 => x"81",
          5502 => x"74",
          5503 => x"53",
          5504 => x"83",
          5505 => x"78",
          5506 => x"8f",
          5507 => x"2e",
          5508 => x"c0",
          5509 => x"52",
          5510 => x"87",
          5511 => x"08",
          5512 => x"2e",
          5513 => x"84",
          5514 => x"38",
          5515 => x"87",
          5516 => x"15",
          5517 => x"70",
          5518 => x"52",
          5519 => x"ff",
          5520 => x"39",
          5521 => x"81",
          5522 => x"ff",
          5523 => x"57",
          5524 => x"90",
          5525 => x"80",
          5526 => x"71",
          5527 => x"78",
          5528 => x"38",
          5529 => x"80",
          5530 => x"80",
          5531 => x"81",
          5532 => x"72",
          5533 => x"0c",
          5534 => x"04",
          5535 => x"60",
          5536 => x"8c",
          5537 => x"33",
          5538 => x"5b",
          5539 => x"74",
          5540 => x"e1",
          5541 => x"f8",
          5542 => x"79",
          5543 => x"78",
          5544 => x"06",
          5545 => x"77",
          5546 => x"87",
          5547 => x"11",
          5548 => x"8c",
          5549 => x"92",
          5550 => x"59",
          5551 => x"85",
          5552 => x"98",
          5553 => x"7d",
          5554 => x"0c",
          5555 => x"08",
          5556 => x"70",
          5557 => x"53",
          5558 => x"2e",
          5559 => x"70",
          5560 => x"33",
          5561 => x"18",
          5562 => x"2a",
          5563 => x"51",
          5564 => x"2e",
          5565 => x"c0",
          5566 => x"52",
          5567 => x"87",
          5568 => x"08",
          5569 => x"2e",
          5570 => x"84",
          5571 => x"38",
          5572 => x"87",
          5573 => x"15",
          5574 => x"70",
          5575 => x"52",
          5576 => x"ff",
          5577 => x"39",
          5578 => x"81",
          5579 => x"80",
          5580 => x"52",
          5581 => x"90",
          5582 => x"80",
          5583 => x"71",
          5584 => x"7a",
          5585 => x"38",
          5586 => x"80",
          5587 => x"80",
          5588 => x"81",
          5589 => x"72",
          5590 => x"0c",
          5591 => x"04",
          5592 => x"7a",
          5593 => x"a3",
          5594 => x"88",
          5595 => x"33",
          5596 => x"56",
          5597 => x"3f",
          5598 => x"08",
          5599 => x"83",
          5600 => x"fe",
          5601 => x"87",
          5602 => x"0c",
          5603 => x"76",
          5604 => x"38",
          5605 => x"93",
          5606 => x"2b",
          5607 => x"8c",
          5608 => x"71",
          5609 => x"38",
          5610 => x"71",
          5611 => x"c6",
          5612 => x"39",
          5613 => x"81",
          5614 => x"06",
          5615 => x"71",
          5616 => x"38",
          5617 => x"8c",
          5618 => x"e8",
          5619 => x"98",
          5620 => x"71",
          5621 => x"73",
          5622 => x"92",
          5623 => x"72",
          5624 => x"06",
          5625 => x"f7",
          5626 => x"80",
          5627 => x"88",
          5628 => x"0c",
          5629 => x"80",
          5630 => x"56",
          5631 => x"56",
          5632 => x"82",
          5633 => x"88",
          5634 => x"fe",
          5635 => x"81",
          5636 => x"33",
          5637 => x"07",
          5638 => x"0c",
          5639 => x"3d",
          5640 => x"3d",
          5641 => x"11",
          5642 => x"33",
          5643 => x"71",
          5644 => x"81",
          5645 => x"72",
          5646 => x"75",
          5647 => x"82",
          5648 => x"52",
          5649 => x"54",
          5650 => x"0d",
          5651 => x"0d",
          5652 => x"05",
          5653 => x"52",
          5654 => x"70",
          5655 => x"34",
          5656 => x"51",
          5657 => x"83",
          5658 => x"ff",
          5659 => x"75",
          5660 => x"72",
          5661 => x"54",
          5662 => x"2a",
          5663 => x"70",
          5664 => x"34",
          5665 => x"51",
          5666 => x"81",
          5667 => x"70",
          5668 => x"70",
          5669 => x"3d",
          5670 => x"3d",
          5671 => x"77",
          5672 => x"70",
          5673 => x"38",
          5674 => x"05",
          5675 => x"70",
          5676 => x"34",
          5677 => x"eb",
          5678 => x"0d",
          5679 => x"0d",
          5680 => x"54",
          5681 => x"72",
          5682 => x"54",
          5683 => x"51",
          5684 => x"84",
          5685 => x"fc",
          5686 => x"77",
          5687 => x"53",
          5688 => x"05",
          5689 => x"70",
          5690 => x"33",
          5691 => x"ff",
          5692 => x"52",
          5693 => x"2e",
          5694 => x"80",
          5695 => x"71",
          5696 => x"0c",
          5697 => x"04",
          5698 => x"74",
          5699 => x"89",
          5700 => x"2e",
          5701 => x"11",
          5702 => x"52",
          5703 => x"70",
          5704 => x"f8",
          5705 => x"0d",
          5706 => x"82",
          5707 => x"04",
          5708 => x"77",
          5709 => x"70",
          5710 => x"33",
          5711 => x"55",
          5712 => x"ff",
          5713 => x"f8",
          5714 => x"72",
          5715 => x"38",
          5716 => x"72",
          5717 => x"b6",
          5718 => x"f8",
          5719 => x"ff",
          5720 => x"80",
          5721 => x"73",
          5722 => x"55",
          5723 => x"f8",
          5724 => x"0d",
          5725 => x"0d",
          5726 => x"0b",
          5727 => x"56",
          5728 => x"2e",
          5729 => x"81",
          5730 => x"08",
          5731 => x"70",
          5732 => x"33",
          5733 => x"e4",
          5734 => x"f8",
          5735 => x"09",
          5736 => x"38",
          5737 => x"08",
          5738 => x"b4",
          5739 => x"a8",
          5740 => x"a0",
          5741 => x"56",
          5742 => x"27",
          5743 => x"16",
          5744 => x"82",
          5745 => x"06",
          5746 => x"54",
          5747 => x"78",
          5748 => x"33",
          5749 => x"3f",
          5750 => x"5a",
          5751 => x"f8",
          5752 => x"0d",
          5753 => x"0d",
          5754 => x"56",
          5755 => x"b4",
          5756 => x"af",
          5757 => x"fe",
          5758 => x"d4",
          5759 => x"82",
          5760 => x"9f",
          5761 => x"74",
          5762 => x"52",
          5763 => x"51",
          5764 => x"82",
          5765 => x"80",
          5766 => x"ff",
          5767 => x"74",
          5768 => x"76",
          5769 => x"0c",
          5770 => x"04",
          5771 => x"7a",
          5772 => x"fe",
          5773 => x"d4",
          5774 => x"82",
          5775 => x"81",
          5776 => x"33",
          5777 => x"2e",
          5778 => x"80",
          5779 => x"17",
          5780 => x"81",
          5781 => x"06",
          5782 => x"84",
          5783 => x"d4",
          5784 => x"b8",
          5785 => x"56",
          5786 => x"82",
          5787 => x"84",
          5788 => x"fb",
          5789 => x"8b",
          5790 => x"52",
          5791 => x"eb",
          5792 => x"85",
          5793 => x"84",
          5794 => x"fb",
          5795 => x"17",
          5796 => x"a0",
          5797 => x"d3",
          5798 => x"08",
          5799 => x"17",
          5800 => x"3f",
          5801 => x"81",
          5802 => x"19",
          5803 => x"53",
          5804 => x"17",
          5805 => x"c4",
          5806 => x"18",
          5807 => x"80",
          5808 => x"33",
          5809 => x"3f",
          5810 => x"08",
          5811 => x"38",
          5812 => x"82",
          5813 => x"8a",
          5814 => x"fb",
          5815 => x"fe",
          5816 => x"08",
          5817 => x"56",
          5818 => x"74",
          5819 => x"38",
          5820 => x"75",
          5821 => x"16",
          5822 => x"53",
          5823 => x"f8",
          5824 => x"0d",
          5825 => x"0d",
          5826 => x"08",
          5827 => x"81",
          5828 => x"df",
          5829 => x"15",
          5830 => x"d7",
          5831 => x"33",
          5832 => x"82",
          5833 => x"38",
          5834 => x"89",
          5835 => x"2e",
          5836 => x"bf",
          5837 => x"2e",
          5838 => x"81",
          5839 => x"81",
          5840 => x"89",
          5841 => x"08",
          5842 => x"52",
          5843 => x"3f",
          5844 => x"08",
          5845 => x"74",
          5846 => x"14",
          5847 => x"81",
          5848 => x"2a",
          5849 => x"05",
          5850 => x"57",
          5851 => x"f5",
          5852 => x"f8",
          5853 => x"38",
          5854 => x"06",
          5855 => x"33",
          5856 => x"78",
          5857 => x"06",
          5858 => x"5c",
          5859 => x"53",
          5860 => x"38",
          5861 => x"06",
          5862 => x"39",
          5863 => x"a8",
          5864 => x"52",
          5865 => x"bd",
          5866 => x"f8",
          5867 => x"38",
          5868 => x"fe",
          5869 => x"b8",
          5870 => x"cf",
          5871 => x"f8",
          5872 => x"ff",
          5873 => x"39",
          5874 => x"a8",
          5875 => x"52",
          5876 => x"91",
          5877 => x"f8",
          5878 => x"76",
          5879 => x"fc",
          5880 => x"b8",
          5881 => x"ba",
          5882 => x"f8",
          5883 => x"06",
          5884 => x"81",
          5885 => x"d4",
          5886 => x"3d",
          5887 => x"3d",
          5888 => x"7e",
          5889 => x"82",
          5890 => x"27",
          5891 => x"76",
          5892 => x"27",
          5893 => x"75",
          5894 => x"79",
          5895 => x"38",
          5896 => x"89",
          5897 => x"2e",
          5898 => x"80",
          5899 => x"2e",
          5900 => x"81",
          5901 => x"81",
          5902 => x"89",
          5903 => x"08",
          5904 => x"52",
          5905 => x"3f",
          5906 => x"08",
          5907 => x"f8",
          5908 => x"38",
          5909 => x"06",
          5910 => x"81",
          5911 => x"06",
          5912 => x"77",
          5913 => x"2e",
          5914 => x"84",
          5915 => x"06",
          5916 => x"06",
          5917 => x"53",
          5918 => x"81",
          5919 => x"34",
          5920 => x"a8",
          5921 => x"52",
          5922 => x"d9",
          5923 => x"f8",
          5924 => x"d4",
          5925 => x"94",
          5926 => x"ff",
          5927 => x"05",
          5928 => x"54",
          5929 => x"38",
          5930 => x"74",
          5931 => x"06",
          5932 => x"07",
          5933 => x"74",
          5934 => x"39",
          5935 => x"a8",
          5936 => x"52",
          5937 => x"9d",
          5938 => x"f8",
          5939 => x"d4",
          5940 => x"d8",
          5941 => x"ff",
          5942 => x"76",
          5943 => x"06",
          5944 => x"05",
          5945 => x"3f",
          5946 => x"87",
          5947 => x"08",
          5948 => x"51",
          5949 => x"82",
          5950 => x"59",
          5951 => x"08",
          5952 => x"f0",
          5953 => x"82",
          5954 => x"06",
          5955 => x"05",
          5956 => x"54",
          5957 => x"3f",
          5958 => x"08",
          5959 => x"74",
          5960 => x"51",
          5961 => x"81",
          5962 => x"34",
          5963 => x"f8",
          5964 => x"0d",
          5965 => x"0d",
          5966 => x"72",
          5967 => x"56",
          5968 => x"27",
          5969 => x"9c",
          5970 => x"9d",
          5971 => x"2e",
          5972 => x"53",
          5973 => x"51",
          5974 => x"82",
          5975 => x"54",
          5976 => x"08",
          5977 => x"93",
          5978 => x"80",
          5979 => x"54",
          5980 => x"82",
          5981 => x"54",
          5982 => x"74",
          5983 => x"fb",
          5984 => x"d4",
          5985 => x"82",
          5986 => x"80",
          5987 => x"38",
          5988 => x"08",
          5989 => x"38",
          5990 => x"08",
          5991 => x"38",
          5992 => x"52",
          5993 => x"d6",
          5994 => x"f8",
          5995 => x"9c",
          5996 => x"11",
          5997 => x"57",
          5998 => x"74",
          5999 => x"81",
          6000 => x"0c",
          6001 => x"81",
          6002 => x"84",
          6003 => x"55",
          6004 => x"ff",
          6005 => x"54",
          6006 => x"f8",
          6007 => x"0d",
          6008 => x"0d",
          6009 => x"08",
          6010 => x"79",
          6011 => x"17",
          6012 => x"80",
          6013 => x"9c",
          6014 => x"26",
          6015 => x"58",
          6016 => x"52",
          6017 => x"fd",
          6018 => x"74",
          6019 => x"08",
          6020 => x"38",
          6021 => x"08",
          6022 => x"f8",
          6023 => x"82",
          6024 => x"17",
          6025 => x"f8",
          6026 => x"c7",
          6027 => x"94",
          6028 => x"56",
          6029 => x"2e",
          6030 => x"77",
          6031 => x"81",
          6032 => x"38",
          6033 => x"9c",
          6034 => x"26",
          6035 => x"56",
          6036 => x"51",
          6037 => x"80",
          6038 => x"f8",
          6039 => x"09",
          6040 => x"38",
          6041 => x"08",
          6042 => x"f8",
          6043 => x"30",
          6044 => x"80",
          6045 => x"07",
          6046 => x"08",
          6047 => x"55",
          6048 => x"ef",
          6049 => x"f8",
          6050 => x"95",
          6051 => x"08",
          6052 => x"27",
          6053 => x"9c",
          6054 => x"89",
          6055 => x"85",
          6056 => x"db",
          6057 => x"81",
          6058 => x"17",
          6059 => x"89",
          6060 => x"75",
          6061 => x"ac",
          6062 => x"7a",
          6063 => x"3f",
          6064 => x"08",
          6065 => x"38",
          6066 => x"d4",
          6067 => x"2e",
          6068 => x"86",
          6069 => x"f8",
          6070 => x"d4",
          6071 => x"70",
          6072 => x"07",
          6073 => x"7c",
          6074 => x"55",
          6075 => x"f8",
          6076 => x"2e",
          6077 => x"ff",
          6078 => x"55",
          6079 => x"ff",
          6080 => x"76",
          6081 => x"3f",
          6082 => x"08",
          6083 => x"08",
          6084 => x"d4",
          6085 => x"80",
          6086 => x"55",
          6087 => x"94",
          6088 => x"2e",
          6089 => x"53",
          6090 => x"51",
          6091 => x"82",
          6092 => x"55",
          6093 => x"75",
          6094 => x"9c",
          6095 => x"05",
          6096 => x"56",
          6097 => x"26",
          6098 => x"15",
          6099 => x"84",
          6100 => x"07",
          6101 => x"18",
          6102 => x"ff",
          6103 => x"2e",
          6104 => x"39",
          6105 => x"39",
          6106 => x"08",
          6107 => x"81",
          6108 => x"74",
          6109 => x"0c",
          6110 => x"04",
          6111 => x"7a",
          6112 => x"f3",
          6113 => x"d4",
          6114 => x"81",
          6115 => x"f8",
          6116 => x"38",
          6117 => x"51",
          6118 => x"82",
          6119 => x"82",
          6120 => x"b4",
          6121 => x"84",
          6122 => x"52",
          6123 => x"52",
          6124 => x"3f",
          6125 => x"39",
          6126 => x"8a",
          6127 => x"75",
          6128 => x"38",
          6129 => x"19",
          6130 => x"81",
          6131 => x"ed",
          6132 => x"d4",
          6133 => x"2e",
          6134 => x"15",
          6135 => x"70",
          6136 => x"07",
          6137 => x"53",
          6138 => x"75",
          6139 => x"0c",
          6140 => x"04",
          6141 => x"7a",
          6142 => x"58",
          6143 => x"f0",
          6144 => x"80",
          6145 => x"9f",
          6146 => x"80",
          6147 => x"90",
          6148 => x"17",
          6149 => x"aa",
          6150 => x"53",
          6151 => x"88",
          6152 => x"08",
          6153 => x"38",
          6154 => x"53",
          6155 => x"17",
          6156 => x"72",
          6157 => x"fe",
          6158 => x"08",
          6159 => x"80",
          6160 => x"16",
          6161 => x"2b",
          6162 => x"75",
          6163 => x"73",
          6164 => x"f5",
          6165 => x"d4",
          6166 => x"82",
          6167 => x"ff",
          6168 => x"81",
          6169 => x"f8",
          6170 => x"38",
          6171 => x"82",
          6172 => x"26",
          6173 => x"58",
          6174 => x"73",
          6175 => x"39",
          6176 => x"51",
          6177 => x"82",
          6178 => x"98",
          6179 => x"94",
          6180 => x"17",
          6181 => x"58",
          6182 => x"9a",
          6183 => x"81",
          6184 => x"74",
          6185 => x"98",
          6186 => x"83",
          6187 => x"b8",
          6188 => x"0c",
          6189 => x"82",
          6190 => x"8a",
          6191 => x"f8",
          6192 => x"70",
          6193 => x"08",
          6194 => x"57",
          6195 => x"0a",
          6196 => x"38",
          6197 => x"15",
          6198 => x"08",
          6199 => x"72",
          6200 => x"cb",
          6201 => x"ff",
          6202 => x"81",
          6203 => x"13",
          6204 => x"94",
          6205 => x"74",
          6206 => x"85",
          6207 => x"22",
          6208 => x"73",
          6209 => x"38",
          6210 => x"8a",
          6211 => x"05",
          6212 => x"06",
          6213 => x"8a",
          6214 => x"73",
          6215 => x"3f",
          6216 => x"08",
          6217 => x"81",
          6218 => x"f8",
          6219 => x"ff",
          6220 => x"82",
          6221 => x"ff",
          6222 => x"38",
          6223 => x"82",
          6224 => x"26",
          6225 => x"7b",
          6226 => x"98",
          6227 => x"55",
          6228 => x"94",
          6229 => x"73",
          6230 => x"3f",
          6231 => x"08",
          6232 => x"82",
          6233 => x"80",
          6234 => x"38",
          6235 => x"d4",
          6236 => x"2e",
          6237 => x"55",
          6238 => x"08",
          6239 => x"38",
          6240 => x"08",
          6241 => x"fb",
          6242 => x"d4",
          6243 => x"38",
          6244 => x"0c",
          6245 => x"51",
          6246 => x"82",
          6247 => x"98",
          6248 => x"90",
          6249 => x"16",
          6250 => x"15",
          6251 => x"74",
          6252 => x"0c",
          6253 => x"04",
          6254 => x"7b",
          6255 => x"5b",
          6256 => x"52",
          6257 => x"ac",
          6258 => x"f8",
          6259 => x"d4",
          6260 => x"ec",
          6261 => x"f8",
          6262 => x"17",
          6263 => x"51",
          6264 => x"82",
          6265 => x"54",
          6266 => x"08",
          6267 => x"82",
          6268 => x"9c",
          6269 => x"33",
          6270 => x"72",
          6271 => x"09",
          6272 => x"38",
          6273 => x"d4",
          6274 => x"72",
          6275 => x"55",
          6276 => x"53",
          6277 => x"8e",
          6278 => x"56",
          6279 => x"09",
          6280 => x"38",
          6281 => x"d4",
          6282 => x"81",
          6283 => x"fd",
          6284 => x"d4",
          6285 => x"82",
          6286 => x"80",
          6287 => x"38",
          6288 => x"09",
          6289 => x"38",
          6290 => x"82",
          6291 => x"8b",
          6292 => x"fd",
          6293 => x"9a",
          6294 => x"eb",
          6295 => x"d4",
          6296 => x"ff",
          6297 => x"70",
          6298 => x"53",
          6299 => x"09",
          6300 => x"38",
          6301 => x"eb",
          6302 => x"d4",
          6303 => x"2b",
          6304 => x"72",
          6305 => x"0c",
          6306 => x"04",
          6307 => x"77",
          6308 => x"ff",
          6309 => x"9a",
          6310 => x"55",
          6311 => x"76",
          6312 => x"53",
          6313 => x"09",
          6314 => x"38",
          6315 => x"52",
          6316 => x"eb",
          6317 => x"3d",
          6318 => x"3d",
          6319 => x"80",
          6320 => x"70",
          6321 => x"81",
          6322 => x"74",
          6323 => x"56",
          6324 => x"70",
          6325 => x"ff",
          6326 => x"51",
          6327 => x"38",
          6328 => x"f8",
          6329 => x"0d",
          6330 => x"0d",
          6331 => x"59",
          6332 => x"5f",
          6333 => x"70",
          6334 => x"19",
          6335 => x"83",
          6336 => x"19",
          6337 => x"51",
          6338 => x"82",
          6339 => x"5b",
          6340 => x"08",
          6341 => x"9c",
          6342 => x"33",
          6343 => x"86",
          6344 => x"82",
          6345 => x"15",
          6346 => x"70",
          6347 => x"58",
          6348 => x"1a",
          6349 => x"f8",
          6350 => x"81",
          6351 => x"81",
          6352 => x"81",
          6353 => x"f8",
          6354 => x"ae",
          6355 => x"06",
          6356 => x"53",
          6357 => x"53",
          6358 => x"82",
          6359 => x"77",
          6360 => x"56",
          6361 => x"09",
          6362 => x"38",
          6363 => x"7f",
          6364 => x"81",
          6365 => x"ef",
          6366 => x"2e",
          6367 => x"81",
          6368 => x"86",
          6369 => x"06",
          6370 => x"80",
          6371 => x"8d",
          6372 => x"81",
          6373 => x"90",
          6374 => x"1d",
          6375 => x"5d",
          6376 => x"09",
          6377 => x"9c",
          6378 => x"33",
          6379 => x"2e",
          6380 => x"81",
          6381 => x"1e",
          6382 => x"52",
          6383 => x"3f",
          6384 => x"08",
          6385 => x"06",
          6386 => x"f8",
          6387 => x"70",
          6388 => x"8d",
          6389 => x"51",
          6390 => x"58",
          6391 => x"80",
          6392 => x"05",
          6393 => x"3f",
          6394 => x"08",
          6395 => x"06",
          6396 => x"2e",
          6397 => x"81",
          6398 => x"c8",
          6399 => x"1a",
          6400 => x"75",
          6401 => x"14",
          6402 => x"75",
          6403 => x"2e",
          6404 => x"b0",
          6405 => x"57",
          6406 => x"c1",
          6407 => x"70",
          6408 => x"81",
          6409 => x"55",
          6410 => x"8e",
          6411 => x"fe",
          6412 => x"73",
          6413 => x"80",
          6414 => x"1c",
          6415 => x"06",
          6416 => x"39",
          6417 => x"72",
          6418 => x"7b",
          6419 => x"51",
          6420 => x"82",
          6421 => x"81",
          6422 => x"72",
          6423 => x"38",
          6424 => x"1a",
          6425 => x"80",
          6426 => x"f8",
          6427 => x"d4",
          6428 => x"82",
          6429 => x"89",
          6430 => x"08",
          6431 => x"86",
          6432 => x"98",
          6433 => x"82",
          6434 => x"90",
          6435 => x"f2",
          6436 => x"70",
          6437 => x"80",
          6438 => x"f6",
          6439 => x"d4",
          6440 => x"82",
          6441 => x"83",
          6442 => x"ff",
          6443 => x"ff",
          6444 => x"0c",
          6445 => x"52",
          6446 => x"a9",
          6447 => x"f8",
          6448 => x"d4",
          6449 => x"85",
          6450 => x"08",
          6451 => x"57",
          6452 => x"84",
          6453 => x"39",
          6454 => x"bf",
          6455 => x"ff",
          6456 => x"73",
          6457 => x"75",
          6458 => x"82",
          6459 => x"83",
          6460 => x"06",
          6461 => x"8f",
          6462 => x"73",
          6463 => x"74",
          6464 => x"81",
          6465 => x"38",
          6466 => x"70",
          6467 => x"81",
          6468 => x"55",
          6469 => x"38",
          6470 => x"70",
          6471 => x"54",
          6472 => x"92",
          6473 => x"33",
          6474 => x"06",
          6475 => x"08",
          6476 => x"58",
          6477 => x"7c",
          6478 => x"06",
          6479 => x"8d",
          6480 => x"7d",
          6481 => x"81",
          6482 => x"38",
          6483 => x"9a",
          6484 => x"e5",
          6485 => x"d4",
          6486 => x"ff",
          6487 => x"74",
          6488 => x"76",
          6489 => x"06",
          6490 => x"05",
          6491 => x"75",
          6492 => x"c7",
          6493 => x"77",
          6494 => x"8f",
          6495 => x"f8",
          6496 => x"ff",
          6497 => x"80",
          6498 => x"77",
          6499 => x"80",
          6500 => x"51",
          6501 => x"3f",
          6502 => x"08",
          6503 => x"70",
          6504 => x"81",
          6505 => x"80",
          6506 => x"74",
          6507 => x"08",
          6508 => x"06",
          6509 => x"75",
          6510 => x"75",
          6511 => x"2e",
          6512 => x"b3",
          6513 => x"5b",
          6514 => x"ff",
          6515 => x"33",
          6516 => x"70",
          6517 => x"55",
          6518 => x"2e",
          6519 => x"80",
          6520 => x"77",
          6521 => x"22",
          6522 => x"8b",
          6523 => x"70",
          6524 => x"51",
          6525 => x"81",
          6526 => x"5c",
          6527 => x"93",
          6528 => x"f9",
          6529 => x"d4",
          6530 => x"ff",
          6531 => x"7e",
          6532 => x"ab",
          6533 => x"06",
          6534 => x"38",
          6535 => x"19",
          6536 => x"08",
          6537 => x"3f",
          6538 => x"08",
          6539 => x"38",
          6540 => x"ff",
          6541 => x"0c",
          6542 => x"51",
          6543 => x"82",
          6544 => x"58",
          6545 => x"08",
          6546 => x"e8",
          6547 => x"d4",
          6548 => x"3d",
          6549 => x"3d",
          6550 => x"08",
          6551 => x"81",
          6552 => x"5d",
          6553 => x"73",
          6554 => x"73",
          6555 => x"70",
          6556 => x"5d",
          6557 => x"8d",
          6558 => x"70",
          6559 => x"22",
          6560 => x"f0",
          6561 => x"a0",
          6562 => x"92",
          6563 => x"5f",
          6564 => x"3f",
          6565 => x"05",
          6566 => x"54",
          6567 => x"82",
          6568 => x"c0",
          6569 => x"34",
          6570 => x"1c",
          6571 => x"58",
          6572 => x"52",
          6573 => x"e2",
          6574 => x"27",
          6575 => x"7a",
          6576 => x"70",
          6577 => x"06",
          6578 => x"80",
          6579 => x"74",
          6580 => x"06",
          6581 => x"55",
          6582 => x"81",
          6583 => x"07",
          6584 => x"71",
          6585 => x"81",
          6586 => x"56",
          6587 => x"2e",
          6588 => x"84",
          6589 => x"56",
          6590 => x"76",
          6591 => x"38",
          6592 => x"55",
          6593 => x"05",
          6594 => x"57",
          6595 => x"bf",
          6596 => x"74",
          6597 => x"87",
          6598 => x"76",
          6599 => x"ff",
          6600 => x"2a",
          6601 => x"74",
          6602 => x"3d",
          6603 => x"54",
          6604 => x"34",
          6605 => x"b5",
          6606 => x"54",
          6607 => x"ad",
          6608 => x"70",
          6609 => x"e3",
          6610 => x"d4",
          6611 => x"2e",
          6612 => x"17",
          6613 => x"2e",
          6614 => x"15",
          6615 => x"55",
          6616 => x"89",
          6617 => x"70",
          6618 => x"d0",
          6619 => x"77",
          6620 => x"54",
          6621 => x"16",
          6622 => x"56",
          6623 => x"8a",
          6624 => x"81",
          6625 => x"58",
          6626 => x"78",
          6627 => x"27",
          6628 => x"51",
          6629 => x"82",
          6630 => x"8b",
          6631 => x"5b",
          6632 => x"27",
          6633 => x"87",
          6634 => x"e4",
          6635 => x"38",
          6636 => x"08",
          6637 => x"f8",
          6638 => x"09",
          6639 => x"df",
          6640 => x"cb",
          6641 => x"1b",
          6642 => x"cb",
          6643 => x"81",
          6644 => x"06",
          6645 => x"81",
          6646 => x"2e",
          6647 => x"52",
          6648 => x"fe",
          6649 => x"82",
          6650 => x"19",
          6651 => x"79",
          6652 => x"3f",
          6653 => x"08",
          6654 => x"f8",
          6655 => x"38",
          6656 => x"78",
          6657 => x"d4",
          6658 => x"2b",
          6659 => x"71",
          6660 => x"79",
          6661 => x"3f",
          6662 => x"08",
          6663 => x"f8",
          6664 => x"38",
          6665 => x"f5",
          6666 => x"d4",
          6667 => x"ff",
          6668 => x"1a",
          6669 => x"51",
          6670 => x"82",
          6671 => x"57",
          6672 => x"08",
          6673 => x"8c",
          6674 => x"1b",
          6675 => x"ff",
          6676 => x"5b",
          6677 => x"34",
          6678 => x"17",
          6679 => x"f8",
          6680 => x"34",
          6681 => x"08",
          6682 => x"51",
          6683 => x"77",
          6684 => x"05",
          6685 => x"73",
          6686 => x"2e",
          6687 => x"10",
          6688 => x"81",
          6689 => x"54",
          6690 => x"c7",
          6691 => x"76",
          6692 => x"b9",
          6693 => x"38",
          6694 => x"54",
          6695 => x"8c",
          6696 => x"38",
          6697 => x"ff",
          6698 => x"74",
          6699 => x"22",
          6700 => x"86",
          6701 => x"c0",
          6702 => x"76",
          6703 => x"83",
          6704 => x"52",
          6705 => x"f7",
          6706 => x"f8",
          6707 => x"d4",
          6708 => x"c9",
          6709 => x"59",
          6710 => x"38",
          6711 => x"52",
          6712 => x"81",
          6713 => x"f8",
          6714 => x"d4",
          6715 => x"38",
          6716 => x"d4",
          6717 => x"9c",
          6718 => x"df",
          6719 => x"53",
          6720 => x"9c",
          6721 => x"df",
          6722 => x"1a",
          6723 => x"33",
          6724 => x"55",
          6725 => x"34",
          6726 => x"1d",
          6727 => x"74",
          6728 => x"0c",
          6729 => x"04",
          6730 => x"78",
          6731 => x"12",
          6732 => x"08",
          6733 => x"55",
          6734 => x"94",
          6735 => x"74",
          6736 => x"3f",
          6737 => x"08",
          6738 => x"f8",
          6739 => x"38",
          6740 => x"52",
          6741 => x"8d",
          6742 => x"f8",
          6743 => x"d4",
          6744 => x"38",
          6745 => x"53",
          6746 => x"81",
          6747 => x"34",
          6748 => x"77",
          6749 => x"82",
          6750 => x"52",
          6751 => x"bf",
          6752 => x"f8",
          6753 => x"d4",
          6754 => x"2e",
          6755 => x"84",
          6756 => x"06",
          6757 => x"54",
          6758 => x"f8",
          6759 => x"0d",
          6760 => x"0d",
          6761 => x"08",
          6762 => x"80",
          6763 => x"34",
          6764 => x"80",
          6765 => x"38",
          6766 => x"ff",
          6767 => x"38",
          6768 => x"7f",
          6769 => x"70",
          6770 => x"5b",
          6771 => x"77",
          6772 => x"38",
          6773 => x"70",
          6774 => x"5b",
          6775 => x"97",
          6776 => x"80",
          6777 => x"ff",
          6778 => x"53",
          6779 => x"26",
          6780 => x"5b",
          6781 => x"76",
          6782 => x"81",
          6783 => x"58",
          6784 => x"b5",
          6785 => x"2b",
          6786 => x"80",
          6787 => x"82",
          6788 => x"83",
          6789 => x"55",
          6790 => x"27",
          6791 => x"76",
          6792 => x"74",
          6793 => x"72",
          6794 => x"97",
          6795 => x"55",
          6796 => x"30",
          6797 => x"78",
          6798 => x"72",
          6799 => x"52",
          6800 => x"80",
          6801 => x"80",
          6802 => x"74",
          6803 => x"55",
          6804 => x"80",
          6805 => x"08",
          6806 => x"70",
          6807 => x"54",
          6808 => x"38",
          6809 => x"80",
          6810 => x"79",
          6811 => x"53",
          6812 => x"05",
          6813 => x"82",
          6814 => x"70",
          6815 => x"5a",
          6816 => x"08",
          6817 => x"81",
          6818 => x"53",
          6819 => x"b7",
          6820 => x"2e",
          6821 => x"84",
          6822 => x"55",
          6823 => x"70",
          6824 => x"07",
          6825 => x"54",
          6826 => x"26",
          6827 => x"80",
          6828 => x"ae",
          6829 => x"05",
          6830 => x"17",
          6831 => x"70",
          6832 => x"34",
          6833 => x"8a",
          6834 => x"b5",
          6835 => x"88",
          6836 => x"0b",
          6837 => x"96",
          6838 => x"72",
          6839 => x"76",
          6840 => x"0b",
          6841 => x"81",
          6842 => x"39",
          6843 => x"1a",
          6844 => x"57",
          6845 => x"80",
          6846 => x"18",
          6847 => x"56",
          6848 => x"bf",
          6849 => x"72",
          6850 => x"38",
          6851 => x"8c",
          6852 => x"53",
          6853 => x"87",
          6854 => x"2a",
          6855 => x"72",
          6856 => x"72",
          6857 => x"72",
          6858 => x"38",
          6859 => x"83",
          6860 => x"56",
          6861 => x"70",
          6862 => x"34",
          6863 => x"15",
          6864 => x"33",
          6865 => x"59",
          6866 => x"38",
          6867 => x"05",
          6868 => x"82",
          6869 => x"1c",
          6870 => x"33",
          6871 => x"85",
          6872 => x"19",
          6873 => x"08",
          6874 => x"33",
          6875 => x"9c",
          6876 => x"11",
          6877 => x"aa",
          6878 => x"f8",
          6879 => x"96",
          6880 => x"87",
          6881 => x"f8",
          6882 => x"23",
          6883 => x"d8",
          6884 => x"d4",
          6885 => x"19",
          6886 => x"0d",
          6887 => x"0d",
          6888 => x"41",
          6889 => x"70",
          6890 => x"55",
          6891 => x"83",
          6892 => x"73",
          6893 => x"92",
          6894 => x"2e",
          6895 => x"98",
          6896 => x"1f",
          6897 => x"81",
          6898 => x"64",
          6899 => x"56",
          6900 => x"2e",
          6901 => x"83",
          6902 => x"73",
          6903 => x"70",
          6904 => x"25",
          6905 => x"51",
          6906 => x"38",
          6907 => x"0c",
          6908 => x"51",
          6909 => x"26",
          6910 => x"80",
          6911 => x"34",
          6912 => x"51",
          6913 => x"82",
          6914 => x"56",
          6915 => x"63",
          6916 => x"8c",
          6917 => x"54",
          6918 => x"3d",
          6919 => x"da",
          6920 => x"d4",
          6921 => x"2e",
          6922 => x"83",
          6923 => x"82",
          6924 => x"27",
          6925 => x"10",
          6926 => x"f8",
          6927 => x"55",
          6928 => x"23",
          6929 => x"82",
          6930 => x"83",
          6931 => x"70",
          6932 => x"30",
          6933 => x"71",
          6934 => x"51",
          6935 => x"73",
          6936 => x"80",
          6937 => x"38",
          6938 => x"26",
          6939 => x"52",
          6940 => x"51",
          6941 => x"82",
          6942 => x"81",
          6943 => x"81",
          6944 => x"d7",
          6945 => x"1a",
          6946 => x"23",
          6947 => x"ff",
          6948 => x"15",
          6949 => x"70",
          6950 => x"57",
          6951 => x"09",
          6952 => x"38",
          6953 => x"80",
          6954 => x"30",
          6955 => x"79",
          6956 => x"54",
          6957 => x"74",
          6958 => x"27",
          6959 => x"78",
          6960 => x"81",
          6961 => x"79",
          6962 => x"ae",
          6963 => x"80",
          6964 => x"82",
          6965 => x"06",
          6966 => x"82",
          6967 => x"73",
          6968 => x"81",
          6969 => x"38",
          6970 => x"73",
          6971 => x"81",
          6972 => x"78",
          6973 => x"80",
          6974 => x"0b",
          6975 => x"58",
          6976 => x"78",
          6977 => x"a0",
          6978 => x"70",
          6979 => x"34",
          6980 => x"8a",
          6981 => x"38",
          6982 => x"54",
          6983 => x"34",
          6984 => x"78",
          6985 => x"38",
          6986 => x"fe",
          6987 => x"22",
          6988 => x"72",
          6989 => x"30",
          6990 => x"51",
          6991 => x"56",
          6992 => x"2e",
          6993 => x"87",
          6994 => x"59",
          6995 => x"78",
          6996 => x"55",
          6997 => x"23",
          6998 => x"86",
          6999 => x"39",
          7000 => x"57",
          7001 => x"80",
          7002 => x"83",
          7003 => x"56",
          7004 => x"a0",
          7005 => x"06",
          7006 => x"1d",
          7007 => x"70",
          7008 => x"5d",
          7009 => x"f2",
          7010 => x"38",
          7011 => x"ff",
          7012 => x"ae",
          7013 => x"06",
          7014 => x"83",
          7015 => x"80",
          7016 => x"79",
          7017 => x"70",
          7018 => x"73",
          7019 => x"38",
          7020 => x"fe",
          7021 => x"19",
          7022 => x"2e",
          7023 => x"15",
          7024 => x"55",
          7025 => x"09",
          7026 => x"38",
          7027 => x"52",
          7028 => x"d5",
          7029 => x"70",
          7030 => x"5f",
          7031 => x"70",
          7032 => x"5f",
          7033 => x"80",
          7034 => x"38",
          7035 => x"96",
          7036 => x"32",
          7037 => x"80",
          7038 => x"54",
          7039 => x"8c",
          7040 => x"2e",
          7041 => x"83",
          7042 => x"39",
          7043 => x"5b",
          7044 => x"83",
          7045 => x"7c",
          7046 => x"30",
          7047 => x"80",
          7048 => x"07",
          7049 => x"55",
          7050 => x"a6",
          7051 => x"2e",
          7052 => x"7c",
          7053 => x"38",
          7054 => x"57",
          7055 => x"81",
          7056 => x"5d",
          7057 => x"7c",
          7058 => x"fc",
          7059 => x"ff",
          7060 => x"ff",
          7061 => x"38",
          7062 => x"57",
          7063 => x"75",
          7064 => x"c2",
          7065 => x"f8",
          7066 => x"ff",
          7067 => x"2a",
          7068 => x"51",
          7069 => x"80",
          7070 => x"75",
          7071 => x"82",
          7072 => x"33",
          7073 => x"ff",
          7074 => x"38",
          7075 => x"73",
          7076 => x"38",
          7077 => x"7f",
          7078 => x"c0",
          7079 => x"a0",
          7080 => x"2a",
          7081 => x"75",
          7082 => x"58",
          7083 => x"75",
          7084 => x"38",
          7085 => x"c6",
          7086 => x"cc",
          7087 => x"f8",
          7088 => x"8a",
          7089 => x"77",
          7090 => x"56",
          7091 => x"bf",
          7092 => x"99",
          7093 => x"7b",
          7094 => x"ff",
          7095 => x"73",
          7096 => x"38",
          7097 => x"e0",
          7098 => x"ff",
          7099 => x"55",
          7100 => x"a0",
          7101 => x"74",
          7102 => x"58",
          7103 => x"a0",
          7104 => x"73",
          7105 => x"09",
          7106 => x"38",
          7107 => x"1f",
          7108 => x"2e",
          7109 => x"88",
          7110 => x"2b",
          7111 => x"5c",
          7112 => x"54",
          7113 => x"8d",
          7114 => x"06",
          7115 => x"2e",
          7116 => x"85",
          7117 => x"07",
          7118 => x"2a",
          7119 => x"51",
          7120 => x"38",
          7121 => x"54",
          7122 => x"85",
          7123 => x"07",
          7124 => x"2a",
          7125 => x"51",
          7126 => x"2e",
          7127 => x"88",
          7128 => x"ab",
          7129 => x"51",
          7130 => x"82",
          7131 => x"ab",
          7132 => x"56",
          7133 => x"08",
          7134 => x"38",
          7135 => x"08",
          7136 => x"81",
          7137 => x"38",
          7138 => x"70",
          7139 => x"82",
          7140 => x"54",
          7141 => x"96",
          7142 => x"06",
          7143 => x"2e",
          7144 => x"ff",
          7145 => x"1f",
          7146 => x"80",
          7147 => x"81",
          7148 => x"bb",
          7149 => x"b7",
          7150 => x"2a",
          7151 => x"51",
          7152 => x"38",
          7153 => x"70",
          7154 => x"81",
          7155 => x"55",
          7156 => x"e1",
          7157 => x"08",
          7158 => x"60",
          7159 => x"52",
          7160 => x"ef",
          7161 => x"f8",
          7162 => x"0c",
          7163 => x"75",
          7164 => x"0c",
          7165 => x"04",
          7166 => x"7c",
          7167 => x"08",
          7168 => x"55",
          7169 => x"59",
          7170 => x"81",
          7171 => x"70",
          7172 => x"33",
          7173 => x"52",
          7174 => x"2e",
          7175 => x"ee",
          7176 => x"2e",
          7177 => x"81",
          7178 => x"33",
          7179 => x"81",
          7180 => x"52",
          7181 => x"26",
          7182 => x"14",
          7183 => x"06",
          7184 => x"52",
          7185 => x"80",
          7186 => x"0b",
          7187 => x"59",
          7188 => x"7a",
          7189 => x"70",
          7190 => x"33",
          7191 => x"05",
          7192 => x"9f",
          7193 => x"53",
          7194 => x"89",
          7195 => x"70",
          7196 => x"54",
          7197 => x"12",
          7198 => x"26",
          7199 => x"12",
          7200 => x"06",
          7201 => x"30",
          7202 => x"51",
          7203 => x"2e",
          7204 => x"85",
          7205 => x"be",
          7206 => x"74",
          7207 => x"30",
          7208 => x"9f",
          7209 => x"2a",
          7210 => x"54",
          7211 => x"2e",
          7212 => x"15",
          7213 => x"55",
          7214 => x"ff",
          7215 => x"39",
          7216 => x"86",
          7217 => x"7c",
          7218 => x"51",
          7219 => x"ec",
          7220 => x"70",
          7221 => x"0c",
          7222 => x"04",
          7223 => x"78",
          7224 => x"83",
          7225 => x"0b",
          7226 => x"79",
          7227 => x"d1",
          7228 => x"55",
          7229 => x"08",
          7230 => x"84",
          7231 => x"ce",
          7232 => x"d4",
          7233 => x"ff",
          7234 => x"83",
          7235 => x"d4",
          7236 => x"81",
          7237 => x"38",
          7238 => x"17",
          7239 => x"74",
          7240 => x"09",
          7241 => x"38",
          7242 => x"81",
          7243 => x"30",
          7244 => x"79",
          7245 => x"54",
          7246 => x"74",
          7247 => x"09",
          7248 => x"38",
          7249 => x"c6",
          7250 => x"ee",
          7251 => x"87",
          7252 => x"f8",
          7253 => x"d4",
          7254 => x"2e",
          7255 => x"53",
          7256 => x"52",
          7257 => x"51",
          7258 => x"82",
          7259 => x"55",
          7260 => x"08",
          7261 => x"38",
          7262 => x"82",
          7263 => x"88",
          7264 => x"f2",
          7265 => x"02",
          7266 => x"cb",
          7267 => x"55",
          7268 => x"60",
          7269 => x"3f",
          7270 => x"08",
          7271 => x"80",
          7272 => x"f8",
          7273 => x"84",
          7274 => x"f8",
          7275 => x"82",
          7276 => x"70",
          7277 => x"8c",
          7278 => x"2e",
          7279 => x"73",
          7280 => x"81",
          7281 => x"33",
          7282 => x"80",
          7283 => x"81",
          7284 => x"c6",
          7285 => x"d4",
          7286 => x"ff",
          7287 => x"06",
          7288 => x"98",
          7289 => x"2e",
          7290 => x"74",
          7291 => x"81",
          7292 => x"8a",
          7293 => x"b4",
          7294 => x"39",
          7295 => x"77",
          7296 => x"81",
          7297 => x"33",
          7298 => x"3f",
          7299 => x"08",
          7300 => x"70",
          7301 => x"55",
          7302 => x"86",
          7303 => x"80",
          7304 => x"74",
          7305 => x"81",
          7306 => x"8a",
          7307 => x"fc",
          7308 => x"53",
          7309 => x"fd",
          7310 => x"d4",
          7311 => x"ff",
          7312 => x"82",
          7313 => x"06",
          7314 => x"8c",
          7315 => x"58",
          7316 => x"fa",
          7317 => x"58",
          7318 => x"2e",
          7319 => x"fe",
          7320 => x"be",
          7321 => x"f8",
          7322 => x"78",
          7323 => x"5a",
          7324 => x"90",
          7325 => x"75",
          7326 => x"38",
          7327 => x"3d",
          7328 => x"70",
          7329 => x"08",
          7330 => x"7a",
          7331 => x"38",
          7332 => x"51",
          7333 => x"82",
          7334 => x"81",
          7335 => x"81",
          7336 => x"38",
          7337 => x"83",
          7338 => x"38",
          7339 => x"84",
          7340 => x"38",
          7341 => x"81",
          7342 => x"38",
          7343 => x"51",
          7344 => x"82",
          7345 => x"83",
          7346 => x"53",
          7347 => x"2e",
          7348 => x"84",
          7349 => x"ce",
          7350 => x"af",
          7351 => x"f8",
          7352 => x"ff",
          7353 => x"8d",
          7354 => x"14",
          7355 => x"3f",
          7356 => x"08",
          7357 => x"15",
          7358 => x"14",
          7359 => x"34",
          7360 => x"33",
          7361 => x"81",
          7362 => x"54",
          7363 => x"72",
          7364 => x"98",
          7365 => x"ff",
          7366 => x"29",
          7367 => x"33",
          7368 => x"72",
          7369 => x"72",
          7370 => x"38",
          7371 => x"06",
          7372 => x"2e",
          7373 => x"56",
          7374 => x"80",
          7375 => x"c9",
          7376 => x"d4",
          7377 => x"82",
          7378 => x"88",
          7379 => x"8f",
          7380 => x"56",
          7381 => x"38",
          7382 => x"51",
          7383 => x"82",
          7384 => x"83",
          7385 => x"55",
          7386 => x"80",
          7387 => x"c9",
          7388 => x"d4",
          7389 => x"80",
          7390 => x"c9",
          7391 => x"d4",
          7392 => x"ff",
          7393 => x"8d",
          7394 => x"2e",
          7395 => x"88",
          7396 => x"14",
          7397 => x"05",
          7398 => x"75",
          7399 => x"38",
          7400 => x"52",
          7401 => x"51",
          7402 => x"3f",
          7403 => x"08",
          7404 => x"f8",
          7405 => x"82",
          7406 => x"d4",
          7407 => x"ff",
          7408 => x"26",
          7409 => x"57",
          7410 => x"f5",
          7411 => x"82",
          7412 => x"f5",
          7413 => x"81",
          7414 => x"8d",
          7415 => x"2e",
          7416 => x"82",
          7417 => x"16",
          7418 => x"16",
          7419 => x"70",
          7420 => x"7a",
          7421 => x"0c",
          7422 => x"83",
          7423 => x"06",
          7424 => x"e2",
          7425 => x"83",
          7426 => x"f8",
          7427 => x"ff",
          7428 => x"56",
          7429 => x"38",
          7430 => x"38",
          7431 => x"51",
          7432 => x"82",
          7433 => x"ac",
          7434 => x"82",
          7435 => x"39",
          7436 => x"80",
          7437 => x"38",
          7438 => x"15",
          7439 => x"53",
          7440 => x"8d",
          7441 => x"15",
          7442 => x"76",
          7443 => x"51",
          7444 => x"13",
          7445 => x"8d",
          7446 => x"15",
          7447 => x"cc",
          7448 => x"94",
          7449 => x"0b",
          7450 => x"ff",
          7451 => x"15",
          7452 => x"2e",
          7453 => x"81",
          7454 => x"e8",
          7455 => x"8b",
          7456 => x"f8",
          7457 => x"ff",
          7458 => x"81",
          7459 => x"06",
          7460 => x"81",
          7461 => x"51",
          7462 => x"82",
          7463 => x"80",
          7464 => x"d4",
          7465 => x"15",
          7466 => x"14",
          7467 => x"3f",
          7468 => x"08",
          7469 => x"06",
          7470 => x"d4",
          7471 => x"81",
          7472 => x"38",
          7473 => x"c6",
          7474 => x"d4",
          7475 => x"8b",
          7476 => x"2e",
          7477 => x"b3",
          7478 => x"14",
          7479 => x"3f",
          7480 => x"08",
          7481 => x"e4",
          7482 => x"81",
          7483 => x"84",
          7484 => x"c6",
          7485 => x"d4",
          7486 => x"15",
          7487 => x"14",
          7488 => x"3f",
          7489 => x"08",
          7490 => x"76",
          7491 => x"ec",
          7492 => x"05",
          7493 => x"ec",
          7494 => x"86",
          7495 => x"ec",
          7496 => x"15",
          7497 => x"98",
          7498 => x"56",
          7499 => x"f8",
          7500 => x"0d",
          7501 => x"0d",
          7502 => x"55",
          7503 => x"ba",
          7504 => x"53",
          7505 => x"b2",
          7506 => x"52",
          7507 => x"aa",
          7508 => x"22",
          7509 => x"57",
          7510 => x"2e",
          7511 => x"9a",
          7512 => x"33",
          7513 => x"8d",
          7514 => x"f8",
          7515 => x"52",
          7516 => x"71",
          7517 => x"55",
          7518 => x"53",
          7519 => x"0c",
          7520 => x"d4",
          7521 => x"3d",
          7522 => x"3d",
          7523 => x"05",
          7524 => x"89",
          7525 => x"52",
          7526 => x"3f",
          7527 => x"0b",
          7528 => x"08",
          7529 => x"82",
          7530 => x"84",
          7531 => x"c0",
          7532 => x"55",
          7533 => x"2e",
          7534 => x"74",
          7535 => x"73",
          7536 => x"38",
          7537 => x"78",
          7538 => x"54",
          7539 => x"92",
          7540 => x"89",
          7541 => x"84",
          7542 => x"a7",
          7543 => x"f8",
          7544 => x"82",
          7545 => x"88",
          7546 => x"ea",
          7547 => x"02",
          7548 => x"eb",
          7549 => x"59",
          7550 => x"80",
          7551 => x"38",
          7552 => x"70",
          7553 => x"cc",
          7554 => x"3d",
          7555 => x"58",
          7556 => x"82",
          7557 => x"55",
          7558 => x"08",
          7559 => x"7a",
          7560 => x"8c",
          7561 => x"56",
          7562 => x"82",
          7563 => x"55",
          7564 => x"08",
          7565 => x"80",
          7566 => x"70",
          7567 => x"57",
          7568 => x"83",
          7569 => x"77",
          7570 => x"73",
          7571 => x"ab",
          7572 => x"2e",
          7573 => x"84",
          7574 => x"06",
          7575 => x"51",
          7576 => x"82",
          7577 => x"55",
          7578 => x"b2",
          7579 => x"06",
          7580 => x"b8",
          7581 => x"2a",
          7582 => x"51",
          7583 => x"2e",
          7584 => x"55",
          7585 => x"77",
          7586 => x"74",
          7587 => x"77",
          7588 => x"81",
          7589 => x"73",
          7590 => x"af",
          7591 => x"7a",
          7592 => x"3f",
          7593 => x"08",
          7594 => x"b2",
          7595 => x"8e",
          7596 => x"b7",
          7597 => x"a0",
          7598 => x"34",
          7599 => x"52",
          7600 => x"c8",
          7601 => x"62",
          7602 => x"c3",
          7603 => x"54",
          7604 => x"15",
          7605 => x"2e",
          7606 => x"7a",
          7607 => x"51",
          7608 => x"75",
          7609 => x"d0",
          7610 => x"c9",
          7611 => x"f8",
          7612 => x"d4",
          7613 => x"ca",
          7614 => x"74",
          7615 => x"02",
          7616 => x"70",
          7617 => x"81",
          7618 => x"56",
          7619 => x"86",
          7620 => x"82",
          7621 => x"81",
          7622 => x"06",
          7623 => x"80",
          7624 => x"75",
          7625 => x"73",
          7626 => x"38",
          7627 => x"92",
          7628 => x"7a",
          7629 => x"3f",
          7630 => x"08",
          7631 => x"90",
          7632 => x"55",
          7633 => x"08",
          7634 => x"77",
          7635 => x"81",
          7636 => x"73",
          7637 => x"38",
          7638 => x"07",
          7639 => x"11",
          7640 => x"0c",
          7641 => x"0c",
          7642 => x"52",
          7643 => x"3f",
          7644 => x"08",
          7645 => x"08",
          7646 => x"63",
          7647 => x"5a",
          7648 => x"82",
          7649 => x"82",
          7650 => x"8c",
          7651 => x"7a",
          7652 => x"17",
          7653 => x"23",
          7654 => x"34",
          7655 => x"1a",
          7656 => x"9c",
          7657 => x"0b",
          7658 => x"77",
          7659 => x"81",
          7660 => x"73",
          7661 => x"8d",
          7662 => x"f8",
          7663 => x"81",
          7664 => x"d4",
          7665 => x"1a",
          7666 => x"22",
          7667 => x"7b",
          7668 => x"a8",
          7669 => x"78",
          7670 => x"3f",
          7671 => x"08",
          7672 => x"f8",
          7673 => x"83",
          7674 => x"82",
          7675 => x"ff",
          7676 => x"06",
          7677 => x"55",
          7678 => x"56",
          7679 => x"76",
          7680 => x"51",
          7681 => x"27",
          7682 => x"70",
          7683 => x"5a",
          7684 => x"76",
          7685 => x"74",
          7686 => x"83",
          7687 => x"73",
          7688 => x"38",
          7689 => x"51",
          7690 => x"82",
          7691 => x"85",
          7692 => x"8e",
          7693 => x"2a",
          7694 => x"08",
          7695 => x"0c",
          7696 => x"79",
          7697 => x"73",
          7698 => x"0c",
          7699 => x"04",
          7700 => x"60",
          7701 => x"40",
          7702 => x"80",
          7703 => x"3d",
          7704 => x"78",
          7705 => x"3f",
          7706 => x"08",
          7707 => x"f8",
          7708 => x"91",
          7709 => x"74",
          7710 => x"38",
          7711 => x"c7",
          7712 => x"33",
          7713 => x"87",
          7714 => x"2e",
          7715 => x"95",
          7716 => x"91",
          7717 => x"56",
          7718 => x"81",
          7719 => x"34",
          7720 => x"a3",
          7721 => x"08",
          7722 => x"31",
          7723 => x"27",
          7724 => x"5c",
          7725 => x"82",
          7726 => x"19",
          7727 => x"ff",
          7728 => x"74",
          7729 => x"7e",
          7730 => x"ff",
          7731 => x"2a",
          7732 => x"79",
          7733 => x"87",
          7734 => x"08",
          7735 => x"98",
          7736 => x"78",
          7737 => x"3f",
          7738 => x"08",
          7739 => x"27",
          7740 => x"74",
          7741 => x"a3",
          7742 => x"1a",
          7743 => x"08",
          7744 => x"c3",
          7745 => x"d4",
          7746 => x"2e",
          7747 => x"82",
          7748 => x"1a",
          7749 => x"59",
          7750 => x"2e",
          7751 => x"77",
          7752 => x"11",
          7753 => x"55",
          7754 => x"85",
          7755 => x"31",
          7756 => x"76",
          7757 => x"81",
          7758 => x"ff",
          7759 => x"82",
          7760 => x"fe",
          7761 => x"83",
          7762 => x"56",
          7763 => x"a0",
          7764 => x"08",
          7765 => x"74",
          7766 => x"38",
          7767 => x"b8",
          7768 => x"16",
          7769 => x"89",
          7770 => x"51",
          7771 => x"3f",
          7772 => x"56",
          7773 => x"9c",
          7774 => x"19",
          7775 => x"06",
          7776 => x"31",
          7777 => x"76",
          7778 => x"7b",
          7779 => x"08",
          7780 => x"c0",
          7781 => x"d4",
          7782 => x"ff",
          7783 => x"94",
          7784 => x"ff",
          7785 => x"05",
          7786 => x"ff",
          7787 => x"7b",
          7788 => x"08",
          7789 => x"76",
          7790 => x"08",
          7791 => x"0c",
          7792 => x"f0",
          7793 => x"75",
          7794 => x"0c",
          7795 => x"04",
          7796 => x"60",
          7797 => x"40",
          7798 => x"80",
          7799 => x"3d",
          7800 => x"77",
          7801 => x"3f",
          7802 => x"08",
          7803 => x"f8",
          7804 => x"91",
          7805 => x"74",
          7806 => x"38",
          7807 => x"be",
          7808 => x"33",
          7809 => x"70",
          7810 => x"56",
          7811 => x"74",
          7812 => x"aa",
          7813 => x"82",
          7814 => x"34",
          7815 => x"9e",
          7816 => x"91",
          7817 => x"56",
          7818 => x"94",
          7819 => x"11",
          7820 => x"76",
          7821 => x"75",
          7822 => x"80",
          7823 => x"38",
          7824 => x"70",
          7825 => x"56",
          7826 => x"81",
          7827 => x"11",
          7828 => x"77",
          7829 => x"5c",
          7830 => x"38",
          7831 => x"88",
          7832 => x"74",
          7833 => x"52",
          7834 => x"18",
          7835 => x"51",
          7836 => x"82",
          7837 => x"55",
          7838 => x"08",
          7839 => x"b1",
          7840 => x"2e",
          7841 => x"74",
          7842 => x"95",
          7843 => x"19",
          7844 => x"08",
          7845 => x"88",
          7846 => x"55",
          7847 => x"9c",
          7848 => x"09",
          7849 => x"38",
          7850 => x"bd",
          7851 => x"d4",
          7852 => x"ed",
          7853 => x"08",
          7854 => x"c0",
          7855 => x"d4",
          7856 => x"2e",
          7857 => x"82",
          7858 => x"1b",
          7859 => x"5a",
          7860 => x"2e",
          7861 => x"78",
          7862 => x"11",
          7863 => x"55",
          7864 => x"85",
          7865 => x"31",
          7866 => x"76",
          7867 => x"81",
          7868 => x"ff",
          7869 => x"82",
          7870 => x"fe",
          7871 => x"b4",
          7872 => x"31",
          7873 => x"79",
          7874 => x"84",
          7875 => x"16",
          7876 => x"89",
          7877 => x"52",
          7878 => x"ff",
          7879 => x"7e",
          7880 => x"83",
          7881 => x"89",
          7882 => x"de",
          7883 => x"08",
          7884 => x"26",
          7885 => x"51",
          7886 => x"3f",
          7887 => x"08",
          7888 => x"7e",
          7889 => x"0c",
          7890 => x"19",
          7891 => x"08",
          7892 => x"84",
          7893 => x"57",
          7894 => x"27",
          7895 => x"56",
          7896 => x"52",
          7897 => x"bc",
          7898 => x"d4",
          7899 => x"b1",
          7900 => x"7c",
          7901 => x"08",
          7902 => x"1f",
          7903 => x"ff",
          7904 => x"7e",
          7905 => x"83",
          7906 => x"76",
          7907 => x"17",
          7908 => x"1e",
          7909 => x"18",
          7910 => x"0c",
          7911 => x"58",
          7912 => x"74",
          7913 => x"38",
          7914 => x"8c",
          7915 => x"8a",
          7916 => x"33",
          7917 => x"55",
          7918 => x"34",
          7919 => x"82",
          7920 => x"90",
          7921 => x"f8",
          7922 => x"8b",
          7923 => x"53",
          7924 => x"f2",
          7925 => x"d4",
          7926 => x"82",
          7927 => x"81",
          7928 => x"16",
          7929 => x"2a",
          7930 => x"51",
          7931 => x"80",
          7932 => x"38",
          7933 => x"52",
          7934 => x"bb",
          7935 => x"d4",
          7936 => x"82",
          7937 => x"80",
          7938 => x"16",
          7939 => x"33",
          7940 => x"55",
          7941 => x"34",
          7942 => x"53",
          7943 => x"08",
          7944 => x"3f",
          7945 => x"52",
          7946 => x"ff",
          7947 => x"82",
          7948 => x"52",
          7949 => x"ff",
          7950 => x"76",
          7951 => x"51",
          7952 => x"3f",
          7953 => x"0b",
          7954 => x"78",
          7955 => x"dc",
          7956 => x"f8",
          7957 => x"33",
          7958 => x"55",
          7959 => x"17",
          7960 => x"d4",
          7961 => x"3d",
          7962 => x"3d",
          7963 => x"52",
          7964 => x"3f",
          7965 => x"08",
          7966 => x"f8",
          7967 => x"86",
          7968 => x"52",
          7969 => x"ad",
          7970 => x"f8",
          7971 => x"d4",
          7972 => x"38",
          7973 => x"08",
          7974 => x"82",
          7975 => x"86",
          7976 => x"ff",
          7977 => x"3d",
          7978 => x"3f",
          7979 => x"0b",
          7980 => x"08",
          7981 => x"82",
          7982 => x"82",
          7983 => x"80",
          7984 => x"d4",
          7985 => x"3d",
          7986 => x"3d",
          7987 => x"94",
          7988 => x"52",
          7989 => x"e9",
          7990 => x"d4",
          7991 => x"82",
          7992 => x"80",
          7993 => x"58",
          7994 => x"3d",
          7995 => x"dd",
          7996 => x"d4",
          7997 => x"82",
          7998 => x"bc",
          7999 => x"c7",
          8000 => x"98",
          8001 => x"73",
          8002 => x"38",
          8003 => x"12",
          8004 => x"39",
          8005 => x"33",
          8006 => x"70",
          8007 => x"55",
          8008 => x"2e",
          8009 => x"7f",
          8010 => x"54",
          8011 => x"82",
          8012 => x"98",
          8013 => x"39",
          8014 => x"08",
          8015 => x"81",
          8016 => x"85",
          8017 => x"d4",
          8018 => x"3d",
          8019 => x"a3",
          8020 => x"e1",
          8021 => x"e1",
          8022 => x"5b",
          8023 => x"80",
          8024 => x"3d",
          8025 => x"52",
          8026 => x"51",
          8027 => x"82",
          8028 => x"57",
          8029 => x"08",
          8030 => x"7b",
          8031 => x"0c",
          8032 => x"11",
          8033 => x"3d",
          8034 => x"80",
          8035 => x"54",
          8036 => x"82",
          8037 => x"52",
          8038 => x"70",
          8039 => x"d4",
          8040 => x"f8",
          8041 => x"d4",
          8042 => x"ef",
          8043 => x"3d",
          8044 => x"51",
          8045 => x"3f",
          8046 => x"08",
          8047 => x"f8",
          8048 => x"38",
          8049 => x"08",
          8050 => x"c9",
          8051 => x"d4",
          8052 => x"d6",
          8053 => x"52",
          8054 => x"98",
          8055 => x"f8",
          8056 => x"d4",
          8057 => x"b3",
          8058 => x"74",
          8059 => x"3f",
          8060 => x"08",
          8061 => x"f8",
          8062 => x"80",
          8063 => x"52",
          8064 => x"cf",
          8065 => x"d4",
          8066 => x"a6",
          8067 => x"74",
          8068 => x"3f",
          8069 => x"08",
          8070 => x"f8",
          8071 => x"c9",
          8072 => x"2e",
          8073 => x"86",
          8074 => x"81",
          8075 => x"81",
          8076 => x"df",
          8077 => x"05",
          8078 => x"d6",
          8079 => x"93",
          8080 => x"82",
          8081 => x"56",
          8082 => x"80",
          8083 => x"02",
          8084 => x"55",
          8085 => x"16",
          8086 => x"56",
          8087 => x"38",
          8088 => x"73",
          8089 => x"99",
          8090 => x"2e",
          8091 => x"16",
          8092 => x"ff",
          8093 => x"3d",
          8094 => x"18",
          8095 => x"58",
          8096 => x"33",
          8097 => x"eb",
          8098 => x"80",
          8099 => x"11",
          8100 => x"74",
          8101 => x"39",
          8102 => x"09",
          8103 => x"38",
          8104 => x"e1",
          8105 => x"55",
          8106 => x"34",
          8107 => x"ec",
          8108 => x"84",
          8109 => x"f0",
          8110 => x"70",
          8111 => x"56",
          8112 => x"76",
          8113 => x"81",
          8114 => x"70",
          8115 => x"56",
          8116 => x"82",
          8117 => x"78",
          8118 => x"80",
          8119 => x"27",
          8120 => x"19",
          8121 => x"7a",
          8122 => x"5c",
          8123 => x"55",
          8124 => x"7a",
          8125 => x"5c",
          8126 => x"2e",
          8127 => x"85",
          8128 => x"97",
          8129 => x"3d",
          8130 => x"19",
          8131 => x"33",
          8132 => x"05",
          8133 => x"78",
          8134 => x"80",
          8135 => x"82",
          8136 => x"80",
          8137 => x"04",
          8138 => x"7b",
          8139 => x"fc",
          8140 => x"53",
          8141 => x"fd",
          8142 => x"f8",
          8143 => x"d4",
          8144 => x"fe",
          8145 => x"33",
          8146 => x"f6",
          8147 => x"08",
          8148 => x"27",
          8149 => x"15",
          8150 => x"2a",
          8151 => x"51",
          8152 => x"83",
          8153 => x"94",
          8154 => x"80",
          8155 => x"0c",
          8156 => x"2e",
          8157 => x"79",
          8158 => x"70",
          8159 => x"51",
          8160 => x"2e",
          8161 => x"52",
          8162 => x"fe",
          8163 => x"82",
          8164 => x"ff",
          8165 => x"70",
          8166 => x"fe",
          8167 => x"82",
          8168 => x"73",
          8169 => x"76",
          8170 => x"06",
          8171 => x"0c",
          8172 => x"98",
          8173 => x"58",
          8174 => x"39",
          8175 => x"54",
          8176 => x"73",
          8177 => x"ff",
          8178 => x"82",
          8179 => x"54",
          8180 => x"08",
          8181 => x"9d",
          8182 => x"f8",
          8183 => x"81",
          8184 => x"d4",
          8185 => x"16",
          8186 => x"16",
          8187 => x"2e",
          8188 => x"76",
          8189 => x"de",
          8190 => x"31",
          8191 => x"18",
          8192 => x"90",
          8193 => x"81",
          8194 => x"06",
          8195 => x"56",
          8196 => x"9b",
          8197 => x"74",
          8198 => x"c5",
          8199 => x"f8",
          8200 => x"d4",
          8201 => x"38",
          8202 => x"08",
          8203 => x"73",
          8204 => x"ff",
          8205 => x"82",
          8206 => x"54",
          8207 => x"bf",
          8208 => x"27",
          8209 => x"53",
          8210 => x"08",
          8211 => x"73",
          8212 => x"ff",
          8213 => x"15",
          8214 => x"16",
          8215 => x"ff",
          8216 => x"80",
          8217 => x"73",
          8218 => x"ff",
          8219 => x"82",
          8220 => x"94",
          8221 => x"91",
          8222 => x"53",
          8223 => x"81",
          8224 => x"34",
          8225 => x"39",
          8226 => x"82",
          8227 => x"05",
          8228 => x"08",
          8229 => x"08",
          8230 => x"38",
          8231 => x"0c",
          8232 => x"80",
          8233 => x"72",
          8234 => x"73",
          8235 => x"53",
          8236 => x"8c",
          8237 => x"16",
          8238 => x"38",
          8239 => x"0c",
          8240 => x"82",
          8241 => x"8b",
          8242 => x"f9",
          8243 => x"56",
          8244 => x"80",
          8245 => x"38",
          8246 => x"3d",
          8247 => x"8a",
          8248 => x"51",
          8249 => x"82",
          8250 => x"55",
          8251 => x"08",
          8252 => x"77",
          8253 => x"52",
          8254 => x"a1",
          8255 => x"f8",
          8256 => x"d4",
          8257 => x"c4",
          8258 => x"33",
          8259 => x"55",
          8260 => x"24",
          8261 => x"16",
          8262 => x"2a",
          8263 => x"51",
          8264 => x"80",
          8265 => x"9c",
          8266 => x"77",
          8267 => x"3f",
          8268 => x"08",
          8269 => x"77",
          8270 => x"22",
          8271 => x"74",
          8272 => x"ff",
          8273 => x"82",
          8274 => x"55",
          8275 => x"09",
          8276 => x"38",
          8277 => x"39",
          8278 => x"84",
          8279 => x"0c",
          8280 => x"82",
          8281 => x"89",
          8282 => x"fc",
          8283 => x"87",
          8284 => x"53",
          8285 => x"e7",
          8286 => x"d4",
          8287 => x"38",
          8288 => x"08",
          8289 => x"3d",
          8290 => x"3d",
          8291 => x"89",
          8292 => x"54",
          8293 => x"54",
          8294 => x"82",
          8295 => x"53",
          8296 => x"08",
          8297 => x"74",
          8298 => x"d4",
          8299 => x"73",
          8300 => x"c0",
          8301 => x"f8",
          8302 => x"cb",
          8303 => x"f8",
          8304 => x"51",
          8305 => x"82",
          8306 => x"53",
          8307 => x"08",
          8308 => x"81",
          8309 => x"80",
          8310 => x"82",
          8311 => x"a7",
          8312 => x"73",
          8313 => x"3f",
          8314 => x"51",
          8315 => x"3f",
          8316 => x"08",
          8317 => x"30",
          8318 => x"9f",
          8319 => x"d4",
          8320 => x"51",
          8321 => x"72",
          8322 => x"0c",
          8323 => x"04",
          8324 => x"66",
          8325 => x"89",
          8326 => x"97",
          8327 => x"de",
          8328 => x"d4",
          8329 => x"82",
          8330 => x"b2",
          8331 => x"75",
          8332 => x"3f",
          8333 => x"08",
          8334 => x"f8",
          8335 => x"02",
          8336 => x"33",
          8337 => x"55",
          8338 => x"25",
          8339 => x"55",
          8340 => x"80",
          8341 => x"76",
          8342 => x"ce",
          8343 => x"82",
          8344 => x"95",
          8345 => x"f0",
          8346 => x"65",
          8347 => x"53",
          8348 => x"05",
          8349 => x"51",
          8350 => x"82",
          8351 => x"5b",
          8352 => x"08",
          8353 => x"7c",
          8354 => x"08",
          8355 => x"fe",
          8356 => x"08",
          8357 => x"55",
          8358 => x"91",
          8359 => x"0c",
          8360 => x"81",
          8361 => x"39",
          8362 => x"c9",
          8363 => x"f8",
          8364 => x"55",
          8365 => x"2e",
          8366 => x"80",
          8367 => x"75",
          8368 => x"52",
          8369 => x"05",
          8370 => x"b9",
          8371 => x"f8",
          8372 => x"cf",
          8373 => x"f8",
          8374 => x"cc",
          8375 => x"f8",
          8376 => x"82",
          8377 => x"07",
          8378 => x"05",
          8379 => x"53",
          8380 => x"9c",
          8381 => x"26",
          8382 => x"f9",
          8383 => x"08",
          8384 => x"08",
          8385 => x"98",
          8386 => x"81",
          8387 => x"58",
          8388 => x"3f",
          8389 => x"08",
          8390 => x"f8",
          8391 => x"38",
          8392 => x"77",
          8393 => x"5d",
          8394 => x"74",
          8395 => x"81",
          8396 => x"b8",
          8397 => x"a9",
          8398 => x"d4",
          8399 => x"ff",
          8400 => x"30",
          8401 => x"1b",
          8402 => x"5b",
          8403 => x"39",
          8404 => x"ff",
          8405 => x"82",
          8406 => x"f0",
          8407 => x"30",
          8408 => x"1b",
          8409 => x"5b",
          8410 => x"83",
          8411 => x"58",
          8412 => x"92",
          8413 => x"0c",
          8414 => x"12",
          8415 => x"33",
          8416 => x"54",
          8417 => x"34",
          8418 => x"f8",
          8419 => x"0d",
          8420 => x"0d",
          8421 => x"fc",
          8422 => x"52",
          8423 => x"3f",
          8424 => x"08",
          8425 => x"f8",
          8426 => x"38",
          8427 => x"56",
          8428 => x"38",
          8429 => x"70",
          8430 => x"81",
          8431 => x"55",
          8432 => x"80",
          8433 => x"38",
          8434 => x"54",
          8435 => x"08",
          8436 => x"38",
          8437 => x"82",
          8438 => x"53",
          8439 => x"52",
          8440 => x"b2",
          8441 => x"d4",
          8442 => x"88",
          8443 => x"80",
          8444 => x"17",
          8445 => x"51",
          8446 => x"3f",
          8447 => x"08",
          8448 => x"81",
          8449 => x"81",
          8450 => x"f8",
          8451 => x"09",
          8452 => x"38",
          8453 => x"39",
          8454 => x"77",
          8455 => x"f8",
          8456 => x"08",
          8457 => x"98",
          8458 => x"82",
          8459 => x"52",
          8460 => x"b2",
          8461 => x"d4",
          8462 => x"94",
          8463 => x"18",
          8464 => x"33",
          8465 => x"54",
          8466 => x"34",
          8467 => x"85",
          8468 => x"18",
          8469 => x"74",
          8470 => x"0c",
          8471 => x"04",
          8472 => x"82",
          8473 => x"ff",
          8474 => x"a3",
          8475 => x"93",
          8476 => x"f8",
          8477 => x"d4",
          8478 => x"f9",
          8479 => x"a3",
          8480 => x"96",
          8481 => x"58",
          8482 => x"82",
          8483 => x"55",
          8484 => x"08",
          8485 => x"02",
          8486 => x"33",
          8487 => x"70",
          8488 => x"55",
          8489 => x"73",
          8490 => x"75",
          8491 => x"80",
          8492 => x"c1",
          8493 => x"da",
          8494 => x"81",
          8495 => x"87",
          8496 => x"b1",
          8497 => x"78",
          8498 => x"87",
          8499 => x"f8",
          8500 => x"2a",
          8501 => x"51",
          8502 => x"80",
          8503 => x"38",
          8504 => x"d4",
          8505 => x"15",
          8506 => x"89",
          8507 => x"82",
          8508 => x"5c",
          8509 => x"3d",
          8510 => x"ff",
          8511 => x"82",
          8512 => x"55",
          8513 => x"08",
          8514 => x"82",
          8515 => x"52",
          8516 => x"bb",
          8517 => x"d4",
          8518 => x"82",
          8519 => x"86",
          8520 => x"80",
          8521 => x"d4",
          8522 => x"2e",
          8523 => x"d4",
          8524 => x"c1",
          8525 => x"c7",
          8526 => x"d4",
          8527 => x"d4",
          8528 => x"70",
          8529 => x"08",
          8530 => x"51",
          8531 => x"80",
          8532 => x"73",
          8533 => x"38",
          8534 => x"52",
          8535 => x"af",
          8536 => x"d4",
          8537 => x"74",
          8538 => x"51",
          8539 => x"3f",
          8540 => x"08",
          8541 => x"d4",
          8542 => x"3d",
          8543 => x"3d",
          8544 => x"9a",
          8545 => x"05",
          8546 => x"51",
          8547 => x"82",
          8548 => x"54",
          8549 => x"08",
          8550 => x"78",
          8551 => x"8e",
          8552 => x"58",
          8553 => x"82",
          8554 => x"54",
          8555 => x"08",
          8556 => x"54",
          8557 => x"82",
          8558 => x"84",
          8559 => x"06",
          8560 => x"02",
          8561 => x"33",
          8562 => x"81",
          8563 => x"86",
          8564 => x"fd",
          8565 => x"74",
          8566 => x"70",
          8567 => x"b0",
          8568 => x"d4",
          8569 => x"55",
          8570 => x"f8",
          8571 => x"87",
          8572 => x"f8",
          8573 => x"09",
          8574 => x"38",
          8575 => x"d4",
          8576 => x"2e",
          8577 => x"86",
          8578 => x"81",
          8579 => x"81",
          8580 => x"d4",
          8581 => x"78",
          8582 => x"e0",
          8583 => x"f8",
          8584 => x"d4",
          8585 => x"9f",
          8586 => x"a0",
          8587 => x"51",
          8588 => x"3f",
          8589 => x"0b",
          8590 => x"78",
          8591 => x"80",
          8592 => x"82",
          8593 => x"52",
          8594 => x"51",
          8595 => x"3f",
          8596 => x"b8",
          8597 => x"ff",
          8598 => x"a0",
          8599 => x"11",
          8600 => x"05",
          8601 => x"b2",
          8602 => x"ae",
          8603 => x"15",
          8604 => x"78",
          8605 => x"53",
          8606 => x"90",
          8607 => x"81",
          8608 => x"34",
          8609 => x"bf",
          8610 => x"d4",
          8611 => x"82",
          8612 => x"b3",
          8613 => x"b2",
          8614 => x"96",
          8615 => x"a3",
          8616 => x"53",
          8617 => x"51",
          8618 => x"3f",
          8619 => x"0b",
          8620 => x"78",
          8621 => x"83",
          8622 => x"51",
          8623 => x"3f",
          8624 => x"08",
          8625 => x"80",
          8626 => x"76",
          8627 => x"e5",
          8628 => x"d4",
          8629 => x"3d",
          8630 => x"3d",
          8631 => x"84",
          8632 => x"94",
          8633 => x"aa",
          8634 => x"05",
          8635 => x"51",
          8636 => x"82",
          8637 => x"55",
          8638 => x"08",
          8639 => x"78",
          8640 => x"08",
          8641 => x"70",
          8642 => x"91",
          8643 => x"f8",
          8644 => x"d4",
          8645 => x"be",
          8646 => x"9f",
          8647 => x"a0",
          8648 => x"55",
          8649 => x"38",
          8650 => x"3d",
          8651 => x"3d",
          8652 => x"51",
          8653 => x"3f",
          8654 => x"52",
          8655 => x"52",
          8656 => x"d6",
          8657 => x"08",
          8658 => x"c8",
          8659 => x"d4",
          8660 => x"82",
          8661 => x"97",
          8662 => x"3d",
          8663 => x"81",
          8664 => x"65",
          8665 => x"2e",
          8666 => x"55",
          8667 => x"82",
          8668 => x"84",
          8669 => x"06",
          8670 => x"73",
          8671 => x"d6",
          8672 => x"f8",
          8673 => x"d4",
          8674 => x"ca",
          8675 => x"93",
          8676 => x"ff",
          8677 => x"8d",
          8678 => x"a1",
          8679 => x"af",
          8680 => x"17",
          8681 => x"33",
          8682 => x"70",
          8683 => x"55",
          8684 => x"38",
          8685 => x"54",
          8686 => x"34",
          8687 => x"0b",
          8688 => x"8b",
          8689 => x"84",
          8690 => x"06",
          8691 => x"73",
          8692 => x"e7",
          8693 => x"2e",
          8694 => x"75",
          8695 => x"ff",
          8696 => x"82",
          8697 => x"52",
          8698 => x"a5",
          8699 => x"55",
          8700 => x"08",
          8701 => x"de",
          8702 => x"f8",
          8703 => x"51",
          8704 => x"3f",
          8705 => x"08",
          8706 => x"11",
          8707 => x"82",
          8708 => x"80",
          8709 => x"16",
          8710 => x"ae",
          8711 => x"06",
          8712 => x"53",
          8713 => x"51",
          8714 => x"3f",
          8715 => x"0b",
          8716 => x"87",
          8717 => x"f8",
          8718 => x"77",
          8719 => x"3f",
          8720 => x"08",
          8721 => x"f8",
          8722 => x"78",
          8723 => x"dc",
          8724 => x"f8",
          8725 => x"82",
          8726 => x"aa",
          8727 => x"ec",
          8728 => x"80",
          8729 => x"02",
          8730 => x"e3",
          8731 => x"57",
          8732 => x"3d",
          8733 => x"97",
          8734 => x"87",
          8735 => x"f8",
          8736 => x"d4",
          8737 => x"cf",
          8738 => x"66",
          8739 => x"d0",
          8740 => x"89",
          8741 => x"f8",
          8742 => x"d4",
          8743 => x"38",
          8744 => x"05",
          8745 => x"06",
          8746 => x"73",
          8747 => x"a7",
          8748 => x"09",
          8749 => x"71",
          8750 => x"06",
          8751 => x"55",
          8752 => x"15",
          8753 => x"81",
          8754 => x"34",
          8755 => x"a2",
          8756 => x"d4",
          8757 => x"74",
          8758 => x"0c",
          8759 => x"04",
          8760 => x"65",
          8761 => x"94",
          8762 => x"52",
          8763 => x"d1",
          8764 => x"d4",
          8765 => x"82",
          8766 => x"80",
          8767 => x"58",
          8768 => x"3d",
          8769 => x"c5",
          8770 => x"d4",
          8771 => x"82",
          8772 => x"b4",
          8773 => x"c7",
          8774 => x"a0",
          8775 => x"55",
          8776 => x"84",
          8777 => x"17",
          8778 => x"2b",
          8779 => x"96",
          8780 => x"9e",
          8781 => x"54",
          8782 => x"15",
          8783 => x"ff",
          8784 => x"82",
          8785 => x"55",
          8786 => x"f8",
          8787 => x"0d",
          8788 => x"0d",
          8789 => x"5a",
          8790 => x"3d",
          8791 => x"9a",
          8792 => x"9f",
          8793 => x"f8",
          8794 => x"f8",
          8795 => x"82",
          8796 => x"07",
          8797 => x"55",
          8798 => x"2e",
          8799 => x"81",
          8800 => x"55",
          8801 => x"2e",
          8802 => x"7b",
          8803 => x"80",
          8804 => x"70",
          8805 => x"ac",
          8806 => x"d4",
          8807 => x"82",
          8808 => x"80",
          8809 => x"52",
          8810 => x"b2",
          8811 => x"d4",
          8812 => x"82",
          8813 => x"bf",
          8814 => x"f8",
          8815 => x"f8",
          8816 => x"59",
          8817 => x"81",
          8818 => x"56",
          8819 => x"33",
          8820 => x"16",
          8821 => x"27",
          8822 => x"56",
          8823 => x"80",
          8824 => x"80",
          8825 => x"ff",
          8826 => x"70",
          8827 => x"56",
          8828 => x"e8",
          8829 => x"76",
          8830 => x"81",
          8831 => x"80",
          8832 => x"57",
          8833 => x"78",
          8834 => x"51",
          8835 => x"2e",
          8836 => x"73",
          8837 => x"38",
          8838 => x"08",
          8839 => x"9f",
          8840 => x"d4",
          8841 => x"82",
          8842 => x"a7",
          8843 => x"33",
          8844 => x"c3",
          8845 => x"2e",
          8846 => x"e4",
          8847 => x"2e",
          8848 => x"56",
          8849 => x"05",
          8850 => x"d6",
          8851 => x"f8",
          8852 => x"76",
          8853 => x"0c",
          8854 => x"04",
          8855 => x"82",
          8856 => x"ff",
          8857 => x"9d",
          8858 => x"97",
          8859 => x"f8",
          8860 => x"f8",
          8861 => x"82",
          8862 => x"82",
          8863 => x"53",
          8864 => x"3d",
          8865 => x"ff",
          8866 => x"73",
          8867 => x"51",
          8868 => x"74",
          8869 => x"38",
          8870 => x"3d",
          8871 => x"90",
          8872 => x"f8",
          8873 => x"ff",
          8874 => x"38",
          8875 => x"08",
          8876 => x"3f",
          8877 => x"82",
          8878 => x"51",
          8879 => x"82",
          8880 => x"83",
          8881 => x"55",
          8882 => x"a3",
          8883 => x"82",
          8884 => x"ff",
          8885 => x"82",
          8886 => x"93",
          8887 => x"75",
          8888 => x"75",
          8889 => x"38",
          8890 => x"76",
          8891 => x"86",
          8892 => x"39",
          8893 => x"27",
          8894 => x"88",
          8895 => x"77",
          8896 => x"59",
          8897 => x"56",
          8898 => x"81",
          8899 => x"81",
          8900 => x"33",
          8901 => x"73",
          8902 => x"fe",
          8903 => x"33",
          8904 => x"73",
          8905 => x"81",
          8906 => x"80",
          8907 => x"02",
          8908 => x"75",
          8909 => x"51",
          8910 => x"2e",
          8911 => x"87",
          8912 => x"56",
          8913 => x"78",
          8914 => x"80",
          8915 => x"70",
          8916 => x"a9",
          8917 => x"d4",
          8918 => x"82",
          8919 => x"80",
          8920 => x"52",
          8921 => x"af",
          8922 => x"d4",
          8923 => x"82",
          8924 => x"8d",
          8925 => x"c4",
          8926 => x"e5",
          8927 => x"c6",
          8928 => x"f8",
          8929 => x"09",
          8930 => x"cc",
          8931 => x"75",
          8932 => x"c4",
          8933 => x"74",
          8934 => x"9c",
          8935 => x"f8",
          8936 => x"d4",
          8937 => x"38",
          8938 => x"d4",
          8939 => x"66",
          8940 => x"89",
          8941 => x"88",
          8942 => x"34",
          8943 => x"52",
          8944 => x"99",
          8945 => x"54",
          8946 => x"15",
          8947 => x"ff",
          8948 => x"82",
          8949 => x"54",
          8950 => x"82",
          8951 => x"9c",
          8952 => x"f2",
          8953 => x"62",
          8954 => x"80",
          8955 => x"93",
          8956 => x"55",
          8957 => x"5e",
          8958 => x"3f",
          8959 => x"08",
          8960 => x"f8",
          8961 => x"38",
          8962 => x"58",
          8963 => x"38",
          8964 => x"97",
          8965 => x"08",
          8966 => x"38",
          8967 => x"70",
          8968 => x"81",
          8969 => x"55",
          8970 => x"87",
          8971 => x"39",
          8972 => x"90",
          8973 => x"82",
          8974 => x"8a",
          8975 => x"89",
          8976 => x"7f",
          8977 => x"56",
          8978 => x"3f",
          8979 => x"06",
          8980 => x"72",
          8981 => x"82",
          8982 => x"05",
          8983 => x"7c",
          8984 => x"55",
          8985 => x"27",
          8986 => x"16",
          8987 => x"83",
          8988 => x"76",
          8989 => x"80",
          8990 => x"79",
          8991 => x"85",
          8992 => x"7f",
          8993 => x"14",
          8994 => x"83",
          8995 => x"82",
          8996 => x"81",
          8997 => x"38",
          8998 => x"08",
          8999 => x"95",
          9000 => x"f8",
          9001 => x"81",
          9002 => x"7b",
          9003 => x"06",
          9004 => x"39",
          9005 => x"56",
          9006 => x"09",
          9007 => x"b9",
          9008 => x"80",
          9009 => x"80",
          9010 => x"78",
          9011 => x"7a",
          9012 => x"38",
          9013 => x"73",
          9014 => x"81",
          9015 => x"ff",
          9016 => x"74",
          9017 => x"ff",
          9018 => x"82",
          9019 => x"58",
          9020 => x"08",
          9021 => x"74",
          9022 => x"16",
          9023 => x"73",
          9024 => x"39",
          9025 => x"7e",
          9026 => x"0c",
          9027 => x"2e",
          9028 => x"88",
          9029 => x"8c",
          9030 => x"1a",
          9031 => x"07",
          9032 => x"1b",
          9033 => x"08",
          9034 => x"16",
          9035 => x"75",
          9036 => x"38",
          9037 => x"94",
          9038 => x"15",
          9039 => x"54",
          9040 => x"34",
          9041 => x"82",
          9042 => x"90",
          9043 => x"e9",
          9044 => x"6d",
          9045 => x"80",
          9046 => x"9d",
          9047 => x"5c",
          9048 => x"3f",
          9049 => x"0b",
          9050 => x"08",
          9051 => x"38",
          9052 => x"08",
          9053 => x"ec",
          9054 => x"08",
          9055 => x"80",
          9056 => x"80",
          9057 => x"d4",
          9058 => x"ff",
          9059 => x"52",
          9060 => x"8e",
          9061 => x"d4",
          9062 => x"ff",
          9063 => x"06",
          9064 => x"56",
          9065 => x"38",
          9066 => x"70",
          9067 => x"55",
          9068 => x"8b",
          9069 => x"3d",
          9070 => x"83",
          9071 => x"ff",
          9072 => x"82",
          9073 => x"99",
          9074 => x"74",
          9075 => x"38",
          9076 => x"80",
          9077 => x"ff",
          9078 => x"55",
          9079 => x"83",
          9080 => x"78",
          9081 => x"38",
          9082 => x"26",
          9083 => x"81",
          9084 => x"8b",
          9085 => x"79",
          9086 => x"80",
          9087 => x"93",
          9088 => x"39",
          9089 => x"6e",
          9090 => x"89",
          9091 => x"48",
          9092 => x"83",
          9093 => x"61",
          9094 => x"25",
          9095 => x"55",
          9096 => x"8a",
          9097 => x"3d",
          9098 => x"81",
          9099 => x"ff",
          9100 => x"81",
          9101 => x"f8",
          9102 => x"38",
          9103 => x"70",
          9104 => x"d4",
          9105 => x"56",
          9106 => x"38",
          9107 => x"55",
          9108 => x"75",
          9109 => x"38",
          9110 => x"70",
          9111 => x"ff",
          9112 => x"83",
          9113 => x"78",
          9114 => x"89",
          9115 => x"81",
          9116 => x"06",
          9117 => x"80",
          9118 => x"77",
          9119 => x"74",
          9120 => x"8d",
          9121 => x"06",
          9122 => x"2e",
          9123 => x"77",
          9124 => x"93",
          9125 => x"74",
          9126 => x"cb",
          9127 => x"7d",
          9128 => x"81",
          9129 => x"38",
          9130 => x"66",
          9131 => x"81",
          9132 => x"b4",
          9133 => x"74",
          9134 => x"38",
          9135 => x"98",
          9136 => x"b4",
          9137 => x"82",
          9138 => x"57",
          9139 => x"80",
          9140 => x"76",
          9141 => x"38",
          9142 => x"51",
          9143 => x"3f",
          9144 => x"08",
          9145 => x"87",
          9146 => x"2a",
          9147 => x"5c",
          9148 => x"d4",
          9149 => x"80",
          9150 => x"44",
          9151 => x"0a",
          9152 => x"ec",
          9153 => x"39",
          9154 => x"66",
          9155 => x"81",
          9156 => x"a4",
          9157 => x"74",
          9158 => x"38",
          9159 => x"98",
          9160 => x"a4",
          9161 => x"82",
          9162 => x"57",
          9163 => x"80",
          9164 => x"76",
          9165 => x"38",
          9166 => x"51",
          9167 => x"3f",
          9168 => x"08",
          9169 => x"57",
          9170 => x"08",
          9171 => x"96",
          9172 => x"82",
          9173 => x"10",
          9174 => x"08",
          9175 => x"72",
          9176 => x"59",
          9177 => x"ff",
          9178 => x"5d",
          9179 => x"44",
          9180 => x"11",
          9181 => x"70",
          9182 => x"71",
          9183 => x"06",
          9184 => x"52",
          9185 => x"40",
          9186 => x"09",
          9187 => x"38",
          9188 => x"18",
          9189 => x"39",
          9190 => x"79",
          9191 => x"70",
          9192 => x"58",
          9193 => x"76",
          9194 => x"38",
          9195 => x"7d",
          9196 => x"70",
          9197 => x"55",
          9198 => x"3f",
          9199 => x"08",
          9200 => x"2e",
          9201 => x"9b",
          9202 => x"f8",
          9203 => x"f5",
          9204 => x"38",
          9205 => x"38",
          9206 => x"59",
          9207 => x"38",
          9208 => x"7d",
          9209 => x"81",
          9210 => x"38",
          9211 => x"0b",
          9212 => x"08",
          9213 => x"78",
          9214 => x"1a",
          9215 => x"c0",
          9216 => x"74",
          9217 => x"39",
          9218 => x"55",
          9219 => x"8f",
          9220 => x"fd",
          9221 => x"d4",
          9222 => x"f5",
          9223 => x"78",
          9224 => x"79",
          9225 => x"80",
          9226 => x"f1",
          9227 => x"39",
          9228 => x"81",
          9229 => x"06",
          9230 => x"55",
          9231 => x"27",
          9232 => x"81",
          9233 => x"56",
          9234 => x"38",
          9235 => x"80",
          9236 => x"ff",
          9237 => x"8b",
          9238 => x"bc",
          9239 => x"ff",
          9240 => x"84",
          9241 => x"1b",
          9242 => x"e1",
          9243 => x"1c",
          9244 => x"ff",
          9245 => x"8e",
          9246 => x"8f",
          9247 => x"0b",
          9248 => x"7d",
          9249 => x"30",
          9250 => x"84",
          9251 => x"51",
          9252 => x"51",
          9253 => x"3f",
          9254 => x"83",
          9255 => x"90",
          9256 => x"ff",
          9257 => x"93",
          9258 => x"8f",
          9259 => x"39",
          9260 => x"1b",
          9261 => x"b3",
          9262 => x"95",
          9263 => x"52",
          9264 => x"ff",
          9265 => x"81",
          9266 => x"1b",
          9267 => x"fd",
          9268 => x"9c",
          9269 => x"8f",
          9270 => x"83",
          9271 => x"06",
          9272 => x"82",
          9273 => x"52",
          9274 => x"51",
          9275 => x"3f",
          9276 => x"1b",
          9277 => x"f3",
          9278 => x"ac",
          9279 => x"8e",
          9280 => x"52",
          9281 => x"ff",
          9282 => x"86",
          9283 => x"51",
          9284 => x"3f",
          9285 => x"80",
          9286 => x"a9",
          9287 => x"1c",
          9288 => x"82",
          9289 => x"80",
          9290 => x"ae",
          9291 => x"b2",
          9292 => x"1b",
          9293 => x"b3",
          9294 => x"ff",
          9295 => x"96",
          9296 => x"8e",
          9297 => x"80",
          9298 => x"34",
          9299 => x"1c",
          9300 => x"82",
          9301 => x"ab",
          9302 => x"8e",
          9303 => x"d4",
          9304 => x"fe",
          9305 => x"59",
          9306 => x"3f",
          9307 => x"53",
          9308 => x"51",
          9309 => x"3f",
          9310 => x"d4",
          9311 => x"e7",
          9312 => x"2e",
          9313 => x"80",
          9314 => x"54",
          9315 => x"53",
          9316 => x"51",
          9317 => x"3f",
          9318 => x"80",
          9319 => x"ff",
          9320 => x"84",
          9321 => x"d2",
          9322 => x"ff",
          9323 => x"86",
          9324 => x"f2",
          9325 => x"1b",
          9326 => x"af",
          9327 => x"52",
          9328 => x"51",
          9329 => x"3f",
          9330 => x"ec",
          9331 => x"8d",
          9332 => x"d4",
          9333 => x"51",
          9334 => x"3f",
          9335 => x"87",
          9336 => x"52",
          9337 => x"89",
          9338 => x"54",
          9339 => x"7a",
          9340 => x"ff",
          9341 => x"65",
          9342 => x"7a",
          9343 => x"bd",
          9344 => x"80",
          9345 => x"2e",
          9346 => x"9a",
          9347 => x"7a",
          9348 => x"d7",
          9349 => x"84",
          9350 => x"8c",
          9351 => x"0a",
          9352 => x"51",
          9353 => x"ff",
          9354 => x"7d",
          9355 => x"38",
          9356 => x"52",
          9357 => x"8c",
          9358 => x"55",
          9359 => x"62",
          9360 => x"74",
          9361 => x"75",
          9362 => x"7e",
          9363 => x"ac",
          9364 => x"f8",
          9365 => x"38",
          9366 => x"82",
          9367 => x"52",
          9368 => x"8c",
          9369 => x"16",
          9370 => x"56",
          9371 => x"38",
          9372 => x"77",
          9373 => x"8d",
          9374 => x"7d",
          9375 => x"38",
          9376 => x"57",
          9377 => x"83",
          9378 => x"76",
          9379 => x"7a",
          9380 => x"ff",
          9381 => x"82",
          9382 => x"81",
          9383 => x"16",
          9384 => x"56",
          9385 => x"38",
          9386 => x"83",
          9387 => x"86",
          9388 => x"ff",
          9389 => x"38",
          9390 => x"82",
          9391 => x"81",
          9392 => x"06",
          9393 => x"fe",
          9394 => x"53",
          9395 => x"51",
          9396 => x"3f",
          9397 => x"52",
          9398 => x"8a",
          9399 => x"be",
          9400 => x"75",
          9401 => x"81",
          9402 => x"0b",
          9403 => x"77",
          9404 => x"75",
          9405 => x"60",
          9406 => x"80",
          9407 => x"75",
          9408 => x"aa",
          9409 => x"85",
          9410 => x"d4",
          9411 => x"2a",
          9412 => x"75",
          9413 => x"82",
          9414 => x"87",
          9415 => x"52",
          9416 => x"51",
          9417 => x"3f",
          9418 => x"ca",
          9419 => x"8a",
          9420 => x"54",
          9421 => x"52",
          9422 => x"86",
          9423 => x"56",
          9424 => x"08",
          9425 => x"53",
          9426 => x"51",
          9427 => x"3f",
          9428 => x"d4",
          9429 => x"38",
          9430 => x"56",
          9431 => x"56",
          9432 => x"d4",
          9433 => x"75",
          9434 => x"0c",
          9435 => x"04",
          9436 => x"7d",
          9437 => x"80",
          9438 => x"05",
          9439 => x"76",
          9440 => x"38",
          9441 => x"11",
          9442 => x"53",
          9443 => x"79",
          9444 => x"3f",
          9445 => x"09",
          9446 => x"38",
          9447 => x"55",
          9448 => x"db",
          9449 => x"70",
          9450 => x"34",
          9451 => x"74",
          9452 => x"81",
          9453 => x"80",
          9454 => x"55",
          9455 => x"76",
          9456 => x"d4",
          9457 => x"3d",
          9458 => x"3d",
          9459 => x"84",
          9460 => x"33",
          9461 => x"8a",
          9462 => x"06",
          9463 => x"52",
          9464 => x"3f",
          9465 => x"56",
          9466 => x"be",
          9467 => x"08",
          9468 => x"05",
          9469 => x"75",
          9470 => x"56",
          9471 => x"a1",
          9472 => x"fc",
          9473 => x"53",
          9474 => x"76",
          9475 => x"c0",
          9476 => x"32",
          9477 => x"72",
          9478 => x"70",
          9479 => x"56",
          9480 => x"18",
          9481 => x"88",
          9482 => x"3d",
          9483 => x"3d",
          9484 => x"11",
          9485 => x"80",
          9486 => x"38",
          9487 => x"05",
          9488 => x"8c",
          9489 => x"08",
          9490 => x"3f",
          9491 => x"08",
          9492 => x"16",
          9493 => x"09",
          9494 => x"38",
          9495 => x"55",
          9496 => x"55",
          9497 => x"f8",
          9498 => x"0d",
          9499 => x"0d",
          9500 => x"cc",
          9501 => x"73",
          9502 => x"c1",
          9503 => x"0c",
          9504 => x"04",
          9505 => x"02",
          9506 => x"33",
          9507 => x"3d",
          9508 => x"54",
          9509 => x"52",
          9510 => x"ae",
          9511 => x"ff",
          9512 => x"3d",
          9513 => x"3d",
          9514 => x"84",
          9515 => x"22",
          9516 => x"52",
          9517 => x"26",
          9518 => x"83",
          9519 => x"52",
          9520 => x"83",
          9521 => x"27",
          9522 => x"b5",
          9523 => x"06",
          9524 => x"80",
          9525 => x"82",
          9526 => x"51",
          9527 => x"9c",
          9528 => x"70",
          9529 => x"06",
          9530 => x"80",
          9531 => x"38",
          9532 => x"c8",
          9533 => x"22",
          9534 => x"39",
          9535 => x"70",
          9536 => x"53",
          9537 => x"d4",
          9538 => x"3d",
          9539 => x"3d",
          9540 => x"05",
          9541 => x"05",
          9542 => x"53",
          9543 => x"70",
          9544 => x"85",
          9545 => x"9a",
          9546 => x"b5",
          9547 => x"06",
          9548 => x"81",
          9549 => x"38",
          9550 => x"c6",
          9551 => x"22",
          9552 => x"82",
          9553 => x"84",
          9554 => x"fb",
          9555 => x"51",
          9556 => x"ff",
          9557 => x"38",
          9558 => x"ff",
          9559 => x"c4",
          9560 => x"ff",
          9561 => x"38",
          9562 => x"56",
          9563 => x"05",
          9564 => x"30",
          9565 => x"72",
          9566 => x"51",
          9567 => x"80",
          9568 => x"70",
          9569 => x"22",
          9570 => x"71",
          9571 => x"70",
          9572 => x"55",
          9573 => x"25",
          9574 => x"73",
          9575 => x"dc",
          9576 => x"29",
          9577 => x"05",
          9578 => x"04",
          9579 => x"10",
          9580 => x"22",
          9581 => x"80",
          9582 => x"75",
          9583 => x"72",
          9584 => x"51",
          9585 => x"12",
          9586 => x"e0",
          9587 => x"39",
          9588 => x"95",
          9589 => x"51",
          9590 => x"12",
          9591 => x"ff",
          9592 => x"85",
          9593 => x"12",
          9594 => x"ff",
          9595 => x"8c",
          9596 => x"f8",
          9597 => x"16",
          9598 => x"39",
          9599 => x"82",
          9600 => x"87",
          9601 => x"00",
          9602 => x"ff",
          9603 => x"ff",
          9604 => x"ff",
          9605 => x"00",
          9606 => x"51",
          9607 => x"d5",
          9608 => x"dc",
          9609 => x"e3",
          9610 => x"ea",
          9611 => x"f1",
          9612 => x"f8",
          9613 => x"ff",
          9614 => x"06",
          9615 => x"0d",
          9616 => x"14",
          9617 => x"1b",
          9618 => x"21",
          9619 => x"27",
          9620 => x"2d",
          9621 => x"33",
          9622 => x"39",
          9623 => x"3f",
          9624 => x"45",
          9625 => x"4b",
          9626 => x"8a",
          9627 => x"90",
          9628 => x"96",
          9629 => x"9c",
          9630 => x"a2",
          9631 => x"80",
          9632 => x"80",
          9633 => x"91",
          9634 => x"e9",
          9635 => x"68",
          9636 => x"55",
          9637 => x"59",
          9638 => x"ba",
          9639 => x"9c",
          9640 => x"32",
          9641 => x"b8",
          9642 => x"3b",
          9643 => x"55",
          9644 => x"91",
          9645 => x"ba",
          9646 => x"59",
          9647 => x"55",
          9648 => x"55",
          9649 => x"b8",
          9650 => x"32",
          9651 => x"ba",
          9652 => x"e9",
          9653 => x"ac",
          9654 => x"ba",
          9655 => x"c6",
          9656 => x"cb",
          9657 => x"d0",
          9658 => x"d5",
          9659 => x"da",
          9660 => x"df",
          9661 => x"e5",
          9662 => x"31",
          9663 => x"1a",
          9664 => x"1a",
          9665 => x"60",
          9666 => x"1a",
          9667 => x"1a",
          9668 => x"1a",
          9669 => x"1a",
          9670 => x"1a",
          9671 => x"1a",
          9672 => x"1a",
          9673 => x"1d",
          9674 => x"1a",
          9675 => x"48",
          9676 => x"78",
          9677 => x"1a",
          9678 => x"1a",
          9679 => x"1a",
          9680 => x"1a",
          9681 => x"1a",
          9682 => x"1a",
          9683 => x"1a",
          9684 => x"1a",
          9685 => x"1a",
          9686 => x"1a",
          9687 => x"1a",
          9688 => x"1a",
          9689 => x"1a",
          9690 => x"1a",
          9691 => x"1a",
          9692 => x"1a",
          9693 => x"1a",
          9694 => x"1a",
          9695 => x"1a",
          9696 => x"1a",
          9697 => x"1a",
          9698 => x"1a",
          9699 => x"1a",
          9700 => x"1a",
          9701 => x"1a",
          9702 => x"1a",
          9703 => x"1a",
          9704 => x"1a",
          9705 => x"1a",
          9706 => x"1a",
          9707 => x"1a",
          9708 => x"1a",
          9709 => x"1a",
          9710 => x"1a",
          9711 => x"1a",
          9712 => x"1a",
          9713 => x"a8",
          9714 => x"1a",
          9715 => x"1a",
          9716 => x"1a",
          9717 => x"1a",
          9718 => x"16",
          9719 => x"1a",
          9720 => x"1a",
          9721 => x"1a",
          9722 => x"1a",
          9723 => x"1a",
          9724 => x"1a",
          9725 => x"1a",
          9726 => x"1a",
          9727 => x"1a",
          9728 => x"1a",
          9729 => x"d8",
          9730 => x"3f",
          9731 => x"af",
          9732 => x"af",
          9733 => x"af",
          9734 => x"1a",
          9735 => x"3f",
          9736 => x"1a",
          9737 => x"1a",
          9738 => x"98",
          9739 => x"1a",
          9740 => x"1a",
          9741 => x"ec",
          9742 => x"f7",
          9743 => x"1a",
          9744 => x"1a",
          9745 => x"11",
          9746 => x"1a",
          9747 => x"1f",
          9748 => x"1a",
          9749 => x"1a",
          9750 => x"16",
          9751 => x"69",
          9752 => x"00",
          9753 => x"63",
          9754 => x"00",
          9755 => x"69",
          9756 => x"00",
          9757 => x"61",
          9758 => x"00",
          9759 => x"65",
          9760 => x"00",
          9761 => x"65",
          9762 => x"00",
          9763 => x"70",
          9764 => x"00",
          9765 => x"66",
          9766 => x"00",
          9767 => x"6d",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"00",
          9776 => x"6c",
          9777 => x"00",
          9778 => x"00",
          9779 => x"74",
          9780 => x"00",
          9781 => x"65",
          9782 => x"00",
          9783 => x"6f",
          9784 => x"00",
          9785 => x"74",
          9786 => x"00",
          9787 => x"73",
          9788 => x"00",
          9789 => x"73",
          9790 => x"00",
          9791 => x"6f",
          9792 => x"00",
          9793 => x"00",
          9794 => x"6b",
          9795 => x"72",
          9796 => x"00",
          9797 => x"65",
          9798 => x"6c",
          9799 => x"72",
          9800 => x"00",
          9801 => x"6b",
          9802 => x"74",
          9803 => x"61",
          9804 => x"00",
          9805 => x"66",
          9806 => x"20",
          9807 => x"6e",
          9808 => x"00",
          9809 => x"70",
          9810 => x"20",
          9811 => x"6e",
          9812 => x"00",
          9813 => x"61",
          9814 => x"20",
          9815 => x"65",
          9816 => x"65",
          9817 => x"00",
          9818 => x"65",
          9819 => x"64",
          9820 => x"65",
          9821 => x"00",
          9822 => x"65",
          9823 => x"72",
          9824 => x"79",
          9825 => x"69",
          9826 => x"2e",
          9827 => x"00",
          9828 => x"65",
          9829 => x"6e",
          9830 => x"20",
          9831 => x"61",
          9832 => x"2e",
          9833 => x"00",
          9834 => x"69",
          9835 => x"72",
          9836 => x"20",
          9837 => x"74",
          9838 => x"65",
          9839 => x"00",
          9840 => x"76",
          9841 => x"75",
          9842 => x"72",
          9843 => x"20",
          9844 => x"61",
          9845 => x"2e",
          9846 => x"00",
          9847 => x"6b",
          9848 => x"74",
          9849 => x"61",
          9850 => x"64",
          9851 => x"00",
          9852 => x"63",
          9853 => x"61",
          9854 => x"6c",
          9855 => x"69",
          9856 => x"79",
          9857 => x"6d",
          9858 => x"75",
          9859 => x"6f",
          9860 => x"69",
          9861 => x"00",
          9862 => x"6d",
          9863 => x"61",
          9864 => x"74",
          9865 => x"00",
          9866 => x"65",
          9867 => x"2c",
          9868 => x"65",
          9869 => x"69",
          9870 => x"63",
          9871 => x"65",
          9872 => x"64",
          9873 => x"00",
          9874 => x"65",
          9875 => x"20",
          9876 => x"6b",
          9877 => x"00",
          9878 => x"75",
          9879 => x"63",
          9880 => x"74",
          9881 => x"6d",
          9882 => x"2e",
          9883 => x"00",
          9884 => x"20",
          9885 => x"79",
          9886 => x"65",
          9887 => x"69",
          9888 => x"2e",
          9889 => x"00",
          9890 => x"61",
          9891 => x"65",
          9892 => x"69",
          9893 => x"72",
          9894 => x"74",
          9895 => x"00",
          9896 => x"63",
          9897 => x"2e",
          9898 => x"00",
          9899 => x"6e",
          9900 => x"20",
          9901 => x"6f",
          9902 => x"00",
          9903 => x"75",
          9904 => x"74",
          9905 => x"25",
          9906 => x"74",
          9907 => x"75",
          9908 => x"74",
          9909 => x"73",
          9910 => x"0a",
          9911 => x"00",
          9912 => x"64",
          9913 => x"00",
          9914 => x"30",
          9915 => x"2c",
          9916 => x"25",
          9917 => x"78",
          9918 => x"3d",
          9919 => x"6c",
          9920 => x"5f",
          9921 => x"3d",
          9922 => x"6c",
          9923 => x"30",
          9924 => x"20",
          9925 => x"6c",
          9926 => x"00",
          9927 => x"6c",
          9928 => x"00",
          9929 => x"00",
          9930 => x"58",
          9931 => x"00",
          9932 => x"20",
          9933 => x"20",
          9934 => x"00",
          9935 => x"58",
          9936 => x"00",
          9937 => x"00",
          9938 => x"00",
          9939 => x"00",
          9940 => x"00",
          9941 => x"20",
          9942 => x"28",
          9943 => x"00",
          9944 => x"31",
          9945 => x"30",
          9946 => x"00",
          9947 => x"30",
          9948 => x"00",
          9949 => x"55",
          9950 => x"65",
          9951 => x"30",
          9952 => x"20",
          9953 => x"25",
          9954 => x"2a",
          9955 => x"00",
          9956 => x"20",
          9957 => x"65",
          9958 => x"70",
          9959 => x"61",
          9960 => x"65",
          9961 => x"00",
          9962 => x"65",
          9963 => x"6e",
          9964 => x"72",
          9965 => x"00",
          9966 => x"20",
          9967 => x"65",
          9968 => x"70",
          9969 => x"00",
          9970 => x"54",
          9971 => x"44",
          9972 => x"74",
          9973 => x"75",
          9974 => x"00",
          9975 => x"54",
          9976 => x"52",
          9977 => x"74",
          9978 => x"75",
          9979 => x"00",
          9980 => x"54",
          9981 => x"58",
          9982 => x"74",
          9983 => x"75",
          9984 => x"00",
          9985 => x"54",
          9986 => x"58",
          9987 => x"74",
          9988 => x"75",
          9989 => x"00",
          9990 => x"54",
          9991 => x"58",
          9992 => x"74",
          9993 => x"75",
          9994 => x"00",
          9995 => x"54",
          9996 => x"58",
          9997 => x"74",
          9998 => x"75",
          9999 => x"00",
         10000 => x"74",
         10001 => x"20",
         10002 => x"74",
         10003 => x"72",
         10004 => x"00",
         10005 => x"62",
         10006 => x"67",
         10007 => x"6d",
         10008 => x"2e",
         10009 => x"00",
         10010 => x"6f",
         10011 => x"63",
         10012 => x"74",
         10013 => x"00",
         10014 => x"2e",
         10015 => x"00",
         10016 => x"00",
         10017 => x"6c",
         10018 => x"74",
         10019 => x"6e",
         10020 => x"61",
         10021 => x"65",
         10022 => x"20",
         10023 => x"64",
         10024 => x"20",
         10025 => x"61",
         10026 => x"69",
         10027 => x"20",
         10028 => x"75",
         10029 => x"79",
         10030 => x"00",
         10031 => x"00",
         10032 => x"61",
         10033 => x"67",
         10034 => x"2e",
         10035 => x"00",
         10036 => x"79",
         10037 => x"2e",
         10038 => x"00",
         10039 => x"70",
         10040 => x"6e",
         10041 => x"2e",
         10042 => x"00",
         10043 => x"6c",
         10044 => x"30",
         10045 => x"2d",
         10046 => x"38",
         10047 => x"25",
         10048 => x"29",
         10049 => x"00",
         10050 => x"70",
         10051 => x"6d",
         10052 => x"00",
         10053 => x"6d",
         10054 => x"74",
         10055 => x"00",
         10056 => x"6c",
         10057 => x"30",
         10058 => x"00",
         10059 => x"00",
         10060 => x"6c",
         10061 => x"30",
         10062 => x"00",
         10063 => x"6c",
         10064 => x"30",
         10065 => x"2d",
         10066 => x"00",
         10067 => x"63",
         10068 => x"6e",
         10069 => x"6f",
         10070 => x"40",
         10071 => x"38",
         10072 => x"2e",
         10073 => x"00",
         10074 => x"6c",
         10075 => x"20",
         10076 => x"65",
         10077 => x"25",
         10078 => x"78",
         10079 => x"2e",
         10080 => x"00",
         10081 => x"6c",
         10082 => x"74",
         10083 => x"65",
         10084 => x"6f",
         10085 => x"28",
         10086 => x"2e",
         10087 => x"00",
         10088 => x"74",
         10089 => x"69",
         10090 => x"61",
         10091 => x"69",
         10092 => x"69",
         10093 => x"2e",
         10094 => x"00",
         10095 => x"64",
         10096 => x"62",
         10097 => x"69",
         10098 => x"2e",
         10099 => x"00",
         10100 => x"00",
         10101 => x"00",
         10102 => x"5c",
         10103 => x"25",
         10104 => x"73",
         10105 => x"00",
         10106 => x"5c",
         10107 => x"25",
         10108 => x"00",
         10109 => x"5c",
         10110 => x"00",
         10111 => x"20",
         10112 => x"6d",
         10113 => x"2e",
         10114 => x"00",
         10115 => x"6f",
         10116 => x"65",
         10117 => x"75",
         10118 => x"64",
         10119 => x"61",
         10120 => x"74",
         10121 => x"6f",
         10122 => x"73",
         10123 => x"6d",
         10124 => x"64",
         10125 => x"00",
         10126 => x"6e",
         10127 => x"2e",
         10128 => x"00",
         10129 => x"62",
         10130 => x"67",
         10131 => x"74",
         10132 => x"75",
         10133 => x"2e",
         10134 => x"00",
         10135 => x"25",
         10136 => x"64",
         10137 => x"3a",
         10138 => x"25",
         10139 => x"64",
         10140 => x"00",
         10141 => x"20",
         10142 => x"66",
         10143 => x"72",
         10144 => x"6f",
         10145 => x"00",
         10146 => x"72",
         10147 => x"53",
         10148 => x"63",
         10149 => x"69",
         10150 => x"00",
         10151 => x"65",
         10152 => x"65",
         10153 => x"6d",
         10154 => x"6d",
         10155 => x"65",
         10156 => x"00",
         10157 => x"20",
         10158 => x"53",
         10159 => x"4d",
         10160 => x"25",
         10161 => x"3a",
         10162 => x"58",
         10163 => x"00",
         10164 => x"20",
         10165 => x"41",
         10166 => x"20",
         10167 => x"25",
         10168 => x"3a",
         10169 => x"58",
         10170 => x"00",
         10171 => x"20",
         10172 => x"4e",
         10173 => x"41",
         10174 => x"25",
         10175 => x"3a",
         10176 => x"58",
         10177 => x"00",
         10178 => x"20",
         10179 => x"4d",
         10180 => x"20",
         10181 => x"25",
         10182 => x"3a",
         10183 => x"58",
         10184 => x"00",
         10185 => x"20",
         10186 => x"20",
         10187 => x"20",
         10188 => x"25",
         10189 => x"3a",
         10190 => x"58",
         10191 => x"00",
         10192 => x"20",
         10193 => x"43",
         10194 => x"20",
         10195 => x"44",
         10196 => x"63",
         10197 => x"3d",
         10198 => x"64",
         10199 => x"00",
         10200 => x"20",
         10201 => x"45",
         10202 => x"20",
         10203 => x"54",
         10204 => x"72",
         10205 => x"3d",
         10206 => x"64",
         10207 => x"00",
         10208 => x"20",
         10209 => x"52",
         10210 => x"52",
         10211 => x"43",
         10212 => x"6e",
         10213 => x"3d",
         10214 => x"64",
         10215 => x"00",
         10216 => x"20",
         10217 => x"48",
         10218 => x"45",
         10219 => x"53",
         10220 => x"00",
         10221 => x"20",
         10222 => x"49",
         10223 => x"00",
         10224 => x"20",
         10225 => x"54",
         10226 => x"00",
         10227 => x"20",
         10228 => x"00",
         10229 => x"20",
         10230 => x"00",
         10231 => x"72",
         10232 => x"65",
         10233 => x"00",
         10234 => x"20",
         10235 => x"20",
         10236 => x"65",
         10237 => x"65",
         10238 => x"72",
         10239 => x"64",
         10240 => x"73",
         10241 => x"25",
         10242 => x"0a",
         10243 => x"00",
         10244 => x"20",
         10245 => x"20",
         10246 => x"6f",
         10247 => x"53",
         10248 => x"74",
         10249 => x"64",
         10250 => x"73",
         10251 => x"25",
         10252 => x"0a",
         10253 => x"00",
         10254 => x"20",
         10255 => x"63",
         10256 => x"74",
         10257 => x"20",
         10258 => x"72",
         10259 => x"20",
         10260 => x"20",
         10261 => x"25",
         10262 => x"0a",
         10263 => x"00",
         10264 => x"63",
         10265 => x"00",
         10266 => x"20",
         10267 => x"20",
         10268 => x"20",
         10269 => x"20",
         10270 => x"20",
         10271 => x"20",
         10272 => x"20",
         10273 => x"25",
         10274 => x"0a",
         10275 => x"00",
         10276 => x"20",
         10277 => x"74",
         10278 => x"43",
         10279 => x"6b",
         10280 => x"65",
         10281 => x"20",
         10282 => x"20",
         10283 => x"25",
         10284 => x"30",
         10285 => x"48",
         10286 => x"00",
         10287 => x"20",
         10288 => x"41",
         10289 => x"6c",
         10290 => x"20",
         10291 => x"71",
         10292 => x"20",
         10293 => x"20",
         10294 => x"25",
         10295 => x"30",
         10296 => x"48",
         10297 => x"00",
         10298 => x"20",
         10299 => x"68",
         10300 => x"65",
         10301 => x"52",
         10302 => x"43",
         10303 => x"6b",
         10304 => x"65",
         10305 => x"25",
         10306 => x"30",
         10307 => x"48",
         10308 => x"00",
         10309 => x"6c",
         10310 => x"00",
         10311 => x"69",
         10312 => x"00",
         10313 => x"78",
         10314 => x"00",
         10315 => x"00",
         10316 => x"6d",
         10317 => x"00",
         10318 => x"6e",
         10319 => x"00",
         10320 => x"9c",
         10321 => x"00",
         10322 => x"02",
         10323 => x"98",
         10324 => x"00",
         10325 => x"03",
         10326 => x"94",
         10327 => x"00",
         10328 => x"04",
         10329 => x"90",
         10330 => x"00",
         10331 => x"05",
         10332 => x"8c",
         10333 => x"00",
         10334 => x"06",
         10335 => x"88",
         10336 => x"00",
         10337 => x"07",
         10338 => x"84",
         10339 => x"00",
         10340 => x"01",
         10341 => x"80",
         10342 => x"00",
         10343 => x"08",
         10344 => x"7c",
         10345 => x"00",
         10346 => x"0b",
         10347 => x"78",
         10348 => x"00",
         10349 => x"09",
         10350 => x"74",
         10351 => x"00",
         10352 => x"0a",
         10353 => x"70",
         10354 => x"00",
         10355 => x"0d",
         10356 => x"6c",
         10357 => x"00",
         10358 => x"0c",
         10359 => x"68",
         10360 => x"00",
         10361 => x"0e",
         10362 => x"64",
         10363 => x"00",
         10364 => x"0f",
         10365 => x"60",
         10366 => x"00",
         10367 => x"0f",
         10368 => x"5c",
         10369 => x"00",
         10370 => x"10",
         10371 => x"58",
         10372 => x"00",
         10373 => x"11",
         10374 => x"54",
         10375 => x"00",
         10376 => x"12",
         10377 => x"50",
         10378 => x"00",
         10379 => x"13",
         10380 => x"4c",
         10381 => x"00",
         10382 => x"14",
         10383 => x"48",
         10384 => x"00",
         10385 => x"15",
         10386 => x"00",
         10387 => x"00",
         10388 => x"00",
         10389 => x"00",
         10390 => x"7e",
         10391 => x"7e",
         10392 => x"7e",
         10393 => x"00",
         10394 => x"7e",
         10395 => x"7e",
         10396 => x"7e",
         10397 => x"00",
         10398 => x"00",
         10399 => x"00",
         10400 => x"00",
         10401 => x"00",
         10402 => x"00",
         10403 => x"00",
         10404 => x"00",
         10405 => x"00",
         10406 => x"00",
         10407 => x"00",
         10408 => x"74",
         10409 => x"00",
         10410 => x"74",
         10411 => x"00",
         10412 => x"00",
         10413 => x"6c",
         10414 => x"25",
         10415 => x"00",
         10416 => x"6c",
         10417 => x"74",
         10418 => x"65",
         10419 => x"20",
         10420 => x"20",
         10421 => x"74",
         10422 => x"20",
         10423 => x"65",
         10424 => x"20",
         10425 => x"2e",
         10426 => x"00",
         10427 => x"6e",
         10428 => x"6f",
         10429 => x"2f",
         10430 => x"61",
         10431 => x"68",
         10432 => x"6f",
         10433 => x"66",
         10434 => x"2c",
         10435 => x"73",
         10436 => x"69",
         10437 => x"00",
         10438 => x"00",
         10439 => x"3c",
         10440 => x"7f",
         10441 => x"00",
         10442 => x"3d",
         10443 => x"00",
         10444 => x"00",
         10445 => x"33",
         10446 => x"00",
         10447 => x"4d",
         10448 => x"53",
         10449 => x"00",
         10450 => x"4e",
         10451 => x"20",
         10452 => x"46",
         10453 => x"32",
         10454 => x"00",
         10455 => x"4e",
         10456 => x"20",
         10457 => x"46",
         10458 => x"20",
         10459 => x"00",
         10460 => x"18",
         10461 => x"00",
         10462 => x"00",
         10463 => x"00",
         10464 => x"07",
         10465 => x"12",
         10466 => x"1c",
         10467 => x"00",
         10468 => x"41",
         10469 => x"80",
         10470 => x"49",
         10471 => x"8f",
         10472 => x"4f",
         10473 => x"55",
         10474 => x"9b",
         10475 => x"9f",
         10476 => x"55",
         10477 => x"a7",
         10478 => x"ab",
         10479 => x"af",
         10480 => x"b3",
         10481 => x"b7",
         10482 => x"bb",
         10483 => x"bf",
         10484 => x"c3",
         10485 => x"c7",
         10486 => x"cb",
         10487 => x"cf",
         10488 => x"d3",
         10489 => x"d7",
         10490 => x"db",
         10491 => x"df",
         10492 => x"e3",
         10493 => x"e7",
         10494 => x"eb",
         10495 => x"ef",
         10496 => x"f3",
         10497 => x"f7",
         10498 => x"fb",
         10499 => x"ff",
         10500 => x"3b",
         10501 => x"2f",
         10502 => x"3a",
         10503 => x"7c",
         10504 => x"00",
         10505 => x"04",
         10506 => x"40",
         10507 => x"00",
         10508 => x"00",
         10509 => x"02",
         10510 => x"08",
         10511 => x"20",
         10512 => x"00",
         10513 => x"fc",
         10514 => x"e2",
         10515 => x"e0",
         10516 => x"e7",
         10517 => x"eb",
         10518 => x"ef",
         10519 => x"ec",
         10520 => x"c5",
         10521 => x"e6",
         10522 => x"f4",
         10523 => x"f2",
         10524 => x"f9",
         10525 => x"d6",
         10526 => x"a2",
         10527 => x"a5",
         10528 => x"92",
         10529 => x"ed",
         10530 => x"fa",
         10531 => x"d1",
         10532 => x"ba",
         10533 => x"10",
         10534 => x"bd",
         10535 => x"a1",
         10536 => x"bb",
         10537 => x"92",
         10538 => x"02",
         10539 => x"61",
         10540 => x"56",
         10541 => x"63",
         10542 => x"57",
         10543 => x"5c",
         10544 => x"10",
         10545 => x"34",
         10546 => x"1c",
         10547 => x"3c",
         10548 => x"5f",
         10549 => x"54",
         10550 => x"66",
         10551 => x"50",
         10552 => x"67",
         10553 => x"64",
         10554 => x"59",
         10555 => x"52",
         10556 => x"6b",
         10557 => x"18",
         10558 => x"88",
         10559 => x"8c",
         10560 => x"80",
         10561 => x"df",
         10562 => x"c0",
         10563 => x"c3",
         10564 => x"c4",
         10565 => x"98",
         10566 => x"b4",
         10567 => x"c6",
         10568 => x"29",
         10569 => x"b1",
         10570 => x"64",
         10571 => x"21",
         10572 => x"48",
         10573 => x"19",
         10574 => x"1a",
         10575 => x"b2",
         10576 => x"a0",
         10577 => x"1a",
         10578 => x"17",
         10579 => x"07",
         10580 => x"01",
         10581 => x"00",
         10582 => x"32",
         10583 => x"39",
         10584 => x"4a",
         10585 => x"79",
         10586 => x"80",
         10587 => x"43",
         10588 => x"82",
         10589 => x"84",
         10590 => x"86",
         10591 => x"87",
         10592 => x"8a",
         10593 => x"8b",
         10594 => x"8e",
         10595 => x"90",
         10596 => x"91",
         10597 => x"94",
         10598 => x"96",
         10599 => x"98",
         10600 => x"3d",
         10601 => x"9c",
         10602 => x"20",
         10603 => x"a0",
         10604 => x"a2",
         10605 => x"a4",
         10606 => x"a6",
         10607 => x"a7",
         10608 => x"aa",
         10609 => x"ac",
         10610 => x"ae",
         10611 => x"af",
         10612 => x"b2",
         10613 => x"b3",
         10614 => x"b5",
         10615 => x"b8",
         10616 => x"ba",
         10617 => x"bc",
         10618 => x"be",
         10619 => x"c0",
         10620 => x"c2",
         10621 => x"c4",
         10622 => x"c4",
         10623 => x"c8",
         10624 => x"ca",
         10625 => x"ca",
         10626 => x"10",
         10627 => x"01",
         10628 => x"de",
         10629 => x"f3",
         10630 => x"f1",
         10631 => x"f4",
         10632 => x"28",
         10633 => x"12",
         10634 => x"09",
         10635 => x"3b",
         10636 => x"3d",
         10637 => x"3f",
         10638 => x"41",
         10639 => x"46",
         10640 => x"53",
         10641 => x"81",
         10642 => x"55",
         10643 => x"8a",
         10644 => x"8f",
         10645 => x"90",
         10646 => x"5d",
         10647 => x"5f",
         10648 => x"61",
         10649 => x"94",
         10650 => x"65",
         10651 => x"67",
         10652 => x"96",
         10653 => x"62",
         10654 => x"6d",
         10655 => x"9c",
         10656 => x"71",
         10657 => x"73",
         10658 => x"9f",
         10659 => x"77",
         10660 => x"79",
         10661 => x"7b",
         10662 => x"64",
         10663 => x"7f",
         10664 => x"81",
         10665 => x"a9",
         10666 => x"85",
         10667 => x"87",
         10668 => x"44",
         10669 => x"b2",
         10670 => x"8d",
         10671 => x"8f",
         10672 => x"91",
         10673 => x"7b",
         10674 => x"fd",
         10675 => x"ff",
         10676 => x"04",
         10677 => x"88",
         10678 => x"8a",
         10679 => x"11",
         10680 => x"02",
         10681 => x"a3",
         10682 => x"08",
         10683 => x"03",
         10684 => x"8e",
         10685 => x"d8",
         10686 => x"f2",
         10687 => x"f9",
         10688 => x"f4",
         10689 => x"f6",
         10690 => x"f7",
         10691 => x"fa",
         10692 => x"30",
         10693 => x"50",
         10694 => x"60",
         10695 => x"8a",
         10696 => x"c1",
         10697 => x"cf",
         10698 => x"c0",
         10699 => x"44",
         10700 => x"26",
         10701 => x"00",
         10702 => x"01",
         10703 => x"00",
         10704 => x"a0",
         10705 => x"00",
         10706 => x"10",
         10707 => x"20",
         10708 => x"30",
         10709 => x"40",
         10710 => x"51",
         10711 => x"59",
         10712 => x"5b",
         10713 => x"5d",
         10714 => x"5f",
         10715 => x"08",
         10716 => x"0e",
         10717 => x"bb",
         10718 => x"c9",
         10719 => x"cb",
         10720 => x"db",
         10721 => x"f9",
         10722 => x"eb",
         10723 => x"fb",
         10724 => x"08",
         10725 => x"08",
         10726 => x"08",
         10727 => x"04",
         10728 => x"b9",
         10729 => x"bc",
         10730 => x"01",
         10731 => x"d0",
         10732 => x"e0",
         10733 => x"e5",
         10734 => x"ec",
         10735 => x"01",
         10736 => x"4e",
         10737 => x"32",
         10738 => x"10",
         10739 => x"01",
         10740 => x"d0",
         10741 => x"30",
         10742 => x"60",
         10743 => x"67",
         10744 => x"75",
         10745 => x"80",
         10746 => x"00",
         10747 => x"41",
         10748 => x"00",
         10749 => x"00",
         10750 => x"5c",
         10751 => x"00",
         10752 => x"00",
         10753 => x"00",
         10754 => x"64",
         10755 => x"00",
         10756 => x"00",
         10757 => x"00",
         10758 => x"6c",
         10759 => x"00",
         10760 => x"00",
         10761 => x"00",
         10762 => x"74",
         10763 => x"00",
         10764 => x"00",
         10765 => x"00",
         10766 => x"7c",
         10767 => x"00",
         10768 => x"00",
         10769 => x"00",
         10770 => x"84",
         10771 => x"00",
         10772 => x"00",
         10773 => x"00",
         10774 => x"8c",
         10775 => x"00",
         10776 => x"00",
         10777 => x"00",
         10778 => x"94",
         10779 => x"00",
         10780 => x"00",
         10781 => x"00",
         10782 => x"9c",
         10783 => x"00",
         10784 => x"00",
         10785 => x"00",
         10786 => x"a4",
         10787 => x"00",
         10788 => x"00",
         10789 => x"00",
         10790 => x"a8",
         10791 => x"00",
         10792 => x"00",
         10793 => x"00",
         10794 => x"ac",
         10795 => x"00",
         10796 => x"00",
         10797 => x"00",
         10798 => x"b0",
         10799 => x"00",
         10800 => x"00",
         10801 => x"00",
         10802 => x"b4",
         10803 => x"00",
         10804 => x"00",
         10805 => x"00",
         10806 => x"b8",
         10807 => x"00",
         10808 => x"00",
         10809 => x"00",
         10810 => x"bc",
         10811 => x"00",
         10812 => x"00",
         10813 => x"00",
         10814 => x"c0",
         10815 => x"00",
         10816 => x"00",
         10817 => x"00",
         10818 => x"c8",
         10819 => x"00",
         10820 => x"00",
         10821 => x"00",
         10822 => x"cc",
         10823 => x"00",
         10824 => x"00",
         10825 => x"00",
         10826 => x"d4",
         10827 => x"00",
         10828 => x"00",
         10829 => x"00",
         10830 => x"dc",
         10831 => x"00",
         10832 => x"00",
         10833 => x"00",
         10834 => x"e4",
         10835 => x"00",
         10836 => x"00",
         10837 => x"00",
         10838 => x"ec",
         10839 => x"00",
         10840 => x"00",
         10841 => x"00",
         10842 => x"f4",
         10843 => x"00",
         10844 => x"00",
         10845 => x"00",
         10846 => x"fc",
         10847 => x"00",
         10848 => x"00",
         10849 => x"00",
         10850 => x"04",
         10851 => x"00",
         10852 => x"00",
         10853 => x"00",
         10854 => x"00",
         10855 => x"00",
         10856 => x"ff",
         10857 => x"00",
         10858 => x"ff",
         10859 => x"00",
         10860 => x"ff",
         10861 => x"00",
         10862 => x"00",
         10863 => x"00",
         10864 => x"ff",
         10865 => x"00",
         10866 => x"00",
         10867 => x"00",
         10868 => x"00",
         10869 => x"00",
         10870 => x"00",
         10871 => x"00",
         10872 => x"00",
         10873 => x"01",
         10874 => x"01",
         10875 => x"01",
         10876 => x"00",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"00",
         10884 => x"00",
         10885 => x"00",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"00",
         10890 => x"00",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"00",
         10895 => x"00",
         10896 => x"00",
         10897 => x"00",
         10898 => x"00",
         10899 => x"00",
         10900 => x"00",
         10901 => x"a0",
         10902 => x"00",
         10903 => x"a8",
         10904 => x"00",
         10905 => x"b0",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"0b",
             2 => x"b9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"82",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a4",
           270 => x"0b",
           271 => x"0b",
           272 => x"c2",
           273 => x"0b",
           274 => x"0b",
           275 => x"e0",
           276 => x"0b",
           277 => x"0b",
           278 => x"80",
           279 => x"0b",
           280 => x"0b",
           281 => x"9e",
           282 => x"0b",
           283 => x"0b",
           284 => x"bd",
           285 => x"0b",
           286 => x"0b",
           287 => x"dd",
           288 => x"0b",
           289 => x"0b",
           290 => x"fd",
           291 => x"0b",
           292 => x"0b",
           293 => x"9d",
           294 => x"0b",
           295 => x"0b",
           296 => x"bd",
           297 => x"0b",
           298 => x"0b",
           299 => x"dd",
           300 => x"0b",
           301 => x"0b",
           302 => x"fd",
           303 => x"0b",
           304 => x"0b",
           305 => x"9d",
           306 => x"0b",
           307 => x"0b",
           308 => x"bd",
           309 => x"0b",
           310 => x"0b",
           311 => x"dd",
           312 => x"0b",
           313 => x"0b",
           314 => x"fd",
           315 => x"0b",
           316 => x"0b",
           317 => x"9d",
           318 => x"0b",
           319 => x"0b",
           320 => x"bd",
           321 => x"0b",
           322 => x"0b",
           323 => x"dd",
           324 => x"0b",
           325 => x"0b",
           326 => x"fd",
           327 => x"0b",
           328 => x"0b",
           329 => x"9d",
           330 => x"0b",
           331 => x"0b",
           332 => x"bd",
           333 => x"0b",
           334 => x"0b",
           335 => x"dd",
           336 => x"0b",
           337 => x"0b",
           338 => x"fd",
           339 => x"0b",
           340 => x"0b",
           341 => x"9d",
           342 => x"0b",
           343 => x"0b",
           344 => x"bd",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"d5",
           386 => x"f7",
           387 => x"d5",
           388 => x"80",
           389 => x"d5",
           390 => x"b2",
           391 => x"84",
           392 => x"90",
           393 => x"84",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"82",
           399 => x"84",
           400 => x"82",
           401 => x"94",
           402 => x"d5",
           403 => x"80",
           404 => x"d5",
           405 => x"c2",
           406 => x"84",
           407 => x"90",
           408 => x"84",
           409 => x"f7",
           410 => x"84",
           411 => x"90",
           412 => x"84",
           413 => x"a6",
           414 => x"84",
           415 => x"90",
           416 => x"84",
           417 => x"2d",
           418 => x"08",
           419 => x"04",
           420 => x"0c",
           421 => x"82",
           422 => x"84",
           423 => x"82",
           424 => x"97",
           425 => x"d5",
           426 => x"80",
           427 => x"d5",
           428 => x"fa",
           429 => x"d5",
           430 => x"80",
           431 => x"d5",
           432 => x"fb",
           433 => x"d5",
           434 => x"80",
           435 => x"d5",
           436 => x"f2",
           437 => x"d5",
           438 => x"80",
           439 => x"d5",
           440 => x"f4",
           441 => x"d5",
           442 => x"80",
           443 => x"d5",
           444 => x"f6",
           445 => x"d5",
           446 => x"80",
           447 => x"d5",
           448 => x"eb",
           449 => x"d5",
           450 => x"80",
           451 => x"d5",
           452 => x"f8",
           453 => x"d5",
           454 => x"80",
           455 => x"d5",
           456 => x"f0",
           457 => x"d5",
           458 => x"80",
           459 => x"d5",
           460 => x"f3",
           461 => x"d5",
           462 => x"80",
           463 => x"d5",
           464 => x"fe",
           465 => x"d5",
           466 => x"80",
           467 => x"d5",
           468 => x"87",
           469 => x"d5",
           470 => x"80",
           471 => x"d5",
           472 => x"f7",
           473 => x"d5",
           474 => x"80",
           475 => x"d5",
           476 => x"81",
           477 => x"d5",
           478 => x"80",
           479 => x"d5",
           480 => x"82",
           481 => x"d5",
           482 => x"80",
           483 => x"d5",
           484 => x"83",
           485 => x"d5",
           486 => x"80",
           487 => x"d5",
           488 => x"8a",
           489 => x"d5",
           490 => x"80",
           491 => x"d5",
           492 => x"88",
           493 => x"d5",
           494 => x"80",
           495 => x"d5",
           496 => x"8d",
           497 => x"d5",
           498 => x"80",
           499 => x"d5",
           500 => x"84",
           501 => x"d5",
           502 => x"80",
           503 => x"d5",
           504 => x"90",
           505 => x"d5",
           506 => x"80",
           507 => x"d5",
           508 => x"91",
           509 => x"d5",
           510 => x"80",
           511 => x"d5",
           512 => x"f9",
           513 => x"d5",
           514 => x"80",
           515 => x"d5",
           516 => x"f9",
           517 => x"d5",
           518 => x"80",
           519 => x"d5",
           520 => x"fa",
           521 => x"d5",
           522 => x"80",
           523 => x"d5",
           524 => x"84",
           525 => x"d5",
           526 => x"80",
           527 => x"d5",
           528 => x"92",
           529 => x"d5",
           530 => x"80",
           531 => x"d5",
           532 => x"94",
           533 => x"d5",
           534 => x"80",
           535 => x"d5",
           536 => x"97",
           537 => x"d5",
           538 => x"80",
           539 => x"d5",
           540 => x"eb",
           541 => x"d5",
           542 => x"80",
           543 => x"d5",
           544 => x"9a",
           545 => x"d5",
           546 => x"80",
           547 => x"d5",
           548 => x"a9",
           549 => x"d5",
           550 => x"80",
           551 => x"d5",
           552 => x"a6",
           553 => x"d5",
           554 => x"80",
           555 => x"d5",
           556 => x"ab",
           557 => x"d5",
           558 => x"80",
           559 => x"d5",
           560 => x"ac",
           561 => x"d5",
           562 => x"80",
           563 => x"d5",
           564 => x"ae",
           565 => x"d5",
           566 => x"80",
           567 => x"d5",
           568 => x"f3",
           569 => x"d5",
           570 => x"80",
           571 => x"d5",
           572 => x"f4",
           573 => x"d5",
           574 => x"80",
           575 => x"d5",
           576 => x"f8",
           577 => x"d5",
           578 => x"80",
           579 => x"d5",
           580 => x"d7",
           581 => x"d5",
           582 => x"80",
           583 => x"d5",
           584 => x"a5",
           585 => x"d5",
           586 => x"80",
           587 => x"d5",
           588 => x"a5",
           589 => x"d5",
           590 => x"80",
           591 => x"d5",
           592 => x"a9",
           593 => x"d5",
           594 => x"80",
           595 => x"d5",
           596 => x"a2",
           597 => x"d5",
           598 => x"80",
           599 => x"04",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"04",
           609 => x"81",
           610 => x"83",
           611 => x"05",
           612 => x"10",
           613 => x"72",
           614 => x"51",
           615 => x"72",
           616 => x"06",
           617 => x"72",
           618 => x"10",
           619 => x"10",
           620 => x"ed",
           621 => x"53",
           622 => x"d4",
           623 => x"f0",
           624 => x"38",
           625 => x"84",
           626 => x"0b",
           627 => x"bc",
           628 => x"51",
           629 => x"04",
           630 => x"84",
           631 => x"d5",
           632 => x"3d",
           633 => x"84",
           634 => x"70",
           635 => x"08",
           636 => x"82",
           637 => x"fc",
           638 => x"82",
           639 => x"88",
           640 => x"82",
           641 => x"52",
           642 => x"3f",
           643 => x"08",
           644 => x"84",
           645 => x"0c",
           646 => x"08",
           647 => x"70",
           648 => x"0c",
           649 => x"3d",
           650 => x"84",
           651 => x"d5",
           652 => x"82",
           653 => x"fb",
           654 => x"d5",
           655 => x"05",
           656 => x"33",
           657 => x"70",
           658 => x"51",
           659 => x"8f",
           660 => x"82",
           661 => x"8c",
           662 => x"83",
           663 => x"80",
           664 => x"84",
           665 => x"0c",
           666 => x"82",
           667 => x"8c",
           668 => x"05",
           669 => x"08",
           670 => x"80",
           671 => x"84",
           672 => x"0c",
           673 => x"08",
           674 => x"82",
           675 => x"fc",
           676 => x"d5",
           677 => x"05",
           678 => x"80",
           679 => x"0b",
           680 => x"08",
           681 => x"25",
           682 => x"82",
           683 => x"90",
           684 => x"a0",
           685 => x"d4",
           686 => x"82",
           687 => x"f8",
           688 => x"82",
           689 => x"f8",
           690 => x"2e",
           691 => x"8d",
           692 => x"82",
           693 => x"f4",
           694 => x"d2",
           695 => x"84",
           696 => x"08",
           697 => x"08",
           698 => x"53",
           699 => x"34",
           700 => x"08",
           701 => x"ff",
           702 => x"84",
           703 => x"0c",
           704 => x"08",
           705 => x"81",
           706 => x"84",
           707 => x"0c",
           708 => x"82",
           709 => x"fc",
           710 => x"80",
           711 => x"d5",
           712 => x"05",
           713 => x"d5",
           714 => x"05",
           715 => x"d5",
           716 => x"05",
           717 => x"f8",
           718 => x"0d",
           719 => x"0c",
           720 => x"84",
           721 => x"d5",
           722 => x"3d",
           723 => x"82",
           724 => x"e5",
           725 => x"d5",
           726 => x"05",
           727 => x"84",
           728 => x"0c",
           729 => x"82",
           730 => x"e8",
           731 => x"d5",
           732 => x"05",
           733 => x"84",
           734 => x"0c",
           735 => x"08",
           736 => x"54",
           737 => x"08",
           738 => x"53",
           739 => x"08",
           740 => x"53",
           741 => x"8d",
           742 => x"f8",
           743 => x"d5",
           744 => x"05",
           745 => x"84",
           746 => x"08",
           747 => x"08",
           748 => x"05",
           749 => x"74",
           750 => x"84",
           751 => x"08",
           752 => x"f8",
           753 => x"3d",
           754 => x"84",
           755 => x"d5",
           756 => x"82",
           757 => x"fb",
           758 => x"d5",
           759 => x"05",
           760 => x"84",
           761 => x"0c",
           762 => x"08",
           763 => x"54",
           764 => x"08",
           765 => x"53",
           766 => x"08",
           767 => x"52",
           768 => x"82",
           769 => x"70",
           770 => x"08",
           771 => x"82",
           772 => x"f8",
           773 => x"82",
           774 => x"51",
           775 => x"0d",
           776 => x"0c",
           777 => x"84",
           778 => x"d5",
           779 => x"3d",
           780 => x"82",
           781 => x"e4",
           782 => x"d5",
           783 => x"05",
           784 => x"0b",
           785 => x"82",
           786 => x"88",
           787 => x"11",
           788 => x"2a",
           789 => x"70",
           790 => x"51",
           791 => x"72",
           792 => x"38",
           793 => x"d5",
           794 => x"05",
           795 => x"39",
           796 => x"08",
           797 => x"53",
           798 => x"72",
           799 => x"08",
           800 => x"72",
           801 => x"53",
           802 => x"95",
           803 => x"d5",
           804 => x"05",
           805 => x"82",
           806 => x"8c",
           807 => x"d5",
           808 => x"05",
           809 => x"06",
           810 => x"80",
           811 => x"38",
           812 => x"08",
           813 => x"53",
           814 => x"81",
           815 => x"d5",
           816 => x"05",
           817 => x"b9",
           818 => x"38",
           819 => x"08",
           820 => x"53",
           821 => x"09",
           822 => x"c5",
           823 => x"84",
           824 => x"33",
           825 => x"70",
           826 => x"51",
           827 => x"38",
           828 => x"08",
           829 => x"70",
           830 => x"81",
           831 => x"06",
           832 => x"53",
           833 => x"99",
           834 => x"84",
           835 => x"22",
           836 => x"07",
           837 => x"82",
           838 => x"e4",
           839 => x"d0",
           840 => x"84",
           841 => x"33",
           842 => x"70",
           843 => x"70",
           844 => x"11",
           845 => x"51",
           846 => x"55",
           847 => x"d5",
           848 => x"05",
           849 => x"84",
           850 => x"33",
           851 => x"84",
           852 => x"33",
           853 => x"11",
           854 => x"72",
           855 => x"08",
           856 => x"82",
           857 => x"e8",
           858 => x"98",
           859 => x"2c",
           860 => x"72",
           861 => x"38",
           862 => x"82",
           863 => x"e8",
           864 => x"d5",
           865 => x"05",
           866 => x"2a",
           867 => x"51",
           868 => x"fd",
           869 => x"d5",
           870 => x"05",
           871 => x"2b",
           872 => x"70",
           873 => x"88",
           874 => x"51",
           875 => x"82",
           876 => x"ec",
           877 => x"b8",
           878 => x"84",
           879 => x"22",
           880 => x"70",
           881 => x"51",
           882 => x"2e",
           883 => x"d5",
           884 => x"05",
           885 => x"2b",
           886 => x"51",
           887 => x"8a",
           888 => x"82",
           889 => x"e8",
           890 => x"d5",
           891 => x"05",
           892 => x"82",
           893 => x"c4",
           894 => x"82",
           895 => x"c4",
           896 => x"d8",
           897 => x"38",
           898 => x"08",
           899 => x"70",
           900 => x"ad",
           901 => x"08",
           902 => x"53",
           903 => x"d5",
           904 => x"05",
           905 => x"07",
           906 => x"82",
           907 => x"e4",
           908 => x"d5",
           909 => x"05",
           910 => x"07",
           911 => x"82",
           912 => x"e4",
           913 => x"a8",
           914 => x"84",
           915 => x"22",
           916 => x"07",
           917 => x"82",
           918 => x"e4",
           919 => x"90",
           920 => x"84",
           921 => x"22",
           922 => x"07",
           923 => x"82",
           924 => x"e4",
           925 => x"f8",
           926 => x"84",
           927 => x"22",
           928 => x"51",
           929 => x"d5",
           930 => x"05",
           931 => x"82",
           932 => x"e8",
           933 => x"d8",
           934 => x"84",
           935 => x"22",
           936 => x"51",
           937 => x"d5",
           938 => x"05",
           939 => x"39",
           940 => x"d5",
           941 => x"05",
           942 => x"84",
           943 => x"22",
           944 => x"53",
           945 => x"84",
           946 => x"23",
           947 => x"82",
           948 => x"f8",
           949 => x"a8",
           950 => x"84",
           951 => x"08",
           952 => x"08",
           953 => x"84",
           954 => x"84",
           955 => x"0c",
           956 => x"53",
           957 => x"84",
           958 => x"34",
           959 => x"08",
           960 => x"ff",
           961 => x"72",
           962 => x"08",
           963 => x"8c",
           964 => x"d5",
           965 => x"05",
           966 => x"84",
           967 => x"08",
           968 => x"d5",
           969 => x"05",
           970 => x"82",
           971 => x"fc",
           972 => x"d5",
           973 => x"05",
           974 => x"2a",
           975 => x"51",
           976 => x"72",
           977 => x"38",
           978 => x"08",
           979 => x"70",
           980 => x"72",
           981 => x"82",
           982 => x"fc",
           983 => x"53",
           984 => x"82",
           985 => x"53",
           986 => x"84",
           987 => x"23",
           988 => x"d5",
           989 => x"05",
           990 => x"8a",
           991 => x"f8",
           992 => x"82",
           993 => x"f4",
           994 => x"d5",
           995 => x"05",
           996 => x"d5",
           997 => x"05",
           998 => x"31",
           999 => x"82",
          1000 => x"ec",
          1001 => x"d8",
          1002 => x"84",
          1003 => x"08",
          1004 => x"08",
          1005 => x"84",
          1006 => x"84",
          1007 => x"0c",
          1008 => x"d5",
          1009 => x"05",
          1010 => x"84",
          1011 => x"22",
          1012 => x"70",
          1013 => x"51",
          1014 => x"80",
          1015 => x"82",
          1016 => x"e8",
          1017 => x"98",
          1018 => x"98",
          1019 => x"d5",
          1020 => x"05",
          1021 => x"a2",
          1022 => x"d4",
          1023 => x"72",
          1024 => x"08",
          1025 => x"99",
          1026 => x"84",
          1027 => x"08",
          1028 => x"3f",
          1029 => x"08",
          1030 => x"d5",
          1031 => x"05",
          1032 => x"84",
          1033 => x"22",
          1034 => x"84",
          1035 => x"22",
          1036 => x"54",
          1037 => x"d5",
          1038 => x"05",
          1039 => x"39",
          1040 => x"08",
          1041 => x"70",
          1042 => x"81",
          1043 => x"53",
          1044 => x"a4",
          1045 => x"84",
          1046 => x"08",
          1047 => x"08",
          1048 => x"84",
          1049 => x"84",
          1050 => x"0c",
          1051 => x"d5",
          1052 => x"05",
          1053 => x"39",
          1054 => x"08",
          1055 => x"82",
          1056 => x"90",
          1057 => x"05",
          1058 => x"08",
          1059 => x"70",
          1060 => x"84",
          1061 => x"0c",
          1062 => x"84",
          1063 => x"08",
          1064 => x"08",
          1065 => x"82",
          1066 => x"fc",
          1067 => x"25",
          1068 => x"d5",
          1069 => x"05",
          1070 => x"07",
          1071 => x"82",
          1072 => x"e4",
          1073 => x"d5",
          1074 => x"05",
          1075 => x"d5",
          1076 => x"05",
          1077 => x"84",
          1078 => x"22",
          1079 => x"06",
          1080 => x"82",
          1081 => x"e4",
          1082 => x"af",
          1083 => x"82",
          1084 => x"f4",
          1085 => x"39",
          1086 => x"08",
          1087 => x"70",
          1088 => x"51",
          1089 => x"d5",
          1090 => x"05",
          1091 => x"0b",
          1092 => x"08",
          1093 => x"90",
          1094 => x"84",
          1095 => x"23",
          1096 => x"08",
          1097 => x"70",
          1098 => x"81",
          1099 => x"53",
          1100 => x"a4",
          1101 => x"84",
          1102 => x"08",
          1103 => x"08",
          1104 => x"84",
          1105 => x"84",
          1106 => x"0c",
          1107 => x"d5",
          1108 => x"05",
          1109 => x"39",
          1110 => x"08",
          1111 => x"82",
          1112 => x"90",
          1113 => x"05",
          1114 => x"08",
          1115 => x"70",
          1116 => x"84",
          1117 => x"0c",
          1118 => x"84",
          1119 => x"08",
          1120 => x"08",
          1121 => x"82",
          1122 => x"e4",
          1123 => x"cf",
          1124 => x"72",
          1125 => x"08",
          1126 => x"82",
          1127 => x"82",
          1128 => x"f0",
          1129 => x"d5",
          1130 => x"05",
          1131 => x"84",
          1132 => x"22",
          1133 => x"08",
          1134 => x"71",
          1135 => x"56",
          1136 => x"9e",
          1137 => x"f8",
          1138 => x"75",
          1139 => x"84",
          1140 => x"08",
          1141 => x"08",
          1142 => x"82",
          1143 => x"f0",
          1144 => x"33",
          1145 => x"73",
          1146 => x"82",
          1147 => x"f0",
          1148 => x"72",
          1149 => x"d5",
          1150 => x"05",
          1151 => x"df",
          1152 => x"53",
          1153 => x"84",
          1154 => x"34",
          1155 => x"d5",
          1156 => x"05",
          1157 => x"33",
          1158 => x"53",
          1159 => x"84",
          1160 => x"34",
          1161 => x"08",
          1162 => x"53",
          1163 => x"08",
          1164 => x"73",
          1165 => x"84",
          1166 => x"08",
          1167 => x"d5",
          1168 => x"05",
          1169 => x"84",
          1170 => x"22",
          1171 => x"d5",
          1172 => x"05",
          1173 => x"a3",
          1174 => x"d4",
          1175 => x"82",
          1176 => x"fc",
          1177 => x"82",
          1178 => x"fc",
          1179 => x"2e",
          1180 => x"b2",
          1181 => x"84",
          1182 => x"08",
          1183 => x"54",
          1184 => x"74",
          1185 => x"51",
          1186 => x"d5",
          1187 => x"05",
          1188 => x"84",
          1189 => x"22",
          1190 => x"51",
          1191 => x"2e",
          1192 => x"d5",
          1193 => x"05",
          1194 => x"51",
          1195 => x"d5",
          1196 => x"05",
          1197 => x"84",
          1198 => x"22",
          1199 => x"70",
          1200 => x"51",
          1201 => x"2e",
          1202 => x"82",
          1203 => x"ec",
          1204 => x"90",
          1205 => x"84",
          1206 => x"0c",
          1207 => x"08",
          1208 => x"90",
          1209 => x"84",
          1210 => x"0c",
          1211 => x"08",
          1212 => x"51",
          1213 => x"2e",
          1214 => x"95",
          1215 => x"84",
          1216 => x"08",
          1217 => x"72",
          1218 => x"08",
          1219 => x"93",
          1220 => x"84",
          1221 => x"08",
          1222 => x"72",
          1223 => x"08",
          1224 => x"82",
          1225 => x"c8",
          1226 => x"d5",
          1227 => x"05",
          1228 => x"84",
          1229 => x"22",
          1230 => x"70",
          1231 => x"51",
          1232 => x"2e",
          1233 => x"82",
          1234 => x"e8",
          1235 => x"98",
          1236 => x"2c",
          1237 => x"08",
          1238 => x"57",
          1239 => x"72",
          1240 => x"38",
          1241 => x"08",
          1242 => x"70",
          1243 => x"53",
          1244 => x"84",
          1245 => x"23",
          1246 => x"d5",
          1247 => x"05",
          1248 => x"d5",
          1249 => x"05",
          1250 => x"31",
          1251 => x"82",
          1252 => x"e8",
          1253 => x"d5",
          1254 => x"05",
          1255 => x"2a",
          1256 => x"51",
          1257 => x"80",
          1258 => x"82",
          1259 => x"e8",
          1260 => x"88",
          1261 => x"2b",
          1262 => x"70",
          1263 => x"51",
          1264 => x"72",
          1265 => x"84",
          1266 => x"22",
          1267 => x"51",
          1268 => x"d5",
          1269 => x"05",
          1270 => x"82",
          1271 => x"fc",
          1272 => x"88",
          1273 => x"2b",
          1274 => x"70",
          1275 => x"51",
          1276 => x"72",
          1277 => x"84",
          1278 => x"22",
          1279 => x"51",
          1280 => x"d5",
          1281 => x"05",
          1282 => x"84",
          1283 => x"22",
          1284 => x"06",
          1285 => x"b0",
          1286 => x"84",
          1287 => x"22",
          1288 => x"54",
          1289 => x"84",
          1290 => x"23",
          1291 => x"70",
          1292 => x"53",
          1293 => x"90",
          1294 => x"84",
          1295 => x"08",
          1296 => x"8a",
          1297 => x"39",
          1298 => x"08",
          1299 => x"70",
          1300 => x"81",
          1301 => x"53",
          1302 => x"91",
          1303 => x"84",
          1304 => x"08",
          1305 => x"8a",
          1306 => x"c7",
          1307 => x"84",
          1308 => x"22",
          1309 => x"70",
          1310 => x"51",
          1311 => x"2e",
          1312 => x"d5",
          1313 => x"05",
          1314 => x"51",
          1315 => x"a3",
          1316 => x"84",
          1317 => x"22",
          1318 => x"70",
          1319 => x"51",
          1320 => x"2e",
          1321 => x"d5",
          1322 => x"05",
          1323 => x"51",
          1324 => x"82",
          1325 => x"e4",
          1326 => x"86",
          1327 => x"06",
          1328 => x"72",
          1329 => x"38",
          1330 => x"08",
          1331 => x"52",
          1332 => x"df",
          1333 => x"84",
          1334 => x"22",
          1335 => x"2e",
          1336 => x"94",
          1337 => x"84",
          1338 => x"08",
          1339 => x"84",
          1340 => x"33",
          1341 => x"3f",
          1342 => x"08",
          1343 => x"70",
          1344 => x"81",
          1345 => x"53",
          1346 => x"b0",
          1347 => x"84",
          1348 => x"22",
          1349 => x"54",
          1350 => x"84",
          1351 => x"23",
          1352 => x"70",
          1353 => x"53",
          1354 => x"90",
          1355 => x"84",
          1356 => x"08",
          1357 => x"88",
          1358 => x"39",
          1359 => x"08",
          1360 => x"70",
          1361 => x"81",
          1362 => x"53",
          1363 => x"b0",
          1364 => x"84",
          1365 => x"33",
          1366 => x"54",
          1367 => x"84",
          1368 => x"34",
          1369 => x"70",
          1370 => x"53",
          1371 => x"90",
          1372 => x"84",
          1373 => x"08",
          1374 => x"88",
          1375 => x"39",
          1376 => x"08",
          1377 => x"70",
          1378 => x"81",
          1379 => x"53",
          1380 => x"82",
          1381 => x"ec",
          1382 => x"11",
          1383 => x"82",
          1384 => x"ec",
          1385 => x"90",
          1386 => x"2c",
          1387 => x"73",
          1388 => x"82",
          1389 => x"88",
          1390 => x"a0",
          1391 => x"3f",
          1392 => x"d5",
          1393 => x"05",
          1394 => x"80",
          1395 => x"81",
          1396 => x"82",
          1397 => x"88",
          1398 => x"82",
          1399 => x"fc",
          1400 => x"87",
          1401 => x"ee",
          1402 => x"84",
          1403 => x"33",
          1404 => x"f3",
          1405 => x"06",
          1406 => x"82",
          1407 => x"f4",
          1408 => x"11",
          1409 => x"82",
          1410 => x"f4",
          1411 => x"83",
          1412 => x"53",
          1413 => x"ff",
          1414 => x"38",
          1415 => x"08",
          1416 => x"52",
          1417 => x"08",
          1418 => x"70",
          1419 => x"d5",
          1420 => x"05",
          1421 => x"82",
          1422 => x"fc",
          1423 => x"86",
          1424 => x"b7",
          1425 => x"84",
          1426 => x"33",
          1427 => x"d3",
          1428 => x"06",
          1429 => x"82",
          1430 => x"f4",
          1431 => x"11",
          1432 => x"82",
          1433 => x"f4",
          1434 => x"83",
          1435 => x"53",
          1436 => x"ff",
          1437 => x"38",
          1438 => x"08",
          1439 => x"52",
          1440 => x"08",
          1441 => x"70",
          1442 => x"86",
          1443 => x"d5",
          1444 => x"05",
          1445 => x"82",
          1446 => x"fc",
          1447 => x"b7",
          1448 => x"84",
          1449 => x"08",
          1450 => x"2e",
          1451 => x"d5",
          1452 => x"05",
          1453 => x"d5",
          1454 => x"05",
          1455 => x"82",
          1456 => x"f0",
          1457 => x"d5",
          1458 => x"05",
          1459 => x"52",
          1460 => x"3f",
          1461 => x"d5",
          1462 => x"05",
          1463 => x"2a",
          1464 => x"51",
          1465 => x"80",
          1466 => x"38",
          1467 => x"08",
          1468 => x"ff",
          1469 => x"72",
          1470 => x"08",
          1471 => x"73",
          1472 => x"90",
          1473 => x"80",
          1474 => x"38",
          1475 => x"08",
          1476 => x"52",
          1477 => x"9b",
          1478 => x"82",
          1479 => x"88",
          1480 => x"82",
          1481 => x"f8",
          1482 => x"85",
          1483 => x"0b",
          1484 => x"08",
          1485 => x"ea",
          1486 => x"d5",
          1487 => x"05",
          1488 => x"a5",
          1489 => x"06",
          1490 => x"0b",
          1491 => x"08",
          1492 => x"80",
          1493 => x"84",
          1494 => x"23",
          1495 => x"d5",
          1496 => x"05",
          1497 => x"82",
          1498 => x"f4",
          1499 => x"80",
          1500 => x"84",
          1501 => x"08",
          1502 => x"84",
          1503 => x"33",
          1504 => x"3f",
          1505 => x"82",
          1506 => x"88",
          1507 => x"11",
          1508 => x"d5",
          1509 => x"05",
          1510 => x"82",
          1511 => x"e0",
          1512 => x"d4",
          1513 => x"3d",
          1514 => x"84",
          1515 => x"d5",
          1516 => x"82",
          1517 => x"fd",
          1518 => x"f0",
          1519 => x"82",
          1520 => x"8c",
          1521 => x"82",
          1522 => x"88",
          1523 => x"e4",
          1524 => x"d4",
          1525 => x"82",
          1526 => x"54",
          1527 => x"82",
          1528 => x"04",
          1529 => x"08",
          1530 => x"84",
          1531 => x"0d",
          1532 => x"d5",
          1533 => x"05",
          1534 => x"dc",
          1535 => x"33",
          1536 => x"70",
          1537 => x"81",
          1538 => x"51",
          1539 => x"80",
          1540 => x"ff",
          1541 => x"84",
          1542 => x"0c",
          1543 => x"82",
          1544 => x"88",
          1545 => x"72",
          1546 => x"84",
          1547 => x"08",
          1548 => x"d5",
          1549 => x"05",
          1550 => x"82",
          1551 => x"fc",
          1552 => x"81",
          1553 => x"72",
          1554 => x"38",
          1555 => x"08",
          1556 => x"08",
          1557 => x"84",
          1558 => x"33",
          1559 => x"08",
          1560 => x"2d",
          1561 => x"08",
          1562 => x"2e",
          1563 => x"ff",
          1564 => x"84",
          1565 => x"0c",
          1566 => x"82",
          1567 => x"82",
          1568 => x"53",
          1569 => x"90",
          1570 => x"72",
          1571 => x"f8",
          1572 => x"80",
          1573 => x"ff",
          1574 => x"84",
          1575 => x"0c",
          1576 => x"08",
          1577 => x"70",
          1578 => x"08",
          1579 => x"53",
          1580 => x"08",
          1581 => x"82",
          1582 => x"87",
          1583 => x"d5",
          1584 => x"82",
          1585 => x"02",
          1586 => x"0c",
          1587 => x"80",
          1588 => x"84",
          1589 => x"0c",
          1590 => x"08",
          1591 => x"85",
          1592 => x"81",
          1593 => x"32",
          1594 => x"51",
          1595 => x"53",
          1596 => x"8d",
          1597 => x"82",
          1598 => x"f4",
          1599 => x"f3",
          1600 => x"84",
          1601 => x"08",
          1602 => x"82",
          1603 => x"88",
          1604 => x"05",
          1605 => x"08",
          1606 => x"53",
          1607 => x"84",
          1608 => x"34",
          1609 => x"06",
          1610 => x"2e",
          1611 => x"d5",
          1612 => x"05",
          1613 => x"84",
          1614 => x"08",
          1615 => x"84",
          1616 => x"33",
          1617 => x"08",
          1618 => x"2d",
          1619 => x"08",
          1620 => x"2e",
          1621 => x"ff",
          1622 => x"84",
          1623 => x"0c",
          1624 => x"82",
          1625 => x"f8",
          1626 => x"82",
          1627 => x"f4",
          1628 => x"82",
          1629 => x"f4",
          1630 => x"d4",
          1631 => x"3d",
          1632 => x"84",
          1633 => x"d5",
          1634 => x"82",
          1635 => x"fe",
          1636 => x"f0",
          1637 => x"82",
          1638 => x"88",
          1639 => x"93",
          1640 => x"f8",
          1641 => x"d4",
          1642 => x"84",
          1643 => x"d5",
          1644 => x"82",
          1645 => x"02",
          1646 => x"0c",
          1647 => x"82",
          1648 => x"8c",
          1649 => x"11",
          1650 => x"2a",
          1651 => x"70",
          1652 => x"51",
          1653 => x"72",
          1654 => x"38",
          1655 => x"d5",
          1656 => x"05",
          1657 => x"39",
          1658 => x"08",
          1659 => x"85",
          1660 => x"82",
          1661 => x"06",
          1662 => x"53",
          1663 => x"80",
          1664 => x"d5",
          1665 => x"05",
          1666 => x"84",
          1667 => x"08",
          1668 => x"14",
          1669 => x"08",
          1670 => x"82",
          1671 => x"8c",
          1672 => x"08",
          1673 => x"84",
          1674 => x"08",
          1675 => x"54",
          1676 => x"73",
          1677 => x"74",
          1678 => x"84",
          1679 => x"08",
          1680 => x"81",
          1681 => x"0c",
          1682 => x"08",
          1683 => x"70",
          1684 => x"08",
          1685 => x"51",
          1686 => x"39",
          1687 => x"08",
          1688 => x"82",
          1689 => x"8c",
          1690 => x"82",
          1691 => x"88",
          1692 => x"81",
          1693 => x"90",
          1694 => x"54",
          1695 => x"82",
          1696 => x"53",
          1697 => x"82",
          1698 => x"8c",
          1699 => x"11",
          1700 => x"8c",
          1701 => x"d5",
          1702 => x"05",
          1703 => x"d5",
          1704 => x"05",
          1705 => x"8a",
          1706 => x"82",
          1707 => x"fc",
          1708 => x"d5",
          1709 => x"05",
          1710 => x"f8",
          1711 => x"0d",
          1712 => x"0c",
          1713 => x"84",
          1714 => x"d5",
          1715 => x"3d",
          1716 => x"84",
          1717 => x"08",
          1718 => x"70",
          1719 => x"81",
          1720 => x"51",
          1721 => x"2e",
          1722 => x"0b",
          1723 => x"08",
          1724 => x"83",
          1725 => x"d5",
          1726 => x"05",
          1727 => x"33",
          1728 => x"70",
          1729 => x"51",
          1730 => x"80",
          1731 => x"38",
          1732 => x"08",
          1733 => x"82",
          1734 => x"88",
          1735 => x"53",
          1736 => x"70",
          1737 => x"51",
          1738 => x"14",
          1739 => x"84",
          1740 => x"08",
          1741 => x"81",
          1742 => x"0c",
          1743 => x"08",
          1744 => x"84",
          1745 => x"82",
          1746 => x"f8",
          1747 => x"51",
          1748 => x"39",
          1749 => x"08",
          1750 => x"85",
          1751 => x"82",
          1752 => x"06",
          1753 => x"52",
          1754 => x"80",
          1755 => x"d5",
          1756 => x"05",
          1757 => x"70",
          1758 => x"84",
          1759 => x"0c",
          1760 => x"d5",
          1761 => x"05",
          1762 => x"82",
          1763 => x"88",
          1764 => x"d5",
          1765 => x"05",
          1766 => x"85",
          1767 => x"a0",
          1768 => x"71",
          1769 => x"ff",
          1770 => x"84",
          1771 => x"0c",
          1772 => x"82",
          1773 => x"88",
          1774 => x"08",
          1775 => x"0c",
          1776 => x"39",
          1777 => x"08",
          1778 => x"82",
          1779 => x"88",
          1780 => x"94",
          1781 => x"52",
          1782 => x"d4",
          1783 => x"82",
          1784 => x"fc",
          1785 => x"82",
          1786 => x"fc",
          1787 => x"25",
          1788 => x"82",
          1789 => x"88",
          1790 => x"d5",
          1791 => x"05",
          1792 => x"84",
          1793 => x"08",
          1794 => x"82",
          1795 => x"f0",
          1796 => x"82",
          1797 => x"fc",
          1798 => x"2e",
          1799 => x"95",
          1800 => x"84",
          1801 => x"08",
          1802 => x"71",
          1803 => x"08",
          1804 => x"93",
          1805 => x"84",
          1806 => x"08",
          1807 => x"71",
          1808 => x"08",
          1809 => x"82",
          1810 => x"f4",
          1811 => x"82",
          1812 => x"ec",
          1813 => x"13",
          1814 => x"82",
          1815 => x"f8",
          1816 => x"39",
          1817 => x"08",
          1818 => x"8c",
          1819 => x"05",
          1820 => x"82",
          1821 => x"fc",
          1822 => x"81",
          1823 => x"82",
          1824 => x"f8",
          1825 => x"51",
          1826 => x"84",
          1827 => x"08",
          1828 => x"0c",
          1829 => x"82",
          1830 => x"04",
          1831 => x"08",
          1832 => x"84",
          1833 => x"0d",
          1834 => x"08",
          1835 => x"82",
          1836 => x"fc",
          1837 => x"d5",
          1838 => x"05",
          1839 => x"84",
          1840 => x"0c",
          1841 => x"08",
          1842 => x"80",
          1843 => x"38",
          1844 => x"08",
          1845 => x"82",
          1846 => x"fc",
          1847 => x"81",
          1848 => x"d5",
          1849 => x"05",
          1850 => x"84",
          1851 => x"08",
          1852 => x"d5",
          1853 => x"05",
          1854 => x"81",
          1855 => x"d5",
          1856 => x"05",
          1857 => x"84",
          1858 => x"08",
          1859 => x"84",
          1860 => x"0c",
          1861 => x"08",
          1862 => x"82",
          1863 => x"90",
          1864 => x"82",
          1865 => x"f8",
          1866 => x"d5",
          1867 => x"05",
          1868 => x"82",
          1869 => x"90",
          1870 => x"d5",
          1871 => x"05",
          1872 => x"82",
          1873 => x"90",
          1874 => x"d5",
          1875 => x"05",
          1876 => x"81",
          1877 => x"d5",
          1878 => x"05",
          1879 => x"82",
          1880 => x"fc",
          1881 => x"d5",
          1882 => x"05",
          1883 => x"82",
          1884 => x"f8",
          1885 => x"d5",
          1886 => x"05",
          1887 => x"84",
          1888 => x"08",
          1889 => x"33",
          1890 => x"ae",
          1891 => x"84",
          1892 => x"08",
          1893 => x"d5",
          1894 => x"05",
          1895 => x"84",
          1896 => x"08",
          1897 => x"d5",
          1898 => x"05",
          1899 => x"84",
          1900 => x"08",
          1901 => x"38",
          1902 => x"08",
          1903 => x"51",
          1904 => x"d5",
          1905 => x"05",
          1906 => x"82",
          1907 => x"f8",
          1908 => x"d5",
          1909 => x"05",
          1910 => x"71",
          1911 => x"d5",
          1912 => x"05",
          1913 => x"82",
          1914 => x"fc",
          1915 => x"ad",
          1916 => x"84",
          1917 => x"08",
          1918 => x"f8",
          1919 => x"3d",
          1920 => x"84",
          1921 => x"d5",
          1922 => x"82",
          1923 => x"fe",
          1924 => x"d5",
          1925 => x"05",
          1926 => x"84",
          1927 => x"0c",
          1928 => x"08",
          1929 => x"52",
          1930 => x"d5",
          1931 => x"05",
          1932 => x"82",
          1933 => x"fc",
          1934 => x"81",
          1935 => x"51",
          1936 => x"83",
          1937 => x"82",
          1938 => x"fc",
          1939 => x"05",
          1940 => x"08",
          1941 => x"82",
          1942 => x"fc",
          1943 => x"d5",
          1944 => x"05",
          1945 => x"82",
          1946 => x"51",
          1947 => x"82",
          1948 => x"04",
          1949 => x"08",
          1950 => x"84",
          1951 => x"0d",
          1952 => x"08",
          1953 => x"82",
          1954 => x"fc",
          1955 => x"d5",
          1956 => x"05",
          1957 => x"33",
          1958 => x"08",
          1959 => x"81",
          1960 => x"84",
          1961 => x"0c",
          1962 => x"08",
          1963 => x"53",
          1964 => x"34",
          1965 => x"08",
          1966 => x"81",
          1967 => x"84",
          1968 => x"0c",
          1969 => x"06",
          1970 => x"2e",
          1971 => x"be",
          1972 => x"84",
          1973 => x"08",
          1974 => x"f8",
          1975 => x"3d",
          1976 => x"84",
          1977 => x"d5",
          1978 => x"82",
          1979 => x"fd",
          1980 => x"d5",
          1981 => x"05",
          1982 => x"84",
          1983 => x"0c",
          1984 => x"08",
          1985 => x"82",
          1986 => x"f8",
          1987 => x"d5",
          1988 => x"05",
          1989 => x"80",
          1990 => x"d5",
          1991 => x"05",
          1992 => x"82",
          1993 => x"90",
          1994 => x"d5",
          1995 => x"05",
          1996 => x"82",
          1997 => x"90",
          1998 => x"d5",
          1999 => x"05",
          2000 => x"ba",
          2001 => x"84",
          2002 => x"08",
          2003 => x"82",
          2004 => x"f8",
          2005 => x"05",
          2006 => x"08",
          2007 => x"82",
          2008 => x"fc",
          2009 => x"52",
          2010 => x"82",
          2011 => x"fc",
          2012 => x"05",
          2013 => x"08",
          2014 => x"ff",
          2015 => x"d5",
          2016 => x"05",
          2017 => x"d4",
          2018 => x"85",
          2019 => x"d5",
          2020 => x"82",
          2021 => x"02",
          2022 => x"0c",
          2023 => x"82",
          2024 => x"90",
          2025 => x"2e",
          2026 => x"82",
          2027 => x"8c",
          2028 => x"71",
          2029 => x"84",
          2030 => x"08",
          2031 => x"d5",
          2032 => x"05",
          2033 => x"84",
          2034 => x"08",
          2035 => x"81",
          2036 => x"54",
          2037 => x"71",
          2038 => x"80",
          2039 => x"d5",
          2040 => x"05",
          2041 => x"33",
          2042 => x"08",
          2043 => x"81",
          2044 => x"84",
          2045 => x"0c",
          2046 => x"06",
          2047 => x"8d",
          2048 => x"82",
          2049 => x"fc",
          2050 => x"9b",
          2051 => x"84",
          2052 => x"08",
          2053 => x"d5",
          2054 => x"05",
          2055 => x"84",
          2056 => x"08",
          2057 => x"38",
          2058 => x"82",
          2059 => x"90",
          2060 => x"2e",
          2061 => x"82",
          2062 => x"88",
          2063 => x"33",
          2064 => x"8d",
          2065 => x"82",
          2066 => x"fc",
          2067 => x"d7",
          2068 => x"84",
          2069 => x"08",
          2070 => x"d5",
          2071 => x"05",
          2072 => x"84",
          2073 => x"08",
          2074 => x"52",
          2075 => x"81",
          2076 => x"84",
          2077 => x"0c",
          2078 => x"d5",
          2079 => x"05",
          2080 => x"82",
          2081 => x"8c",
          2082 => x"33",
          2083 => x"70",
          2084 => x"08",
          2085 => x"53",
          2086 => x"53",
          2087 => x"0b",
          2088 => x"08",
          2089 => x"82",
          2090 => x"fc",
          2091 => x"d4",
          2092 => x"3d",
          2093 => x"84",
          2094 => x"d5",
          2095 => x"82",
          2096 => x"fa",
          2097 => x"d5",
          2098 => x"05",
          2099 => x"d5",
          2100 => x"05",
          2101 => x"8d",
          2102 => x"f8",
          2103 => x"d5",
          2104 => x"05",
          2105 => x"84",
          2106 => x"08",
          2107 => x"53",
          2108 => x"e3",
          2109 => x"d4",
          2110 => x"82",
          2111 => x"fc",
          2112 => x"82",
          2113 => x"fc",
          2114 => x"38",
          2115 => x"d5",
          2116 => x"05",
          2117 => x"82",
          2118 => x"fc",
          2119 => x"d5",
          2120 => x"05",
          2121 => x"80",
          2122 => x"d5",
          2123 => x"05",
          2124 => x"d5",
          2125 => x"05",
          2126 => x"d5",
          2127 => x"05",
          2128 => x"a2",
          2129 => x"f8",
          2130 => x"d5",
          2131 => x"05",
          2132 => x"d5",
          2133 => x"05",
          2134 => x"f8",
          2135 => x"0d",
          2136 => x"0c",
          2137 => x"84",
          2138 => x"d5",
          2139 => x"3d",
          2140 => x"84",
          2141 => x"08",
          2142 => x"08",
          2143 => x"82",
          2144 => x"8c",
          2145 => x"38",
          2146 => x"d5",
          2147 => x"05",
          2148 => x"39",
          2149 => x"08",
          2150 => x"52",
          2151 => x"d5",
          2152 => x"05",
          2153 => x"82",
          2154 => x"f8",
          2155 => x"81",
          2156 => x"51",
          2157 => x"9f",
          2158 => x"84",
          2159 => x"08",
          2160 => x"d5",
          2161 => x"05",
          2162 => x"84",
          2163 => x"08",
          2164 => x"38",
          2165 => x"82",
          2166 => x"f8",
          2167 => x"05",
          2168 => x"08",
          2169 => x"82",
          2170 => x"f8",
          2171 => x"d5",
          2172 => x"05",
          2173 => x"82",
          2174 => x"fc",
          2175 => x"82",
          2176 => x"fc",
          2177 => x"d4",
          2178 => x"3d",
          2179 => x"84",
          2180 => x"d5",
          2181 => x"82",
          2182 => x"fe",
          2183 => x"d5",
          2184 => x"05",
          2185 => x"84",
          2186 => x"0c",
          2187 => x"08",
          2188 => x"80",
          2189 => x"38",
          2190 => x"08",
          2191 => x"81",
          2192 => x"84",
          2193 => x"0c",
          2194 => x"08",
          2195 => x"ff",
          2196 => x"84",
          2197 => x"0c",
          2198 => x"08",
          2199 => x"80",
          2200 => x"82",
          2201 => x"8c",
          2202 => x"70",
          2203 => x"08",
          2204 => x"52",
          2205 => x"34",
          2206 => x"08",
          2207 => x"81",
          2208 => x"84",
          2209 => x"0c",
          2210 => x"82",
          2211 => x"88",
          2212 => x"82",
          2213 => x"51",
          2214 => x"82",
          2215 => x"04",
          2216 => x"08",
          2217 => x"84",
          2218 => x"0d",
          2219 => x"d5",
          2220 => x"05",
          2221 => x"84",
          2222 => x"08",
          2223 => x"38",
          2224 => x"08",
          2225 => x"30",
          2226 => x"08",
          2227 => x"80",
          2228 => x"84",
          2229 => x"0c",
          2230 => x"08",
          2231 => x"8a",
          2232 => x"82",
          2233 => x"f4",
          2234 => x"d5",
          2235 => x"05",
          2236 => x"84",
          2237 => x"0c",
          2238 => x"08",
          2239 => x"80",
          2240 => x"82",
          2241 => x"8c",
          2242 => x"82",
          2243 => x"8c",
          2244 => x"0b",
          2245 => x"08",
          2246 => x"82",
          2247 => x"fc",
          2248 => x"38",
          2249 => x"d5",
          2250 => x"05",
          2251 => x"84",
          2252 => x"08",
          2253 => x"08",
          2254 => x"80",
          2255 => x"84",
          2256 => x"08",
          2257 => x"84",
          2258 => x"08",
          2259 => x"3f",
          2260 => x"08",
          2261 => x"84",
          2262 => x"0c",
          2263 => x"84",
          2264 => x"08",
          2265 => x"38",
          2266 => x"08",
          2267 => x"30",
          2268 => x"08",
          2269 => x"82",
          2270 => x"f8",
          2271 => x"82",
          2272 => x"54",
          2273 => x"82",
          2274 => x"04",
          2275 => x"08",
          2276 => x"84",
          2277 => x"0d",
          2278 => x"d5",
          2279 => x"05",
          2280 => x"84",
          2281 => x"08",
          2282 => x"38",
          2283 => x"08",
          2284 => x"30",
          2285 => x"08",
          2286 => x"81",
          2287 => x"84",
          2288 => x"0c",
          2289 => x"08",
          2290 => x"80",
          2291 => x"82",
          2292 => x"8c",
          2293 => x"82",
          2294 => x"8c",
          2295 => x"53",
          2296 => x"08",
          2297 => x"52",
          2298 => x"08",
          2299 => x"51",
          2300 => x"82",
          2301 => x"70",
          2302 => x"08",
          2303 => x"54",
          2304 => x"08",
          2305 => x"80",
          2306 => x"82",
          2307 => x"f8",
          2308 => x"82",
          2309 => x"f8",
          2310 => x"d5",
          2311 => x"05",
          2312 => x"d4",
          2313 => x"87",
          2314 => x"d5",
          2315 => x"82",
          2316 => x"02",
          2317 => x"0c",
          2318 => x"80",
          2319 => x"84",
          2320 => x"08",
          2321 => x"84",
          2322 => x"08",
          2323 => x"3f",
          2324 => x"08",
          2325 => x"f8",
          2326 => x"3d",
          2327 => x"84",
          2328 => x"d5",
          2329 => x"82",
          2330 => x"fd",
          2331 => x"53",
          2332 => x"08",
          2333 => x"52",
          2334 => x"08",
          2335 => x"51",
          2336 => x"d4",
          2337 => x"82",
          2338 => x"54",
          2339 => x"82",
          2340 => x"04",
          2341 => x"08",
          2342 => x"84",
          2343 => x"0d",
          2344 => x"d5",
          2345 => x"05",
          2346 => x"82",
          2347 => x"f8",
          2348 => x"d5",
          2349 => x"05",
          2350 => x"84",
          2351 => x"08",
          2352 => x"82",
          2353 => x"fc",
          2354 => x"2e",
          2355 => x"0b",
          2356 => x"08",
          2357 => x"24",
          2358 => x"d5",
          2359 => x"05",
          2360 => x"d5",
          2361 => x"05",
          2362 => x"84",
          2363 => x"08",
          2364 => x"84",
          2365 => x"0c",
          2366 => x"82",
          2367 => x"fc",
          2368 => x"2e",
          2369 => x"82",
          2370 => x"8c",
          2371 => x"d5",
          2372 => x"05",
          2373 => x"38",
          2374 => x"08",
          2375 => x"82",
          2376 => x"8c",
          2377 => x"82",
          2378 => x"88",
          2379 => x"d5",
          2380 => x"05",
          2381 => x"84",
          2382 => x"08",
          2383 => x"84",
          2384 => x"0c",
          2385 => x"08",
          2386 => x"81",
          2387 => x"84",
          2388 => x"0c",
          2389 => x"08",
          2390 => x"81",
          2391 => x"84",
          2392 => x"0c",
          2393 => x"82",
          2394 => x"90",
          2395 => x"2e",
          2396 => x"d5",
          2397 => x"05",
          2398 => x"d5",
          2399 => x"05",
          2400 => x"39",
          2401 => x"08",
          2402 => x"70",
          2403 => x"08",
          2404 => x"51",
          2405 => x"08",
          2406 => x"82",
          2407 => x"85",
          2408 => x"d5",
          2409 => x"82",
          2410 => x"02",
          2411 => x"0c",
          2412 => x"80",
          2413 => x"84",
          2414 => x"34",
          2415 => x"08",
          2416 => x"53",
          2417 => x"82",
          2418 => x"88",
          2419 => x"08",
          2420 => x"33",
          2421 => x"d5",
          2422 => x"05",
          2423 => x"ff",
          2424 => x"a0",
          2425 => x"06",
          2426 => x"d5",
          2427 => x"05",
          2428 => x"81",
          2429 => x"53",
          2430 => x"d5",
          2431 => x"05",
          2432 => x"ad",
          2433 => x"06",
          2434 => x"0b",
          2435 => x"08",
          2436 => x"82",
          2437 => x"88",
          2438 => x"08",
          2439 => x"0c",
          2440 => x"53",
          2441 => x"d5",
          2442 => x"05",
          2443 => x"84",
          2444 => x"33",
          2445 => x"2e",
          2446 => x"81",
          2447 => x"d5",
          2448 => x"05",
          2449 => x"81",
          2450 => x"70",
          2451 => x"72",
          2452 => x"84",
          2453 => x"34",
          2454 => x"08",
          2455 => x"82",
          2456 => x"e8",
          2457 => x"d5",
          2458 => x"05",
          2459 => x"2e",
          2460 => x"d5",
          2461 => x"05",
          2462 => x"2e",
          2463 => x"cd",
          2464 => x"82",
          2465 => x"f4",
          2466 => x"d5",
          2467 => x"05",
          2468 => x"81",
          2469 => x"70",
          2470 => x"72",
          2471 => x"84",
          2472 => x"34",
          2473 => x"82",
          2474 => x"84",
          2475 => x"34",
          2476 => x"08",
          2477 => x"70",
          2478 => x"71",
          2479 => x"51",
          2480 => x"82",
          2481 => x"f8",
          2482 => x"fe",
          2483 => x"84",
          2484 => x"33",
          2485 => x"26",
          2486 => x"0b",
          2487 => x"08",
          2488 => x"83",
          2489 => x"d5",
          2490 => x"05",
          2491 => x"73",
          2492 => x"82",
          2493 => x"f8",
          2494 => x"72",
          2495 => x"38",
          2496 => x"0b",
          2497 => x"08",
          2498 => x"82",
          2499 => x"0b",
          2500 => x"08",
          2501 => x"b2",
          2502 => x"84",
          2503 => x"33",
          2504 => x"27",
          2505 => x"d5",
          2506 => x"05",
          2507 => x"b9",
          2508 => x"8d",
          2509 => x"82",
          2510 => x"ec",
          2511 => x"a5",
          2512 => x"82",
          2513 => x"f4",
          2514 => x"0b",
          2515 => x"08",
          2516 => x"82",
          2517 => x"f8",
          2518 => x"a0",
          2519 => x"cf",
          2520 => x"84",
          2521 => x"33",
          2522 => x"73",
          2523 => x"82",
          2524 => x"f8",
          2525 => x"11",
          2526 => x"82",
          2527 => x"f8",
          2528 => x"d5",
          2529 => x"05",
          2530 => x"51",
          2531 => x"d5",
          2532 => x"05",
          2533 => x"84",
          2534 => x"33",
          2535 => x"27",
          2536 => x"d5",
          2537 => x"05",
          2538 => x"51",
          2539 => x"d5",
          2540 => x"05",
          2541 => x"84",
          2542 => x"33",
          2543 => x"26",
          2544 => x"0b",
          2545 => x"08",
          2546 => x"81",
          2547 => x"d5",
          2548 => x"05",
          2549 => x"84",
          2550 => x"33",
          2551 => x"74",
          2552 => x"80",
          2553 => x"84",
          2554 => x"0c",
          2555 => x"82",
          2556 => x"f4",
          2557 => x"82",
          2558 => x"fc",
          2559 => x"82",
          2560 => x"f8",
          2561 => x"12",
          2562 => x"08",
          2563 => x"82",
          2564 => x"88",
          2565 => x"08",
          2566 => x"0c",
          2567 => x"51",
          2568 => x"72",
          2569 => x"84",
          2570 => x"34",
          2571 => x"82",
          2572 => x"f0",
          2573 => x"72",
          2574 => x"38",
          2575 => x"08",
          2576 => x"30",
          2577 => x"08",
          2578 => x"82",
          2579 => x"8c",
          2580 => x"d5",
          2581 => x"05",
          2582 => x"53",
          2583 => x"d5",
          2584 => x"05",
          2585 => x"84",
          2586 => x"08",
          2587 => x"0c",
          2588 => x"82",
          2589 => x"04",
          2590 => x"08",
          2591 => x"84",
          2592 => x"0d",
          2593 => x"d5",
          2594 => x"05",
          2595 => x"84",
          2596 => x"08",
          2597 => x"0c",
          2598 => x"08",
          2599 => x"70",
          2600 => x"72",
          2601 => x"82",
          2602 => x"f8",
          2603 => x"81",
          2604 => x"72",
          2605 => x"81",
          2606 => x"82",
          2607 => x"88",
          2608 => x"08",
          2609 => x"0c",
          2610 => x"82",
          2611 => x"f8",
          2612 => x"72",
          2613 => x"81",
          2614 => x"81",
          2615 => x"84",
          2616 => x"34",
          2617 => x"08",
          2618 => x"70",
          2619 => x"71",
          2620 => x"51",
          2621 => x"82",
          2622 => x"f8",
          2623 => x"d5",
          2624 => x"05",
          2625 => x"b0",
          2626 => x"06",
          2627 => x"82",
          2628 => x"88",
          2629 => x"08",
          2630 => x"0c",
          2631 => x"53",
          2632 => x"d5",
          2633 => x"05",
          2634 => x"84",
          2635 => x"33",
          2636 => x"08",
          2637 => x"82",
          2638 => x"e8",
          2639 => x"e2",
          2640 => x"82",
          2641 => x"e8",
          2642 => x"f8",
          2643 => x"80",
          2644 => x"0b",
          2645 => x"08",
          2646 => x"82",
          2647 => x"88",
          2648 => x"08",
          2649 => x"0c",
          2650 => x"53",
          2651 => x"d5",
          2652 => x"05",
          2653 => x"39",
          2654 => x"d5",
          2655 => x"05",
          2656 => x"84",
          2657 => x"08",
          2658 => x"05",
          2659 => x"08",
          2660 => x"33",
          2661 => x"08",
          2662 => x"80",
          2663 => x"d5",
          2664 => x"05",
          2665 => x"a0",
          2666 => x"81",
          2667 => x"84",
          2668 => x"0c",
          2669 => x"82",
          2670 => x"f8",
          2671 => x"af",
          2672 => x"38",
          2673 => x"08",
          2674 => x"53",
          2675 => x"83",
          2676 => x"80",
          2677 => x"84",
          2678 => x"0c",
          2679 => x"88",
          2680 => x"84",
          2681 => x"34",
          2682 => x"d5",
          2683 => x"05",
          2684 => x"73",
          2685 => x"82",
          2686 => x"f8",
          2687 => x"72",
          2688 => x"38",
          2689 => x"0b",
          2690 => x"08",
          2691 => x"82",
          2692 => x"0b",
          2693 => x"08",
          2694 => x"80",
          2695 => x"84",
          2696 => x"0c",
          2697 => x"08",
          2698 => x"53",
          2699 => x"81",
          2700 => x"d5",
          2701 => x"05",
          2702 => x"e0",
          2703 => x"38",
          2704 => x"08",
          2705 => x"e0",
          2706 => x"72",
          2707 => x"08",
          2708 => x"82",
          2709 => x"f8",
          2710 => x"11",
          2711 => x"82",
          2712 => x"f8",
          2713 => x"d5",
          2714 => x"05",
          2715 => x"73",
          2716 => x"82",
          2717 => x"f8",
          2718 => x"11",
          2719 => x"82",
          2720 => x"f8",
          2721 => x"d5",
          2722 => x"05",
          2723 => x"89",
          2724 => x"80",
          2725 => x"84",
          2726 => x"0c",
          2727 => x"82",
          2728 => x"f8",
          2729 => x"d5",
          2730 => x"05",
          2731 => x"72",
          2732 => x"38",
          2733 => x"d5",
          2734 => x"05",
          2735 => x"39",
          2736 => x"08",
          2737 => x"70",
          2738 => x"08",
          2739 => x"29",
          2740 => x"08",
          2741 => x"70",
          2742 => x"84",
          2743 => x"0c",
          2744 => x"08",
          2745 => x"70",
          2746 => x"71",
          2747 => x"51",
          2748 => x"53",
          2749 => x"d5",
          2750 => x"05",
          2751 => x"39",
          2752 => x"08",
          2753 => x"53",
          2754 => x"90",
          2755 => x"84",
          2756 => x"08",
          2757 => x"84",
          2758 => x"0c",
          2759 => x"08",
          2760 => x"82",
          2761 => x"fc",
          2762 => x"0c",
          2763 => x"82",
          2764 => x"ec",
          2765 => x"d5",
          2766 => x"05",
          2767 => x"f8",
          2768 => x"0d",
          2769 => x"0c",
          2770 => x"0d",
          2771 => x"70",
          2772 => x"74",
          2773 => x"df",
          2774 => x"77",
          2775 => x"85",
          2776 => x"80",
          2777 => x"33",
          2778 => x"2e",
          2779 => x"86",
          2780 => x"55",
          2781 => x"57",
          2782 => x"82",
          2783 => x"70",
          2784 => x"e5",
          2785 => x"d4",
          2786 => x"d4",
          2787 => x"75",
          2788 => x"52",
          2789 => x"3f",
          2790 => x"08",
          2791 => x"16",
          2792 => x"81",
          2793 => x"38",
          2794 => x"81",
          2795 => x"54",
          2796 => x"c4",
          2797 => x"73",
          2798 => x"0c",
          2799 => x"04",
          2800 => x"73",
          2801 => x"26",
          2802 => x"71",
          2803 => x"ac",
          2804 => x"71",
          2805 => x"b2",
          2806 => x"80",
          2807 => x"94",
          2808 => x"39",
          2809 => x"51",
          2810 => x"82",
          2811 => x"80",
          2812 => x"b2",
          2813 => x"e4",
          2814 => x"d4",
          2815 => x"39",
          2816 => x"51",
          2817 => x"82",
          2818 => x"80",
          2819 => x"b3",
          2820 => x"c8",
          2821 => x"a8",
          2822 => x"39",
          2823 => x"51",
          2824 => x"b3",
          2825 => x"39",
          2826 => x"51",
          2827 => x"b4",
          2828 => x"39",
          2829 => x"51",
          2830 => x"b4",
          2831 => x"39",
          2832 => x"51",
          2833 => x"b4",
          2834 => x"39",
          2835 => x"51",
          2836 => x"b5",
          2837 => x"39",
          2838 => x"51",
          2839 => x"83",
          2840 => x"fb",
          2841 => x"79",
          2842 => x"87",
          2843 => x"38",
          2844 => x"87",
          2845 => x"90",
          2846 => x"52",
          2847 => x"af",
          2848 => x"f8",
          2849 => x"51",
          2850 => x"82",
          2851 => x"54",
          2852 => x"52",
          2853 => x"51",
          2854 => x"3f",
          2855 => x"04",
          2856 => x"66",
          2857 => x"80",
          2858 => x"5b",
          2859 => x"78",
          2860 => x"07",
          2861 => x"57",
          2862 => x"56",
          2863 => x"26",
          2864 => x"56",
          2865 => x"70",
          2866 => x"51",
          2867 => x"74",
          2868 => x"81",
          2869 => x"8c",
          2870 => x"56",
          2871 => x"3f",
          2872 => x"08",
          2873 => x"f8",
          2874 => x"82",
          2875 => x"87",
          2876 => x"0c",
          2877 => x"08",
          2878 => x"d4",
          2879 => x"80",
          2880 => x"75",
          2881 => x"c9",
          2882 => x"f8",
          2883 => x"d4",
          2884 => x"38",
          2885 => x"80",
          2886 => x"74",
          2887 => x"59",
          2888 => x"96",
          2889 => x"51",
          2890 => x"3f",
          2891 => x"78",
          2892 => x"7b",
          2893 => x"2a",
          2894 => x"57",
          2895 => x"80",
          2896 => x"82",
          2897 => x"87",
          2898 => x"08",
          2899 => x"fe",
          2900 => x"56",
          2901 => x"f8",
          2902 => x"0d",
          2903 => x"0d",
          2904 => x"05",
          2905 => x"59",
          2906 => x"80",
          2907 => x"7b",
          2908 => x"3f",
          2909 => x"08",
          2910 => x"77",
          2911 => x"38",
          2912 => x"bf",
          2913 => x"82",
          2914 => x"82",
          2915 => x"82",
          2916 => x"82",
          2917 => x"54",
          2918 => x"08",
          2919 => x"d8",
          2920 => x"b5",
          2921 => x"b8",
          2922 => x"f0",
          2923 => x"55",
          2924 => x"d4",
          2925 => x"52",
          2926 => x"2d",
          2927 => x"08",
          2928 => x"79",
          2929 => x"d4",
          2930 => x"3d",
          2931 => x"3d",
          2932 => x"63",
          2933 => x"80",
          2934 => x"73",
          2935 => x"41",
          2936 => x"5e",
          2937 => x"52",
          2938 => x"51",
          2939 => x"3f",
          2940 => x"51",
          2941 => x"3f",
          2942 => x"79",
          2943 => x"38",
          2944 => x"89",
          2945 => x"2e",
          2946 => x"c6",
          2947 => x"53",
          2948 => x"8e",
          2949 => x"52",
          2950 => x"51",
          2951 => x"3f",
          2952 => x"b6",
          2953 => x"b7",
          2954 => x"15",
          2955 => x"39",
          2956 => x"72",
          2957 => x"38",
          2958 => x"82",
          2959 => x"ff",
          2960 => x"89",
          2961 => x"b0",
          2962 => x"8d",
          2963 => x"55",
          2964 => x"18",
          2965 => x"27",
          2966 => x"33",
          2967 => x"bc",
          2968 => x"f5",
          2969 => x"82",
          2970 => x"ff",
          2971 => x"81",
          2972 => x"f0",
          2973 => x"a0",
          2974 => x"3f",
          2975 => x"82",
          2976 => x"ff",
          2977 => x"80",
          2978 => x"27",
          2979 => x"74",
          2980 => x"55",
          2981 => x"72",
          2982 => x"38",
          2983 => x"53",
          2984 => x"83",
          2985 => x"75",
          2986 => x"81",
          2987 => x"53",
          2988 => x"90",
          2989 => x"fe",
          2990 => x"82",
          2991 => x"52",
          2992 => x"39",
          2993 => x"08",
          2994 => x"d5",
          2995 => x"15",
          2996 => x"39",
          2997 => x"51",
          2998 => x"78",
          2999 => x"5c",
          3000 => x"3f",
          3001 => x"08",
          3002 => x"98",
          3003 => x"76",
          3004 => x"81",
          3005 => x"9d",
          3006 => x"d4",
          3007 => x"2b",
          3008 => x"70",
          3009 => x"30",
          3010 => x"70",
          3011 => x"07",
          3012 => x"06",
          3013 => x"59",
          3014 => x"80",
          3015 => x"38",
          3016 => x"09",
          3017 => x"38",
          3018 => x"39",
          3019 => x"72",
          3020 => x"b2",
          3021 => x"72",
          3022 => x"0c",
          3023 => x"04",
          3024 => x"02",
          3025 => x"82",
          3026 => x"82",
          3027 => x"55",
          3028 => x"3f",
          3029 => x"22",
          3030 => x"3f",
          3031 => x"54",
          3032 => x"53",
          3033 => x"33",
          3034 => x"f4",
          3035 => x"e9",
          3036 => x"2e",
          3037 => x"ca",
          3038 => x"0d",
          3039 => x"0d",
          3040 => x"80",
          3041 => x"b2",
          3042 => x"99",
          3043 => x"b7",
          3044 => x"95",
          3045 => x"98",
          3046 => x"81",
          3047 => x"06",
          3048 => x"80",
          3049 => x"81",
          3050 => x"3f",
          3051 => x"51",
          3052 => x"80",
          3053 => x"3f",
          3054 => x"70",
          3055 => x"52",
          3056 => x"92",
          3057 => x"98",
          3058 => x"b7",
          3059 => x"d9",
          3060 => x"98",
          3061 => x"83",
          3062 => x"06",
          3063 => x"80",
          3064 => x"81",
          3065 => x"3f",
          3066 => x"51",
          3067 => x"80",
          3068 => x"3f",
          3069 => x"70",
          3070 => x"52",
          3071 => x"92",
          3072 => x"98",
          3073 => x"b7",
          3074 => x"9d",
          3075 => x"97",
          3076 => x"85",
          3077 => x"06",
          3078 => x"80",
          3079 => x"81",
          3080 => x"3f",
          3081 => x"51",
          3082 => x"80",
          3083 => x"3f",
          3084 => x"70",
          3085 => x"52",
          3086 => x"92",
          3087 => x"97",
          3088 => x"b8",
          3089 => x"e1",
          3090 => x"97",
          3091 => x"87",
          3092 => x"06",
          3093 => x"80",
          3094 => x"81",
          3095 => x"3f",
          3096 => x"51",
          3097 => x"80",
          3098 => x"3f",
          3099 => x"70",
          3100 => x"52",
          3101 => x"92",
          3102 => x"97",
          3103 => x"b8",
          3104 => x"a5",
          3105 => x"97",
          3106 => x"b6",
          3107 => x"0d",
          3108 => x"0d",
          3109 => x"05",
          3110 => x"70",
          3111 => x"80",
          3112 => x"e2",
          3113 => x"0b",
          3114 => x"33",
          3115 => x"38",
          3116 => x"b8",
          3117 => x"ec",
          3118 => x"8a",
          3119 => x"d4",
          3120 => x"70",
          3121 => x"08",
          3122 => x"82",
          3123 => x"51",
          3124 => x"0b",
          3125 => x"34",
          3126 => x"cf",
          3127 => x"73",
          3128 => x"81",
          3129 => x"82",
          3130 => x"74",
          3131 => x"81",
          3132 => x"82",
          3133 => x"80",
          3134 => x"82",
          3135 => x"51",
          3136 => x"91",
          3137 => x"88",
          3138 => x"df",
          3139 => x"0b",
          3140 => x"f4",
          3141 => x"82",
          3142 => x"54",
          3143 => x"09",
          3144 => x"38",
          3145 => x"53",
          3146 => x"51",
          3147 => x"80",
          3148 => x"f8",
          3149 => x"0d",
          3150 => x"0d",
          3151 => x"5e",
          3152 => x"ec",
          3153 => x"81",
          3154 => x"80",
          3155 => x"82",
          3156 => x"81",
          3157 => x"78",
          3158 => x"81",
          3159 => x"97",
          3160 => x"53",
          3161 => x"52",
          3162 => x"fa",
          3163 => x"78",
          3164 => x"a4",
          3165 => x"93",
          3166 => x"f8",
          3167 => x"88",
          3168 => x"84",
          3169 => x"39",
          3170 => x"5e",
          3171 => x"51",
          3172 => x"3f",
          3173 => x"47",
          3174 => x"52",
          3175 => x"f1",
          3176 => x"ff",
          3177 => x"f3",
          3178 => x"d4",
          3179 => x"2b",
          3180 => x"51",
          3181 => x"c2",
          3182 => x"38",
          3183 => x"24",
          3184 => x"bd",
          3185 => x"38",
          3186 => x"90",
          3187 => x"2e",
          3188 => x"78",
          3189 => x"da",
          3190 => x"39",
          3191 => x"2e",
          3192 => x"78",
          3193 => x"85",
          3194 => x"bf",
          3195 => x"38",
          3196 => x"78",
          3197 => x"89",
          3198 => x"80",
          3199 => x"38",
          3200 => x"2e",
          3201 => x"78",
          3202 => x"89",
          3203 => x"a1",
          3204 => x"83",
          3205 => x"38",
          3206 => x"24",
          3207 => x"81",
          3208 => x"ed",
          3209 => x"39",
          3210 => x"2e",
          3211 => x"8a",
          3212 => x"3d",
          3213 => x"53",
          3214 => x"51",
          3215 => x"82",
          3216 => x"80",
          3217 => x"38",
          3218 => x"fc",
          3219 => x"84",
          3220 => x"a4",
          3221 => x"f8",
          3222 => x"fe",
          3223 => x"3d",
          3224 => x"53",
          3225 => x"51",
          3226 => x"82",
          3227 => x"86",
          3228 => x"f8",
          3229 => x"b9",
          3230 => x"ae",
          3231 => x"64",
          3232 => x"7b",
          3233 => x"38",
          3234 => x"7a",
          3235 => x"5c",
          3236 => x"26",
          3237 => x"db",
          3238 => x"ff",
          3239 => x"ff",
          3240 => x"eb",
          3241 => x"d4",
          3242 => x"2e",
          3243 => x"b5",
          3244 => x"11",
          3245 => x"05",
          3246 => x"3f",
          3247 => x"08",
          3248 => x"c8",
          3249 => x"fe",
          3250 => x"ff",
          3251 => x"eb",
          3252 => x"d4",
          3253 => x"2e",
          3254 => x"82",
          3255 => x"ff",
          3256 => x"64",
          3257 => x"27",
          3258 => x"62",
          3259 => x"81",
          3260 => x"79",
          3261 => x"05",
          3262 => x"b5",
          3263 => x"11",
          3264 => x"05",
          3265 => x"3f",
          3266 => x"08",
          3267 => x"fc",
          3268 => x"fe",
          3269 => x"ff",
          3270 => x"ea",
          3271 => x"d4",
          3272 => x"2e",
          3273 => x"b5",
          3274 => x"11",
          3275 => x"05",
          3276 => x"3f",
          3277 => x"08",
          3278 => x"d0",
          3279 => x"dc",
          3280 => x"95",
          3281 => x"79",
          3282 => x"38",
          3283 => x"7b",
          3284 => x"5b",
          3285 => x"92",
          3286 => x"7a",
          3287 => x"53",
          3288 => x"b9",
          3289 => x"ac",
          3290 => x"1a",
          3291 => x"44",
          3292 => x"8a",
          3293 => x"3f",
          3294 => x"b5",
          3295 => x"11",
          3296 => x"05",
          3297 => x"3f",
          3298 => x"08",
          3299 => x"82",
          3300 => x"59",
          3301 => x"89",
          3302 => x"9c",
          3303 => x"cd",
          3304 => x"e5",
          3305 => x"80",
          3306 => x"82",
          3307 => x"45",
          3308 => x"d3",
          3309 => x"78",
          3310 => x"38",
          3311 => x"08",
          3312 => x"82",
          3313 => x"59",
          3314 => x"88",
          3315 => x"b4",
          3316 => x"39",
          3317 => x"33",
          3318 => x"2e",
          3319 => x"d3",
          3320 => x"89",
          3321 => x"cc",
          3322 => x"05",
          3323 => x"fe",
          3324 => x"ff",
          3325 => x"e8",
          3326 => x"d4",
          3327 => x"de",
          3328 => x"e4",
          3329 => x"80",
          3330 => x"82",
          3331 => x"44",
          3332 => x"82",
          3333 => x"59",
          3334 => x"88",
          3335 => x"a8",
          3336 => x"39",
          3337 => x"33",
          3338 => x"2e",
          3339 => x"d3",
          3340 => x"aa",
          3341 => x"e7",
          3342 => x"80",
          3343 => x"82",
          3344 => x"44",
          3345 => x"d3",
          3346 => x"78",
          3347 => x"38",
          3348 => x"08",
          3349 => x"82",
          3350 => x"88",
          3351 => x"3d",
          3352 => x"53",
          3353 => x"51",
          3354 => x"82",
          3355 => x"80",
          3356 => x"80",
          3357 => x"7a",
          3358 => x"38",
          3359 => x"90",
          3360 => x"70",
          3361 => x"2a",
          3362 => x"51",
          3363 => x"78",
          3364 => x"38",
          3365 => x"83",
          3366 => x"82",
          3367 => x"c6",
          3368 => x"55",
          3369 => x"53",
          3370 => x"51",
          3371 => x"82",
          3372 => x"87",
          3373 => x"3d",
          3374 => x"53",
          3375 => x"51",
          3376 => x"82",
          3377 => x"80",
          3378 => x"38",
          3379 => x"fc",
          3380 => x"84",
          3381 => x"a0",
          3382 => x"f8",
          3383 => x"a4",
          3384 => x"02",
          3385 => x"33",
          3386 => x"81",
          3387 => x"3d",
          3388 => x"53",
          3389 => x"51",
          3390 => x"82",
          3391 => x"e1",
          3392 => x"39",
          3393 => x"54",
          3394 => x"a0",
          3395 => x"c9",
          3396 => x"d8",
          3397 => x"f8",
          3398 => x"ff",
          3399 => x"79",
          3400 => x"59",
          3401 => x"f8",
          3402 => x"79",
          3403 => x"b5",
          3404 => x"11",
          3405 => x"05",
          3406 => x"3f",
          3407 => x"08",
          3408 => x"38",
          3409 => x"80",
          3410 => x"79",
          3411 => x"05",
          3412 => x"39",
          3413 => x"51",
          3414 => x"ff",
          3415 => x"3d",
          3416 => x"53",
          3417 => x"51",
          3418 => x"82",
          3419 => x"80",
          3420 => x"38",
          3421 => x"f0",
          3422 => x"84",
          3423 => x"a7",
          3424 => x"f8",
          3425 => x"a6",
          3426 => x"02",
          3427 => x"22",
          3428 => x"05",
          3429 => x"42",
          3430 => x"f0",
          3431 => x"84",
          3432 => x"83",
          3433 => x"f8",
          3434 => x"f7",
          3435 => x"70",
          3436 => x"82",
          3437 => x"ff",
          3438 => x"82",
          3439 => x"53",
          3440 => x"79",
          3441 => x"e6",
          3442 => x"79",
          3443 => x"ae",
          3444 => x"38",
          3445 => x"87",
          3446 => x"05",
          3447 => x"b5",
          3448 => x"11",
          3449 => x"05",
          3450 => x"3f",
          3451 => x"08",
          3452 => x"38",
          3453 => x"80",
          3454 => x"79",
          3455 => x"5b",
          3456 => x"ff",
          3457 => x"ba",
          3458 => x"d8",
          3459 => x"39",
          3460 => x"f4",
          3461 => x"84",
          3462 => x"8b",
          3463 => x"f8",
          3464 => x"f6",
          3465 => x"3d",
          3466 => x"53",
          3467 => x"51",
          3468 => x"82",
          3469 => x"80",
          3470 => x"61",
          3471 => x"59",
          3472 => x"42",
          3473 => x"f0",
          3474 => x"84",
          3475 => x"d7",
          3476 => x"f8",
          3477 => x"f6",
          3478 => x"70",
          3479 => x"82",
          3480 => x"ff",
          3481 => x"82",
          3482 => x"53",
          3483 => x"79",
          3484 => x"ba",
          3485 => x"79",
          3486 => x"ae",
          3487 => x"38",
          3488 => x"9b",
          3489 => x"fe",
          3490 => x"ff",
          3491 => x"de",
          3492 => x"d4",
          3493 => x"2e",
          3494 => x"61",
          3495 => x"61",
          3496 => x"ff",
          3497 => x"ba",
          3498 => x"b8",
          3499 => x"39",
          3500 => x"80",
          3501 => x"84",
          3502 => x"bc",
          3503 => x"f8",
          3504 => x"f5",
          3505 => x"52",
          3506 => x"51",
          3507 => x"3f",
          3508 => x"04",
          3509 => x"80",
          3510 => x"84",
          3511 => x"98",
          3512 => x"f8",
          3513 => x"f5",
          3514 => x"52",
          3515 => x"51",
          3516 => x"3f",
          3517 => x"2d",
          3518 => x"08",
          3519 => x"8c",
          3520 => x"f8",
          3521 => x"bb",
          3522 => x"a5",
          3523 => x"fc",
          3524 => x"a0",
          3525 => x"3f",
          3526 => x"3f",
          3527 => x"82",
          3528 => x"c1",
          3529 => x"59",
          3530 => x"92",
          3531 => x"dc",
          3532 => x"33",
          3533 => x"2e",
          3534 => x"80",
          3535 => x"51",
          3536 => x"82",
          3537 => x"5d",
          3538 => x"08",
          3539 => x"92",
          3540 => x"f8",
          3541 => x"3d",
          3542 => x"51",
          3543 => x"82",
          3544 => x"60",
          3545 => x"5c",
          3546 => x"81",
          3547 => x"d4",
          3548 => x"cd",
          3549 => x"d4",
          3550 => x"26",
          3551 => x"81",
          3552 => x"2e",
          3553 => x"82",
          3554 => x"7a",
          3555 => x"38",
          3556 => x"7a",
          3557 => x"38",
          3558 => x"82",
          3559 => x"7b",
          3560 => x"d4",
          3561 => x"82",
          3562 => x"b5",
          3563 => x"05",
          3564 => x"8d",
          3565 => x"7b",
          3566 => x"ff",
          3567 => x"cd",
          3568 => x"39",
          3569 => x"bb",
          3570 => x"53",
          3571 => x"52",
          3572 => x"b0",
          3573 => x"a6",
          3574 => x"39",
          3575 => x"53",
          3576 => x"52",
          3577 => x"b0",
          3578 => x"a6",
          3579 => x"d3",
          3580 => x"d5",
          3581 => x"56",
          3582 => x"54",
          3583 => x"53",
          3584 => x"52",
          3585 => x"b0",
          3586 => x"d1",
          3587 => x"f8",
          3588 => x"f8",
          3589 => x"30",
          3590 => x"80",
          3591 => x"5b",
          3592 => x"7a",
          3593 => x"38",
          3594 => x"7a",
          3595 => x"80",
          3596 => x"81",
          3597 => x"ff",
          3598 => x"7a",
          3599 => x"7f",
          3600 => x"81",
          3601 => x"78",
          3602 => x"ff",
          3603 => x"06",
          3604 => x"bb",
          3605 => x"bf",
          3606 => x"51",
          3607 => x"f2",
          3608 => x"bc",
          3609 => x"be",
          3610 => x"a0",
          3611 => x"0d",
          3612 => x"d5",
          3613 => x"c0",
          3614 => x"53",
          3615 => x"52",
          3616 => x"ab",
          3617 => x"f8",
          3618 => x"87",
          3619 => x"08",
          3620 => x"84",
          3621 => x"51",
          3622 => x"72",
          3623 => x"08",
          3624 => x"94",
          3625 => x"c0",
          3626 => x"53",
          3627 => x"52",
          3628 => x"fb",
          3629 => x"f8",
          3630 => x"87",
          3631 => x"08",
          3632 => x"84",
          3633 => x"51",
          3634 => x"72",
          3635 => x"08",
          3636 => x"94",
          3637 => x"80",
          3638 => x"c0",
          3639 => x"8c",
          3640 => x"87",
          3641 => x"0c",
          3642 => x"53",
          3643 => x"84",
          3644 => x"05",
          3645 => x"bf",
          3646 => x"27",
          3647 => x"80",
          3648 => x"de",
          3649 => x"73",
          3650 => x"55",
          3651 => x"ff",
          3652 => x"ee",
          3653 => x"a4",
          3654 => x"90",
          3655 => x"84",
          3656 => x"34",
          3657 => x"3d",
          3658 => x"e0",
          3659 => x"f0",
          3660 => x"f0",
          3661 => x"be",
          3662 => x"3f",
          3663 => x"51",
          3664 => x"3f",
          3665 => x"51",
          3666 => x"3f",
          3667 => x"51",
          3668 => x"81",
          3669 => x"3f",
          3670 => x"80",
          3671 => x"0d",
          3672 => x"53",
          3673 => x"52",
          3674 => x"82",
          3675 => x"81",
          3676 => x"07",
          3677 => x"52",
          3678 => x"e8",
          3679 => x"d4",
          3680 => x"3d",
          3681 => x"3d",
          3682 => x"08",
          3683 => x"73",
          3684 => x"74",
          3685 => x"38",
          3686 => x"70",
          3687 => x"81",
          3688 => x"81",
          3689 => x"39",
          3690 => x"70",
          3691 => x"81",
          3692 => x"81",
          3693 => x"54",
          3694 => x"81",
          3695 => x"06",
          3696 => x"39",
          3697 => x"80",
          3698 => x"54",
          3699 => x"83",
          3700 => x"70",
          3701 => x"38",
          3702 => x"98",
          3703 => x"52",
          3704 => x"52",
          3705 => x"2e",
          3706 => x"54",
          3707 => x"84",
          3708 => x"38",
          3709 => x"52",
          3710 => x"2e",
          3711 => x"83",
          3712 => x"70",
          3713 => x"30",
          3714 => x"76",
          3715 => x"51",
          3716 => x"88",
          3717 => x"70",
          3718 => x"34",
          3719 => x"72",
          3720 => x"d4",
          3721 => x"3d",
          3722 => x"3d",
          3723 => x"72",
          3724 => x"91",
          3725 => x"fc",
          3726 => x"51",
          3727 => x"82",
          3728 => x"85",
          3729 => x"83",
          3730 => x"72",
          3731 => x"0c",
          3732 => x"04",
          3733 => x"76",
          3734 => x"ff",
          3735 => x"81",
          3736 => x"26",
          3737 => x"83",
          3738 => x"05",
          3739 => x"70",
          3740 => x"8a",
          3741 => x"33",
          3742 => x"70",
          3743 => x"fe",
          3744 => x"33",
          3745 => x"70",
          3746 => x"f2",
          3747 => x"33",
          3748 => x"70",
          3749 => x"e6",
          3750 => x"22",
          3751 => x"74",
          3752 => x"80",
          3753 => x"13",
          3754 => x"52",
          3755 => x"26",
          3756 => x"81",
          3757 => x"98",
          3758 => x"22",
          3759 => x"bc",
          3760 => x"33",
          3761 => x"b8",
          3762 => x"33",
          3763 => x"b4",
          3764 => x"33",
          3765 => x"b0",
          3766 => x"33",
          3767 => x"ac",
          3768 => x"33",
          3769 => x"a8",
          3770 => x"c0",
          3771 => x"73",
          3772 => x"a0",
          3773 => x"87",
          3774 => x"0c",
          3775 => x"82",
          3776 => x"86",
          3777 => x"f3",
          3778 => x"5b",
          3779 => x"9c",
          3780 => x"0c",
          3781 => x"bc",
          3782 => x"7b",
          3783 => x"98",
          3784 => x"79",
          3785 => x"87",
          3786 => x"08",
          3787 => x"1c",
          3788 => x"98",
          3789 => x"79",
          3790 => x"87",
          3791 => x"08",
          3792 => x"1c",
          3793 => x"98",
          3794 => x"79",
          3795 => x"87",
          3796 => x"08",
          3797 => x"1c",
          3798 => x"98",
          3799 => x"79",
          3800 => x"80",
          3801 => x"83",
          3802 => x"59",
          3803 => x"ff",
          3804 => x"1b",
          3805 => x"1b",
          3806 => x"1b",
          3807 => x"1b",
          3808 => x"1b",
          3809 => x"83",
          3810 => x"52",
          3811 => x"51",
          3812 => x"3f",
          3813 => x"04",
          3814 => x"02",
          3815 => x"82",
          3816 => x"70",
          3817 => x"58",
          3818 => x"c0",
          3819 => x"75",
          3820 => x"38",
          3821 => x"94",
          3822 => x"70",
          3823 => x"81",
          3824 => x"52",
          3825 => x"8c",
          3826 => x"2a",
          3827 => x"51",
          3828 => x"38",
          3829 => x"70",
          3830 => x"51",
          3831 => x"8d",
          3832 => x"2a",
          3833 => x"51",
          3834 => x"be",
          3835 => x"ff",
          3836 => x"c0",
          3837 => x"70",
          3838 => x"38",
          3839 => x"90",
          3840 => x"0c",
          3841 => x"f8",
          3842 => x"0d",
          3843 => x"0d",
          3844 => x"33",
          3845 => x"9f",
          3846 => x"52",
          3847 => x"98",
          3848 => x"0d",
          3849 => x"0d",
          3850 => x"33",
          3851 => x"2e",
          3852 => x"87",
          3853 => x"8d",
          3854 => x"82",
          3855 => x"70",
          3856 => x"58",
          3857 => x"94",
          3858 => x"80",
          3859 => x"87",
          3860 => x"53",
          3861 => x"96",
          3862 => x"06",
          3863 => x"72",
          3864 => x"38",
          3865 => x"70",
          3866 => x"53",
          3867 => x"74",
          3868 => x"81",
          3869 => x"72",
          3870 => x"38",
          3871 => x"70",
          3872 => x"53",
          3873 => x"38",
          3874 => x"06",
          3875 => x"94",
          3876 => x"80",
          3877 => x"87",
          3878 => x"54",
          3879 => x"80",
          3880 => x"f8",
          3881 => x"0d",
          3882 => x"0d",
          3883 => x"74",
          3884 => x"ff",
          3885 => x"57",
          3886 => x"80",
          3887 => x"81",
          3888 => x"15",
          3889 => x"33",
          3890 => x"06",
          3891 => x"58",
          3892 => x"84",
          3893 => x"2e",
          3894 => x"c0",
          3895 => x"70",
          3896 => x"2a",
          3897 => x"53",
          3898 => x"80",
          3899 => x"71",
          3900 => x"81",
          3901 => x"70",
          3902 => x"81",
          3903 => x"06",
          3904 => x"80",
          3905 => x"71",
          3906 => x"81",
          3907 => x"70",
          3908 => x"74",
          3909 => x"51",
          3910 => x"80",
          3911 => x"2e",
          3912 => x"c0",
          3913 => x"77",
          3914 => x"17",
          3915 => x"81",
          3916 => x"53",
          3917 => x"86",
          3918 => x"d4",
          3919 => x"3d",
          3920 => x"3d",
          3921 => x"98",
          3922 => x"ff",
          3923 => x"87",
          3924 => x"51",
          3925 => x"86",
          3926 => x"94",
          3927 => x"08",
          3928 => x"70",
          3929 => x"51",
          3930 => x"2e",
          3931 => x"81",
          3932 => x"87",
          3933 => x"52",
          3934 => x"86",
          3935 => x"94",
          3936 => x"08",
          3937 => x"06",
          3938 => x"0c",
          3939 => x"0d",
          3940 => x"3f",
          3941 => x"08",
          3942 => x"82",
          3943 => x"04",
          3944 => x"82",
          3945 => x"70",
          3946 => x"52",
          3947 => x"94",
          3948 => x"80",
          3949 => x"87",
          3950 => x"52",
          3951 => x"82",
          3952 => x"06",
          3953 => x"ff",
          3954 => x"2e",
          3955 => x"81",
          3956 => x"87",
          3957 => x"52",
          3958 => x"86",
          3959 => x"94",
          3960 => x"08",
          3961 => x"70",
          3962 => x"53",
          3963 => x"d4",
          3964 => x"3d",
          3965 => x"3d",
          3966 => x"9e",
          3967 => x"9c",
          3968 => x"51",
          3969 => x"2e",
          3970 => x"87",
          3971 => x"08",
          3972 => x"0c",
          3973 => x"a8",
          3974 => x"a0",
          3975 => x"9e",
          3976 => x"d3",
          3977 => x"c0",
          3978 => x"82",
          3979 => x"87",
          3980 => x"08",
          3981 => x"0c",
          3982 => x"a0",
          3983 => x"b0",
          3984 => x"9e",
          3985 => x"d3",
          3986 => x"c0",
          3987 => x"82",
          3988 => x"87",
          3989 => x"08",
          3990 => x"0c",
          3991 => x"b8",
          3992 => x"c0",
          3993 => x"9e",
          3994 => x"d3",
          3995 => x"c0",
          3996 => x"82",
          3997 => x"87",
          3998 => x"08",
          3999 => x"0c",
          4000 => x"80",
          4001 => x"82",
          4002 => x"87",
          4003 => x"08",
          4004 => x"0c",
          4005 => x"88",
          4006 => x"d8",
          4007 => x"9e",
          4008 => x"d3",
          4009 => x"0b",
          4010 => x"34",
          4011 => x"c0",
          4012 => x"70",
          4013 => x"06",
          4014 => x"70",
          4015 => x"38",
          4016 => x"82",
          4017 => x"80",
          4018 => x"9e",
          4019 => x"88",
          4020 => x"51",
          4021 => x"80",
          4022 => x"81",
          4023 => x"d3",
          4024 => x"0b",
          4025 => x"90",
          4026 => x"80",
          4027 => x"52",
          4028 => x"2e",
          4029 => x"52",
          4030 => x"e3",
          4031 => x"87",
          4032 => x"08",
          4033 => x"80",
          4034 => x"52",
          4035 => x"83",
          4036 => x"71",
          4037 => x"34",
          4038 => x"c0",
          4039 => x"70",
          4040 => x"06",
          4041 => x"70",
          4042 => x"38",
          4043 => x"82",
          4044 => x"80",
          4045 => x"9e",
          4046 => x"90",
          4047 => x"51",
          4048 => x"80",
          4049 => x"81",
          4050 => x"d3",
          4051 => x"0b",
          4052 => x"90",
          4053 => x"80",
          4054 => x"52",
          4055 => x"2e",
          4056 => x"52",
          4057 => x"e7",
          4058 => x"87",
          4059 => x"08",
          4060 => x"80",
          4061 => x"52",
          4062 => x"83",
          4063 => x"71",
          4064 => x"34",
          4065 => x"c0",
          4066 => x"70",
          4067 => x"06",
          4068 => x"70",
          4069 => x"38",
          4070 => x"82",
          4071 => x"80",
          4072 => x"9e",
          4073 => x"80",
          4074 => x"51",
          4075 => x"80",
          4076 => x"81",
          4077 => x"d3",
          4078 => x"0b",
          4079 => x"90",
          4080 => x"80",
          4081 => x"52",
          4082 => x"83",
          4083 => x"71",
          4084 => x"34",
          4085 => x"90",
          4086 => x"80",
          4087 => x"2a",
          4088 => x"70",
          4089 => x"34",
          4090 => x"c0",
          4091 => x"70",
          4092 => x"51",
          4093 => x"80",
          4094 => x"81",
          4095 => x"d3",
          4096 => x"c0",
          4097 => x"70",
          4098 => x"70",
          4099 => x"51",
          4100 => x"d3",
          4101 => x"0b",
          4102 => x"90",
          4103 => x"06",
          4104 => x"70",
          4105 => x"38",
          4106 => x"82",
          4107 => x"87",
          4108 => x"08",
          4109 => x"51",
          4110 => x"d3",
          4111 => x"3d",
          4112 => x"3d",
          4113 => x"f4",
          4114 => x"8d",
          4115 => x"e0",
          4116 => x"80",
          4117 => x"82",
          4118 => x"ff",
          4119 => x"82",
          4120 => x"ff",
          4121 => x"82",
          4122 => x"54",
          4123 => x"94",
          4124 => x"bc",
          4125 => x"c0",
          4126 => x"52",
          4127 => x"51",
          4128 => x"3f",
          4129 => x"33",
          4130 => x"2e",
          4131 => x"d3",
          4132 => x"d3",
          4133 => x"54",
          4134 => x"d0",
          4135 => x"b9",
          4136 => x"e4",
          4137 => x"80",
          4138 => x"82",
          4139 => x"82",
          4140 => x"11",
          4141 => x"bd",
          4142 => x"92",
          4143 => x"d3",
          4144 => x"73",
          4145 => x"38",
          4146 => x"08",
          4147 => x"08",
          4148 => x"82",
          4149 => x"ff",
          4150 => x"82",
          4151 => x"54",
          4152 => x"94",
          4153 => x"ac",
          4154 => x"b0",
          4155 => x"52",
          4156 => x"51",
          4157 => x"3f",
          4158 => x"33",
          4159 => x"2e",
          4160 => x"d3",
          4161 => x"82",
          4162 => x"ff",
          4163 => x"82",
          4164 => x"54",
          4165 => x"8e",
          4166 => x"f0",
          4167 => x"be",
          4168 => x"91",
          4169 => x"d3",
          4170 => x"73",
          4171 => x"38",
          4172 => x"33",
          4173 => x"80",
          4174 => x"9d",
          4175 => x"e1",
          4176 => x"80",
          4177 => x"82",
          4178 => x"ff",
          4179 => x"82",
          4180 => x"54",
          4181 => x"89",
          4182 => x"b4",
          4183 => x"84",
          4184 => x"e8",
          4185 => x"80",
          4186 => x"82",
          4187 => x"ff",
          4188 => x"82",
          4189 => x"54",
          4190 => x"89",
          4191 => x"cc",
          4192 => x"e0",
          4193 => x"ea",
          4194 => x"80",
          4195 => x"82",
          4196 => x"ff",
          4197 => x"82",
          4198 => x"ff",
          4199 => x"82",
          4200 => x"52",
          4201 => x"51",
          4202 => x"3f",
          4203 => x"08",
          4204 => x"90",
          4205 => x"a1",
          4206 => x"cc",
          4207 => x"c0",
          4208 => x"90",
          4209 => x"c0",
          4210 => x"ac",
          4211 => x"d3",
          4212 => x"82",
          4213 => x"ff",
          4214 => x"82",
          4215 => x"56",
          4216 => x"52",
          4217 => x"c7",
          4218 => x"f8",
          4219 => x"c0",
          4220 => x"31",
          4221 => x"d4",
          4222 => x"82",
          4223 => x"ff",
          4224 => x"82",
          4225 => x"54",
          4226 => x"a9",
          4227 => x"d8",
          4228 => x"84",
          4229 => x"51",
          4230 => x"82",
          4231 => x"bd",
          4232 => x"76",
          4233 => x"54",
          4234 => x"08",
          4235 => x"bc",
          4236 => x"a5",
          4237 => x"e2",
          4238 => x"80",
          4239 => x"82",
          4240 => x"56",
          4241 => x"52",
          4242 => x"e3",
          4243 => x"f8",
          4244 => x"c0",
          4245 => x"31",
          4246 => x"d4",
          4247 => x"82",
          4248 => x"ff",
          4249 => x"8a",
          4250 => x"9a",
          4251 => x"0d",
          4252 => x"0d",
          4253 => x"33",
          4254 => x"71",
          4255 => x"38",
          4256 => x"82",
          4257 => x"52",
          4258 => x"82",
          4259 => x"9d",
          4260 => x"9c",
          4261 => x"82",
          4262 => x"91",
          4263 => x"ac",
          4264 => x"82",
          4265 => x"85",
          4266 => x"b8",
          4267 => x"a9",
          4268 => x"0d",
          4269 => x"80",
          4270 => x"0b",
          4271 => x"84",
          4272 => x"d3",
          4273 => x"c0",
          4274 => x"04",
          4275 => x"76",
          4276 => x"98",
          4277 => x"2b",
          4278 => x"72",
          4279 => x"82",
          4280 => x"51",
          4281 => x"80",
          4282 => x"c4",
          4283 => x"53",
          4284 => x"9c",
          4285 => x"c0",
          4286 => x"02",
          4287 => x"05",
          4288 => x"52",
          4289 => x"72",
          4290 => x"06",
          4291 => x"53",
          4292 => x"f8",
          4293 => x"0d",
          4294 => x"0d",
          4295 => x"05",
          4296 => x"71",
          4297 => x"54",
          4298 => x"b1",
          4299 => x"dc",
          4300 => x"51",
          4301 => x"3f",
          4302 => x"08",
          4303 => x"ff",
          4304 => x"82",
          4305 => x"52",
          4306 => x"ac",
          4307 => x"33",
          4308 => x"72",
          4309 => x"81",
          4310 => x"cc",
          4311 => x"ff",
          4312 => x"74",
          4313 => x"3d",
          4314 => x"3d",
          4315 => x"84",
          4316 => x"33",
          4317 => x"bb",
          4318 => x"d4",
          4319 => x"84",
          4320 => x"f8",
          4321 => x"51",
          4322 => x"58",
          4323 => x"2e",
          4324 => x"51",
          4325 => x"82",
          4326 => x"70",
          4327 => x"d3",
          4328 => x"19",
          4329 => x"56",
          4330 => x"3f",
          4331 => x"08",
          4332 => x"d4",
          4333 => x"84",
          4334 => x"f8",
          4335 => x"51",
          4336 => x"80",
          4337 => x"75",
          4338 => x"74",
          4339 => x"96",
          4340 => x"d0",
          4341 => x"55",
          4342 => x"d0",
          4343 => x"ff",
          4344 => x"75",
          4345 => x"80",
          4346 => x"d0",
          4347 => x"2e",
          4348 => x"d4",
          4349 => x"75",
          4350 => x"38",
          4351 => x"33",
          4352 => x"38",
          4353 => x"05",
          4354 => x"78",
          4355 => x"80",
          4356 => x"82",
          4357 => x"52",
          4358 => x"a0",
          4359 => x"d4",
          4360 => x"80",
          4361 => x"8c",
          4362 => x"fd",
          4363 => x"d3",
          4364 => x"54",
          4365 => x"71",
          4366 => x"38",
          4367 => x"d1",
          4368 => x"0c",
          4369 => x"14",
          4370 => x"80",
          4371 => x"80",
          4372 => x"d0",
          4373 => x"cc",
          4374 => x"80",
          4375 => x"71",
          4376 => x"87",
          4377 => x"cc",
          4378 => x"a5",
          4379 => x"82",
          4380 => x"85",
          4381 => x"dc",
          4382 => x"57",
          4383 => x"d4",
          4384 => x"80",
          4385 => x"82",
          4386 => x"80",
          4387 => x"d4",
          4388 => x"80",
          4389 => x"3d",
          4390 => x"81",
          4391 => x"82",
          4392 => x"80",
          4393 => x"75",
          4394 => x"da",
          4395 => x"f8",
          4396 => x"0b",
          4397 => x"08",
          4398 => x"82",
          4399 => x"ff",
          4400 => x"55",
          4401 => x"34",
          4402 => x"52",
          4403 => x"c5",
          4404 => x"ff",
          4405 => x"74",
          4406 => x"81",
          4407 => x"38",
          4408 => x"04",
          4409 => x"aa",
          4410 => x"3d",
          4411 => x"81",
          4412 => x"80",
          4413 => x"cc",
          4414 => x"f4",
          4415 => x"d4",
          4416 => x"95",
          4417 => x"82",
          4418 => x"54",
          4419 => x"52",
          4420 => x"52",
          4421 => x"d9",
          4422 => x"f8",
          4423 => x"a5",
          4424 => x"ff",
          4425 => x"82",
          4426 => x"81",
          4427 => x"80",
          4428 => x"f8",
          4429 => x"38",
          4430 => x"08",
          4431 => x"17",
          4432 => x"74",
          4433 => x"70",
          4434 => x"07",
          4435 => x"55",
          4436 => x"2e",
          4437 => x"ff",
          4438 => x"d4",
          4439 => x"11",
          4440 => x"80",
          4441 => x"82",
          4442 => x"80",
          4443 => x"82",
          4444 => x"ff",
          4445 => x"78",
          4446 => x"81",
          4447 => x"75",
          4448 => x"ff",
          4449 => x"79",
          4450 => x"fa",
          4451 => x"08",
          4452 => x"f8",
          4453 => x"80",
          4454 => x"d4",
          4455 => x"3d",
          4456 => x"3d",
          4457 => x"71",
          4458 => x"33",
          4459 => x"58",
          4460 => x"09",
          4461 => x"38",
          4462 => x"05",
          4463 => x"27",
          4464 => x"17",
          4465 => x"71",
          4466 => x"55",
          4467 => x"09",
          4468 => x"38",
          4469 => x"ea",
          4470 => x"73",
          4471 => x"d4",
          4472 => x"08",
          4473 => x"b0",
          4474 => x"d4",
          4475 => x"79",
          4476 => x"51",
          4477 => x"3f",
          4478 => x"08",
          4479 => x"84",
          4480 => x"74",
          4481 => x"38",
          4482 => x"88",
          4483 => x"fc",
          4484 => x"39",
          4485 => x"8c",
          4486 => x"53",
          4487 => x"c4",
          4488 => x"d4",
          4489 => x"2e",
          4490 => x"1b",
          4491 => x"77",
          4492 => x"3f",
          4493 => x"08",
          4494 => x"55",
          4495 => x"74",
          4496 => x"81",
          4497 => x"ff",
          4498 => x"82",
          4499 => x"8b",
          4500 => x"73",
          4501 => x"0c",
          4502 => x"04",
          4503 => x"b0",
          4504 => x"3d",
          4505 => x"08",
          4506 => x"80",
          4507 => x"34",
          4508 => x"33",
          4509 => x"08",
          4510 => x"81",
          4511 => x"82",
          4512 => x"55",
          4513 => x"38",
          4514 => x"80",
          4515 => x"38",
          4516 => x"06",
          4517 => x"80",
          4518 => x"38",
          4519 => x"87",
          4520 => x"f8",
          4521 => x"cc",
          4522 => x"f8",
          4523 => x"81",
          4524 => x"53",
          4525 => x"d4",
          4526 => x"80",
          4527 => x"82",
          4528 => x"80",
          4529 => x"82",
          4530 => x"ff",
          4531 => x"80",
          4532 => x"d4",
          4533 => x"82",
          4534 => x"53",
          4535 => x"90",
          4536 => x"54",
          4537 => x"3f",
          4538 => x"08",
          4539 => x"f8",
          4540 => x"09",
          4541 => x"d0",
          4542 => x"f8",
          4543 => x"ae",
          4544 => x"d4",
          4545 => x"80",
          4546 => x"f8",
          4547 => x"38",
          4548 => x"08",
          4549 => x"17",
          4550 => x"74",
          4551 => x"74",
          4552 => x"52",
          4553 => x"c2",
          4554 => x"70",
          4555 => x"5c",
          4556 => x"27",
          4557 => x"5b",
          4558 => x"09",
          4559 => x"97",
          4560 => x"75",
          4561 => x"34",
          4562 => x"82",
          4563 => x"80",
          4564 => x"f9",
          4565 => x"3d",
          4566 => x"3f",
          4567 => x"08",
          4568 => x"98",
          4569 => x"78",
          4570 => x"38",
          4571 => x"06",
          4572 => x"33",
          4573 => x"70",
          4574 => x"ec",
          4575 => x"98",
          4576 => x"2c",
          4577 => x"05",
          4578 => x"82",
          4579 => x"70",
          4580 => x"33",
          4581 => x"51",
          4582 => x"59",
          4583 => x"56",
          4584 => x"80",
          4585 => x"74",
          4586 => x"74",
          4587 => x"29",
          4588 => x"05",
          4589 => x"51",
          4590 => x"24",
          4591 => x"76",
          4592 => x"77",
          4593 => x"3f",
          4594 => x"08",
          4595 => x"54",
          4596 => x"d7",
          4597 => x"ec",
          4598 => x"56",
          4599 => x"81",
          4600 => x"81",
          4601 => x"70",
          4602 => x"81",
          4603 => x"51",
          4604 => x"26",
          4605 => x"53",
          4606 => x"51",
          4607 => x"82",
          4608 => x"81",
          4609 => x"73",
          4610 => x"39",
          4611 => x"80",
          4612 => x"38",
          4613 => x"74",
          4614 => x"34",
          4615 => x"70",
          4616 => x"ec",
          4617 => x"98",
          4618 => x"2c",
          4619 => x"70",
          4620 => x"c2",
          4621 => x"5e",
          4622 => x"57",
          4623 => x"74",
          4624 => x"81",
          4625 => x"38",
          4626 => x"14",
          4627 => x"80",
          4628 => x"b4",
          4629 => x"82",
          4630 => x"92",
          4631 => x"ec",
          4632 => x"82",
          4633 => x"78",
          4634 => x"75",
          4635 => x"54",
          4636 => x"fd",
          4637 => x"84",
          4638 => x"fc",
          4639 => x"08",
          4640 => x"bc",
          4641 => x"7e",
          4642 => x"38",
          4643 => x"33",
          4644 => x"27",
          4645 => x"98",
          4646 => x"2c",
          4647 => x"75",
          4648 => x"74",
          4649 => x"33",
          4650 => x"74",
          4651 => x"29",
          4652 => x"05",
          4653 => x"82",
          4654 => x"56",
          4655 => x"39",
          4656 => x"33",
          4657 => x"54",
          4658 => x"bc",
          4659 => x"54",
          4660 => x"74",
          4661 => x"b8",
          4662 => x"7e",
          4663 => x"81",
          4664 => x"82",
          4665 => x"82",
          4666 => x"70",
          4667 => x"29",
          4668 => x"05",
          4669 => x"82",
          4670 => x"5a",
          4671 => x"74",
          4672 => x"38",
          4673 => x"08",
          4674 => x"70",
          4675 => x"ff",
          4676 => x"74",
          4677 => x"29",
          4678 => x"05",
          4679 => x"82",
          4680 => x"56",
          4681 => x"75",
          4682 => x"82",
          4683 => x"70",
          4684 => x"98",
          4685 => x"b8",
          4686 => x"56",
          4687 => x"25",
          4688 => x"82",
          4689 => x"52",
          4690 => x"a0",
          4691 => x"81",
          4692 => x"81",
          4693 => x"70",
          4694 => x"ec",
          4695 => x"51",
          4696 => x"24",
          4697 => x"ee",
          4698 => x"34",
          4699 => x"1b",
          4700 => x"bc",
          4701 => x"82",
          4702 => x"f3",
          4703 => x"fd",
          4704 => x"bc",
          4705 => x"ff",
          4706 => x"73",
          4707 => x"c6",
          4708 => x"b8",
          4709 => x"54",
          4710 => x"b8",
          4711 => x"54",
          4712 => x"bc",
          4713 => x"dc",
          4714 => x"51",
          4715 => x"3f",
          4716 => x"33",
          4717 => x"70",
          4718 => x"ec",
          4719 => x"51",
          4720 => x"74",
          4721 => x"74",
          4722 => x"14",
          4723 => x"82",
          4724 => x"52",
          4725 => x"ff",
          4726 => x"74",
          4727 => x"29",
          4728 => x"05",
          4729 => x"82",
          4730 => x"58",
          4731 => x"75",
          4732 => x"82",
          4733 => x"52",
          4734 => x"9f",
          4735 => x"ec",
          4736 => x"98",
          4737 => x"2c",
          4738 => x"33",
          4739 => x"57",
          4740 => x"fa",
          4741 => x"f0",
          4742 => x"88",
          4743 => x"93",
          4744 => x"80",
          4745 => x"80",
          4746 => x"98",
          4747 => x"b8",
          4748 => x"55",
          4749 => x"de",
          4750 => x"39",
          4751 => x"33",
          4752 => x"80",
          4753 => x"f0",
          4754 => x"8a",
          4755 => x"e3",
          4756 => x"b8",
          4757 => x"f6",
          4758 => x"d4",
          4759 => x"ff",
          4760 => x"96",
          4761 => x"b8",
          4762 => x"80",
          4763 => x"81",
          4764 => x"79",
          4765 => x"3f",
          4766 => x"7a",
          4767 => x"82",
          4768 => x"80",
          4769 => x"b8",
          4770 => x"d4",
          4771 => x"3d",
          4772 => x"ec",
          4773 => x"73",
          4774 => x"ba",
          4775 => x"dc",
          4776 => x"51",
          4777 => x"3f",
          4778 => x"33",
          4779 => x"73",
          4780 => x"34",
          4781 => x"06",
          4782 => x"82",
          4783 => x"82",
          4784 => x"55",
          4785 => x"2e",
          4786 => x"ff",
          4787 => x"82",
          4788 => x"74",
          4789 => x"98",
          4790 => x"ff",
          4791 => x"55",
          4792 => x"ad",
          4793 => x"54",
          4794 => x"74",
          4795 => x"dc",
          4796 => x"33",
          4797 => x"bb",
          4798 => x"80",
          4799 => x"80",
          4800 => x"98",
          4801 => x"b8",
          4802 => x"55",
          4803 => x"d5",
          4804 => x"dc",
          4805 => x"51",
          4806 => x"3f",
          4807 => x"33",
          4808 => x"70",
          4809 => x"ec",
          4810 => x"51",
          4811 => x"74",
          4812 => x"38",
          4813 => x"08",
          4814 => x"ff",
          4815 => x"74",
          4816 => x"29",
          4817 => x"05",
          4818 => x"82",
          4819 => x"58",
          4820 => x"75",
          4821 => x"f7",
          4822 => x"ec",
          4823 => x"81",
          4824 => x"ec",
          4825 => x"56",
          4826 => x"27",
          4827 => x"82",
          4828 => x"52",
          4829 => x"73",
          4830 => x"34",
          4831 => x"33",
          4832 => x"9c",
          4833 => x"ec",
          4834 => x"81",
          4835 => x"ec",
          4836 => x"56",
          4837 => x"26",
          4838 => x"ba",
          4839 => x"bc",
          4840 => x"82",
          4841 => x"ee",
          4842 => x"0b",
          4843 => x"34",
          4844 => x"ec",
          4845 => x"9e",
          4846 => x"38",
          4847 => x"08",
          4848 => x"2e",
          4849 => x"51",
          4850 => x"3f",
          4851 => x"08",
          4852 => x"34",
          4853 => x"08",
          4854 => x"81",
          4855 => x"52",
          4856 => x"a6",
          4857 => x"5b",
          4858 => x"7a",
          4859 => x"d3",
          4860 => x"11",
          4861 => x"74",
          4862 => x"38",
          4863 => x"a4",
          4864 => x"d4",
          4865 => x"ec",
          4866 => x"d4",
          4867 => x"ff",
          4868 => x"53",
          4869 => x"51",
          4870 => x"3f",
          4871 => x"80",
          4872 => x"08",
          4873 => x"2e",
          4874 => x"74",
          4875 => x"d6",
          4876 => x"7a",
          4877 => x"81",
          4878 => x"82",
          4879 => x"55",
          4880 => x"a4",
          4881 => x"ff",
          4882 => x"82",
          4883 => x"82",
          4884 => x"82",
          4885 => x"81",
          4886 => x"05",
          4887 => x"79",
          4888 => x"82",
          4889 => x"39",
          4890 => x"82",
          4891 => x"70",
          4892 => x"74",
          4893 => x"38",
          4894 => x"a3",
          4895 => x"d4",
          4896 => x"ec",
          4897 => x"d4",
          4898 => x"ff",
          4899 => x"53",
          4900 => x"51",
          4901 => x"3f",
          4902 => x"73",
          4903 => x"5b",
          4904 => x"82",
          4905 => x"74",
          4906 => x"ec",
          4907 => x"ec",
          4908 => x"79",
          4909 => x"3f",
          4910 => x"82",
          4911 => x"70",
          4912 => x"82",
          4913 => x"59",
          4914 => x"77",
          4915 => x"38",
          4916 => x"08",
          4917 => x"54",
          4918 => x"bc",
          4919 => x"70",
          4920 => x"ff",
          4921 => x"f4",
          4922 => x"ec",
          4923 => x"73",
          4924 => x"e2",
          4925 => x"dc",
          4926 => x"51",
          4927 => x"3f",
          4928 => x"33",
          4929 => x"73",
          4930 => x"34",
          4931 => x"f9",
          4932 => x"ff",
          4933 => x"d4",
          4934 => x"80",
          4935 => x"ec",
          4936 => x"80",
          4937 => x"86",
          4938 => x"ff",
          4939 => x"82",
          4940 => x"54",
          4941 => x"74",
          4942 => x"76",
          4943 => x"82",
          4944 => x"54",
          4945 => x"34",
          4946 => x"34",
          4947 => x"08",
          4948 => x"15",
          4949 => x"15",
          4950 => x"f0",
          4951 => x"ec",
          4952 => x"fe",
          4953 => x"70",
          4954 => x"06",
          4955 => x"58",
          4956 => x"74",
          4957 => x"73",
          4958 => x"82",
          4959 => x"70",
          4960 => x"d4",
          4961 => x"f8",
          4962 => x"55",
          4963 => x"34",
          4964 => x"34",
          4965 => x"04",
          4966 => x"73",
          4967 => x"84",
          4968 => x"38",
          4969 => x"2a",
          4970 => x"83",
          4971 => x"51",
          4972 => x"82",
          4973 => x"83",
          4974 => x"f9",
          4975 => x"a6",
          4976 => x"84",
          4977 => x"22",
          4978 => x"d4",
          4979 => x"83",
          4980 => x"74",
          4981 => x"11",
          4982 => x"12",
          4983 => x"2b",
          4984 => x"05",
          4985 => x"71",
          4986 => x"06",
          4987 => x"2a",
          4988 => x"59",
          4989 => x"57",
          4990 => x"71",
          4991 => x"81",
          4992 => x"d4",
          4993 => x"75",
          4994 => x"54",
          4995 => x"34",
          4996 => x"34",
          4997 => x"08",
          4998 => x"33",
          4999 => x"71",
          5000 => x"70",
          5001 => x"ff",
          5002 => x"52",
          5003 => x"05",
          5004 => x"ff",
          5005 => x"2a",
          5006 => x"71",
          5007 => x"72",
          5008 => x"53",
          5009 => x"34",
          5010 => x"08",
          5011 => x"76",
          5012 => x"17",
          5013 => x"0d",
          5014 => x"0d",
          5015 => x"08",
          5016 => x"9e",
          5017 => x"83",
          5018 => x"86",
          5019 => x"12",
          5020 => x"2b",
          5021 => x"07",
          5022 => x"52",
          5023 => x"05",
          5024 => x"85",
          5025 => x"88",
          5026 => x"88",
          5027 => x"56",
          5028 => x"13",
          5029 => x"13",
          5030 => x"f0",
          5031 => x"84",
          5032 => x"12",
          5033 => x"2b",
          5034 => x"07",
          5035 => x"52",
          5036 => x"12",
          5037 => x"33",
          5038 => x"07",
          5039 => x"54",
          5040 => x"70",
          5041 => x"73",
          5042 => x"82",
          5043 => x"13",
          5044 => x"12",
          5045 => x"2b",
          5046 => x"ff",
          5047 => x"88",
          5048 => x"53",
          5049 => x"73",
          5050 => x"14",
          5051 => x"0d",
          5052 => x"0d",
          5053 => x"22",
          5054 => x"08",
          5055 => x"71",
          5056 => x"81",
          5057 => x"88",
          5058 => x"88",
          5059 => x"33",
          5060 => x"71",
          5061 => x"90",
          5062 => x"5f",
          5063 => x"5a",
          5064 => x"54",
          5065 => x"80",
          5066 => x"51",
          5067 => x"82",
          5068 => x"70",
          5069 => x"81",
          5070 => x"8b",
          5071 => x"2b",
          5072 => x"70",
          5073 => x"33",
          5074 => x"07",
          5075 => x"8f",
          5076 => x"51",
          5077 => x"53",
          5078 => x"72",
          5079 => x"2a",
          5080 => x"82",
          5081 => x"83",
          5082 => x"d4",
          5083 => x"16",
          5084 => x"12",
          5085 => x"2b",
          5086 => x"07",
          5087 => x"55",
          5088 => x"33",
          5089 => x"71",
          5090 => x"70",
          5091 => x"06",
          5092 => x"57",
          5093 => x"52",
          5094 => x"71",
          5095 => x"88",
          5096 => x"fb",
          5097 => x"d4",
          5098 => x"84",
          5099 => x"22",
          5100 => x"72",
          5101 => x"33",
          5102 => x"71",
          5103 => x"83",
          5104 => x"5b",
          5105 => x"52",
          5106 => x"33",
          5107 => x"71",
          5108 => x"02",
          5109 => x"05",
          5110 => x"70",
          5111 => x"51",
          5112 => x"71",
          5113 => x"81",
          5114 => x"d4",
          5115 => x"15",
          5116 => x"12",
          5117 => x"2b",
          5118 => x"07",
          5119 => x"52",
          5120 => x"12",
          5121 => x"33",
          5122 => x"07",
          5123 => x"54",
          5124 => x"70",
          5125 => x"72",
          5126 => x"82",
          5127 => x"14",
          5128 => x"83",
          5129 => x"88",
          5130 => x"d4",
          5131 => x"54",
          5132 => x"04",
          5133 => x"7b",
          5134 => x"08",
          5135 => x"70",
          5136 => x"06",
          5137 => x"53",
          5138 => x"82",
          5139 => x"76",
          5140 => x"11",
          5141 => x"83",
          5142 => x"8b",
          5143 => x"2b",
          5144 => x"70",
          5145 => x"33",
          5146 => x"71",
          5147 => x"53",
          5148 => x"53",
          5149 => x"59",
          5150 => x"25",
          5151 => x"80",
          5152 => x"51",
          5153 => x"81",
          5154 => x"14",
          5155 => x"33",
          5156 => x"71",
          5157 => x"76",
          5158 => x"2a",
          5159 => x"58",
          5160 => x"14",
          5161 => x"ff",
          5162 => x"87",
          5163 => x"d4",
          5164 => x"19",
          5165 => x"85",
          5166 => x"88",
          5167 => x"88",
          5168 => x"5b",
          5169 => x"84",
          5170 => x"85",
          5171 => x"d4",
          5172 => x"53",
          5173 => x"14",
          5174 => x"87",
          5175 => x"d4",
          5176 => x"76",
          5177 => x"75",
          5178 => x"82",
          5179 => x"18",
          5180 => x"12",
          5181 => x"2b",
          5182 => x"80",
          5183 => x"88",
          5184 => x"55",
          5185 => x"74",
          5186 => x"15",
          5187 => x"0d",
          5188 => x"0d",
          5189 => x"d4",
          5190 => x"38",
          5191 => x"71",
          5192 => x"38",
          5193 => x"8c",
          5194 => x"0d",
          5195 => x"0d",
          5196 => x"58",
          5197 => x"82",
          5198 => x"83",
          5199 => x"82",
          5200 => x"84",
          5201 => x"12",
          5202 => x"2b",
          5203 => x"59",
          5204 => x"81",
          5205 => x"75",
          5206 => x"cb",
          5207 => x"29",
          5208 => x"81",
          5209 => x"88",
          5210 => x"81",
          5211 => x"79",
          5212 => x"ff",
          5213 => x"7f",
          5214 => x"51",
          5215 => x"77",
          5216 => x"38",
          5217 => x"85",
          5218 => x"5a",
          5219 => x"33",
          5220 => x"71",
          5221 => x"57",
          5222 => x"38",
          5223 => x"ff",
          5224 => x"7a",
          5225 => x"80",
          5226 => x"82",
          5227 => x"11",
          5228 => x"12",
          5229 => x"2b",
          5230 => x"ff",
          5231 => x"52",
          5232 => x"55",
          5233 => x"83",
          5234 => x"80",
          5235 => x"26",
          5236 => x"74",
          5237 => x"2e",
          5238 => x"77",
          5239 => x"81",
          5240 => x"75",
          5241 => x"3f",
          5242 => x"82",
          5243 => x"79",
          5244 => x"f7",
          5245 => x"d4",
          5246 => x"1c",
          5247 => x"87",
          5248 => x"8b",
          5249 => x"2b",
          5250 => x"5e",
          5251 => x"7a",
          5252 => x"ff",
          5253 => x"88",
          5254 => x"56",
          5255 => x"15",
          5256 => x"ff",
          5257 => x"85",
          5258 => x"d4",
          5259 => x"83",
          5260 => x"72",
          5261 => x"33",
          5262 => x"71",
          5263 => x"70",
          5264 => x"5b",
          5265 => x"56",
          5266 => x"19",
          5267 => x"19",
          5268 => x"f0",
          5269 => x"84",
          5270 => x"12",
          5271 => x"2b",
          5272 => x"07",
          5273 => x"55",
          5274 => x"78",
          5275 => x"76",
          5276 => x"82",
          5277 => x"70",
          5278 => x"84",
          5279 => x"12",
          5280 => x"2b",
          5281 => x"2a",
          5282 => x"52",
          5283 => x"84",
          5284 => x"85",
          5285 => x"d4",
          5286 => x"84",
          5287 => x"82",
          5288 => x"8d",
          5289 => x"fe",
          5290 => x"52",
          5291 => x"08",
          5292 => x"db",
          5293 => x"71",
          5294 => x"38",
          5295 => x"ed",
          5296 => x"f8",
          5297 => x"82",
          5298 => x"84",
          5299 => x"ee",
          5300 => x"66",
          5301 => x"70",
          5302 => x"d4",
          5303 => x"2e",
          5304 => x"84",
          5305 => x"3f",
          5306 => x"7e",
          5307 => x"3f",
          5308 => x"08",
          5309 => x"39",
          5310 => x"7b",
          5311 => x"3f",
          5312 => x"ba",
          5313 => x"f5",
          5314 => x"d4",
          5315 => x"ff",
          5316 => x"d4",
          5317 => x"71",
          5318 => x"70",
          5319 => x"06",
          5320 => x"73",
          5321 => x"81",
          5322 => x"88",
          5323 => x"75",
          5324 => x"ff",
          5325 => x"88",
          5326 => x"73",
          5327 => x"70",
          5328 => x"33",
          5329 => x"07",
          5330 => x"53",
          5331 => x"48",
          5332 => x"54",
          5333 => x"56",
          5334 => x"80",
          5335 => x"76",
          5336 => x"06",
          5337 => x"83",
          5338 => x"42",
          5339 => x"33",
          5340 => x"71",
          5341 => x"70",
          5342 => x"70",
          5343 => x"33",
          5344 => x"71",
          5345 => x"53",
          5346 => x"56",
          5347 => x"25",
          5348 => x"75",
          5349 => x"ff",
          5350 => x"54",
          5351 => x"81",
          5352 => x"18",
          5353 => x"2e",
          5354 => x"8f",
          5355 => x"f6",
          5356 => x"83",
          5357 => x"58",
          5358 => x"7f",
          5359 => x"74",
          5360 => x"78",
          5361 => x"3f",
          5362 => x"7f",
          5363 => x"75",
          5364 => x"38",
          5365 => x"11",
          5366 => x"33",
          5367 => x"07",
          5368 => x"f4",
          5369 => x"52",
          5370 => x"b7",
          5371 => x"f8",
          5372 => x"ff",
          5373 => x"7c",
          5374 => x"2b",
          5375 => x"08",
          5376 => x"53",
          5377 => x"91",
          5378 => x"d4",
          5379 => x"84",
          5380 => x"ff",
          5381 => x"5c",
          5382 => x"60",
          5383 => x"74",
          5384 => x"38",
          5385 => x"c9",
          5386 => x"f0",
          5387 => x"11",
          5388 => x"33",
          5389 => x"07",
          5390 => x"f4",
          5391 => x"52",
          5392 => x"df",
          5393 => x"f8",
          5394 => x"ff",
          5395 => x"7c",
          5396 => x"2b",
          5397 => x"08",
          5398 => x"53",
          5399 => x"90",
          5400 => x"d4",
          5401 => x"84",
          5402 => x"05",
          5403 => x"73",
          5404 => x"06",
          5405 => x"7b",
          5406 => x"f9",
          5407 => x"d4",
          5408 => x"82",
          5409 => x"80",
          5410 => x"7d",
          5411 => x"82",
          5412 => x"51",
          5413 => x"3f",
          5414 => x"98",
          5415 => x"7a",
          5416 => x"38",
          5417 => x"52",
          5418 => x"8f",
          5419 => x"83",
          5420 => x"f0",
          5421 => x"05",
          5422 => x"3f",
          5423 => x"82",
          5424 => x"94",
          5425 => x"fc",
          5426 => x"77",
          5427 => x"54",
          5428 => x"82",
          5429 => x"55",
          5430 => x"08",
          5431 => x"38",
          5432 => x"52",
          5433 => x"08",
          5434 => x"a6",
          5435 => x"d4",
          5436 => x"3d",
          5437 => x"3d",
          5438 => x"05",
          5439 => x"52",
          5440 => x"87",
          5441 => x"f4",
          5442 => x"71",
          5443 => x"0c",
          5444 => x"04",
          5445 => x"02",
          5446 => x"02",
          5447 => x"05",
          5448 => x"83",
          5449 => x"26",
          5450 => x"72",
          5451 => x"c0",
          5452 => x"53",
          5453 => x"74",
          5454 => x"38",
          5455 => x"73",
          5456 => x"c0",
          5457 => x"51",
          5458 => x"85",
          5459 => x"98",
          5460 => x"52",
          5461 => x"82",
          5462 => x"70",
          5463 => x"38",
          5464 => x"8c",
          5465 => x"ec",
          5466 => x"fc",
          5467 => x"52",
          5468 => x"87",
          5469 => x"08",
          5470 => x"2e",
          5471 => x"82",
          5472 => x"34",
          5473 => x"13",
          5474 => x"82",
          5475 => x"86",
          5476 => x"f3",
          5477 => x"62",
          5478 => x"05",
          5479 => x"57",
          5480 => x"83",
          5481 => x"fe",
          5482 => x"d4",
          5483 => x"06",
          5484 => x"71",
          5485 => x"71",
          5486 => x"2b",
          5487 => x"80",
          5488 => x"92",
          5489 => x"c0",
          5490 => x"41",
          5491 => x"5a",
          5492 => x"87",
          5493 => x"0c",
          5494 => x"84",
          5495 => x"08",
          5496 => x"70",
          5497 => x"53",
          5498 => x"2e",
          5499 => x"08",
          5500 => x"70",
          5501 => x"34",
          5502 => x"80",
          5503 => x"53",
          5504 => x"2e",
          5505 => x"53",
          5506 => x"26",
          5507 => x"80",
          5508 => x"87",
          5509 => x"08",
          5510 => x"38",
          5511 => x"8c",
          5512 => x"80",
          5513 => x"78",
          5514 => x"99",
          5515 => x"0c",
          5516 => x"8c",
          5517 => x"08",
          5518 => x"51",
          5519 => x"38",
          5520 => x"8d",
          5521 => x"17",
          5522 => x"81",
          5523 => x"53",
          5524 => x"2e",
          5525 => x"fc",
          5526 => x"52",
          5527 => x"7d",
          5528 => x"ed",
          5529 => x"80",
          5530 => x"71",
          5531 => x"38",
          5532 => x"53",
          5533 => x"f8",
          5534 => x"0d",
          5535 => x"0d",
          5536 => x"02",
          5537 => x"05",
          5538 => x"58",
          5539 => x"80",
          5540 => x"fc",
          5541 => x"d4",
          5542 => x"06",
          5543 => x"71",
          5544 => x"81",
          5545 => x"38",
          5546 => x"2b",
          5547 => x"80",
          5548 => x"92",
          5549 => x"c0",
          5550 => x"40",
          5551 => x"5a",
          5552 => x"c0",
          5553 => x"76",
          5554 => x"76",
          5555 => x"75",
          5556 => x"2a",
          5557 => x"51",
          5558 => x"80",
          5559 => x"7a",
          5560 => x"5c",
          5561 => x"81",
          5562 => x"81",
          5563 => x"06",
          5564 => x"80",
          5565 => x"87",
          5566 => x"08",
          5567 => x"38",
          5568 => x"8c",
          5569 => x"80",
          5570 => x"77",
          5571 => x"99",
          5572 => x"0c",
          5573 => x"8c",
          5574 => x"08",
          5575 => x"51",
          5576 => x"38",
          5577 => x"8d",
          5578 => x"70",
          5579 => x"84",
          5580 => x"5b",
          5581 => x"2e",
          5582 => x"fc",
          5583 => x"52",
          5584 => x"7d",
          5585 => x"f8",
          5586 => x"80",
          5587 => x"71",
          5588 => x"38",
          5589 => x"53",
          5590 => x"f8",
          5591 => x"0d",
          5592 => x"0d",
          5593 => x"05",
          5594 => x"02",
          5595 => x"05",
          5596 => x"54",
          5597 => x"fe",
          5598 => x"f8",
          5599 => x"53",
          5600 => x"80",
          5601 => x"0b",
          5602 => x"8c",
          5603 => x"71",
          5604 => x"dc",
          5605 => x"24",
          5606 => x"84",
          5607 => x"92",
          5608 => x"54",
          5609 => x"8d",
          5610 => x"39",
          5611 => x"80",
          5612 => x"cb",
          5613 => x"70",
          5614 => x"81",
          5615 => x"52",
          5616 => x"8a",
          5617 => x"98",
          5618 => x"71",
          5619 => x"c0",
          5620 => x"52",
          5621 => x"81",
          5622 => x"c0",
          5623 => x"53",
          5624 => x"82",
          5625 => x"71",
          5626 => x"39",
          5627 => x"39",
          5628 => x"77",
          5629 => x"81",
          5630 => x"72",
          5631 => x"84",
          5632 => x"73",
          5633 => x"0c",
          5634 => x"04",
          5635 => x"74",
          5636 => x"71",
          5637 => x"2b",
          5638 => x"f8",
          5639 => x"84",
          5640 => x"fd",
          5641 => x"83",
          5642 => x"12",
          5643 => x"2b",
          5644 => x"07",
          5645 => x"70",
          5646 => x"2b",
          5647 => x"07",
          5648 => x"0c",
          5649 => x"56",
          5650 => x"3d",
          5651 => x"3d",
          5652 => x"84",
          5653 => x"22",
          5654 => x"72",
          5655 => x"54",
          5656 => x"2a",
          5657 => x"34",
          5658 => x"04",
          5659 => x"73",
          5660 => x"70",
          5661 => x"05",
          5662 => x"88",
          5663 => x"72",
          5664 => x"54",
          5665 => x"2a",
          5666 => x"70",
          5667 => x"34",
          5668 => x"51",
          5669 => x"83",
          5670 => x"fe",
          5671 => x"75",
          5672 => x"51",
          5673 => x"92",
          5674 => x"81",
          5675 => x"73",
          5676 => x"55",
          5677 => x"51",
          5678 => x"3d",
          5679 => x"3d",
          5680 => x"76",
          5681 => x"72",
          5682 => x"05",
          5683 => x"11",
          5684 => x"38",
          5685 => x"04",
          5686 => x"78",
          5687 => x"56",
          5688 => x"81",
          5689 => x"74",
          5690 => x"56",
          5691 => x"31",
          5692 => x"52",
          5693 => x"80",
          5694 => x"71",
          5695 => x"38",
          5696 => x"f8",
          5697 => x"0d",
          5698 => x"0d",
          5699 => x"51",
          5700 => x"73",
          5701 => x"81",
          5702 => x"33",
          5703 => x"38",
          5704 => x"d4",
          5705 => x"3d",
          5706 => x"0b",
          5707 => x"0c",
          5708 => x"0d",
          5709 => x"70",
          5710 => x"52",
          5711 => x"55",
          5712 => x"3f",
          5713 => x"d4",
          5714 => x"38",
          5715 => x"98",
          5716 => x"52",
          5717 => x"f7",
          5718 => x"d4",
          5719 => x"ff",
          5720 => x"72",
          5721 => x"38",
          5722 => x"72",
          5723 => x"d4",
          5724 => x"3d",
          5725 => x"3d",
          5726 => x"80",
          5727 => x"33",
          5728 => x"7a",
          5729 => x"38",
          5730 => x"16",
          5731 => x"16",
          5732 => x"17",
          5733 => x"f9",
          5734 => x"d4",
          5735 => x"2e",
          5736 => x"b7",
          5737 => x"f8",
          5738 => x"34",
          5739 => x"70",
          5740 => x"31",
          5741 => x"59",
          5742 => x"77",
          5743 => x"82",
          5744 => x"74",
          5745 => x"81",
          5746 => x"81",
          5747 => x"53",
          5748 => x"16",
          5749 => x"a5",
          5750 => x"81",
          5751 => x"d4",
          5752 => x"3d",
          5753 => x"3d",
          5754 => x"56",
          5755 => x"74",
          5756 => x"2e",
          5757 => x"51",
          5758 => x"82",
          5759 => x"57",
          5760 => x"08",
          5761 => x"54",
          5762 => x"16",
          5763 => x"33",
          5764 => x"3f",
          5765 => x"08",
          5766 => x"38",
          5767 => x"57",
          5768 => x"0c",
          5769 => x"f8",
          5770 => x"0d",
          5771 => x"0d",
          5772 => x"57",
          5773 => x"82",
          5774 => x"58",
          5775 => x"08",
          5776 => x"76",
          5777 => x"83",
          5778 => x"06",
          5779 => x"84",
          5780 => x"78",
          5781 => x"81",
          5782 => x"38",
          5783 => x"82",
          5784 => x"52",
          5785 => x"52",
          5786 => x"3f",
          5787 => x"52",
          5788 => x"51",
          5789 => x"84",
          5790 => x"d2",
          5791 => x"fb",
          5792 => x"8a",
          5793 => x"52",
          5794 => x"51",
          5795 => x"94",
          5796 => x"84",
          5797 => x"fb",
          5798 => x"17",
          5799 => x"a4",
          5800 => x"c8",
          5801 => x"08",
          5802 => x"b4",
          5803 => x"55",
          5804 => x"81",
          5805 => x"f7",
          5806 => x"84",
          5807 => x"53",
          5808 => x"17",
          5809 => x"99",
          5810 => x"f8",
          5811 => x"83",
          5812 => x"77",
          5813 => x"0c",
          5814 => x"04",
          5815 => x"77",
          5816 => x"12",
          5817 => x"55",
          5818 => x"56",
          5819 => x"8d",
          5820 => x"22",
          5821 => x"b0",
          5822 => x"57",
          5823 => x"d4",
          5824 => x"3d",
          5825 => x"3d",
          5826 => x"70",
          5827 => x"57",
          5828 => x"81",
          5829 => x"9c",
          5830 => x"81",
          5831 => x"74",
          5832 => x"72",
          5833 => x"f5",
          5834 => x"24",
          5835 => x"81",
          5836 => x"81",
          5837 => x"83",
          5838 => x"38",
          5839 => x"76",
          5840 => x"70",
          5841 => x"16",
          5842 => x"74",
          5843 => x"96",
          5844 => x"f8",
          5845 => x"38",
          5846 => x"06",
          5847 => x"33",
          5848 => x"89",
          5849 => x"08",
          5850 => x"54",
          5851 => x"fc",
          5852 => x"d4",
          5853 => x"fe",
          5854 => x"ff",
          5855 => x"11",
          5856 => x"2b",
          5857 => x"81",
          5858 => x"2a",
          5859 => x"51",
          5860 => x"e2",
          5861 => x"ff",
          5862 => x"da",
          5863 => x"2a",
          5864 => x"05",
          5865 => x"fc",
          5866 => x"d4",
          5867 => x"c6",
          5868 => x"83",
          5869 => x"05",
          5870 => x"f8",
          5871 => x"d4",
          5872 => x"ff",
          5873 => x"ae",
          5874 => x"2a",
          5875 => x"05",
          5876 => x"fc",
          5877 => x"d4",
          5878 => x"38",
          5879 => x"83",
          5880 => x"05",
          5881 => x"f8",
          5882 => x"d4",
          5883 => x"0a",
          5884 => x"39",
          5885 => x"82",
          5886 => x"89",
          5887 => x"f8",
          5888 => x"7c",
          5889 => x"56",
          5890 => x"77",
          5891 => x"38",
          5892 => x"08",
          5893 => x"38",
          5894 => x"72",
          5895 => x"9d",
          5896 => x"24",
          5897 => x"81",
          5898 => x"82",
          5899 => x"83",
          5900 => x"38",
          5901 => x"76",
          5902 => x"70",
          5903 => x"18",
          5904 => x"76",
          5905 => x"9e",
          5906 => x"f8",
          5907 => x"d4",
          5908 => x"d9",
          5909 => x"ff",
          5910 => x"05",
          5911 => x"81",
          5912 => x"54",
          5913 => x"80",
          5914 => x"77",
          5915 => x"f0",
          5916 => x"8f",
          5917 => x"51",
          5918 => x"34",
          5919 => x"17",
          5920 => x"2a",
          5921 => x"05",
          5922 => x"fa",
          5923 => x"d4",
          5924 => x"82",
          5925 => x"81",
          5926 => x"83",
          5927 => x"b8",
          5928 => x"2a",
          5929 => x"8f",
          5930 => x"2a",
          5931 => x"f0",
          5932 => x"06",
          5933 => x"72",
          5934 => x"ec",
          5935 => x"2a",
          5936 => x"05",
          5937 => x"fa",
          5938 => x"d4",
          5939 => x"82",
          5940 => x"80",
          5941 => x"83",
          5942 => x"52",
          5943 => x"fe",
          5944 => x"b8",
          5945 => x"e6",
          5946 => x"76",
          5947 => x"17",
          5948 => x"75",
          5949 => x"3f",
          5950 => x"08",
          5951 => x"f8",
          5952 => x"77",
          5953 => x"77",
          5954 => x"fc",
          5955 => x"b8",
          5956 => x"51",
          5957 => x"8b",
          5958 => x"f8",
          5959 => x"06",
          5960 => x"72",
          5961 => x"3f",
          5962 => x"17",
          5963 => x"d4",
          5964 => x"3d",
          5965 => x"3d",
          5966 => x"7e",
          5967 => x"56",
          5968 => x"75",
          5969 => x"74",
          5970 => x"27",
          5971 => x"80",
          5972 => x"ff",
          5973 => x"75",
          5974 => x"3f",
          5975 => x"08",
          5976 => x"f8",
          5977 => x"38",
          5978 => x"54",
          5979 => x"81",
          5980 => x"39",
          5981 => x"08",
          5982 => x"39",
          5983 => x"51",
          5984 => x"82",
          5985 => x"58",
          5986 => x"08",
          5987 => x"c7",
          5988 => x"f8",
          5989 => x"d2",
          5990 => x"f8",
          5991 => x"cf",
          5992 => x"74",
          5993 => x"fc",
          5994 => x"d4",
          5995 => x"38",
          5996 => x"fe",
          5997 => x"08",
          5998 => x"74",
          5999 => x"38",
          6000 => x"17",
          6001 => x"33",
          6002 => x"73",
          6003 => x"77",
          6004 => x"26",
          6005 => x"80",
          6006 => x"d4",
          6007 => x"3d",
          6008 => x"3d",
          6009 => x"71",
          6010 => x"5b",
          6011 => x"90",
          6012 => x"77",
          6013 => x"38",
          6014 => x"78",
          6015 => x"81",
          6016 => x"79",
          6017 => x"f9",
          6018 => x"55",
          6019 => x"f8",
          6020 => x"e0",
          6021 => x"f8",
          6022 => x"d4",
          6023 => x"2e",
          6024 => x"9c",
          6025 => x"d4",
          6026 => x"82",
          6027 => x"58",
          6028 => x"70",
          6029 => x"80",
          6030 => x"38",
          6031 => x"09",
          6032 => x"e2",
          6033 => x"56",
          6034 => x"76",
          6035 => x"82",
          6036 => x"7a",
          6037 => x"3f",
          6038 => x"d4",
          6039 => x"2e",
          6040 => x"86",
          6041 => x"f8",
          6042 => x"d4",
          6043 => x"70",
          6044 => x"07",
          6045 => x"7c",
          6046 => x"f8",
          6047 => x"51",
          6048 => x"81",
          6049 => x"d4",
          6050 => x"2e",
          6051 => x"17",
          6052 => x"74",
          6053 => x"73",
          6054 => x"27",
          6055 => x"58",
          6056 => x"80",
          6057 => x"56",
          6058 => x"9c",
          6059 => x"26",
          6060 => x"56",
          6061 => x"81",
          6062 => x"52",
          6063 => x"c6",
          6064 => x"f8",
          6065 => x"b8",
          6066 => x"82",
          6067 => x"81",
          6068 => x"06",
          6069 => x"d4",
          6070 => x"82",
          6071 => x"09",
          6072 => x"72",
          6073 => x"70",
          6074 => x"51",
          6075 => x"80",
          6076 => x"78",
          6077 => x"06",
          6078 => x"73",
          6079 => x"39",
          6080 => x"52",
          6081 => x"f7",
          6082 => x"f8",
          6083 => x"f8",
          6084 => x"82",
          6085 => x"07",
          6086 => x"55",
          6087 => x"2e",
          6088 => x"80",
          6089 => x"75",
          6090 => x"76",
          6091 => x"3f",
          6092 => x"08",
          6093 => x"38",
          6094 => x"0c",
          6095 => x"fe",
          6096 => x"08",
          6097 => x"74",
          6098 => x"ff",
          6099 => x"0c",
          6100 => x"81",
          6101 => x"84",
          6102 => x"39",
          6103 => x"81",
          6104 => x"8c",
          6105 => x"8c",
          6106 => x"f8",
          6107 => x"39",
          6108 => x"55",
          6109 => x"f8",
          6110 => x"0d",
          6111 => x"0d",
          6112 => x"55",
          6113 => x"82",
          6114 => x"58",
          6115 => x"d4",
          6116 => x"d8",
          6117 => x"74",
          6118 => x"3f",
          6119 => x"08",
          6120 => x"08",
          6121 => x"59",
          6122 => x"77",
          6123 => x"70",
          6124 => x"8a",
          6125 => x"84",
          6126 => x"56",
          6127 => x"58",
          6128 => x"97",
          6129 => x"75",
          6130 => x"52",
          6131 => x"51",
          6132 => x"82",
          6133 => x"80",
          6134 => x"8a",
          6135 => x"32",
          6136 => x"72",
          6137 => x"2a",
          6138 => x"56",
          6139 => x"f8",
          6140 => x"0d",
          6141 => x"0d",
          6142 => x"08",
          6143 => x"74",
          6144 => x"26",
          6145 => x"74",
          6146 => x"72",
          6147 => x"74",
          6148 => x"88",
          6149 => x"73",
          6150 => x"33",
          6151 => x"27",
          6152 => x"16",
          6153 => x"9b",
          6154 => x"2a",
          6155 => x"88",
          6156 => x"58",
          6157 => x"80",
          6158 => x"16",
          6159 => x"0c",
          6160 => x"8a",
          6161 => x"89",
          6162 => x"72",
          6163 => x"38",
          6164 => x"51",
          6165 => x"82",
          6166 => x"54",
          6167 => x"08",
          6168 => x"38",
          6169 => x"d4",
          6170 => x"8b",
          6171 => x"08",
          6172 => x"08",
          6173 => x"82",
          6174 => x"74",
          6175 => x"cb",
          6176 => x"75",
          6177 => x"3f",
          6178 => x"08",
          6179 => x"73",
          6180 => x"98",
          6181 => x"82",
          6182 => x"2e",
          6183 => x"39",
          6184 => x"39",
          6185 => x"13",
          6186 => x"74",
          6187 => x"16",
          6188 => x"18",
          6189 => x"77",
          6190 => x"0c",
          6191 => x"04",
          6192 => x"7a",
          6193 => x"12",
          6194 => x"59",
          6195 => x"80",
          6196 => x"86",
          6197 => x"98",
          6198 => x"14",
          6199 => x"55",
          6200 => x"81",
          6201 => x"83",
          6202 => x"77",
          6203 => x"81",
          6204 => x"0c",
          6205 => x"55",
          6206 => x"76",
          6207 => x"17",
          6208 => x"74",
          6209 => x"9b",
          6210 => x"39",
          6211 => x"ff",
          6212 => x"2a",
          6213 => x"81",
          6214 => x"52",
          6215 => x"e6",
          6216 => x"f8",
          6217 => x"55",
          6218 => x"d4",
          6219 => x"80",
          6220 => x"55",
          6221 => x"08",
          6222 => x"f4",
          6223 => x"08",
          6224 => x"08",
          6225 => x"38",
          6226 => x"77",
          6227 => x"84",
          6228 => x"39",
          6229 => x"52",
          6230 => x"86",
          6231 => x"f8",
          6232 => x"55",
          6233 => x"08",
          6234 => x"c4",
          6235 => x"82",
          6236 => x"81",
          6237 => x"81",
          6238 => x"f8",
          6239 => x"b0",
          6240 => x"f8",
          6241 => x"51",
          6242 => x"82",
          6243 => x"a0",
          6244 => x"15",
          6245 => x"75",
          6246 => x"3f",
          6247 => x"08",
          6248 => x"76",
          6249 => x"77",
          6250 => x"9c",
          6251 => x"55",
          6252 => x"f8",
          6253 => x"0d",
          6254 => x"0d",
          6255 => x"08",
          6256 => x"80",
          6257 => x"fc",
          6258 => x"d4",
          6259 => x"82",
          6260 => x"80",
          6261 => x"d4",
          6262 => x"98",
          6263 => x"78",
          6264 => x"3f",
          6265 => x"08",
          6266 => x"f8",
          6267 => x"38",
          6268 => x"08",
          6269 => x"70",
          6270 => x"58",
          6271 => x"2e",
          6272 => x"83",
          6273 => x"82",
          6274 => x"55",
          6275 => x"81",
          6276 => x"07",
          6277 => x"2e",
          6278 => x"16",
          6279 => x"2e",
          6280 => x"88",
          6281 => x"82",
          6282 => x"56",
          6283 => x"51",
          6284 => x"82",
          6285 => x"54",
          6286 => x"08",
          6287 => x"9b",
          6288 => x"2e",
          6289 => x"83",
          6290 => x"73",
          6291 => x"0c",
          6292 => x"04",
          6293 => x"76",
          6294 => x"54",
          6295 => x"82",
          6296 => x"83",
          6297 => x"76",
          6298 => x"53",
          6299 => x"2e",
          6300 => x"90",
          6301 => x"51",
          6302 => x"82",
          6303 => x"90",
          6304 => x"53",
          6305 => x"f8",
          6306 => x"0d",
          6307 => x"0d",
          6308 => x"83",
          6309 => x"54",
          6310 => x"55",
          6311 => x"3f",
          6312 => x"51",
          6313 => x"2e",
          6314 => x"8b",
          6315 => x"2a",
          6316 => x"51",
          6317 => x"86",
          6318 => x"fd",
          6319 => x"54",
          6320 => x"53",
          6321 => x"71",
          6322 => x"05",
          6323 => x"05",
          6324 => x"05",
          6325 => x"06",
          6326 => x"51",
          6327 => x"e4",
          6328 => x"d4",
          6329 => x"3d",
          6330 => x"3d",
          6331 => x"40",
          6332 => x"08",
          6333 => x"ff",
          6334 => x"98",
          6335 => x"2e",
          6336 => x"98",
          6337 => x"7d",
          6338 => x"3f",
          6339 => x"08",
          6340 => x"f8",
          6341 => x"38",
          6342 => x"70",
          6343 => x"73",
          6344 => x"5b",
          6345 => x"8b",
          6346 => x"06",
          6347 => x"06",
          6348 => x"86",
          6349 => x"d4",
          6350 => x"73",
          6351 => x"09",
          6352 => x"38",
          6353 => x"d4",
          6354 => x"73",
          6355 => x"81",
          6356 => x"81",
          6357 => x"07",
          6358 => x"38",
          6359 => x"08",
          6360 => x"54",
          6361 => x"2e",
          6362 => x"83",
          6363 => x"75",
          6364 => x"38",
          6365 => x"81",
          6366 => x"8f",
          6367 => x"06",
          6368 => x"73",
          6369 => x"81",
          6370 => x"72",
          6371 => x"38",
          6372 => x"74",
          6373 => x"70",
          6374 => x"ac",
          6375 => x"5d",
          6376 => x"2e",
          6377 => x"81",
          6378 => x"15",
          6379 => x"73",
          6380 => x"06",
          6381 => x"8c",
          6382 => x"16",
          6383 => x"cc",
          6384 => x"f8",
          6385 => x"ff",
          6386 => x"80",
          6387 => x"33",
          6388 => x"06",
          6389 => x"05",
          6390 => x"7b",
          6391 => x"c7",
          6392 => x"75",
          6393 => x"a4",
          6394 => x"f8",
          6395 => x"ff",
          6396 => x"80",
          6397 => x"73",
          6398 => x"80",
          6399 => x"10",
          6400 => x"53",
          6401 => x"81",
          6402 => x"39",
          6403 => x"ff",
          6404 => x"06",
          6405 => x"17",
          6406 => x"27",
          6407 => x"33",
          6408 => x"70",
          6409 => x"54",
          6410 => x"2e",
          6411 => x"81",
          6412 => x"38",
          6413 => x"53",
          6414 => x"ff",
          6415 => x"ff",
          6416 => x"84",
          6417 => x"53",
          6418 => x"39",
          6419 => x"74",
          6420 => x"3f",
          6421 => x"08",
          6422 => x"53",
          6423 => x"a7",
          6424 => x"ac",
          6425 => x"39",
          6426 => x"51",
          6427 => x"82",
          6428 => x"5b",
          6429 => x"08",
          6430 => x"19",
          6431 => x"38",
          6432 => x"0b",
          6433 => x"7a",
          6434 => x"0c",
          6435 => x"04",
          6436 => x"60",
          6437 => x"59",
          6438 => x"51",
          6439 => x"82",
          6440 => x"58",
          6441 => x"08",
          6442 => x"81",
          6443 => x"5c",
          6444 => x"1a",
          6445 => x"08",
          6446 => x"ea",
          6447 => x"d4",
          6448 => x"82",
          6449 => x"83",
          6450 => x"19",
          6451 => x"57",
          6452 => x"38",
          6453 => x"f6",
          6454 => x"33",
          6455 => x"81",
          6456 => x"54",
          6457 => x"34",
          6458 => x"2e",
          6459 => x"74",
          6460 => x"81",
          6461 => x"74",
          6462 => x"38",
          6463 => x"38",
          6464 => x"09",
          6465 => x"f7",
          6466 => x"33",
          6467 => x"70",
          6468 => x"55",
          6469 => x"a1",
          6470 => x"2a",
          6471 => x"51",
          6472 => x"2e",
          6473 => x"17",
          6474 => x"bf",
          6475 => x"1c",
          6476 => x"0c",
          6477 => x"75",
          6478 => x"81",
          6479 => x"38",
          6480 => x"56",
          6481 => x"09",
          6482 => x"ac",
          6483 => x"08",
          6484 => x"5d",
          6485 => x"82",
          6486 => x"83",
          6487 => x"55",
          6488 => x"38",
          6489 => x"bf",
          6490 => x"f3",
          6491 => x"81",
          6492 => x"82",
          6493 => x"33",
          6494 => x"e5",
          6495 => x"d4",
          6496 => x"ff",
          6497 => x"79",
          6498 => x"38",
          6499 => x"26",
          6500 => x"75",
          6501 => x"b4",
          6502 => x"f8",
          6503 => x"1e",
          6504 => x"55",
          6505 => x"55",
          6506 => x"3f",
          6507 => x"f8",
          6508 => x"81",
          6509 => x"38",
          6510 => x"39",
          6511 => x"ff",
          6512 => x"06",
          6513 => x"1b",
          6514 => x"27",
          6515 => x"76",
          6516 => x"2a",
          6517 => x"51",
          6518 => x"80",
          6519 => x"73",
          6520 => x"38",
          6521 => x"70",
          6522 => x"73",
          6523 => x"1c",
          6524 => x"06",
          6525 => x"39",
          6526 => x"73",
          6527 => x"7b",
          6528 => x"51",
          6529 => x"82",
          6530 => x"81",
          6531 => x"73",
          6532 => x"38",
          6533 => x"81",
          6534 => x"95",
          6535 => x"a0",
          6536 => x"19",
          6537 => x"b0",
          6538 => x"f8",
          6539 => x"9e",
          6540 => x"5c",
          6541 => x"1a",
          6542 => x"78",
          6543 => x"3f",
          6544 => x"08",
          6545 => x"f8",
          6546 => x"fc",
          6547 => x"82",
          6548 => x"90",
          6549 => x"ee",
          6550 => x"70",
          6551 => x"33",
          6552 => x"56",
          6553 => x"55",
          6554 => x"38",
          6555 => x"08",
          6556 => x"56",
          6557 => x"2e",
          6558 => x"1d",
          6559 => x"70",
          6560 => x"5d",
          6561 => x"53",
          6562 => x"53",
          6563 => x"53",
          6564 => x"87",
          6565 => x"cb",
          6566 => x"06",
          6567 => x"2e",
          6568 => x"80",
          6569 => x"1b",
          6570 => x"8c",
          6571 => x"56",
          6572 => x"7d",
          6573 => x"e3",
          6574 => x"7b",
          6575 => x"38",
          6576 => x"22",
          6577 => x"ff",
          6578 => x"73",
          6579 => x"38",
          6580 => x"ff",
          6581 => x"59",
          6582 => x"74",
          6583 => x"10",
          6584 => x"2a",
          6585 => x"70",
          6586 => x"56",
          6587 => x"80",
          6588 => x"75",
          6589 => x"32",
          6590 => x"57",
          6591 => x"db",
          6592 => x"75",
          6593 => x"84",
          6594 => x"57",
          6595 => x"07",
          6596 => x"b9",
          6597 => x"38",
          6598 => x"73",
          6599 => x"16",
          6600 => x"84",
          6601 => x"56",
          6602 => x"94",
          6603 => x"17",
          6604 => x"74",
          6605 => x"27",
          6606 => x"33",
          6607 => x"2e",
          6608 => x"19",
          6609 => x"54",
          6610 => x"82",
          6611 => x"80",
          6612 => x"ff",
          6613 => x"74",
          6614 => x"81",
          6615 => x"15",
          6616 => x"27",
          6617 => x"19",
          6618 => x"54",
          6619 => x"3d",
          6620 => x"05",
          6621 => x"81",
          6622 => x"a0",
          6623 => x"26",
          6624 => x"17",
          6625 => x"33",
          6626 => x"75",
          6627 => x"75",
          6628 => x"79",
          6629 => x"3f",
          6630 => x"08",
          6631 => x"1b",
          6632 => x"7b",
          6633 => x"38",
          6634 => x"80",
          6635 => x"f0",
          6636 => x"f8",
          6637 => x"d4",
          6638 => x"2e",
          6639 => x"82",
          6640 => x"80",
          6641 => x"ab",
          6642 => x"80",
          6643 => x"70",
          6644 => x"81",
          6645 => x"5e",
          6646 => x"80",
          6647 => x"8d",
          6648 => x"51",
          6649 => x"3f",
          6650 => x"08",
          6651 => x"52",
          6652 => x"c5",
          6653 => x"f8",
          6654 => x"d4",
          6655 => x"9e",
          6656 => x"59",
          6657 => x"81",
          6658 => x"85",
          6659 => x"08",
          6660 => x"54",
          6661 => x"dd",
          6662 => x"f8",
          6663 => x"d4",
          6664 => x"fa",
          6665 => x"51",
          6666 => x"82",
          6667 => x"81",
          6668 => x"98",
          6669 => x"7b",
          6670 => x"3f",
          6671 => x"08",
          6672 => x"f8",
          6673 => x"38",
          6674 => x"9c",
          6675 => x"81",
          6676 => x"57",
          6677 => x"17",
          6678 => x"8b",
          6679 => x"d4",
          6680 => x"17",
          6681 => x"f8",
          6682 => x"16",
          6683 => x"3f",
          6684 => x"f3",
          6685 => x"55",
          6686 => x"ff",
          6687 => x"74",
          6688 => x"22",
          6689 => x"51",
          6690 => x"82",
          6691 => x"33",
          6692 => x"df",
          6693 => x"85",
          6694 => x"ff",
          6695 => x"57",
          6696 => x"d4",
          6697 => x"ff",
          6698 => x"38",
          6699 => x"70",
          6700 => x"73",
          6701 => x"80",
          6702 => x"77",
          6703 => x"0b",
          6704 => x"80",
          6705 => x"ef",
          6706 => x"d4",
          6707 => x"82",
          6708 => x"80",
          6709 => x"19",
          6710 => x"d7",
          6711 => x"08",
          6712 => x"e2",
          6713 => x"d4",
          6714 => x"82",
          6715 => x"ae",
          6716 => x"82",
          6717 => x"52",
          6718 => x"51",
          6719 => x"8b",
          6720 => x"52",
          6721 => x"51",
          6722 => x"9c",
          6723 => x"1b",
          6724 => x"55",
          6725 => x"16",
          6726 => x"83",
          6727 => x"55",
          6728 => x"f8",
          6729 => x"0d",
          6730 => x"0d",
          6731 => x"90",
          6732 => x"13",
          6733 => x"57",
          6734 => x"2e",
          6735 => x"52",
          6736 => x"b1",
          6737 => x"f8",
          6738 => x"d4",
          6739 => x"c9",
          6740 => x"08",
          6741 => x"e1",
          6742 => x"d4",
          6743 => x"82",
          6744 => x"ab",
          6745 => x"08",
          6746 => x"34",
          6747 => x"17",
          6748 => x"08",
          6749 => x"38",
          6750 => x"08",
          6751 => x"ee",
          6752 => x"d4",
          6753 => x"82",
          6754 => x"80",
          6755 => x"73",
          6756 => x"81",
          6757 => x"82",
          6758 => x"d4",
          6759 => x"3d",
          6760 => x"3d",
          6761 => x"71",
          6762 => x"5c",
          6763 => x"19",
          6764 => x"08",
          6765 => x"e2",
          6766 => x"08",
          6767 => x"bb",
          6768 => x"71",
          6769 => x"08",
          6770 => x"57",
          6771 => x"72",
          6772 => x"9d",
          6773 => x"14",
          6774 => x"1b",
          6775 => x"7a",
          6776 => x"d0",
          6777 => x"83",
          6778 => x"51",
          6779 => x"ff",
          6780 => x"74",
          6781 => x"39",
          6782 => x"11",
          6783 => x"31",
          6784 => x"83",
          6785 => x"90",
          6786 => x"51",
          6787 => x"3f",
          6788 => x"08",
          6789 => x"06",
          6790 => x"75",
          6791 => x"81",
          6792 => x"38",
          6793 => x"53",
          6794 => x"74",
          6795 => x"82",
          6796 => x"74",
          6797 => x"70",
          6798 => x"25",
          6799 => x"07",
          6800 => x"73",
          6801 => x"38",
          6802 => x"39",
          6803 => x"81",
          6804 => x"57",
          6805 => x"1d",
          6806 => x"11",
          6807 => x"54",
          6808 => x"f1",
          6809 => x"70",
          6810 => x"30",
          6811 => x"51",
          6812 => x"94",
          6813 => x"0b",
          6814 => x"80",
          6815 => x"58",
          6816 => x"1c",
          6817 => x"33",
          6818 => x"56",
          6819 => x"2e",
          6820 => x"85",
          6821 => x"06",
          6822 => x"e5",
          6823 => x"32",
          6824 => x"72",
          6825 => x"51",
          6826 => x"8b",
          6827 => x"72",
          6828 => x"38",
          6829 => x"81",
          6830 => x"81",
          6831 => x"76",
          6832 => x"58",
          6833 => x"57",
          6834 => x"ff",
          6835 => x"17",
          6836 => x"80",
          6837 => x"34",
          6838 => x"53",
          6839 => x"38",
          6840 => x"bf",
          6841 => x"34",
          6842 => x"e1",
          6843 => x"89",
          6844 => x"5a",
          6845 => x"2e",
          6846 => x"96",
          6847 => x"55",
          6848 => x"ff",
          6849 => x"55",
          6850 => x"aa",
          6851 => x"08",
          6852 => x"51",
          6853 => x"27",
          6854 => x"84",
          6855 => x"39",
          6856 => x"53",
          6857 => x"53",
          6858 => x"8a",
          6859 => x"70",
          6860 => x"06",
          6861 => x"76",
          6862 => x"58",
          6863 => x"81",
          6864 => x"71",
          6865 => x"55",
          6866 => x"b5",
          6867 => x"94",
          6868 => x"0b",
          6869 => x"9c",
          6870 => x"11",
          6871 => x"72",
          6872 => x"89",
          6873 => x"1c",
          6874 => x"13",
          6875 => x"34",
          6876 => x"9c",
          6877 => x"d9",
          6878 => x"d4",
          6879 => x"0c",
          6880 => x"d9",
          6881 => x"d4",
          6882 => x"19",
          6883 => x"51",
          6884 => x"82",
          6885 => x"84",
          6886 => x"3d",
          6887 => x"3d",
          6888 => x"08",
          6889 => x"64",
          6890 => x"55",
          6891 => x"2e",
          6892 => x"55",
          6893 => x"2e",
          6894 => x"80",
          6895 => x"7f",
          6896 => x"88",
          6897 => x"39",
          6898 => x"80",
          6899 => x"56",
          6900 => x"af",
          6901 => x"06",
          6902 => x"56",
          6903 => x"32",
          6904 => x"80",
          6905 => x"51",
          6906 => x"dc",
          6907 => x"1f",
          6908 => x"33",
          6909 => x"9f",
          6910 => x"ff",
          6911 => x"1f",
          6912 => x"7d",
          6913 => x"3f",
          6914 => x"08",
          6915 => x"39",
          6916 => x"08",
          6917 => x"5b",
          6918 => x"92",
          6919 => x"51",
          6920 => x"82",
          6921 => x"ff",
          6922 => x"38",
          6923 => x"0b",
          6924 => x"08",
          6925 => x"78",
          6926 => x"d4",
          6927 => x"2a",
          6928 => x"75",
          6929 => x"59",
          6930 => x"08",
          6931 => x"06",
          6932 => x"70",
          6933 => x"27",
          6934 => x"07",
          6935 => x"56",
          6936 => x"75",
          6937 => x"ae",
          6938 => x"ff",
          6939 => x"75",
          6940 => x"9c",
          6941 => x"3f",
          6942 => x"08",
          6943 => x"78",
          6944 => x"81",
          6945 => x"10",
          6946 => x"74",
          6947 => x"59",
          6948 => x"81",
          6949 => x"61",
          6950 => x"56",
          6951 => x"2e",
          6952 => x"83",
          6953 => x"73",
          6954 => x"70",
          6955 => x"25",
          6956 => x"51",
          6957 => x"38",
          6958 => x"76",
          6959 => x"57",
          6960 => x"09",
          6961 => x"38",
          6962 => x"73",
          6963 => x"38",
          6964 => x"78",
          6965 => x"81",
          6966 => x"38",
          6967 => x"54",
          6968 => x"09",
          6969 => x"c1",
          6970 => x"54",
          6971 => x"09",
          6972 => x"38",
          6973 => x"54",
          6974 => x"80",
          6975 => x"56",
          6976 => x"78",
          6977 => x"38",
          6978 => x"75",
          6979 => x"57",
          6980 => x"58",
          6981 => x"e9",
          6982 => x"07",
          6983 => x"1f",
          6984 => x"39",
          6985 => x"a8",
          6986 => x"1a",
          6987 => x"74",
          6988 => x"71",
          6989 => x"70",
          6990 => x"2a",
          6991 => x"58",
          6992 => x"ae",
          6993 => x"73",
          6994 => x"19",
          6995 => x"38",
          6996 => x"11",
          6997 => x"74",
          6998 => x"38",
          6999 => x"90",
          7000 => x"07",
          7001 => x"39",
          7002 => x"70",
          7003 => x"06",
          7004 => x"73",
          7005 => x"81",
          7006 => x"81",
          7007 => x"1b",
          7008 => x"55",
          7009 => x"2e",
          7010 => x"8f",
          7011 => x"ff",
          7012 => x"73",
          7013 => x"81",
          7014 => x"76",
          7015 => x"78",
          7016 => x"38",
          7017 => x"05",
          7018 => x"54",
          7019 => x"9d",
          7020 => x"1a",
          7021 => x"ff",
          7022 => x"80",
          7023 => x"fe",
          7024 => x"55",
          7025 => x"2e",
          7026 => x"eb",
          7027 => x"a0",
          7028 => x"51",
          7029 => x"80",
          7030 => x"88",
          7031 => x"1a",
          7032 => x"1f",
          7033 => x"75",
          7034 => x"94",
          7035 => x"2e",
          7036 => x"ae",
          7037 => x"70",
          7038 => x"51",
          7039 => x"2e",
          7040 => x"80",
          7041 => x"76",
          7042 => x"d1",
          7043 => x"73",
          7044 => x"26",
          7045 => x"5b",
          7046 => x"70",
          7047 => x"07",
          7048 => x"7e",
          7049 => x"55",
          7050 => x"2e",
          7051 => x"8b",
          7052 => x"38",
          7053 => x"8b",
          7054 => x"07",
          7055 => x"26",
          7056 => x"78",
          7057 => x"8b",
          7058 => x"81",
          7059 => x"5f",
          7060 => x"80",
          7061 => x"af",
          7062 => x"07",
          7063 => x"52",
          7064 => x"cc",
          7065 => x"d4",
          7066 => x"ff",
          7067 => x"87",
          7068 => x"06",
          7069 => x"73",
          7070 => x"38",
          7071 => x"06",
          7072 => x"11",
          7073 => x"81",
          7074 => x"a4",
          7075 => x"54",
          7076 => x"8a",
          7077 => x"07",
          7078 => x"fe",
          7079 => x"18",
          7080 => x"88",
          7081 => x"73",
          7082 => x"18",
          7083 => x"39",
          7084 => x"92",
          7085 => x"82",
          7086 => x"d4",
          7087 => x"d4",
          7088 => x"2e",
          7089 => x"df",
          7090 => x"58",
          7091 => x"ff",
          7092 => x"73",
          7093 => x"38",
          7094 => x"5c",
          7095 => x"54",
          7096 => x"8e",
          7097 => x"07",
          7098 => x"83",
          7099 => x"58",
          7100 => x"18",
          7101 => x"75",
          7102 => x"18",
          7103 => x"39",
          7104 => x"54",
          7105 => x"2e",
          7106 => x"86",
          7107 => x"a0",
          7108 => x"88",
          7109 => x"06",
          7110 => x"82",
          7111 => x"06",
          7112 => x"06",
          7113 => x"2e",
          7114 => x"83",
          7115 => x"83",
          7116 => x"06",
          7117 => x"82",
          7118 => x"81",
          7119 => x"06",
          7120 => x"9f",
          7121 => x"06",
          7122 => x"2e",
          7123 => x"90",
          7124 => x"82",
          7125 => x"06",
          7126 => x"80",
          7127 => x"76",
          7128 => x"76",
          7129 => x"7d",
          7130 => x"3f",
          7131 => x"08",
          7132 => x"56",
          7133 => x"f8",
          7134 => x"be",
          7135 => x"f8",
          7136 => x"09",
          7137 => x"e8",
          7138 => x"2a",
          7139 => x"76",
          7140 => x"51",
          7141 => x"2e",
          7142 => x"81",
          7143 => x"80",
          7144 => x"38",
          7145 => x"ab",
          7146 => x"56",
          7147 => x"74",
          7148 => x"73",
          7149 => x"56",
          7150 => x"82",
          7151 => x"06",
          7152 => x"ac",
          7153 => x"33",
          7154 => x"70",
          7155 => x"55",
          7156 => x"2e",
          7157 => x"1e",
          7158 => x"06",
          7159 => x"05",
          7160 => x"e4",
          7161 => x"d4",
          7162 => x"1f",
          7163 => x"39",
          7164 => x"f8",
          7165 => x"0d",
          7166 => x"0d",
          7167 => x"7b",
          7168 => x"73",
          7169 => x"55",
          7170 => x"2e",
          7171 => x"75",
          7172 => x"57",
          7173 => x"26",
          7174 => x"ba",
          7175 => x"70",
          7176 => x"ba",
          7177 => x"06",
          7178 => x"73",
          7179 => x"70",
          7180 => x"51",
          7181 => x"89",
          7182 => x"82",
          7183 => x"ff",
          7184 => x"56",
          7185 => x"2e",
          7186 => x"80",
          7187 => x"f0",
          7188 => x"08",
          7189 => x"76",
          7190 => x"58",
          7191 => x"81",
          7192 => x"ff",
          7193 => x"53",
          7194 => x"26",
          7195 => x"13",
          7196 => x"06",
          7197 => x"9f",
          7198 => x"99",
          7199 => x"e0",
          7200 => x"ff",
          7201 => x"72",
          7202 => x"2a",
          7203 => x"72",
          7204 => x"06",
          7205 => x"ff",
          7206 => x"30",
          7207 => x"70",
          7208 => x"07",
          7209 => x"9f",
          7210 => x"54",
          7211 => x"80",
          7212 => x"81",
          7213 => x"59",
          7214 => x"25",
          7215 => x"8b",
          7216 => x"24",
          7217 => x"76",
          7218 => x"78",
          7219 => x"82",
          7220 => x"51",
          7221 => x"f8",
          7222 => x"0d",
          7223 => x"0d",
          7224 => x"0b",
          7225 => x"ff",
          7226 => x"0c",
          7227 => x"51",
          7228 => x"84",
          7229 => x"f8",
          7230 => x"38",
          7231 => x"51",
          7232 => x"82",
          7233 => x"83",
          7234 => x"54",
          7235 => x"82",
          7236 => x"09",
          7237 => x"e3",
          7238 => x"b8",
          7239 => x"57",
          7240 => x"2e",
          7241 => x"83",
          7242 => x"74",
          7243 => x"70",
          7244 => x"25",
          7245 => x"51",
          7246 => x"38",
          7247 => x"2e",
          7248 => x"b5",
          7249 => x"82",
          7250 => x"80",
          7251 => x"cf",
          7252 => x"d4",
          7253 => x"82",
          7254 => x"80",
          7255 => x"85",
          7256 => x"b4",
          7257 => x"16",
          7258 => x"3f",
          7259 => x"08",
          7260 => x"f8",
          7261 => x"83",
          7262 => x"74",
          7263 => x"0c",
          7264 => x"04",
          7265 => x"61",
          7266 => x"80",
          7267 => x"58",
          7268 => x"0c",
          7269 => x"e1",
          7270 => x"f8",
          7271 => x"56",
          7272 => x"d4",
          7273 => x"87",
          7274 => x"d4",
          7275 => x"29",
          7276 => x"05",
          7277 => x"53",
          7278 => x"80",
          7279 => x"38",
          7280 => x"76",
          7281 => x"74",
          7282 => x"72",
          7283 => x"38",
          7284 => x"51",
          7285 => x"82",
          7286 => x"81",
          7287 => x"81",
          7288 => x"72",
          7289 => x"80",
          7290 => x"38",
          7291 => x"70",
          7292 => x"53",
          7293 => x"86",
          7294 => x"af",
          7295 => x"34",
          7296 => x"34",
          7297 => x"14",
          7298 => x"88",
          7299 => x"f8",
          7300 => x"06",
          7301 => x"54",
          7302 => x"72",
          7303 => x"76",
          7304 => x"38",
          7305 => x"70",
          7306 => x"53",
          7307 => x"85",
          7308 => x"70",
          7309 => x"5b",
          7310 => x"82",
          7311 => x"81",
          7312 => x"76",
          7313 => x"81",
          7314 => x"38",
          7315 => x"56",
          7316 => x"83",
          7317 => x"70",
          7318 => x"80",
          7319 => x"83",
          7320 => x"cb",
          7321 => x"d4",
          7322 => x"76",
          7323 => x"05",
          7324 => x"16",
          7325 => x"56",
          7326 => x"d7",
          7327 => x"8d",
          7328 => x"72",
          7329 => x"54",
          7330 => x"57",
          7331 => x"95",
          7332 => x"73",
          7333 => x"3f",
          7334 => x"08",
          7335 => x"57",
          7336 => x"89",
          7337 => x"56",
          7338 => x"d7",
          7339 => x"76",
          7340 => x"f9",
          7341 => x"76",
          7342 => x"f1",
          7343 => x"14",
          7344 => x"3f",
          7345 => x"08",
          7346 => x"06",
          7347 => x"80",
          7348 => x"06",
          7349 => x"80",
          7350 => x"ca",
          7351 => x"d4",
          7352 => x"ff",
          7353 => x"77",
          7354 => x"dc",
          7355 => x"b3",
          7356 => x"f8",
          7357 => x"a0",
          7358 => x"c8",
          7359 => x"15",
          7360 => x"14",
          7361 => x"70",
          7362 => x"51",
          7363 => x"56",
          7364 => x"84",
          7365 => x"81",
          7366 => x"71",
          7367 => x"16",
          7368 => x"53",
          7369 => x"23",
          7370 => x"8b",
          7371 => x"73",
          7372 => x"80",
          7373 => x"8d",
          7374 => x"39",
          7375 => x"51",
          7376 => x"82",
          7377 => x"53",
          7378 => x"08",
          7379 => x"72",
          7380 => x"8d",
          7381 => x"d5",
          7382 => x"14",
          7383 => x"3f",
          7384 => x"08",
          7385 => x"06",
          7386 => x"38",
          7387 => x"51",
          7388 => x"82",
          7389 => x"55",
          7390 => x"51",
          7391 => x"82",
          7392 => x"83",
          7393 => x"53",
          7394 => x"80",
          7395 => x"38",
          7396 => x"78",
          7397 => x"2a",
          7398 => x"78",
          7399 => x"8d",
          7400 => x"22",
          7401 => x"31",
          7402 => x"83",
          7403 => x"f8",
          7404 => x"d4",
          7405 => x"2e",
          7406 => x"82",
          7407 => x"80",
          7408 => x"f5",
          7409 => x"83",
          7410 => x"ff",
          7411 => x"38",
          7412 => x"9f",
          7413 => x"38",
          7414 => x"39",
          7415 => x"80",
          7416 => x"38",
          7417 => x"9c",
          7418 => x"a4",
          7419 => x"1c",
          7420 => x"0c",
          7421 => x"17",
          7422 => x"76",
          7423 => x"81",
          7424 => x"80",
          7425 => x"c8",
          7426 => x"d4",
          7427 => x"ff",
          7428 => x"8d",
          7429 => x"95",
          7430 => x"91",
          7431 => x"14",
          7432 => x"3f",
          7433 => x"08",
          7434 => x"74",
          7435 => x"a2",
          7436 => x"79",
          7437 => x"f5",
          7438 => x"ac",
          7439 => x"15",
          7440 => x"2e",
          7441 => x"10",
          7442 => x"2a",
          7443 => x"05",
          7444 => x"ff",
          7445 => x"53",
          7446 => x"a0",
          7447 => x"81",
          7448 => x"0b",
          7449 => x"ff",
          7450 => x"0c",
          7451 => x"84",
          7452 => x"83",
          7453 => x"06",
          7454 => x"80",
          7455 => x"c7",
          7456 => x"d4",
          7457 => x"ff",
          7458 => x"72",
          7459 => x"81",
          7460 => x"38",
          7461 => x"73",
          7462 => x"3f",
          7463 => x"08",
          7464 => x"82",
          7465 => x"84",
          7466 => x"b6",
          7467 => x"dc",
          7468 => x"f8",
          7469 => x"ff",
          7470 => x"82",
          7471 => x"09",
          7472 => x"c8",
          7473 => x"51",
          7474 => x"82",
          7475 => x"84",
          7476 => x"d2",
          7477 => x"06",
          7478 => x"9c",
          7479 => x"c3",
          7480 => x"f8",
          7481 => x"85",
          7482 => x"09",
          7483 => x"38",
          7484 => x"51",
          7485 => x"82",
          7486 => x"94",
          7487 => x"a4",
          7488 => x"9f",
          7489 => x"f8",
          7490 => x"0c",
          7491 => x"82",
          7492 => x"81",
          7493 => x"82",
          7494 => x"72",
          7495 => x"82",
          7496 => x"8c",
          7497 => x"0b",
          7498 => x"80",
          7499 => x"d4",
          7500 => x"3d",
          7501 => x"3d",
          7502 => x"89",
          7503 => x"2e",
          7504 => x"08",
          7505 => x"2e",
          7506 => x"33",
          7507 => x"2e",
          7508 => x"13",
          7509 => x"22",
          7510 => x"76",
          7511 => x"06",
          7512 => x"13",
          7513 => x"bf",
          7514 => x"d4",
          7515 => x"06",
          7516 => x"38",
          7517 => x"54",
          7518 => x"80",
          7519 => x"71",
          7520 => x"82",
          7521 => x"87",
          7522 => x"fa",
          7523 => x"ab",
          7524 => x"58",
          7525 => x"05",
          7526 => x"dd",
          7527 => x"80",
          7528 => x"f8",
          7529 => x"38",
          7530 => x"08",
          7531 => x"ec",
          7532 => x"08",
          7533 => x"80",
          7534 => x"80",
          7535 => x"54",
          7536 => x"84",
          7537 => x"34",
          7538 => x"75",
          7539 => x"2e",
          7540 => x"53",
          7541 => x"53",
          7542 => x"f7",
          7543 => x"d4",
          7544 => x"73",
          7545 => x"0c",
          7546 => x"04",
          7547 => x"68",
          7548 => x"80",
          7549 => x"59",
          7550 => x"78",
          7551 => x"c8",
          7552 => x"06",
          7553 => x"3d",
          7554 => x"9a",
          7555 => x"52",
          7556 => x"3f",
          7557 => x"08",
          7558 => x"f8",
          7559 => x"38",
          7560 => x"52",
          7561 => x"52",
          7562 => x"3f",
          7563 => x"08",
          7564 => x"f8",
          7565 => x"02",
          7566 => x"33",
          7567 => x"55",
          7568 => x"25",
          7569 => x"55",
          7570 => x"54",
          7571 => x"81",
          7572 => x"80",
          7573 => x"74",
          7574 => x"81",
          7575 => x"75",
          7576 => x"3f",
          7577 => x"08",
          7578 => x"02",
          7579 => x"91",
          7580 => x"81",
          7581 => x"82",
          7582 => x"06",
          7583 => x"80",
          7584 => x"88",
          7585 => x"39",
          7586 => x"58",
          7587 => x"38",
          7588 => x"70",
          7589 => x"54",
          7590 => x"81",
          7591 => x"52",
          7592 => x"b0",
          7593 => x"f8",
          7594 => x"88",
          7595 => x"62",
          7596 => x"c3",
          7597 => x"54",
          7598 => x"15",
          7599 => x"62",
          7600 => x"d7",
          7601 => x"52",
          7602 => x"51",
          7603 => x"7a",
          7604 => x"83",
          7605 => x"80",
          7606 => x"38",
          7607 => x"08",
          7608 => x"53",
          7609 => x"3d",
          7610 => x"cc",
          7611 => x"d4",
          7612 => x"82",
          7613 => x"82",
          7614 => x"39",
          7615 => x"38",
          7616 => x"33",
          7617 => x"70",
          7618 => x"55",
          7619 => x"2e",
          7620 => x"55",
          7621 => x"77",
          7622 => x"81",
          7623 => x"73",
          7624 => x"38",
          7625 => x"54",
          7626 => x"a0",
          7627 => x"82",
          7628 => x"52",
          7629 => x"ae",
          7630 => x"f8",
          7631 => x"18",
          7632 => x"55",
          7633 => x"f8",
          7634 => x"38",
          7635 => x"70",
          7636 => x"54",
          7637 => x"86",
          7638 => x"c0",
          7639 => x"b4",
          7640 => x"1b",
          7641 => x"1b",
          7642 => x"70",
          7643 => x"e4",
          7644 => x"f8",
          7645 => x"f8",
          7646 => x"0c",
          7647 => x"52",
          7648 => x"3f",
          7649 => x"08",
          7650 => x"08",
          7651 => x"77",
          7652 => x"86",
          7653 => x"1a",
          7654 => x"1a",
          7655 => x"91",
          7656 => x"0b",
          7657 => x"80",
          7658 => x"0c",
          7659 => x"70",
          7660 => x"54",
          7661 => x"81",
          7662 => x"d4",
          7663 => x"2e",
          7664 => x"82",
          7665 => x"94",
          7666 => x"17",
          7667 => x"2b",
          7668 => x"57",
          7669 => x"52",
          7670 => x"aa",
          7671 => x"f8",
          7672 => x"d4",
          7673 => x"26",
          7674 => x"55",
          7675 => x"08",
          7676 => x"81",
          7677 => x"79",
          7678 => x"31",
          7679 => x"70",
          7680 => x"25",
          7681 => x"76",
          7682 => x"81",
          7683 => x"55",
          7684 => x"38",
          7685 => x"0c",
          7686 => x"75",
          7687 => x"54",
          7688 => x"a2",
          7689 => x"7a",
          7690 => x"3f",
          7691 => x"08",
          7692 => x"55",
          7693 => x"89",
          7694 => x"f8",
          7695 => x"1a",
          7696 => x"80",
          7697 => x"54",
          7698 => x"f8",
          7699 => x"0d",
          7700 => x"0d",
          7701 => x"64",
          7702 => x"59",
          7703 => x"90",
          7704 => x"52",
          7705 => x"ce",
          7706 => x"f8",
          7707 => x"d4",
          7708 => x"38",
          7709 => x"55",
          7710 => x"86",
          7711 => x"82",
          7712 => x"19",
          7713 => x"55",
          7714 => x"80",
          7715 => x"38",
          7716 => x"0b",
          7717 => x"82",
          7718 => x"39",
          7719 => x"1a",
          7720 => x"82",
          7721 => x"19",
          7722 => x"08",
          7723 => x"7c",
          7724 => x"74",
          7725 => x"2e",
          7726 => x"94",
          7727 => x"83",
          7728 => x"56",
          7729 => x"38",
          7730 => x"22",
          7731 => x"89",
          7732 => x"55",
          7733 => x"75",
          7734 => x"19",
          7735 => x"39",
          7736 => x"52",
          7737 => x"9e",
          7738 => x"f8",
          7739 => x"75",
          7740 => x"38",
          7741 => x"ff",
          7742 => x"98",
          7743 => x"19",
          7744 => x"51",
          7745 => x"82",
          7746 => x"80",
          7747 => x"38",
          7748 => x"08",
          7749 => x"2a",
          7750 => x"80",
          7751 => x"38",
          7752 => x"8a",
          7753 => x"5c",
          7754 => x"27",
          7755 => x"7a",
          7756 => x"54",
          7757 => x"52",
          7758 => x"51",
          7759 => x"3f",
          7760 => x"08",
          7761 => x"7e",
          7762 => x"56",
          7763 => x"2e",
          7764 => x"16",
          7765 => x"55",
          7766 => x"95",
          7767 => x"53",
          7768 => x"b4",
          7769 => x"31",
          7770 => x"05",
          7771 => x"ab",
          7772 => x"2b",
          7773 => x"76",
          7774 => x"94",
          7775 => x"ff",
          7776 => x"71",
          7777 => x"7b",
          7778 => x"38",
          7779 => x"19",
          7780 => x"51",
          7781 => x"82",
          7782 => x"fd",
          7783 => x"53",
          7784 => x"83",
          7785 => x"b8",
          7786 => x"51",
          7787 => x"3f",
          7788 => x"7e",
          7789 => x"0c",
          7790 => x"1b",
          7791 => x"1c",
          7792 => x"fd",
          7793 => x"56",
          7794 => x"f8",
          7795 => x"0d",
          7796 => x"0d",
          7797 => x"64",
          7798 => x"58",
          7799 => x"90",
          7800 => x"52",
          7801 => x"ce",
          7802 => x"f8",
          7803 => x"d4",
          7804 => x"38",
          7805 => x"55",
          7806 => x"86",
          7807 => x"83",
          7808 => x"18",
          7809 => x"2a",
          7810 => x"51",
          7811 => x"56",
          7812 => x"83",
          7813 => x"39",
          7814 => x"19",
          7815 => x"83",
          7816 => x"0b",
          7817 => x"81",
          7818 => x"39",
          7819 => x"7c",
          7820 => x"74",
          7821 => x"38",
          7822 => x"7b",
          7823 => x"f2",
          7824 => x"08",
          7825 => x"06",
          7826 => x"82",
          7827 => x"8a",
          7828 => x"05",
          7829 => x"06",
          7830 => x"bf",
          7831 => x"38",
          7832 => x"55",
          7833 => x"7a",
          7834 => x"98",
          7835 => x"77",
          7836 => x"3f",
          7837 => x"08",
          7838 => x"f8",
          7839 => x"82",
          7840 => x"81",
          7841 => x"38",
          7842 => x"ff",
          7843 => x"98",
          7844 => x"18",
          7845 => x"74",
          7846 => x"7e",
          7847 => x"08",
          7848 => x"2e",
          7849 => x"8e",
          7850 => x"ff",
          7851 => x"82",
          7852 => x"fe",
          7853 => x"18",
          7854 => x"51",
          7855 => x"82",
          7856 => x"80",
          7857 => x"38",
          7858 => x"08",
          7859 => x"2a",
          7860 => x"80",
          7861 => x"38",
          7862 => x"8a",
          7863 => x"5b",
          7864 => x"27",
          7865 => x"7b",
          7866 => x"54",
          7867 => x"52",
          7868 => x"51",
          7869 => x"3f",
          7870 => x"08",
          7871 => x"7e",
          7872 => x"78",
          7873 => x"74",
          7874 => x"38",
          7875 => x"b4",
          7876 => x"31",
          7877 => x"05",
          7878 => x"51",
          7879 => x"3f",
          7880 => x"0b",
          7881 => x"78",
          7882 => x"80",
          7883 => x"18",
          7884 => x"08",
          7885 => x"7e",
          7886 => x"ba",
          7887 => x"f8",
          7888 => x"38",
          7889 => x"12",
          7890 => x"9c",
          7891 => x"18",
          7892 => x"06",
          7893 => x"31",
          7894 => x"76",
          7895 => x"7b",
          7896 => x"08",
          7897 => x"ff",
          7898 => x"82",
          7899 => x"fd",
          7900 => x"53",
          7901 => x"18",
          7902 => x"06",
          7903 => x"51",
          7904 => x"3f",
          7905 => x"0b",
          7906 => x"7b",
          7907 => x"08",
          7908 => x"76",
          7909 => x"08",
          7910 => x"1c",
          7911 => x"08",
          7912 => x"5c",
          7913 => x"83",
          7914 => x"74",
          7915 => x"fd",
          7916 => x"18",
          7917 => x"07",
          7918 => x"19",
          7919 => x"75",
          7920 => x"0c",
          7921 => x"04",
          7922 => x"7a",
          7923 => x"05",
          7924 => x"56",
          7925 => x"82",
          7926 => x"57",
          7927 => x"08",
          7928 => x"90",
          7929 => x"86",
          7930 => x"06",
          7931 => x"73",
          7932 => x"ee",
          7933 => x"08",
          7934 => x"ff",
          7935 => x"82",
          7936 => x"57",
          7937 => x"08",
          7938 => x"a4",
          7939 => x"11",
          7940 => x"55",
          7941 => x"16",
          7942 => x"08",
          7943 => x"75",
          7944 => x"e9",
          7945 => x"08",
          7946 => x"51",
          7947 => x"3f",
          7948 => x"0a",
          7949 => x"51",
          7950 => x"3f",
          7951 => x"15",
          7952 => x"8a",
          7953 => x"81",
          7954 => x"34",
          7955 => x"bb",
          7956 => x"d4",
          7957 => x"17",
          7958 => x"06",
          7959 => x"90",
          7960 => x"82",
          7961 => x"8a",
          7962 => x"fc",
          7963 => x"70",
          7964 => x"d4",
          7965 => x"f8",
          7966 => x"d4",
          7967 => x"38",
          7968 => x"05",
          7969 => x"f1",
          7970 => x"d4",
          7971 => x"82",
          7972 => x"87",
          7973 => x"f8",
          7974 => x"72",
          7975 => x"0c",
          7976 => x"04",
          7977 => x"84",
          7978 => x"cd",
          7979 => x"80",
          7980 => x"f8",
          7981 => x"38",
          7982 => x"08",
          7983 => x"34",
          7984 => x"82",
          7985 => x"83",
          7986 => x"ee",
          7987 => x"53",
          7988 => x"05",
          7989 => x"51",
          7990 => x"82",
          7991 => x"55",
          7992 => x"08",
          7993 => x"76",
          7994 => x"94",
          7995 => x"51",
          7996 => x"82",
          7997 => x"55",
          7998 => x"08",
          7999 => x"80",
          8000 => x"70",
          8001 => x"56",
          8002 => x"89",
          8003 => x"98",
          8004 => x"b2",
          8005 => x"05",
          8006 => x"2a",
          8007 => x"51",
          8008 => x"80",
          8009 => x"76",
          8010 => x"52",
          8011 => x"3f",
          8012 => x"08",
          8013 => x"8e",
          8014 => x"f8",
          8015 => x"09",
          8016 => x"38",
          8017 => x"82",
          8018 => x"94",
          8019 => x"ff",
          8020 => x"80",
          8021 => x"80",
          8022 => x"5b",
          8023 => x"34",
          8024 => x"df",
          8025 => x"05",
          8026 => x"3d",
          8027 => x"3f",
          8028 => x"08",
          8029 => x"f8",
          8030 => x"38",
          8031 => x"3d",
          8032 => x"98",
          8033 => x"d8",
          8034 => x"58",
          8035 => x"08",
          8036 => x"2e",
          8037 => x"a0",
          8038 => x"3d",
          8039 => x"c4",
          8040 => x"d4",
          8041 => x"82",
          8042 => x"82",
          8043 => x"d9",
          8044 => x"7b",
          8045 => x"ae",
          8046 => x"f8",
          8047 => x"d4",
          8048 => x"d8",
          8049 => x"3d",
          8050 => x"51",
          8051 => x"82",
          8052 => x"80",
          8053 => x"76",
          8054 => x"c4",
          8055 => x"d4",
          8056 => x"82",
          8057 => x"82",
          8058 => x"52",
          8059 => x"fa",
          8060 => x"f8",
          8061 => x"d4",
          8062 => x"38",
          8063 => x"08",
          8064 => x"c8",
          8065 => x"82",
          8066 => x"2e",
          8067 => x"52",
          8068 => x"ac",
          8069 => x"f8",
          8070 => x"d4",
          8071 => x"2e",
          8072 => x"84",
          8073 => x"06",
          8074 => x"57",
          8075 => x"76",
          8076 => x"80",
          8077 => x"b8",
          8078 => x"51",
          8079 => x"76",
          8080 => x"11",
          8081 => x"51",
          8082 => x"73",
          8083 => x"38",
          8084 => x"05",
          8085 => x"81",
          8086 => x"56",
          8087 => x"f5",
          8088 => x"54",
          8089 => x"81",
          8090 => x"80",
          8091 => x"78",
          8092 => x"55",
          8093 => x"e1",
          8094 => x"ff",
          8095 => x"58",
          8096 => x"74",
          8097 => x"75",
          8098 => x"18",
          8099 => x"08",
          8100 => x"af",
          8101 => x"f4",
          8102 => x"2e",
          8103 => x"8d",
          8104 => x"80",
          8105 => x"11",
          8106 => x"74",
          8107 => x"82",
          8108 => x"70",
          8109 => x"c6",
          8110 => x"08",
          8111 => x"5c",
          8112 => x"73",
          8113 => x"38",
          8114 => x"1a",
          8115 => x"55",
          8116 => x"38",
          8117 => x"73",
          8118 => x"38",
          8119 => x"76",
          8120 => x"74",
          8121 => x"33",
          8122 => x"05",
          8123 => x"15",
          8124 => x"ba",
          8125 => x"05",
          8126 => x"ff",
          8127 => x"06",
          8128 => x"57",
          8129 => x"e0",
          8130 => x"81",
          8131 => x"73",
          8132 => x"81",
          8133 => x"7a",
          8134 => x"38",
          8135 => x"76",
          8136 => x"0c",
          8137 => x"0d",
          8138 => x"0d",
          8139 => x"3d",
          8140 => x"71",
          8141 => x"eb",
          8142 => x"d4",
          8143 => x"82",
          8144 => x"82",
          8145 => x"15",
          8146 => x"82",
          8147 => x"15",
          8148 => x"76",
          8149 => x"90",
          8150 => x"81",
          8151 => x"06",
          8152 => x"72",
          8153 => x"56",
          8154 => x"54",
          8155 => x"17",
          8156 => x"78",
          8157 => x"38",
          8158 => x"22",
          8159 => x"59",
          8160 => x"78",
          8161 => x"76",
          8162 => x"51",
          8163 => x"3f",
          8164 => x"08",
          8165 => x"54",
          8166 => x"53",
          8167 => x"3f",
          8168 => x"08",
          8169 => x"38",
          8170 => x"75",
          8171 => x"18",
          8172 => x"31",
          8173 => x"57",
          8174 => x"b2",
          8175 => x"08",
          8176 => x"38",
          8177 => x"51",
          8178 => x"3f",
          8179 => x"08",
          8180 => x"f8",
          8181 => x"81",
          8182 => x"d4",
          8183 => x"2e",
          8184 => x"82",
          8185 => x"88",
          8186 => x"98",
          8187 => x"80",
          8188 => x"38",
          8189 => x"80",
          8190 => x"77",
          8191 => x"08",
          8192 => x"0c",
          8193 => x"70",
          8194 => x"81",
          8195 => x"5a",
          8196 => x"2e",
          8197 => x"52",
          8198 => x"bb",
          8199 => x"d4",
          8200 => x"82",
          8201 => x"95",
          8202 => x"f8",
          8203 => x"39",
          8204 => x"51",
          8205 => x"3f",
          8206 => x"08",
          8207 => x"2e",
          8208 => x"74",
          8209 => x"79",
          8210 => x"14",
          8211 => x"38",
          8212 => x"0c",
          8213 => x"94",
          8214 => x"94",
          8215 => x"83",
          8216 => x"72",
          8217 => x"38",
          8218 => x"51",
          8219 => x"3f",
          8220 => x"08",
          8221 => x"0b",
          8222 => x"82",
          8223 => x"39",
          8224 => x"16",
          8225 => x"bb",
          8226 => x"2a",
          8227 => x"08",
          8228 => x"15",
          8229 => x"15",
          8230 => x"90",
          8231 => x"16",
          8232 => x"33",
          8233 => x"53",
          8234 => x"34",
          8235 => x"06",
          8236 => x"2e",
          8237 => x"9c",
          8238 => x"85",
          8239 => x"16",
          8240 => x"72",
          8241 => x"0c",
          8242 => x"04",
          8243 => x"79",
          8244 => x"75",
          8245 => x"8b",
          8246 => x"89",
          8247 => x"52",
          8248 => x"05",
          8249 => x"3f",
          8250 => x"08",
          8251 => x"f8",
          8252 => x"38",
          8253 => x"7a",
          8254 => x"d5",
          8255 => x"d4",
          8256 => x"82",
          8257 => x"80",
          8258 => x"16",
          8259 => x"2b",
          8260 => x"74",
          8261 => x"86",
          8262 => x"84",
          8263 => x"06",
          8264 => x"73",
          8265 => x"38",
          8266 => x"52",
          8267 => x"a4",
          8268 => x"f8",
          8269 => x"0c",
          8270 => x"14",
          8271 => x"23",
          8272 => x"51",
          8273 => x"3f",
          8274 => x"08",
          8275 => x"2e",
          8276 => x"85",
          8277 => x"86",
          8278 => x"2e",
          8279 => x"76",
          8280 => x"73",
          8281 => x"0c",
          8282 => x"04",
          8283 => x"76",
          8284 => x"05",
          8285 => x"53",
          8286 => x"82",
          8287 => x"87",
          8288 => x"f8",
          8289 => x"86",
          8290 => x"fb",
          8291 => x"79",
          8292 => x"05",
          8293 => x"56",
          8294 => x"3f",
          8295 => x"08",
          8296 => x"f8",
          8297 => x"38",
          8298 => x"82",
          8299 => x"52",
          8300 => x"bc",
          8301 => x"d4",
          8302 => x"80",
          8303 => x"d4",
          8304 => x"73",
          8305 => x"3f",
          8306 => x"08",
          8307 => x"f8",
          8308 => x"09",
          8309 => x"38",
          8310 => x"39",
          8311 => x"08",
          8312 => x"52",
          8313 => x"ba",
          8314 => x"73",
          8315 => x"d0",
          8316 => x"f8",
          8317 => x"70",
          8318 => x"07",
          8319 => x"82",
          8320 => x"06",
          8321 => x"54",
          8322 => x"f8",
          8323 => x"0d",
          8324 => x"0d",
          8325 => x"53",
          8326 => x"53",
          8327 => x"56",
          8328 => x"82",
          8329 => x"55",
          8330 => x"08",
          8331 => x"52",
          8332 => x"ea",
          8333 => x"f8",
          8334 => x"d4",
          8335 => x"38",
          8336 => x"05",
          8337 => x"2b",
          8338 => x"80",
          8339 => x"86",
          8340 => x"76",
          8341 => x"38",
          8342 => x"51",
          8343 => x"74",
          8344 => x"0c",
          8345 => x"04",
          8346 => x"63",
          8347 => x"80",
          8348 => x"ec",
          8349 => x"3d",
          8350 => x"3f",
          8351 => x"08",
          8352 => x"f8",
          8353 => x"38",
          8354 => x"73",
          8355 => x"08",
          8356 => x"13",
          8357 => x"58",
          8358 => x"26",
          8359 => x"7c",
          8360 => x"39",
          8361 => x"ce",
          8362 => x"81",
          8363 => x"d4",
          8364 => x"33",
          8365 => x"81",
          8366 => x"06",
          8367 => x"82",
          8368 => x"76",
          8369 => x"f0",
          8370 => x"b0",
          8371 => x"d4",
          8372 => x"2e",
          8373 => x"d4",
          8374 => x"2e",
          8375 => x"d4",
          8376 => x"70",
          8377 => x"08",
          8378 => x"7a",
          8379 => x"7f",
          8380 => x"54",
          8381 => x"77",
          8382 => x"80",
          8383 => x"15",
          8384 => x"f8",
          8385 => x"75",
          8386 => x"52",
          8387 => x"52",
          8388 => x"d2",
          8389 => x"f8",
          8390 => x"d4",
          8391 => x"d6",
          8392 => x"33",
          8393 => x"1a",
          8394 => x"54",
          8395 => x"09",
          8396 => x"38",
          8397 => x"ff",
          8398 => x"82",
          8399 => x"83",
          8400 => x"70",
          8401 => x"25",
          8402 => x"59",
          8403 => x"9b",
          8404 => x"51",
          8405 => x"3f",
          8406 => x"08",
          8407 => x"70",
          8408 => x"25",
          8409 => x"59",
          8410 => x"75",
          8411 => x"7a",
          8412 => x"ff",
          8413 => x"7c",
          8414 => x"94",
          8415 => x"11",
          8416 => x"56",
          8417 => x"15",
          8418 => x"d4",
          8419 => x"3d",
          8420 => x"3d",
          8421 => x"3d",
          8422 => x"70",
          8423 => x"96",
          8424 => x"f8",
          8425 => x"d4",
          8426 => x"aa",
          8427 => x"33",
          8428 => x"a2",
          8429 => x"33",
          8430 => x"70",
          8431 => x"55",
          8432 => x"73",
          8433 => x"90",
          8434 => x"08",
          8435 => x"18",
          8436 => x"82",
          8437 => x"38",
          8438 => x"08",
          8439 => x"08",
          8440 => x"ff",
          8441 => x"82",
          8442 => x"74",
          8443 => x"56",
          8444 => x"98",
          8445 => x"76",
          8446 => x"8a",
          8447 => x"f8",
          8448 => x"09",
          8449 => x"38",
          8450 => x"d4",
          8451 => x"2e",
          8452 => x"85",
          8453 => x"a4",
          8454 => x"38",
          8455 => x"d4",
          8456 => x"15",
          8457 => x"38",
          8458 => x"53",
          8459 => x"08",
          8460 => x"ff",
          8461 => x"82",
          8462 => x"56",
          8463 => x"8c",
          8464 => x"17",
          8465 => x"07",
          8466 => x"18",
          8467 => x"2e",
          8468 => x"91",
          8469 => x"55",
          8470 => x"f8",
          8471 => x"0d",
          8472 => x"0d",
          8473 => x"3d",
          8474 => x"52",
          8475 => x"da",
          8476 => x"d4",
          8477 => x"82",
          8478 => x"81",
          8479 => x"46",
          8480 => x"52",
          8481 => x"52",
          8482 => x"3f",
          8483 => x"08",
          8484 => x"f8",
          8485 => x"38",
          8486 => x"05",
          8487 => x"2a",
          8488 => x"51",
          8489 => x"55",
          8490 => x"38",
          8491 => x"54",
          8492 => x"81",
          8493 => x"80",
          8494 => x"70",
          8495 => x"54",
          8496 => x"81",
          8497 => x"52",
          8498 => x"bb",
          8499 => x"d4",
          8500 => x"84",
          8501 => x"06",
          8502 => x"73",
          8503 => x"d6",
          8504 => x"82",
          8505 => x"98",
          8506 => x"81",
          8507 => x"5a",
          8508 => x"08",
          8509 => x"8a",
          8510 => x"54",
          8511 => x"3f",
          8512 => x"08",
          8513 => x"f8",
          8514 => x"38",
          8515 => x"08",
          8516 => x"ff",
          8517 => x"82",
          8518 => x"55",
          8519 => x"08",
          8520 => x"55",
          8521 => x"82",
          8522 => x"84",
          8523 => x"82",
          8524 => x"80",
          8525 => x"51",
          8526 => x"82",
          8527 => x"82",
          8528 => x"30",
          8529 => x"f8",
          8530 => x"25",
          8531 => x"75",
          8532 => x"38",
          8533 => x"90",
          8534 => x"75",
          8535 => x"ff",
          8536 => x"82",
          8537 => x"55",
          8538 => x"78",
          8539 => x"bd",
          8540 => x"f8",
          8541 => x"82",
          8542 => x"a2",
          8543 => x"e8",
          8544 => x"53",
          8545 => x"bc",
          8546 => x"3d",
          8547 => x"3f",
          8548 => x"08",
          8549 => x"f8",
          8550 => x"38",
          8551 => x"52",
          8552 => x"52",
          8553 => x"3f",
          8554 => x"08",
          8555 => x"f8",
          8556 => x"88",
          8557 => x"39",
          8558 => x"08",
          8559 => x"81",
          8560 => x"38",
          8561 => x"05",
          8562 => x"2a",
          8563 => x"55",
          8564 => x"81",
          8565 => x"5a",
          8566 => x"3d",
          8567 => x"ff",
          8568 => x"82",
          8569 => x"75",
          8570 => x"d4",
          8571 => x"38",
          8572 => x"d4",
          8573 => x"2e",
          8574 => x"83",
          8575 => x"82",
          8576 => x"ff",
          8577 => x"06",
          8578 => x"54",
          8579 => x"73",
          8580 => x"82",
          8581 => x"52",
          8582 => x"b2",
          8583 => x"d4",
          8584 => x"82",
          8585 => x"81",
          8586 => x"53",
          8587 => x"19",
          8588 => x"8a",
          8589 => x"ae",
          8590 => x"34",
          8591 => x"0b",
          8592 => x"34",
          8593 => x"0a",
          8594 => x"19",
          8595 => x"9c",
          8596 => x"78",
          8597 => x"51",
          8598 => x"3f",
          8599 => x"b8",
          8600 => x"d8",
          8601 => x"a4",
          8602 => x"54",
          8603 => x"d9",
          8604 => x"53",
          8605 => x"11",
          8606 => x"b8",
          8607 => x"54",
          8608 => x"15",
          8609 => x"ff",
          8610 => x"82",
          8611 => x"54",
          8612 => x"08",
          8613 => x"88",
          8614 => x"64",
          8615 => x"ff",
          8616 => x"75",
          8617 => x"78",
          8618 => x"e1",
          8619 => x"90",
          8620 => x"34",
          8621 => x"0b",
          8622 => x"78",
          8623 => x"ed",
          8624 => x"f8",
          8625 => x"39",
          8626 => x"52",
          8627 => x"ac",
          8628 => x"82",
          8629 => x"9a",
          8630 => x"d8",
          8631 => x"3d",
          8632 => x"d2",
          8633 => x"53",
          8634 => x"fc",
          8635 => x"3d",
          8636 => x"3f",
          8637 => x"08",
          8638 => x"f8",
          8639 => x"38",
          8640 => x"3d",
          8641 => x"3d",
          8642 => x"c9",
          8643 => x"d4",
          8644 => x"82",
          8645 => x"82",
          8646 => x"81",
          8647 => x"81",
          8648 => x"86",
          8649 => x"af",
          8650 => x"a5",
          8651 => x"aa",
          8652 => x"05",
          8653 => x"e3",
          8654 => x"77",
          8655 => x"70",
          8656 => x"a2",
          8657 => x"3d",
          8658 => x"51",
          8659 => x"82",
          8660 => x"55",
          8661 => x"08",
          8662 => x"a1",
          8663 => x"09",
          8664 => x"38",
          8665 => x"08",
          8666 => x"88",
          8667 => x"39",
          8668 => x"08",
          8669 => x"81",
          8670 => x"38",
          8671 => x"bd",
          8672 => x"d4",
          8673 => x"82",
          8674 => x"81",
          8675 => x"56",
          8676 => x"3d",
          8677 => x"52",
          8678 => x"ff",
          8679 => x"02",
          8680 => x"8b",
          8681 => x"16",
          8682 => x"2a",
          8683 => x"51",
          8684 => x"89",
          8685 => x"07",
          8686 => x"17",
          8687 => x"81",
          8688 => x"34",
          8689 => x"70",
          8690 => x"81",
          8691 => x"55",
          8692 => x"80",
          8693 => x"64",
          8694 => x"38",
          8695 => x"51",
          8696 => x"3f",
          8697 => x"08",
          8698 => x"ff",
          8699 => x"82",
          8700 => x"f8",
          8701 => x"80",
          8702 => x"d4",
          8703 => x"78",
          8704 => x"e2",
          8705 => x"f8",
          8706 => x"d8",
          8707 => x"55",
          8708 => x"08",
          8709 => x"81",
          8710 => x"73",
          8711 => x"81",
          8712 => x"63",
          8713 => x"76",
          8714 => x"e1",
          8715 => x"81",
          8716 => x"34",
          8717 => x"d4",
          8718 => x"38",
          8719 => x"e9",
          8720 => x"f8",
          8721 => x"d4",
          8722 => x"38",
          8723 => x"a3",
          8724 => x"d4",
          8725 => x"74",
          8726 => x"0c",
          8727 => x"04",
          8728 => x"02",
          8729 => x"33",
          8730 => x"80",
          8731 => x"57",
          8732 => x"96",
          8733 => x"52",
          8734 => x"d2",
          8735 => x"d4",
          8736 => x"82",
          8737 => x"80",
          8738 => x"5a",
          8739 => x"3d",
          8740 => x"c6",
          8741 => x"d4",
          8742 => x"82",
          8743 => x"b8",
          8744 => x"cf",
          8745 => x"a0",
          8746 => x"55",
          8747 => x"75",
          8748 => x"71",
          8749 => x"33",
          8750 => x"74",
          8751 => x"57",
          8752 => x"8b",
          8753 => x"54",
          8754 => x"15",
          8755 => x"ff",
          8756 => x"82",
          8757 => x"55",
          8758 => x"f8",
          8759 => x"0d",
          8760 => x"0d",
          8761 => x"53",
          8762 => x"05",
          8763 => x"51",
          8764 => x"82",
          8765 => x"55",
          8766 => x"08",
          8767 => x"76",
          8768 => x"94",
          8769 => x"51",
          8770 => x"82",
          8771 => x"55",
          8772 => x"08",
          8773 => x"80",
          8774 => x"81",
          8775 => x"86",
          8776 => x"38",
          8777 => x"86",
          8778 => x"90",
          8779 => x"54",
          8780 => x"ff",
          8781 => x"76",
          8782 => x"83",
          8783 => x"51",
          8784 => x"3f",
          8785 => x"08",
          8786 => x"d4",
          8787 => x"3d",
          8788 => x"3d",
          8789 => x"5c",
          8790 => x"99",
          8791 => x"52",
          8792 => x"d0",
          8793 => x"d4",
          8794 => x"d4",
          8795 => x"70",
          8796 => x"08",
          8797 => x"51",
          8798 => x"80",
          8799 => x"38",
          8800 => x"06",
          8801 => x"80",
          8802 => x"38",
          8803 => x"5f",
          8804 => x"3d",
          8805 => x"ff",
          8806 => x"82",
          8807 => x"57",
          8808 => x"08",
          8809 => x"74",
          8810 => x"ff",
          8811 => x"82",
          8812 => x"57",
          8813 => x"08",
          8814 => x"d4",
          8815 => x"d4",
          8816 => x"5b",
          8817 => x"18",
          8818 => x"18",
          8819 => x"74",
          8820 => x"81",
          8821 => x"78",
          8822 => x"8b",
          8823 => x"54",
          8824 => x"75",
          8825 => x"38",
          8826 => x"1b",
          8827 => x"55",
          8828 => x"2e",
          8829 => x"39",
          8830 => x"09",
          8831 => x"38",
          8832 => x"80",
          8833 => x"70",
          8834 => x"25",
          8835 => x"80",
          8836 => x"38",
          8837 => x"bc",
          8838 => x"11",
          8839 => x"ff",
          8840 => x"82",
          8841 => x"57",
          8842 => x"08",
          8843 => x"70",
          8844 => x"80",
          8845 => x"83",
          8846 => x"80",
          8847 => x"84",
          8848 => x"a7",
          8849 => x"b8",
          8850 => x"9b",
          8851 => x"d4",
          8852 => x"0c",
          8853 => x"f8",
          8854 => x"0d",
          8855 => x"0d",
          8856 => x"3d",
          8857 => x"52",
          8858 => x"ce",
          8859 => x"d4",
          8860 => x"d4",
          8861 => x"54",
          8862 => x"08",
          8863 => x"8b",
          8864 => x"8a",
          8865 => x"58",
          8866 => x"3f",
          8867 => x"33",
          8868 => x"9f",
          8869 => x"86",
          8870 => x"9d",
          8871 => x"9d",
          8872 => x"d4",
          8873 => x"ff",
          8874 => x"c4",
          8875 => x"f8",
          8876 => x"98",
          8877 => x"52",
          8878 => x"08",
          8879 => x"3f",
          8880 => x"08",
          8881 => x"06",
          8882 => x"2e",
          8883 => x"52",
          8884 => x"51",
          8885 => x"3f",
          8886 => x"08",
          8887 => x"ff",
          8888 => x"38",
          8889 => x"88",
          8890 => x"8a",
          8891 => x"38",
          8892 => x"e7",
          8893 => x"75",
          8894 => x"74",
          8895 => x"73",
          8896 => x"05",
          8897 => x"16",
          8898 => x"70",
          8899 => x"34",
          8900 => x"70",
          8901 => x"56",
          8902 => x"fe",
          8903 => x"3d",
          8904 => x"55",
          8905 => x"2e",
          8906 => x"75",
          8907 => x"38",
          8908 => x"55",
          8909 => x"33",
          8910 => x"a0",
          8911 => x"06",
          8912 => x"16",
          8913 => x"38",
          8914 => x"42",
          8915 => x"3d",
          8916 => x"ff",
          8917 => x"82",
          8918 => x"54",
          8919 => x"08",
          8920 => x"81",
          8921 => x"ff",
          8922 => x"82",
          8923 => x"54",
          8924 => x"08",
          8925 => x"80",
          8926 => x"54",
          8927 => x"80",
          8928 => x"d4",
          8929 => x"2e",
          8930 => x"80",
          8931 => x"54",
          8932 => x"80",
          8933 => x"52",
          8934 => x"ac",
          8935 => x"d4",
          8936 => x"82",
          8937 => x"b1",
          8938 => x"82",
          8939 => x"52",
          8940 => x"9a",
          8941 => x"54",
          8942 => x"15",
          8943 => x"77",
          8944 => x"ff",
          8945 => x"78",
          8946 => x"83",
          8947 => x"51",
          8948 => x"3f",
          8949 => x"08",
          8950 => x"74",
          8951 => x"0c",
          8952 => x"04",
          8953 => x"60",
          8954 => x"05",
          8955 => x"33",
          8956 => x"05",
          8957 => x"40",
          8958 => x"ba",
          8959 => x"f8",
          8960 => x"d4",
          8961 => x"bd",
          8962 => x"33",
          8963 => x"b5",
          8964 => x"2e",
          8965 => x"1a",
          8966 => x"90",
          8967 => x"33",
          8968 => x"70",
          8969 => x"55",
          8970 => x"38",
          8971 => x"97",
          8972 => x"82",
          8973 => x"58",
          8974 => x"7e",
          8975 => x"70",
          8976 => x"55",
          8977 => x"56",
          8978 => x"e3",
          8979 => x"7d",
          8980 => x"70",
          8981 => x"2a",
          8982 => x"08",
          8983 => x"08",
          8984 => x"5d",
          8985 => x"77",
          8986 => x"9c",
          8987 => x"26",
          8988 => x"57",
          8989 => x"59",
          8990 => x"52",
          8991 => x"9d",
          8992 => x"15",
          8993 => x"9c",
          8994 => x"26",
          8995 => x"55",
          8996 => x"08",
          8997 => x"99",
          8998 => x"f8",
          8999 => x"ff",
          9000 => x"d4",
          9001 => x"38",
          9002 => x"75",
          9003 => x"81",
          9004 => x"93",
          9005 => x"80",
          9006 => x"2e",
          9007 => x"ff",
          9008 => x"58",
          9009 => x"7d",
          9010 => x"38",
          9011 => x"55",
          9012 => x"b4",
          9013 => x"56",
          9014 => x"09",
          9015 => x"38",
          9016 => x"53",
          9017 => x"51",
          9018 => x"3f",
          9019 => x"08",
          9020 => x"f8",
          9021 => x"38",
          9022 => x"ff",
          9023 => x"5c",
          9024 => x"84",
          9025 => x"5c",
          9026 => x"12",
          9027 => x"80",
          9028 => x"78",
          9029 => x"7c",
          9030 => x"90",
          9031 => x"c0",
          9032 => x"90",
          9033 => x"15",
          9034 => x"94",
          9035 => x"54",
          9036 => x"91",
          9037 => x"31",
          9038 => x"84",
          9039 => x"07",
          9040 => x"16",
          9041 => x"73",
          9042 => x"0c",
          9043 => x"04",
          9044 => x"6b",
          9045 => x"05",
          9046 => x"33",
          9047 => x"5a",
          9048 => x"95",
          9049 => x"80",
          9050 => x"f8",
          9051 => x"f8",
          9052 => x"f8",
          9053 => x"82",
          9054 => x"70",
          9055 => x"74",
          9056 => x"38",
          9057 => x"82",
          9058 => x"81",
          9059 => x"81",
          9060 => x"ff",
          9061 => x"82",
          9062 => x"81",
          9063 => x"81",
          9064 => x"83",
          9065 => x"c0",
          9066 => x"2a",
          9067 => x"51",
          9068 => x"74",
          9069 => x"99",
          9070 => x"53",
          9071 => x"51",
          9072 => x"3f",
          9073 => x"08",
          9074 => x"55",
          9075 => x"92",
          9076 => x"80",
          9077 => x"38",
          9078 => x"06",
          9079 => x"2e",
          9080 => x"48",
          9081 => x"87",
          9082 => x"79",
          9083 => x"78",
          9084 => x"26",
          9085 => x"19",
          9086 => x"74",
          9087 => x"38",
          9088 => x"e4",
          9089 => x"2a",
          9090 => x"70",
          9091 => x"59",
          9092 => x"7a",
          9093 => x"56",
          9094 => x"80",
          9095 => x"51",
          9096 => x"74",
          9097 => x"99",
          9098 => x"53",
          9099 => x"51",
          9100 => x"3f",
          9101 => x"d4",
          9102 => x"ac",
          9103 => x"2a",
          9104 => x"82",
          9105 => x"43",
          9106 => x"83",
          9107 => x"66",
          9108 => x"60",
          9109 => x"90",
          9110 => x"31",
          9111 => x"80",
          9112 => x"8a",
          9113 => x"56",
          9114 => x"26",
          9115 => x"77",
          9116 => x"81",
          9117 => x"74",
          9118 => x"38",
          9119 => x"55",
          9120 => x"83",
          9121 => x"81",
          9122 => x"80",
          9123 => x"38",
          9124 => x"55",
          9125 => x"5e",
          9126 => x"89",
          9127 => x"5a",
          9128 => x"09",
          9129 => x"e1",
          9130 => x"38",
          9131 => x"57",
          9132 => x"c8",
          9133 => x"5a",
          9134 => x"9d",
          9135 => x"26",
          9136 => x"c8",
          9137 => x"10",
          9138 => x"22",
          9139 => x"74",
          9140 => x"38",
          9141 => x"ee",
          9142 => x"66",
          9143 => x"cf",
          9144 => x"f8",
          9145 => x"84",
          9146 => x"89",
          9147 => x"a0",
          9148 => x"82",
          9149 => x"fc",
          9150 => x"56",
          9151 => x"f0",
          9152 => x"80",
          9153 => x"d3",
          9154 => x"38",
          9155 => x"57",
          9156 => x"c8",
          9157 => x"5a",
          9158 => x"9d",
          9159 => x"26",
          9160 => x"c8",
          9161 => x"10",
          9162 => x"22",
          9163 => x"74",
          9164 => x"38",
          9165 => x"ee",
          9166 => x"66",
          9167 => x"ef",
          9168 => x"f8",
          9169 => x"05",
          9170 => x"f8",
          9171 => x"26",
          9172 => x"0b",
          9173 => x"08",
          9174 => x"f8",
          9175 => x"11",
          9176 => x"05",
          9177 => x"83",
          9178 => x"2a",
          9179 => x"a0",
          9180 => x"7d",
          9181 => x"69",
          9182 => x"05",
          9183 => x"72",
          9184 => x"5c",
          9185 => x"59",
          9186 => x"2e",
          9187 => x"89",
          9188 => x"60",
          9189 => x"84",
          9190 => x"5d",
          9191 => x"18",
          9192 => x"68",
          9193 => x"74",
          9194 => x"af",
          9195 => x"31",
          9196 => x"53",
          9197 => x"52",
          9198 => x"f3",
          9199 => x"f8",
          9200 => x"83",
          9201 => x"06",
          9202 => x"d4",
          9203 => x"ff",
          9204 => x"dd",
          9205 => x"83",
          9206 => x"2a",
          9207 => x"be",
          9208 => x"39",
          9209 => x"09",
          9210 => x"c5",
          9211 => x"f5",
          9212 => x"f8",
          9213 => x"38",
          9214 => x"79",
          9215 => x"80",
          9216 => x"38",
          9217 => x"96",
          9218 => x"06",
          9219 => x"2e",
          9220 => x"5e",
          9221 => x"82",
          9222 => x"9f",
          9223 => x"38",
          9224 => x"38",
          9225 => x"81",
          9226 => x"fc",
          9227 => x"ab",
          9228 => x"7d",
          9229 => x"81",
          9230 => x"7d",
          9231 => x"78",
          9232 => x"74",
          9233 => x"8e",
          9234 => x"9c",
          9235 => x"53",
          9236 => x"51",
          9237 => x"3f",
          9238 => x"c6",
          9239 => x"51",
          9240 => x"3f",
          9241 => x"8b",
          9242 => x"8f",
          9243 => x"8d",
          9244 => x"83",
          9245 => x"52",
          9246 => x"ff",
          9247 => x"81",
          9248 => x"34",
          9249 => x"70",
          9250 => x"2a",
          9251 => x"54",
          9252 => x"1b",
          9253 => x"b6",
          9254 => x"74",
          9255 => x"26",
          9256 => x"83",
          9257 => x"52",
          9258 => x"ff",
          9259 => x"8a",
          9260 => x"a0",
          9261 => x"8f",
          9262 => x"0b",
          9263 => x"bf",
          9264 => x"51",
          9265 => x"3f",
          9266 => x"9a",
          9267 => x"8e",
          9268 => x"52",
          9269 => x"ff",
          9270 => x"7d",
          9271 => x"81",
          9272 => x"38",
          9273 => x"0a",
          9274 => x"1b",
          9275 => x"fc",
          9276 => x"a4",
          9277 => x"8e",
          9278 => x"52",
          9279 => x"ff",
          9280 => x"81",
          9281 => x"51",
          9282 => x"3f",
          9283 => x"1b",
          9284 => x"ba",
          9285 => x"0b",
          9286 => x"34",
          9287 => x"c2",
          9288 => x"53",
          9289 => x"52",
          9290 => x"51",
          9291 => x"88",
          9292 => x"a7",
          9293 => x"8e",
          9294 => x"83",
          9295 => x"52",
          9296 => x"ff",
          9297 => x"ff",
          9298 => x"1c",
          9299 => x"a6",
          9300 => x"53",
          9301 => x"52",
          9302 => x"ff",
          9303 => x"82",
          9304 => x"83",
          9305 => x"52",
          9306 => x"e2",
          9307 => x"60",
          9308 => x"7e",
          9309 => x"85",
          9310 => x"82",
          9311 => x"83",
          9312 => x"83",
          9313 => x"06",
          9314 => x"75",
          9315 => x"05",
          9316 => x"7e",
          9317 => x"e5",
          9318 => x"53",
          9319 => x"51",
          9320 => x"3f",
          9321 => x"a4",
          9322 => x"51",
          9323 => x"3f",
          9324 => x"e4",
          9325 => x"e4",
          9326 => x"8d",
          9327 => x"18",
          9328 => x"1b",
          9329 => x"a4",
          9330 => x"83",
          9331 => x"ff",
          9332 => x"82",
          9333 => x"78",
          9334 => x"f2",
          9335 => x"60",
          9336 => x"7a",
          9337 => x"ff",
          9338 => x"75",
          9339 => x"53",
          9340 => x"51",
          9341 => x"3f",
          9342 => x"52",
          9343 => x"8d",
          9344 => x"56",
          9345 => x"83",
          9346 => x"06",
          9347 => x"52",
          9348 => x"8c",
          9349 => x"52",
          9350 => x"ff",
          9351 => x"f0",
          9352 => x"1b",
          9353 => x"87",
          9354 => x"55",
          9355 => x"83",
          9356 => x"74",
          9357 => x"ff",
          9358 => x"7c",
          9359 => x"74",
          9360 => x"38",
          9361 => x"54",
          9362 => x"52",
          9363 => x"88",
          9364 => x"d4",
          9365 => x"87",
          9366 => x"53",
          9367 => x"08",
          9368 => x"ff",
          9369 => x"76",
          9370 => x"31",
          9371 => x"cd",
          9372 => x"58",
          9373 => x"ff",
          9374 => x"55",
          9375 => x"83",
          9376 => x"61",
          9377 => x"26",
          9378 => x"57",
          9379 => x"53",
          9380 => x"51",
          9381 => x"3f",
          9382 => x"08",
          9383 => x"76",
          9384 => x"31",
          9385 => x"db",
          9386 => x"7d",
          9387 => x"38",
          9388 => x"83",
          9389 => x"8a",
          9390 => x"7d",
          9391 => x"38",
          9392 => x"81",
          9393 => x"80",
          9394 => x"80",
          9395 => x"7a",
          9396 => x"ea",
          9397 => x"d5",
          9398 => x"ff",
          9399 => x"83",
          9400 => x"77",
          9401 => x"0b",
          9402 => x"81",
          9403 => x"34",
          9404 => x"34",
          9405 => x"34",
          9406 => x"56",
          9407 => x"52",
          9408 => x"a2",
          9409 => x"0b",
          9410 => x"82",
          9411 => x"82",
          9412 => x"56",
          9413 => x"34",
          9414 => x"08",
          9415 => x"60",
          9416 => x"1b",
          9417 => x"c4",
          9418 => x"83",
          9419 => x"ff",
          9420 => x"81",
          9421 => x"7a",
          9422 => x"ff",
          9423 => x"81",
          9424 => x"f8",
          9425 => x"80",
          9426 => x"7e",
          9427 => x"91",
          9428 => x"82",
          9429 => x"90",
          9430 => x"8e",
          9431 => x"81",
          9432 => x"82",
          9433 => x"56",
          9434 => x"f8",
          9435 => x"0d",
          9436 => x"0d",
          9437 => x"59",
          9438 => x"ff",
          9439 => x"57",
          9440 => x"b4",
          9441 => x"f8",
          9442 => x"81",
          9443 => x"52",
          9444 => x"bd",
          9445 => x"2e",
          9446 => x"9c",
          9447 => x"33",
          9448 => x"2e",
          9449 => x"76",
          9450 => x"58",
          9451 => x"57",
          9452 => x"09",
          9453 => x"38",
          9454 => x"78",
          9455 => x"38",
          9456 => x"82",
          9457 => x"8d",
          9458 => x"f7",
          9459 => x"02",
          9460 => x"05",
          9461 => x"77",
          9462 => x"81",
          9463 => x"8d",
          9464 => x"e7",
          9465 => x"08",
          9466 => x"24",
          9467 => x"17",
          9468 => x"8c",
          9469 => x"77",
          9470 => x"16",
          9471 => x"25",
          9472 => x"3d",
          9473 => x"75",
          9474 => x"52",
          9475 => x"cb",
          9476 => x"76",
          9477 => x"70",
          9478 => x"2a",
          9479 => x"51",
          9480 => x"84",
          9481 => x"19",
          9482 => x"8b",
          9483 => x"f9",
          9484 => x"84",
          9485 => x"56",
          9486 => x"a7",
          9487 => x"fc",
          9488 => x"53",
          9489 => x"75",
          9490 => x"85",
          9491 => x"f8",
          9492 => x"84",
          9493 => x"2e",
          9494 => x"87",
          9495 => x"08",
          9496 => x"ff",
          9497 => x"d4",
          9498 => x"3d",
          9499 => x"3d",
          9500 => x"80",
          9501 => x"52",
          9502 => x"88",
          9503 => x"74",
          9504 => x"0d",
          9505 => x"0d",
          9506 => x"05",
          9507 => x"86",
          9508 => x"54",
          9509 => x"73",
          9510 => x"fe",
          9511 => x"51",
          9512 => x"98",
          9513 => x"fd",
          9514 => x"02",
          9515 => x"05",
          9516 => x"80",
          9517 => x"ff",
          9518 => x"72",
          9519 => x"06",
          9520 => x"39",
          9521 => x"73",
          9522 => x"83",
          9523 => x"81",
          9524 => x"70",
          9525 => x"38",
          9526 => x"22",
          9527 => x"2e",
          9528 => x"12",
          9529 => x"ff",
          9530 => x"71",
          9531 => x"8d",
          9532 => x"82",
          9533 => x"70",
          9534 => x"e1",
          9535 => x"12",
          9536 => x"06",
          9537 => x"82",
          9538 => x"85",
          9539 => x"fe",
          9540 => x"92",
          9541 => x"84",
          9542 => x"22",
          9543 => x"53",
          9544 => x"26",
          9545 => x"53",
          9546 => x"83",
          9547 => x"81",
          9548 => x"70",
          9549 => x"8b",
          9550 => x"82",
          9551 => x"70",
          9552 => x"72",
          9553 => x"0c",
          9554 => x"04",
          9555 => x"77",
          9556 => x"ff",
          9557 => x"a7",
          9558 => x"ff",
          9559 => x"ca",
          9560 => x"9f",
          9561 => x"85",
          9562 => x"b8",
          9563 => x"82",
          9564 => x"70",
          9565 => x"25",
          9566 => x"07",
          9567 => x"70",
          9568 => x"75",
          9569 => x"57",
          9570 => x"2a",
          9571 => x"06",
          9572 => x"52",
          9573 => x"71",
          9574 => x"38",
          9575 => x"80",
          9576 => x"84",
          9577 => x"d4",
          9578 => x"08",
          9579 => x"31",
          9580 => x"70",
          9581 => x"51",
          9582 => x"71",
          9583 => x"06",
          9584 => x"51",
          9585 => x"f0",
          9586 => x"39",
          9587 => x"9a",
          9588 => x"51",
          9589 => x"12",
          9590 => x"88",
          9591 => x"39",
          9592 => x"51",
          9593 => x"a0",
          9594 => x"83",
          9595 => x"52",
          9596 => x"fe",
          9597 => x"10",
          9598 => x"f1",
          9599 => x"70",
          9600 => x"0c",
          9601 => x"04",
          9602 => x"ff",
          9603 => x"ff",
          9604 => x"00",
          9605 => x"ff",
          9606 => x"2c",
          9607 => x"2b",
          9608 => x"2b",
          9609 => x"2b",
          9610 => x"2b",
          9611 => x"2b",
          9612 => x"2b",
          9613 => x"2b",
          9614 => x"2c",
          9615 => x"2c",
          9616 => x"2c",
          9617 => x"2c",
          9618 => x"2c",
          9619 => x"2c",
          9620 => x"2c",
          9621 => x"2c",
          9622 => x"2c",
          9623 => x"2c",
          9624 => x"2c",
          9625 => x"2c",
          9626 => x"42",
          9627 => x"42",
          9628 => x"42",
          9629 => x"42",
          9630 => x"42",
          9631 => x"48",
          9632 => x"49",
          9633 => x"4a",
          9634 => x"4c",
          9635 => x"49",
          9636 => x"47",
          9637 => x"4b",
          9638 => x"4c",
          9639 => x"4b",
          9640 => x"4c",
          9641 => x"4b",
          9642 => x"4a",
          9643 => x"47",
          9644 => x"4a",
          9645 => x"4a",
          9646 => x"4b",
          9647 => x"47",
          9648 => x"47",
          9649 => x"4b",
          9650 => x"4c",
          9651 => x"4c",
          9652 => x"4c",
          9653 => x"95",
          9654 => x"95",
          9655 => x"95",
          9656 => x"95",
          9657 => x"95",
          9658 => x"95",
          9659 => x"95",
          9660 => x"95",
          9661 => x"95",
          9662 => x"0e",
          9663 => x"17",
          9664 => x"17",
          9665 => x"0e",
          9666 => x"17",
          9667 => x"17",
          9668 => x"17",
          9669 => x"17",
          9670 => x"17",
          9671 => x"17",
          9672 => x"17",
          9673 => x"0e",
          9674 => x"17",
          9675 => x"0e",
          9676 => x"0e",
          9677 => x"17",
          9678 => x"17",
          9679 => x"17",
          9680 => x"17",
          9681 => x"17",
          9682 => x"17",
          9683 => x"17",
          9684 => x"17",
          9685 => x"17",
          9686 => x"17",
          9687 => x"17",
          9688 => x"17",
          9689 => x"17",
          9690 => x"17",
          9691 => x"17",
          9692 => x"17",
          9693 => x"17",
          9694 => x"17",
          9695 => x"17",
          9696 => x"17",
          9697 => x"17",
          9698 => x"17",
          9699 => x"17",
          9700 => x"17",
          9701 => x"17",
          9702 => x"17",
          9703 => x"17",
          9704 => x"17",
          9705 => x"17",
          9706 => x"17",
          9707 => x"17",
          9708 => x"17",
          9709 => x"17",
          9710 => x"17",
          9711 => x"17",
          9712 => x"17",
          9713 => x"0f",
          9714 => x"17",
          9715 => x"17",
          9716 => x"17",
          9717 => x"17",
          9718 => x"11",
          9719 => x"17",
          9720 => x"17",
          9721 => x"17",
          9722 => x"17",
          9723 => x"17",
          9724 => x"17",
          9725 => x"17",
          9726 => x"17",
          9727 => x"17",
          9728 => x"17",
          9729 => x"0e",
          9730 => x"10",
          9731 => x"0e",
          9732 => x"0e",
          9733 => x"0e",
          9734 => x"17",
          9735 => x"10",
          9736 => x"17",
          9737 => x"17",
          9738 => x"0e",
          9739 => x"17",
          9740 => x"17",
          9741 => x"10",
          9742 => x"10",
          9743 => x"17",
          9744 => x"17",
          9745 => x"0f",
          9746 => x"17",
          9747 => x"11",
          9748 => x"17",
          9749 => x"17",
          9750 => x"11",
          9751 => x"6e",
          9752 => x"00",
          9753 => x"6f",
          9754 => x"00",
          9755 => x"6e",
          9756 => x"00",
          9757 => x"6f",
          9758 => x"00",
          9759 => x"78",
          9760 => x"00",
          9761 => x"6c",
          9762 => x"00",
          9763 => x"6f",
          9764 => x"00",
          9765 => x"69",
          9766 => x"00",
          9767 => x"75",
          9768 => x"00",
          9769 => x"62",
          9770 => x"68",
          9771 => x"77",
          9772 => x"64",
          9773 => x"65",
          9774 => x"64",
          9775 => x"65",
          9776 => x"6c",
          9777 => x"00",
          9778 => x"70",
          9779 => x"73",
          9780 => x"74",
          9781 => x"73",
          9782 => x"00",
          9783 => x"66",
          9784 => x"00",
          9785 => x"73",
          9786 => x"00",
          9787 => x"61",
          9788 => x"00",
          9789 => x"61",
          9790 => x"00",
          9791 => x"6c",
          9792 => x"00",
          9793 => x"00",
          9794 => x"73",
          9795 => x"72",
          9796 => x"00",
          9797 => x"74",
          9798 => x"61",
          9799 => x"72",
          9800 => x"2e",
          9801 => x"73",
          9802 => x"6f",
          9803 => x"65",
          9804 => x"2e",
          9805 => x"20",
          9806 => x"65",
          9807 => x"75",
          9808 => x"00",
          9809 => x"20",
          9810 => x"68",
          9811 => x"75",
          9812 => x"00",
          9813 => x"76",
          9814 => x"64",
          9815 => x"6c",
          9816 => x"6d",
          9817 => x"00",
          9818 => x"63",
          9819 => x"20",
          9820 => x"69",
          9821 => x"00",
          9822 => x"6c",
          9823 => x"6c",
          9824 => x"64",
          9825 => x"78",
          9826 => x"73",
          9827 => x"00",
          9828 => x"6c",
          9829 => x"61",
          9830 => x"65",
          9831 => x"76",
          9832 => x"64",
          9833 => x"00",
          9834 => x"20",
          9835 => x"77",
          9836 => x"65",
          9837 => x"6f",
          9838 => x"74",
          9839 => x"00",
          9840 => x"69",
          9841 => x"6e",
          9842 => x"65",
          9843 => x"73",
          9844 => x"76",
          9845 => x"64",
          9846 => x"00",
          9847 => x"73",
          9848 => x"6f",
          9849 => x"6e",
          9850 => x"65",
          9851 => x"00",
          9852 => x"20",
          9853 => x"70",
          9854 => x"62",
          9855 => x"66",
          9856 => x"73",
          9857 => x"65",
          9858 => x"6f",
          9859 => x"20",
          9860 => x"64",
          9861 => x"2e",
          9862 => x"72",
          9863 => x"20",
          9864 => x"72",
          9865 => x"2e",
          9866 => x"6d",
          9867 => x"74",
          9868 => x"70",
          9869 => x"74",
          9870 => x"20",
          9871 => x"63",
          9872 => x"65",
          9873 => x"00",
          9874 => x"6c",
          9875 => x"73",
          9876 => x"63",
          9877 => x"2e",
          9878 => x"73",
          9879 => x"69",
          9880 => x"6e",
          9881 => x"65",
          9882 => x"79",
          9883 => x"00",
          9884 => x"6f",
          9885 => x"6e",
          9886 => x"70",
          9887 => x"66",
          9888 => x"73",
          9889 => x"00",
          9890 => x"72",
          9891 => x"74",
          9892 => x"20",
          9893 => x"6f",
          9894 => x"63",
          9895 => x"00",
          9896 => x"63",
          9897 => x"73",
          9898 => x"00",
          9899 => x"6b",
          9900 => x"6e",
          9901 => x"72",
          9902 => x"00",
          9903 => x"6c",
          9904 => x"79",
          9905 => x"20",
          9906 => x"61",
          9907 => x"6c",
          9908 => x"79",
          9909 => x"2f",
          9910 => x"2e",
          9911 => x"00",
          9912 => x"61",
          9913 => x"00",
          9914 => x"25",
          9915 => x"78",
          9916 => x"3d",
          9917 => x"6c",
          9918 => x"32",
          9919 => x"38",
          9920 => x"20",
          9921 => x"42",
          9922 => x"38",
          9923 => x"25",
          9924 => x"78",
          9925 => x"38",
          9926 => x"00",
          9927 => x"38",
          9928 => x"00",
          9929 => x"20",
          9930 => x"34",
          9931 => x"00",
          9932 => x"20",
          9933 => x"20",
          9934 => x"00",
          9935 => x"32",
          9936 => x"00",
          9937 => x"00",
          9938 => x"00",
          9939 => x"00",
          9940 => x"53",
          9941 => x"2a",
          9942 => x"20",
          9943 => x"00",
          9944 => x"2f",
          9945 => x"32",
          9946 => x"00",
          9947 => x"2e",
          9948 => x"00",
          9949 => x"50",
          9950 => x"72",
          9951 => x"25",
          9952 => x"29",
          9953 => x"20",
          9954 => x"2a",
          9955 => x"00",
          9956 => x"55",
          9957 => x"74",
          9958 => x"75",
          9959 => x"48",
          9960 => x"6c",
          9961 => x"00",
          9962 => x"6d",
          9963 => x"69",
          9964 => x"72",
          9965 => x"74",
          9966 => x"32",
          9967 => x"74",
          9968 => x"75",
          9969 => x"00",
          9970 => x"43",
          9971 => x"52",
          9972 => x"6e",
          9973 => x"72",
          9974 => x"00",
          9975 => x"43",
          9976 => x"57",
          9977 => x"6e",
          9978 => x"72",
          9979 => x"00",
          9980 => x"52",
          9981 => x"52",
          9982 => x"6e",
          9983 => x"72",
          9984 => x"00",
          9985 => x"52",
          9986 => x"54",
          9987 => x"6e",
          9988 => x"72",
          9989 => x"00",
          9990 => x"52",
          9991 => x"52",
          9992 => x"6e",
          9993 => x"72",
          9994 => x"00",
          9995 => x"52",
          9996 => x"54",
          9997 => x"6e",
          9998 => x"72",
          9999 => x"00",
         10000 => x"74",
         10001 => x"67",
         10002 => x"20",
         10003 => x"65",
         10004 => x"2e",
         10005 => x"61",
         10006 => x"6e",
         10007 => x"69",
         10008 => x"2e",
         10009 => x"00",
         10010 => x"74",
         10011 => x"65",
         10012 => x"61",
         10013 => x"00",
         10014 => x"53",
         10015 => x"74",
         10016 => x"00",
         10017 => x"69",
         10018 => x"20",
         10019 => x"69",
         10020 => x"69",
         10021 => x"73",
         10022 => x"64",
         10023 => x"72",
         10024 => x"2c",
         10025 => x"65",
         10026 => x"20",
         10027 => x"74",
         10028 => x"6e",
         10029 => x"6c",
         10030 => x"00",
         10031 => x"00",
         10032 => x"65",
         10033 => x"6e",
         10034 => x"2e",
         10035 => x"00",
         10036 => x"70",
         10037 => x"67",
         10038 => x"00",
         10039 => x"6d",
         10040 => x"69",
         10041 => x"2e",
         10042 => x"00",
         10043 => x"38",
         10044 => x"25",
         10045 => x"29",
         10046 => x"30",
         10047 => x"28",
         10048 => x"78",
         10049 => x"00",
         10050 => x"6d",
         10051 => x"65",
         10052 => x"79",
         10053 => x"6f",
         10054 => x"65",
         10055 => x"00",
         10056 => x"38",
         10057 => x"25",
         10058 => x"2d",
         10059 => x"3f",
         10060 => x"38",
         10061 => x"25",
         10062 => x"2d",
         10063 => x"38",
         10064 => x"25",
         10065 => x"58",
         10066 => x"00",
         10067 => x"65",
         10068 => x"69",
         10069 => x"63",
         10070 => x"20",
         10071 => x"30",
         10072 => x"20",
         10073 => x"0a",
         10074 => x"6c",
         10075 => x"67",
         10076 => x"64",
         10077 => x"20",
         10078 => x"6c",
         10079 => x"2e",
         10080 => x"00",
         10081 => x"6c",
         10082 => x"65",
         10083 => x"6e",
         10084 => x"63",
         10085 => x"20",
         10086 => x"29",
         10087 => x"00",
         10088 => x"73",
         10089 => x"74",
         10090 => x"20",
         10091 => x"6c",
         10092 => x"74",
         10093 => x"2e",
         10094 => x"00",
         10095 => x"6c",
         10096 => x"65",
         10097 => x"74",
         10098 => x"2e",
         10099 => x"00",
         10100 => x"55",
         10101 => x"6e",
         10102 => x"3a",
         10103 => x"5c",
         10104 => x"25",
         10105 => x"00",
         10106 => x"3a",
         10107 => x"5c",
         10108 => x"00",
         10109 => x"3a",
         10110 => x"00",
         10111 => x"64",
         10112 => x"6d",
         10113 => x"64",
         10114 => x"00",
         10115 => x"6d",
         10116 => x"20",
         10117 => x"61",
         10118 => x"65",
         10119 => x"63",
         10120 => x"6f",
         10121 => x"72",
         10122 => x"73",
         10123 => x"6f",
         10124 => x"6e",
         10125 => x"00",
         10126 => x"6e",
         10127 => x"67",
         10128 => x"00",
         10129 => x"61",
         10130 => x"6e",
         10131 => x"6e",
         10132 => x"72",
         10133 => x"73",
         10134 => x"00",
         10135 => x"2f",
         10136 => x"25",
         10137 => x"64",
         10138 => x"3a",
         10139 => x"25",
         10140 => x"0a",
         10141 => x"43",
         10142 => x"6e",
         10143 => x"75",
         10144 => x"69",
         10145 => x"00",
         10146 => x"66",
         10147 => x"20",
         10148 => x"20",
         10149 => x"66",
         10150 => x"00",
         10151 => x"44",
         10152 => x"63",
         10153 => x"69",
         10154 => x"65",
         10155 => x"74",
         10156 => x"00",
         10157 => x"20",
         10158 => x"20",
         10159 => x"41",
         10160 => x"28",
         10161 => x"58",
         10162 => x"38",
         10163 => x"0a",
         10164 => x"20",
         10165 => x"52",
         10166 => x"20",
         10167 => x"28",
         10168 => x"58",
         10169 => x"38",
         10170 => x"0a",
         10171 => x"20",
         10172 => x"53",
         10173 => x"52",
         10174 => x"28",
         10175 => x"58",
         10176 => x"38",
         10177 => x"0a",
         10178 => x"20",
         10179 => x"41",
         10180 => x"20",
         10181 => x"28",
         10182 => x"58",
         10183 => x"38",
         10184 => x"0a",
         10185 => x"20",
         10186 => x"4d",
         10187 => x"20",
         10188 => x"28",
         10189 => x"58",
         10190 => x"38",
         10191 => x"0a",
         10192 => x"20",
         10193 => x"20",
         10194 => x"44",
         10195 => x"28",
         10196 => x"69",
         10197 => x"20",
         10198 => x"32",
         10199 => x"0a",
         10200 => x"20",
         10201 => x"4d",
         10202 => x"20",
         10203 => x"28",
         10204 => x"65",
         10205 => x"20",
         10206 => x"32",
         10207 => x"0a",
         10208 => x"20",
         10209 => x"54",
         10210 => x"54",
         10211 => x"28",
         10212 => x"6e",
         10213 => x"73",
         10214 => x"32",
         10215 => x"0a",
         10216 => x"20",
         10217 => x"53",
         10218 => x"4e",
         10219 => x"55",
         10220 => x"00",
         10221 => x"20",
         10222 => x"20",
         10223 => x"00",
         10224 => x"20",
         10225 => x"43",
         10226 => x"00",
         10227 => x"20",
         10228 => x"32",
         10229 => x"20",
         10230 => x"49",
         10231 => x"64",
         10232 => x"73",
         10233 => x"00",
         10234 => x"20",
         10235 => x"55",
         10236 => x"73",
         10237 => x"56",
         10238 => x"6f",
         10239 => x"64",
         10240 => x"73",
         10241 => x"20",
         10242 => x"58",
         10243 => x"00",
         10244 => x"20",
         10245 => x"55",
         10246 => x"6d",
         10247 => x"20",
         10248 => x"72",
         10249 => x"64",
         10250 => x"73",
         10251 => x"20",
         10252 => x"58",
         10253 => x"00",
         10254 => x"20",
         10255 => x"61",
         10256 => x"53",
         10257 => x"74",
         10258 => x"64",
         10259 => x"73",
         10260 => x"20",
         10261 => x"20",
         10262 => x"58",
         10263 => x"00",
         10264 => x"73",
         10265 => x"00",
         10266 => x"20",
         10267 => x"55",
         10268 => x"20",
         10269 => x"20",
         10270 => x"20",
         10271 => x"20",
         10272 => x"20",
         10273 => x"20",
         10274 => x"58",
         10275 => x"00",
         10276 => x"20",
         10277 => x"73",
         10278 => x"20",
         10279 => x"63",
         10280 => x"72",
         10281 => x"20",
         10282 => x"20",
         10283 => x"20",
         10284 => x"25",
         10285 => x"4d",
         10286 => x"00",
         10287 => x"20",
         10288 => x"52",
         10289 => x"43",
         10290 => x"6b",
         10291 => x"65",
         10292 => x"20",
         10293 => x"20",
         10294 => x"20",
         10295 => x"25",
         10296 => x"4d",
         10297 => x"00",
         10298 => x"20",
         10299 => x"73",
         10300 => x"6e",
         10301 => x"44",
         10302 => x"20",
         10303 => x"63",
         10304 => x"72",
         10305 => x"20",
         10306 => x"25",
         10307 => x"4d",
         10308 => x"00",
         10309 => x"61",
         10310 => x"00",
         10311 => x"64",
         10312 => x"00",
         10313 => x"65",
         10314 => x"00",
         10315 => x"4f",
         10316 => x"4f",
         10317 => x"00",
         10318 => x"6b",
         10319 => x"6e",
         10320 => x"a2",
         10321 => x"00",
         10322 => x"00",
         10323 => x"a2",
         10324 => x"00",
         10325 => x"00",
         10326 => x"a2",
         10327 => x"00",
         10328 => x"00",
         10329 => x"a2",
         10330 => x"00",
         10331 => x"00",
         10332 => x"a2",
         10333 => x"00",
         10334 => x"00",
         10335 => x"a2",
         10336 => x"00",
         10337 => x"00",
         10338 => x"a2",
         10339 => x"00",
         10340 => x"00",
         10341 => x"a2",
         10342 => x"00",
         10343 => x"00",
         10344 => x"a2",
         10345 => x"00",
         10346 => x"00",
         10347 => x"a2",
         10348 => x"00",
         10349 => x"00",
         10350 => x"a2",
         10351 => x"00",
         10352 => x"00",
         10353 => x"a2",
         10354 => x"00",
         10355 => x"00",
         10356 => x"a2",
         10357 => x"00",
         10358 => x"00",
         10359 => x"a2",
         10360 => x"00",
         10361 => x"00",
         10362 => x"a2",
         10363 => x"00",
         10364 => x"00",
         10365 => x"a2",
         10366 => x"00",
         10367 => x"00",
         10368 => x"a2",
         10369 => x"00",
         10370 => x"00",
         10371 => x"a2",
         10372 => x"00",
         10373 => x"00",
         10374 => x"a2",
         10375 => x"00",
         10376 => x"00",
         10377 => x"a2",
         10378 => x"00",
         10379 => x"00",
         10380 => x"a2",
         10381 => x"00",
         10382 => x"00",
         10383 => x"a2",
         10384 => x"00",
         10385 => x"00",
         10386 => x"44",
         10387 => x"43",
         10388 => x"42",
         10389 => x"41",
         10390 => x"36",
         10391 => x"35",
         10392 => x"34",
         10393 => x"46",
         10394 => x"33",
         10395 => x"32",
         10396 => x"31",
         10397 => x"00",
         10398 => x"00",
         10399 => x"00",
         10400 => x"00",
         10401 => x"00",
         10402 => x"00",
         10403 => x"00",
         10404 => x"00",
         10405 => x"00",
         10406 => x"00",
         10407 => x"00",
         10408 => x"73",
         10409 => x"79",
         10410 => x"73",
         10411 => x"00",
         10412 => x"00",
         10413 => x"34",
         10414 => x"20",
         10415 => x"00",
         10416 => x"69",
         10417 => x"20",
         10418 => x"72",
         10419 => x"74",
         10420 => x"65",
         10421 => x"73",
         10422 => x"79",
         10423 => x"6c",
         10424 => x"6f",
         10425 => x"46",
         10426 => x"00",
         10427 => x"6e",
         10428 => x"20",
         10429 => x"6e",
         10430 => x"65",
         10431 => x"20",
         10432 => x"74",
         10433 => x"20",
         10434 => x"65",
         10435 => x"69",
         10436 => x"6c",
         10437 => x"2e",
         10438 => x"00",
         10439 => x"3a",
         10440 => x"7c",
         10441 => x"00",
         10442 => x"3b",
         10443 => x"00",
         10444 => x"54",
         10445 => x"54",
         10446 => x"00",
         10447 => x"90",
         10448 => x"4f",
         10449 => x"30",
         10450 => x"20",
         10451 => x"45",
         10452 => x"20",
         10453 => x"33",
         10454 => x"20",
         10455 => x"20",
         10456 => x"45",
         10457 => x"20",
         10458 => x"20",
         10459 => x"20",
         10460 => x"a3",
         10461 => x"00",
         10462 => x"00",
         10463 => x"00",
         10464 => x"05",
         10465 => x"10",
         10466 => x"18",
         10467 => x"00",
         10468 => x"45",
         10469 => x"8f",
         10470 => x"45",
         10471 => x"8e",
         10472 => x"92",
         10473 => x"55",
         10474 => x"9a",
         10475 => x"9e",
         10476 => x"4f",
         10477 => x"a6",
         10478 => x"aa",
         10479 => x"ae",
         10480 => x"b2",
         10481 => x"b6",
         10482 => x"ba",
         10483 => x"be",
         10484 => x"c2",
         10485 => x"c6",
         10486 => x"ca",
         10487 => x"ce",
         10488 => x"d2",
         10489 => x"d6",
         10490 => x"da",
         10491 => x"de",
         10492 => x"e2",
         10493 => x"e6",
         10494 => x"ea",
         10495 => x"ee",
         10496 => x"f2",
         10497 => x"f6",
         10498 => x"fa",
         10499 => x"fe",
         10500 => x"2c",
         10501 => x"5d",
         10502 => x"2a",
         10503 => x"3f",
         10504 => x"00",
         10505 => x"00",
         10506 => x"00",
         10507 => x"02",
         10508 => x"00",
         10509 => x"00",
         10510 => x"00",
         10511 => x"00",
         10512 => x"00",
         10513 => x"00",
         10514 => x"00",
         10515 => x"00",
         10516 => x"00",
         10517 => x"00",
         10518 => x"00",
         10519 => x"00",
         10520 => x"00",
         10521 => x"00",
         10522 => x"00",
         10523 => x"00",
         10524 => x"00",
         10525 => x"00",
         10526 => x"00",
         10527 => x"00",
         10528 => x"01",
         10529 => x"00",
         10530 => x"00",
         10531 => x"00",
         10532 => x"00",
         10533 => x"23",
         10534 => x"00",
         10535 => x"00",
         10536 => x"00",
         10537 => x"25",
         10538 => x"25",
         10539 => x"25",
         10540 => x"25",
         10541 => x"25",
         10542 => x"25",
         10543 => x"25",
         10544 => x"25",
         10545 => x"25",
         10546 => x"25",
         10547 => x"25",
         10548 => x"25",
         10549 => x"25",
         10550 => x"25",
         10551 => x"25",
         10552 => x"25",
         10553 => x"25",
         10554 => x"25",
         10555 => x"25",
         10556 => x"25",
         10557 => x"25",
         10558 => x"25",
         10559 => x"25",
         10560 => x"25",
         10561 => x"00",
         10562 => x"03",
         10563 => x"03",
         10564 => x"03",
         10565 => x"03",
         10566 => x"03",
         10567 => x"03",
         10568 => x"22",
         10569 => x"00",
         10570 => x"22",
         10571 => x"23",
         10572 => x"22",
         10573 => x"22",
         10574 => x"22",
         10575 => x"00",
         10576 => x"00",
         10577 => x"03",
         10578 => x"03",
         10579 => x"03",
         10580 => x"00",
         10581 => x"01",
         10582 => x"01",
         10583 => x"01",
         10584 => x"01",
         10585 => x"01",
         10586 => x"01",
         10587 => x"02",
         10588 => x"01",
         10589 => x"01",
         10590 => x"01",
         10591 => x"01",
         10592 => x"01",
         10593 => x"01",
         10594 => x"01",
         10595 => x"01",
         10596 => x"01",
         10597 => x"01",
         10598 => x"01",
         10599 => x"01",
         10600 => x"02",
         10601 => x"01",
         10602 => x"02",
         10603 => x"01",
         10604 => x"01",
         10605 => x"01",
         10606 => x"01",
         10607 => x"01",
         10608 => x"01",
         10609 => x"01",
         10610 => x"01",
         10611 => x"01",
         10612 => x"01",
         10613 => x"01",
         10614 => x"01",
         10615 => x"01",
         10616 => x"01",
         10617 => x"01",
         10618 => x"01",
         10619 => x"01",
         10620 => x"01",
         10621 => x"01",
         10622 => x"01",
         10623 => x"01",
         10624 => x"01",
         10625 => x"01",
         10626 => x"01",
         10627 => x"00",
         10628 => x"01",
         10629 => x"01",
         10630 => x"01",
         10631 => x"01",
         10632 => x"01",
         10633 => x"01",
         10634 => x"00",
         10635 => x"02",
         10636 => x"02",
         10637 => x"02",
         10638 => x"02",
         10639 => x"02",
         10640 => x"02",
         10641 => x"01",
         10642 => x"02",
         10643 => x"01",
         10644 => x"01",
         10645 => x"01",
         10646 => x"02",
         10647 => x"02",
         10648 => x"02",
         10649 => x"01",
         10650 => x"02",
         10651 => x"02",
         10652 => x"01",
         10653 => x"2c",
         10654 => x"02",
         10655 => x"01",
         10656 => x"02",
         10657 => x"02",
         10658 => x"01",
         10659 => x"02",
         10660 => x"02",
         10661 => x"02",
         10662 => x"2c",
         10663 => x"02",
         10664 => x"02",
         10665 => x"01",
         10666 => x"02",
         10667 => x"02",
         10668 => x"02",
         10669 => x"01",
         10670 => x"02",
         10671 => x"02",
         10672 => x"02",
         10673 => x"03",
         10674 => x"03",
         10675 => x"03",
         10676 => x"00",
         10677 => x"03",
         10678 => x"03",
         10679 => x"03",
         10680 => x"00",
         10681 => x"03",
         10682 => x"03",
         10683 => x"00",
         10684 => x"03",
         10685 => x"03",
         10686 => x"03",
         10687 => x"03",
         10688 => x"03",
         10689 => x"03",
         10690 => x"03",
         10691 => x"03",
         10692 => x"04",
         10693 => x"04",
         10694 => x"04",
         10695 => x"04",
         10696 => x"04",
         10697 => x"04",
         10698 => x"04",
         10699 => x"01",
         10700 => x"04",
         10701 => x"00",
         10702 => x"00",
         10703 => x"1e",
         10704 => x"1e",
         10705 => x"1f",
         10706 => x"1f",
         10707 => x"1f",
         10708 => x"1f",
         10709 => x"1f",
         10710 => x"1f",
         10711 => x"1f",
         10712 => x"1f",
         10713 => x"1f",
         10714 => x"1f",
         10715 => x"06",
         10716 => x"00",
         10717 => x"1f",
         10718 => x"1f",
         10719 => x"1f",
         10720 => x"1f",
         10721 => x"1f",
         10722 => x"1f",
         10723 => x"1f",
         10724 => x"06",
         10725 => x"06",
         10726 => x"06",
         10727 => x"00",
         10728 => x"1f",
         10729 => x"1f",
         10730 => x"00",
         10731 => x"1f",
         10732 => x"1f",
         10733 => x"1f",
         10734 => x"1f",
         10735 => x"00",
         10736 => x"21",
         10737 => x"21",
         10738 => x"02",
         10739 => x"00",
         10740 => x"24",
         10741 => x"2c",
         10742 => x"2c",
         10743 => x"2c",
         10744 => x"2c",
         10745 => x"2c",
         10746 => x"2d",
         10747 => x"ff",
         10748 => x"00",
         10749 => x"00",
         10750 => x"98",
         10751 => x"01",
         10752 => x"00",
         10753 => x"00",
         10754 => x"98",
         10755 => x"01",
         10756 => x"00",
         10757 => x"00",
         10758 => x"98",
         10759 => x"03",
         10760 => x"00",
         10761 => x"00",
         10762 => x"98",
         10763 => x"03",
         10764 => x"00",
         10765 => x"00",
         10766 => x"98",
         10767 => x"03",
         10768 => x"00",
         10769 => x"00",
         10770 => x"98",
         10771 => x"04",
         10772 => x"00",
         10773 => x"00",
         10774 => x"98",
         10775 => x"04",
         10776 => x"00",
         10777 => x"00",
         10778 => x"98",
         10779 => x"04",
         10780 => x"00",
         10781 => x"00",
         10782 => x"98",
         10783 => x"04",
         10784 => x"00",
         10785 => x"00",
         10786 => x"98",
         10787 => x"04",
         10788 => x"00",
         10789 => x"00",
         10790 => x"98",
         10791 => x"04",
         10792 => x"00",
         10793 => x"00",
         10794 => x"98",
         10795 => x"04",
         10796 => x"00",
         10797 => x"00",
         10798 => x"98",
         10799 => x"05",
         10800 => x"00",
         10801 => x"00",
         10802 => x"98",
         10803 => x"05",
         10804 => x"00",
         10805 => x"00",
         10806 => x"98",
         10807 => x"05",
         10808 => x"00",
         10809 => x"00",
         10810 => x"98",
         10811 => x"05",
         10812 => x"00",
         10813 => x"00",
         10814 => x"98",
         10815 => x"07",
         10816 => x"00",
         10817 => x"00",
         10818 => x"98",
         10819 => x"07",
         10820 => x"00",
         10821 => x"00",
         10822 => x"98",
         10823 => x"08",
         10824 => x"00",
         10825 => x"00",
         10826 => x"98",
         10827 => x"08",
         10828 => x"00",
         10829 => x"00",
         10830 => x"98",
         10831 => x"08",
         10832 => x"00",
         10833 => x"00",
         10834 => x"98",
         10835 => x"08",
         10836 => x"00",
         10837 => x"00",
         10838 => x"98",
         10839 => x"09",
         10840 => x"00",
         10841 => x"00",
         10842 => x"98",
         10843 => x"09",
         10844 => x"00",
         10845 => x"00",
         10846 => x"98",
         10847 => x"09",
         10848 => x"00",
         10849 => x"00",
         10850 => x"99",
         10851 => x"09",
         10852 => x"00",
         10853 => x"00",
         10854 => x"00",
         10855 => x"00",
         10856 => x"7f",
         10857 => x"00",
         10858 => x"7f",
         10859 => x"00",
         10860 => x"7f",
         10861 => x"00",
         10862 => x"00",
         10863 => x"00",
         10864 => x"ff",
         10865 => x"00",
         10866 => x"00",
         10867 => x"78",
         10868 => x"00",
         10869 => x"e1",
         10870 => x"e1",
         10871 => x"e1",
         10872 => x"00",
         10873 => x"01",
         10874 => x"01",
         10875 => x"10",
         10876 => x"00",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"00",
         10884 => x"00",
         10885 => x"00",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"00",
         10890 => x"00",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"00",
         10895 => x"00",
         10896 => x"00",
         10897 => x"00",
         10898 => x"00",
         10899 => x"00",
         10900 => x"00",
         10901 => x"a2",
         10902 => x"00",
         10903 => x"a2",
         10904 => x"00",
         10905 => x"a2",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"85",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"80",
           387 => x"82",
           388 => x"84",
           389 => x"82",
           390 => x"b3",
           391 => x"d5",
           392 => x"80",
           393 => x"d5",
           394 => x"e3",
           395 => x"84",
           396 => x"90",
           397 => x"84",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"82",
           403 => x"84",
           404 => x"82",
           405 => x"b1",
           406 => x"d5",
           407 => x"80",
           408 => x"d5",
           409 => x"d0",
           410 => x"d5",
           411 => x"80",
           412 => x"d5",
           413 => x"cb",
           414 => x"d5",
           415 => x"80",
           416 => x"d5",
           417 => x"d8",
           418 => x"84",
           419 => x"90",
           420 => x"84",
           421 => x"2d",
           422 => x"08",
           423 => x"04",
           424 => x"0c",
           425 => x"82",
           426 => x"84",
           427 => x"82",
           428 => x"80",
           429 => x"82",
           430 => x"84",
           431 => x"82",
           432 => x"80",
           433 => x"82",
           434 => x"84",
           435 => x"82",
           436 => x"80",
           437 => x"82",
           438 => x"84",
           439 => x"82",
           440 => x"80",
           441 => x"82",
           442 => x"84",
           443 => x"82",
           444 => x"80",
           445 => x"82",
           446 => x"84",
           447 => x"82",
           448 => x"81",
           449 => x"82",
           450 => x"84",
           451 => x"82",
           452 => x"81",
           453 => x"82",
           454 => x"84",
           455 => x"82",
           456 => x"81",
           457 => x"82",
           458 => x"84",
           459 => x"82",
           460 => x"81",
           461 => x"82",
           462 => x"84",
           463 => x"82",
           464 => x"81",
           465 => x"82",
           466 => x"84",
           467 => x"82",
           468 => x"82",
           469 => x"82",
           470 => x"84",
           471 => x"82",
           472 => x"81",
           473 => x"82",
           474 => x"84",
           475 => x"82",
           476 => x"82",
           477 => x"82",
           478 => x"84",
           479 => x"82",
           480 => x"82",
           481 => x"82",
           482 => x"84",
           483 => x"82",
           484 => x"82",
           485 => x"82",
           486 => x"84",
           487 => x"82",
           488 => x"82",
           489 => x"82",
           490 => x"84",
           491 => x"82",
           492 => x"82",
           493 => x"82",
           494 => x"84",
           495 => x"82",
           496 => x"82",
           497 => x"82",
           498 => x"84",
           499 => x"82",
           500 => x"82",
           501 => x"82",
           502 => x"84",
           503 => x"82",
           504 => x"82",
           505 => x"82",
           506 => x"84",
           507 => x"82",
           508 => x"82",
           509 => x"82",
           510 => x"84",
           511 => x"82",
           512 => x"81",
           513 => x"82",
           514 => x"84",
           515 => x"82",
           516 => x"81",
           517 => x"82",
           518 => x"84",
           519 => x"82",
           520 => x"81",
           521 => x"82",
           522 => x"84",
           523 => x"82",
           524 => x"82",
           525 => x"82",
           526 => x"84",
           527 => x"82",
           528 => x"82",
           529 => x"82",
           530 => x"84",
           531 => x"82",
           532 => x"82",
           533 => x"82",
           534 => x"84",
           535 => x"82",
           536 => x"82",
           537 => x"82",
           538 => x"84",
           539 => x"82",
           540 => x"81",
           541 => x"82",
           542 => x"84",
           543 => x"82",
           544 => x"82",
           545 => x"82",
           546 => x"84",
           547 => x"82",
           548 => x"82",
           549 => x"82",
           550 => x"84",
           551 => x"82",
           552 => x"82",
           553 => x"82",
           554 => x"84",
           555 => x"82",
           556 => x"81",
           557 => x"82",
           558 => x"84",
           559 => x"82",
           560 => x"81",
           561 => x"82",
           562 => x"84",
           563 => x"82",
           564 => x"81",
           565 => x"82",
           566 => x"84",
           567 => x"82",
           568 => x"80",
           569 => x"82",
           570 => x"84",
           571 => x"82",
           572 => x"80",
           573 => x"82",
           574 => x"84",
           575 => x"82",
           576 => x"80",
           577 => x"82",
           578 => x"84",
           579 => x"82",
           580 => x"80",
           581 => x"82",
           582 => x"84",
           583 => x"82",
           584 => x"81",
           585 => x"82",
           586 => x"84",
           587 => x"82",
           588 => x"81",
           589 => x"82",
           590 => x"84",
           591 => x"82",
           592 => x"81",
           593 => x"82",
           594 => x"84",
           595 => x"82",
           596 => x"81",
           597 => x"82",
           598 => x"84",
           599 => x"3c",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"51",
           609 => x"73",
           610 => x"73",
           611 => x"81",
           612 => x"10",
           613 => x"07",
           614 => x"0c",
           615 => x"72",
           616 => x"81",
           617 => x"09",
           618 => x"71",
           619 => x"0a",
           620 => x"72",
           621 => x"51",
           622 => x"82",
           623 => x"82",
           624 => x"8e",
           625 => x"70",
           626 => x"0c",
           627 => x"93",
           628 => x"81",
           629 => x"ec",
           630 => x"d5",
           631 => x"82",
           632 => x"fb",
           633 => x"d5",
           634 => x"05",
           635 => x"84",
           636 => x"0c",
           637 => x"08",
           638 => x"54",
           639 => x"08",
           640 => x"53",
           641 => x"08",
           642 => x"9a",
           643 => x"f8",
           644 => x"d5",
           645 => x"05",
           646 => x"84",
           647 => x"08",
           648 => x"f8",
           649 => x"87",
           650 => x"d5",
           651 => x"82",
           652 => x"02",
           653 => x"0c",
           654 => x"82",
           655 => x"90",
           656 => x"11",
           657 => x"32",
           658 => x"51",
           659 => x"71",
           660 => x"0b",
           661 => x"08",
           662 => x"25",
           663 => x"39",
           664 => x"d5",
           665 => x"05",
           666 => x"39",
           667 => x"08",
           668 => x"ff",
           669 => x"84",
           670 => x"0c",
           671 => x"d5",
           672 => x"05",
           673 => x"84",
           674 => x"08",
           675 => x"08",
           676 => x"82",
           677 => x"f8",
           678 => x"2e",
           679 => x"80",
           680 => x"84",
           681 => x"08",
           682 => x"38",
           683 => x"08",
           684 => x"51",
           685 => x"82",
           686 => x"70",
           687 => x"08",
           688 => x"52",
           689 => x"08",
           690 => x"ff",
           691 => x"06",
           692 => x"0b",
           693 => x"08",
           694 => x"80",
           695 => x"d5",
           696 => x"05",
           697 => x"84",
           698 => x"08",
           699 => x"73",
           700 => x"84",
           701 => x"08",
           702 => x"d5",
           703 => x"05",
           704 => x"84",
           705 => x"08",
           706 => x"d5",
           707 => x"05",
           708 => x"39",
           709 => x"08",
           710 => x"52",
           711 => x"82",
           712 => x"88",
           713 => x"82",
           714 => x"f4",
           715 => x"82",
           716 => x"f4",
           717 => x"d4",
           718 => x"3d",
           719 => x"84",
           720 => x"d5",
           721 => x"82",
           722 => x"f4",
           723 => x"0b",
           724 => x"08",
           725 => x"82",
           726 => x"88",
           727 => x"d5",
           728 => x"05",
           729 => x"0b",
           730 => x"08",
           731 => x"82",
           732 => x"90",
           733 => x"d5",
           734 => x"05",
           735 => x"84",
           736 => x"08",
           737 => x"84",
           738 => x"08",
           739 => x"84",
           740 => x"70",
           741 => x"81",
           742 => x"d4",
           743 => x"82",
           744 => x"dc",
           745 => x"d5",
           746 => x"05",
           747 => x"84",
           748 => x"08",
           749 => x"80",
           750 => x"d5",
           751 => x"05",
           752 => x"d4",
           753 => x"8e",
           754 => x"d5",
           755 => x"82",
           756 => x"02",
           757 => x"0c",
           758 => x"82",
           759 => x"90",
           760 => x"d5",
           761 => x"05",
           762 => x"84",
           763 => x"08",
           764 => x"84",
           765 => x"08",
           766 => x"84",
           767 => x"08",
           768 => x"3f",
           769 => x"08",
           770 => x"84",
           771 => x"0c",
           772 => x"08",
           773 => x"70",
           774 => x"0c",
           775 => x"3d",
           776 => x"84",
           777 => x"d5",
           778 => x"82",
           779 => x"ed",
           780 => x"0b",
           781 => x"08",
           782 => x"82",
           783 => x"88",
           784 => x"80",
           785 => x"0c",
           786 => x"08",
           787 => x"85",
           788 => x"81",
           789 => x"32",
           790 => x"51",
           791 => x"53",
           792 => x"8d",
           793 => x"82",
           794 => x"e0",
           795 => x"ac",
           796 => x"84",
           797 => x"08",
           798 => x"53",
           799 => x"84",
           800 => x"34",
           801 => x"06",
           802 => x"2e",
           803 => x"82",
           804 => x"8c",
           805 => x"05",
           806 => x"08",
           807 => x"82",
           808 => x"e4",
           809 => x"81",
           810 => x"72",
           811 => x"8b",
           812 => x"84",
           813 => x"33",
           814 => x"27",
           815 => x"82",
           816 => x"f8",
           817 => x"72",
           818 => x"ee",
           819 => x"84",
           820 => x"33",
           821 => x"2e",
           822 => x"80",
           823 => x"d5",
           824 => x"05",
           825 => x"2b",
           826 => x"51",
           827 => x"b2",
           828 => x"84",
           829 => x"22",
           830 => x"70",
           831 => x"81",
           832 => x"51",
           833 => x"2e",
           834 => x"d5",
           835 => x"05",
           836 => x"80",
           837 => x"72",
           838 => x"08",
           839 => x"fe",
           840 => x"d5",
           841 => x"05",
           842 => x"2b",
           843 => x"70",
           844 => x"72",
           845 => x"51",
           846 => x"51",
           847 => x"82",
           848 => x"e8",
           849 => x"d5",
           850 => x"05",
           851 => x"d5",
           852 => x"05",
           853 => x"d0",
           854 => x"53",
           855 => x"84",
           856 => x"34",
           857 => x"08",
           858 => x"70",
           859 => x"98",
           860 => x"53",
           861 => x"8b",
           862 => x"0b",
           863 => x"08",
           864 => x"82",
           865 => x"e4",
           866 => x"83",
           867 => x"06",
           868 => x"72",
           869 => x"82",
           870 => x"e8",
           871 => x"88",
           872 => x"2b",
           873 => x"70",
           874 => x"51",
           875 => x"72",
           876 => x"08",
           877 => x"fd",
           878 => x"d5",
           879 => x"05",
           880 => x"2a",
           881 => x"51",
           882 => x"80",
           883 => x"82",
           884 => x"e8",
           885 => x"98",
           886 => x"2c",
           887 => x"72",
           888 => x"0b",
           889 => x"08",
           890 => x"82",
           891 => x"f8",
           892 => x"11",
           893 => x"08",
           894 => x"53",
           895 => x"08",
           896 => x"80",
           897 => x"94",
           898 => x"84",
           899 => x"08",
           900 => x"82",
           901 => x"70",
           902 => x"51",
           903 => x"82",
           904 => x"e4",
           905 => x"90",
           906 => x"72",
           907 => x"08",
           908 => x"82",
           909 => x"e4",
           910 => x"a0",
           911 => x"72",
           912 => x"08",
           913 => x"fc",
           914 => x"d5",
           915 => x"05",
           916 => x"80",
           917 => x"72",
           918 => x"08",
           919 => x"fc",
           920 => x"d5",
           921 => x"05",
           922 => x"c0",
           923 => x"72",
           924 => x"08",
           925 => x"fb",
           926 => x"d5",
           927 => x"05",
           928 => x"07",
           929 => x"82",
           930 => x"e4",
           931 => x"0b",
           932 => x"08",
           933 => x"fb",
           934 => x"d5",
           935 => x"05",
           936 => x"07",
           937 => x"82",
           938 => x"e4",
           939 => x"c1",
           940 => x"82",
           941 => x"fc",
           942 => x"d5",
           943 => x"05",
           944 => x"51",
           945 => x"d5",
           946 => x"05",
           947 => x"0b",
           948 => x"08",
           949 => x"8d",
           950 => x"d5",
           951 => x"05",
           952 => x"84",
           953 => x"08",
           954 => x"d5",
           955 => x"05",
           956 => x"51",
           957 => x"d5",
           958 => x"05",
           959 => x"84",
           960 => x"22",
           961 => x"53",
           962 => x"84",
           963 => x"23",
           964 => x"82",
           965 => x"90",
           966 => x"d5",
           967 => x"05",
           968 => x"82",
           969 => x"90",
           970 => x"08",
           971 => x"08",
           972 => x"82",
           973 => x"e4",
           974 => x"83",
           975 => x"06",
           976 => x"53",
           977 => x"ab",
           978 => x"84",
           979 => x"33",
           980 => x"53",
           981 => x"53",
           982 => x"08",
           983 => x"52",
           984 => x"3f",
           985 => x"08",
           986 => x"d5",
           987 => x"05",
           988 => x"82",
           989 => x"fc",
           990 => x"9d",
           991 => x"d4",
           992 => x"72",
           993 => x"08",
           994 => x"82",
           995 => x"ec",
           996 => x"82",
           997 => x"f4",
           998 => x"71",
           999 => x"72",
          1000 => x"08",
          1001 => x"8b",
          1002 => x"d5",
          1003 => x"05",
          1004 => x"84",
          1005 => x"08",
          1006 => x"d5",
          1007 => x"05",
          1008 => x"82",
          1009 => x"fc",
          1010 => x"d5",
          1011 => x"05",
          1012 => x"2a",
          1013 => x"51",
          1014 => x"72",
          1015 => x"38",
          1016 => x"08",
          1017 => x"70",
          1018 => x"72",
          1019 => x"82",
          1020 => x"fc",
          1021 => x"53",
          1022 => x"82",
          1023 => x"53",
          1024 => x"84",
          1025 => x"23",
          1026 => x"d5",
          1027 => x"05",
          1028 => x"f3",
          1029 => x"f8",
          1030 => x"82",
          1031 => x"f4",
          1032 => x"d5",
          1033 => x"05",
          1034 => x"d5",
          1035 => x"05",
          1036 => x"31",
          1037 => x"82",
          1038 => x"ec",
          1039 => x"c1",
          1040 => x"84",
          1041 => x"22",
          1042 => x"70",
          1043 => x"51",
          1044 => x"2e",
          1045 => x"d5",
          1046 => x"05",
          1047 => x"84",
          1048 => x"08",
          1049 => x"d5",
          1050 => x"05",
          1051 => x"82",
          1052 => x"dc",
          1053 => x"a2",
          1054 => x"84",
          1055 => x"08",
          1056 => x"08",
          1057 => x"84",
          1058 => x"84",
          1059 => x"0c",
          1060 => x"d5",
          1061 => x"05",
          1062 => x"d5",
          1063 => x"05",
          1064 => x"84",
          1065 => x"0c",
          1066 => x"08",
          1067 => x"80",
          1068 => x"82",
          1069 => x"e4",
          1070 => x"82",
          1071 => x"72",
          1072 => x"08",
          1073 => x"82",
          1074 => x"fc",
          1075 => x"82",
          1076 => x"fc",
          1077 => x"d5",
          1078 => x"05",
          1079 => x"bf",
          1080 => x"72",
          1081 => x"08",
          1082 => x"81",
          1083 => x"0b",
          1084 => x"08",
          1085 => x"a9",
          1086 => x"84",
          1087 => x"22",
          1088 => x"07",
          1089 => x"82",
          1090 => x"e4",
          1091 => x"f8",
          1092 => x"84",
          1093 => x"34",
          1094 => x"d5",
          1095 => x"05",
          1096 => x"84",
          1097 => x"22",
          1098 => x"70",
          1099 => x"51",
          1100 => x"2e",
          1101 => x"d5",
          1102 => x"05",
          1103 => x"84",
          1104 => x"08",
          1105 => x"d5",
          1106 => x"05",
          1107 => x"82",
          1108 => x"d8",
          1109 => x"a2",
          1110 => x"84",
          1111 => x"08",
          1112 => x"08",
          1113 => x"84",
          1114 => x"84",
          1115 => x"0c",
          1116 => x"d5",
          1117 => x"05",
          1118 => x"d5",
          1119 => x"05",
          1120 => x"84",
          1121 => x"0c",
          1122 => x"08",
          1123 => x"70",
          1124 => x"53",
          1125 => x"84",
          1126 => x"23",
          1127 => x"0b",
          1128 => x"08",
          1129 => x"82",
          1130 => x"f0",
          1131 => x"d5",
          1132 => x"05",
          1133 => x"84",
          1134 => x"08",
          1135 => x"54",
          1136 => x"a5",
          1137 => x"d4",
          1138 => x"72",
          1139 => x"d5",
          1140 => x"05",
          1141 => x"84",
          1142 => x"0c",
          1143 => x"08",
          1144 => x"70",
          1145 => x"89",
          1146 => x"38",
          1147 => x"08",
          1148 => x"53",
          1149 => x"82",
          1150 => x"f8",
          1151 => x"15",
          1152 => x"51",
          1153 => x"d5",
          1154 => x"05",
          1155 => x"82",
          1156 => x"f0",
          1157 => x"72",
          1158 => x"51",
          1159 => x"d5",
          1160 => x"05",
          1161 => x"84",
          1162 => x"08",
          1163 => x"84",
          1164 => x"33",
          1165 => x"d5",
          1166 => x"05",
          1167 => x"82",
          1168 => x"f0",
          1169 => x"d5",
          1170 => x"05",
          1171 => x"82",
          1172 => x"fc",
          1173 => x"53",
          1174 => x"82",
          1175 => x"70",
          1176 => x"08",
          1177 => x"53",
          1178 => x"08",
          1179 => x"80",
          1180 => x"fe",
          1181 => x"d5",
          1182 => x"05",
          1183 => x"88",
          1184 => x"54",
          1185 => x"31",
          1186 => x"82",
          1187 => x"fc",
          1188 => x"d5",
          1189 => x"05",
          1190 => x"06",
          1191 => x"80",
          1192 => x"82",
          1193 => x"ec",
          1194 => x"11",
          1195 => x"82",
          1196 => x"ec",
          1197 => x"d5",
          1198 => x"05",
          1199 => x"2a",
          1200 => x"51",
          1201 => x"80",
          1202 => x"38",
          1203 => x"08",
          1204 => x"70",
          1205 => x"d5",
          1206 => x"05",
          1207 => x"84",
          1208 => x"08",
          1209 => x"d5",
          1210 => x"05",
          1211 => x"84",
          1212 => x"22",
          1213 => x"90",
          1214 => x"06",
          1215 => x"d5",
          1216 => x"05",
          1217 => x"53",
          1218 => x"84",
          1219 => x"23",
          1220 => x"d5",
          1221 => x"05",
          1222 => x"53",
          1223 => x"84",
          1224 => x"23",
          1225 => x"08",
          1226 => x"82",
          1227 => x"ec",
          1228 => x"d5",
          1229 => x"05",
          1230 => x"2a",
          1231 => x"51",
          1232 => x"80",
          1233 => x"38",
          1234 => x"08",
          1235 => x"70",
          1236 => x"98",
          1237 => x"84",
          1238 => x"33",
          1239 => x"53",
          1240 => x"97",
          1241 => x"84",
          1242 => x"22",
          1243 => x"51",
          1244 => x"d5",
          1245 => x"05",
          1246 => x"82",
          1247 => x"e8",
          1248 => x"82",
          1249 => x"fc",
          1250 => x"71",
          1251 => x"72",
          1252 => x"08",
          1253 => x"82",
          1254 => x"e4",
          1255 => x"83",
          1256 => x"06",
          1257 => x"72",
          1258 => x"38",
          1259 => x"08",
          1260 => x"70",
          1261 => x"90",
          1262 => x"2c",
          1263 => x"51",
          1264 => x"53",
          1265 => x"d5",
          1266 => x"05",
          1267 => x"31",
          1268 => x"82",
          1269 => x"ec",
          1270 => x"39",
          1271 => x"08",
          1272 => x"70",
          1273 => x"90",
          1274 => x"2c",
          1275 => x"51",
          1276 => x"53",
          1277 => x"d5",
          1278 => x"05",
          1279 => x"31",
          1280 => x"82",
          1281 => x"ec",
          1282 => x"d5",
          1283 => x"05",
          1284 => x"80",
          1285 => x"72",
          1286 => x"d5",
          1287 => x"05",
          1288 => x"54",
          1289 => x"d5",
          1290 => x"05",
          1291 => x"2b",
          1292 => x"51",
          1293 => x"25",
          1294 => x"d5",
          1295 => x"05",
          1296 => x"51",
          1297 => x"d2",
          1298 => x"84",
          1299 => x"22",
          1300 => x"70",
          1301 => x"51",
          1302 => x"2e",
          1303 => x"d5",
          1304 => x"05",
          1305 => x"51",
          1306 => x"80",
          1307 => x"d5",
          1308 => x"05",
          1309 => x"2a",
          1310 => x"51",
          1311 => x"80",
          1312 => x"82",
          1313 => x"88",
          1314 => x"ab",
          1315 => x"3f",
          1316 => x"d5",
          1317 => x"05",
          1318 => x"2a",
          1319 => x"51",
          1320 => x"80",
          1321 => x"82",
          1322 => x"88",
          1323 => x"a0",
          1324 => x"3f",
          1325 => x"08",
          1326 => x"70",
          1327 => x"81",
          1328 => x"53",
          1329 => x"b1",
          1330 => x"84",
          1331 => x"08",
          1332 => x"89",
          1333 => x"d5",
          1334 => x"05",
          1335 => x"90",
          1336 => x"06",
          1337 => x"d5",
          1338 => x"05",
          1339 => x"d5",
          1340 => x"05",
          1341 => x"bc",
          1342 => x"84",
          1343 => x"22",
          1344 => x"70",
          1345 => x"51",
          1346 => x"2e",
          1347 => x"d5",
          1348 => x"05",
          1349 => x"54",
          1350 => x"d5",
          1351 => x"05",
          1352 => x"2b",
          1353 => x"51",
          1354 => x"25",
          1355 => x"d5",
          1356 => x"05",
          1357 => x"51",
          1358 => x"d2",
          1359 => x"84",
          1360 => x"22",
          1361 => x"70",
          1362 => x"51",
          1363 => x"2e",
          1364 => x"d5",
          1365 => x"05",
          1366 => x"54",
          1367 => x"d5",
          1368 => x"05",
          1369 => x"2b",
          1370 => x"51",
          1371 => x"25",
          1372 => x"d5",
          1373 => x"05",
          1374 => x"51",
          1375 => x"d2",
          1376 => x"84",
          1377 => x"22",
          1378 => x"70",
          1379 => x"51",
          1380 => x"38",
          1381 => x"08",
          1382 => x"ff",
          1383 => x"72",
          1384 => x"08",
          1385 => x"73",
          1386 => x"90",
          1387 => x"80",
          1388 => x"38",
          1389 => x"08",
          1390 => x"52",
          1391 => x"f4",
          1392 => x"82",
          1393 => x"f8",
          1394 => x"72",
          1395 => x"09",
          1396 => x"38",
          1397 => x"08",
          1398 => x"52",
          1399 => x"08",
          1400 => x"51",
          1401 => x"81",
          1402 => x"d5",
          1403 => x"05",
          1404 => x"80",
          1405 => x"81",
          1406 => x"38",
          1407 => x"08",
          1408 => x"ff",
          1409 => x"72",
          1410 => x"08",
          1411 => x"72",
          1412 => x"06",
          1413 => x"ff",
          1414 => x"bb",
          1415 => x"84",
          1416 => x"08",
          1417 => x"84",
          1418 => x"08",
          1419 => x"82",
          1420 => x"fc",
          1421 => x"05",
          1422 => x"08",
          1423 => x"53",
          1424 => x"ff",
          1425 => x"d5",
          1426 => x"05",
          1427 => x"80",
          1428 => x"81",
          1429 => x"38",
          1430 => x"08",
          1431 => x"ff",
          1432 => x"72",
          1433 => x"08",
          1434 => x"72",
          1435 => x"06",
          1436 => x"ff",
          1437 => x"df",
          1438 => x"84",
          1439 => x"08",
          1440 => x"84",
          1441 => x"08",
          1442 => x"53",
          1443 => x"82",
          1444 => x"fc",
          1445 => x"05",
          1446 => x"08",
          1447 => x"ff",
          1448 => x"d5",
          1449 => x"05",
          1450 => x"88",
          1451 => x"82",
          1452 => x"88",
          1453 => x"82",
          1454 => x"f0",
          1455 => x"05",
          1456 => x"08",
          1457 => x"82",
          1458 => x"f0",
          1459 => x"33",
          1460 => x"e0",
          1461 => x"82",
          1462 => x"e4",
          1463 => x"87",
          1464 => x"06",
          1465 => x"72",
          1466 => x"c3",
          1467 => x"84",
          1468 => x"22",
          1469 => x"54",
          1470 => x"84",
          1471 => x"23",
          1472 => x"70",
          1473 => x"53",
          1474 => x"a3",
          1475 => x"84",
          1476 => x"08",
          1477 => x"85",
          1478 => x"39",
          1479 => x"08",
          1480 => x"52",
          1481 => x"08",
          1482 => x"51",
          1483 => x"80",
          1484 => x"84",
          1485 => x"23",
          1486 => x"82",
          1487 => x"f8",
          1488 => x"72",
          1489 => x"81",
          1490 => x"81",
          1491 => x"84",
          1492 => x"23",
          1493 => x"d5",
          1494 => x"05",
          1495 => x"82",
          1496 => x"e8",
          1497 => x"0b",
          1498 => x"08",
          1499 => x"ea",
          1500 => x"d5",
          1501 => x"05",
          1502 => x"d5",
          1503 => x"05",
          1504 => x"b0",
          1505 => x"39",
          1506 => x"08",
          1507 => x"8c",
          1508 => x"82",
          1509 => x"e0",
          1510 => x"53",
          1511 => x"08",
          1512 => x"82",
          1513 => x"95",
          1514 => x"d5",
          1515 => x"82",
          1516 => x"02",
          1517 => x"0c",
          1518 => x"82",
          1519 => x"53",
          1520 => x"08",
          1521 => x"52",
          1522 => x"08",
          1523 => x"51",
          1524 => x"82",
          1525 => x"70",
          1526 => x"0c",
          1527 => x"0d",
          1528 => x"0c",
          1529 => x"84",
          1530 => x"d5",
          1531 => x"3d",
          1532 => x"82",
          1533 => x"f8",
          1534 => x"f0",
          1535 => x"11",
          1536 => x"2a",
          1537 => x"70",
          1538 => x"51",
          1539 => x"72",
          1540 => x"38",
          1541 => x"d5",
          1542 => x"05",
          1543 => x"39",
          1544 => x"08",
          1545 => x"53",
          1546 => x"d5",
          1547 => x"05",
          1548 => x"82",
          1549 => x"88",
          1550 => x"72",
          1551 => x"08",
          1552 => x"72",
          1553 => x"53",
          1554 => x"b0",
          1555 => x"dc",
          1556 => x"dc",
          1557 => x"d5",
          1558 => x"05",
          1559 => x"11",
          1560 => x"72",
          1561 => x"f8",
          1562 => x"80",
          1563 => x"38",
          1564 => x"d5",
          1565 => x"05",
          1566 => x"39",
          1567 => x"08",
          1568 => x"08",
          1569 => x"51",
          1570 => x"53",
          1571 => x"d4",
          1572 => x"72",
          1573 => x"38",
          1574 => x"d5",
          1575 => x"05",
          1576 => x"84",
          1577 => x"08",
          1578 => x"84",
          1579 => x"0c",
          1580 => x"84",
          1581 => x"08",
          1582 => x"0c",
          1583 => x"82",
          1584 => x"04",
          1585 => x"08",
          1586 => x"84",
          1587 => x"0d",
          1588 => x"d5",
          1589 => x"05",
          1590 => x"84",
          1591 => x"08",
          1592 => x"70",
          1593 => x"81",
          1594 => x"06",
          1595 => x"51",
          1596 => x"2e",
          1597 => x"0b",
          1598 => x"08",
          1599 => x"80",
          1600 => x"d5",
          1601 => x"05",
          1602 => x"33",
          1603 => x"08",
          1604 => x"81",
          1605 => x"84",
          1606 => x"0c",
          1607 => x"d5",
          1608 => x"05",
          1609 => x"ff",
          1610 => x"80",
          1611 => x"82",
          1612 => x"8c",
          1613 => x"d5",
          1614 => x"05",
          1615 => x"d5",
          1616 => x"05",
          1617 => x"11",
          1618 => x"72",
          1619 => x"f8",
          1620 => x"80",
          1621 => x"38",
          1622 => x"d5",
          1623 => x"05",
          1624 => x"39",
          1625 => x"08",
          1626 => x"70",
          1627 => x"08",
          1628 => x"53",
          1629 => x"08",
          1630 => x"82",
          1631 => x"87",
          1632 => x"d5",
          1633 => x"82",
          1634 => x"02",
          1635 => x"0c",
          1636 => x"82",
          1637 => x"52",
          1638 => x"08",
          1639 => x"51",
          1640 => x"d4",
          1641 => x"82",
          1642 => x"53",
          1643 => x"82",
          1644 => x"04",
          1645 => x"08",
          1646 => x"84",
          1647 => x"0d",
          1648 => x"08",
          1649 => x"85",
          1650 => x"81",
          1651 => x"32",
          1652 => x"51",
          1653 => x"53",
          1654 => x"8d",
          1655 => x"82",
          1656 => x"fc",
          1657 => x"cb",
          1658 => x"84",
          1659 => x"08",
          1660 => x"70",
          1661 => x"81",
          1662 => x"51",
          1663 => x"2e",
          1664 => x"82",
          1665 => x"8c",
          1666 => x"d5",
          1667 => x"05",
          1668 => x"8c",
          1669 => x"14",
          1670 => x"38",
          1671 => x"08",
          1672 => x"70",
          1673 => x"d5",
          1674 => x"05",
          1675 => x"54",
          1676 => x"34",
          1677 => x"05",
          1678 => x"d5",
          1679 => x"05",
          1680 => x"08",
          1681 => x"12",
          1682 => x"84",
          1683 => x"08",
          1684 => x"84",
          1685 => x"0c",
          1686 => x"d7",
          1687 => x"84",
          1688 => x"08",
          1689 => x"08",
          1690 => x"53",
          1691 => x"08",
          1692 => x"70",
          1693 => x"53",
          1694 => x"51",
          1695 => x"2d",
          1696 => x"08",
          1697 => x"38",
          1698 => x"08",
          1699 => x"8c",
          1700 => x"05",
          1701 => x"82",
          1702 => x"88",
          1703 => x"82",
          1704 => x"fc",
          1705 => x"53",
          1706 => x"0b",
          1707 => x"08",
          1708 => x"82",
          1709 => x"fc",
          1710 => x"d4",
          1711 => x"3d",
          1712 => x"84",
          1713 => x"d5",
          1714 => x"82",
          1715 => x"f9",
          1716 => x"d5",
          1717 => x"05",
          1718 => x"33",
          1719 => x"70",
          1720 => x"51",
          1721 => x"80",
          1722 => x"ff",
          1723 => x"84",
          1724 => x"0c",
          1725 => x"82",
          1726 => x"88",
          1727 => x"11",
          1728 => x"2a",
          1729 => x"51",
          1730 => x"71",
          1731 => x"c5",
          1732 => x"84",
          1733 => x"08",
          1734 => x"08",
          1735 => x"53",
          1736 => x"33",
          1737 => x"06",
          1738 => x"85",
          1739 => x"d5",
          1740 => x"05",
          1741 => x"08",
          1742 => x"12",
          1743 => x"84",
          1744 => x"08",
          1745 => x"70",
          1746 => x"08",
          1747 => x"51",
          1748 => x"b6",
          1749 => x"84",
          1750 => x"08",
          1751 => x"70",
          1752 => x"81",
          1753 => x"51",
          1754 => x"2e",
          1755 => x"82",
          1756 => x"88",
          1757 => x"08",
          1758 => x"d5",
          1759 => x"05",
          1760 => x"82",
          1761 => x"fc",
          1762 => x"38",
          1763 => x"08",
          1764 => x"82",
          1765 => x"88",
          1766 => x"53",
          1767 => x"70",
          1768 => x"52",
          1769 => x"34",
          1770 => x"d5",
          1771 => x"05",
          1772 => x"39",
          1773 => x"08",
          1774 => x"70",
          1775 => x"71",
          1776 => x"a1",
          1777 => x"84",
          1778 => x"08",
          1779 => x"08",
          1780 => x"52",
          1781 => x"51",
          1782 => x"82",
          1783 => x"70",
          1784 => x"08",
          1785 => x"52",
          1786 => x"08",
          1787 => x"80",
          1788 => x"38",
          1789 => x"08",
          1790 => x"82",
          1791 => x"f4",
          1792 => x"d5",
          1793 => x"05",
          1794 => x"33",
          1795 => x"08",
          1796 => x"52",
          1797 => x"08",
          1798 => x"ff",
          1799 => x"06",
          1800 => x"d5",
          1801 => x"05",
          1802 => x"52",
          1803 => x"84",
          1804 => x"34",
          1805 => x"d5",
          1806 => x"05",
          1807 => x"52",
          1808 => x"84",
          1809 => x"34",
          1810 => x"08",
          1811 => x"52",
          1812 => x"08",
          1813 => x"85",
          1814 => x"0b",
          1815 => x"08",
          1816 => x"a6",
          1817 => x"84",
          1818 => x"08",
          1819 => x"81",
          1820 => x"0c",
          1821 => x"08",
          1822 => x"70",
          1823 => x"70",
          1824 => x"08",
          1825 => x"51",
          1826 => x"d5",
          1827 => x"05",
          1828 => x"f8",
          1829 => x"0d",
          1830 => x"0c",
          1831 => x"84",
          1832 => x"d5",
          1833 => x"3d",
          1834 => x"84",
          1835 => x"08",
          1836 => x"08",
          1837 => x"82",
          1838 => x"8c",
          1839 => x"d5",
          1840 => x"05",
          1841 => x"84",
          1842 => x"08",
          1843 => x"a2",
          1844 => x"84",
          1845 => x"08",
          1846 => x"08",
          1847 => x"26",
          1848 => x"82",
          1849 => x"f8",
          1850 => x"d5",
          1851 => x"05",
          1852 => x"82",
          1853 => x"fc",
          1854 => x"27",
          1855 => x"82",
          1856 => x"fc",
          1857 => x"d5",
          1858 => x"05",
          1859 => x"d5",
          1860 => x"05",
          1861 => x"84",
          1862 => x"08",
          1863 => x"08",
          1864 => x"05",
          1865 => x"08",
          1866 => x"82",
          1867 => x"90",
          1868 => x"05",
          1869 => x"08",
          1870 => x"82",
          1871 => x"90",
          1872 => x"05",
          1873 => x"08",
          1874 => x"82",
          1875 => x"90",
          1876 => x"2e",
          1877 => x"82",
          1878 => x"fc",
          1879 => x"05",
          1880 => x"08",
          1881 => x"82",
          1882 => x"f8",
          1883 => x"05",
          1884 => x"08",
          1885 => x"82",
          1886 => x"fc",
          1887 => x"d5",
          1888 => x"05",
          1889 => x"71",
          1890 => x"ff",
          1891 => x"d5",
          1892 => x"05",
          1893 => x"82",
          1894 => x"90",
          1895 => x"d5",
          1896 => x"05",
          1897 => x"82",
          1898 => x"90",
          1899 => x"d5",
          1900 => x"05",
          1901 => x"ba",
          1902 => x"84",
          1903 => x"08",
          1904 => x"82",
          1905 => x"f8",
          1906 => x"05",
          1907 => x"08",
          1908 => x"82",
          1909 => x"fc",
          1910 => x"52",
          1911 => x"82",
          1912 => x"fc",
          1913 => x"05",
          1914 => x"08",
          1915 => x"ff",
          1916 => x"d5",
          1917 => x"05",
          1918 => x"d4",
          1919 => x"85",
          1920 => x"d5",
          1921 => x"82",
          1922 => x"02",
          1923 => x"0c",
          1924 => x"82",
          1925 => x"88",
          1926 => x"d5",
          1927 => x"05",
          1928 => x"84",
          1929 => x"08",
          1930 => x"82",
          1931 => x"fc",
          1932 => x"05",
          1933 => x"08",
          1934 => x"70",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"39",
          1938 => x"08",
          1939 => x"ff",
          1940 => x"84",
          1941 => x"0c",
          1942 => x"08",
          1943 => x"82",
          1944 => x"88",
          1945 => x"70",
          1946 => x"0c",
          1947 => x"0d",
          1948 => x"0c",
          1949 => x"84",
          1950 => x"d5",
          1951 => x"3d",
          1952 => x"84",
          1953 => x"08",
          1954 => x"08",
          1955 => x"82",
          1956 => x"8c",
          1957 => x"71",
          1958 => x"84",
          1959 => x"08",
          1960 => x"d5",
          1961 => x"05",
          1962 => x"84",
          1963 => x"08",
          1964 => x"72",
          1965 => x"84",
          1966 => x"08",
          1967 => x"d5",
          1968 => x"05",
          1969 => x"ff",
          1970 => x"80",
          1971 => x"ff",
          1972 => x"d5",
          1973 => x"05",
          1974 => x"d4",
          1975 => x"84",
          1976 => x"d5",
          1977 => x"82",
          1978 => x"02",
          1979 => x"0c",
          1980 => x"82",
          1981 => x"88",
          1982 => x"d5",
          1983 => x"05",
          1984 => x"84",
          1985 => x"08",
          1986 => x"08",
          1987 => x"82",
          1988 => x"90",
          1989 => x"2e",
          1990 => x"82",
          1991 => x"90",
          1992 => x"05",
          1993 => x"08",
          1994 => x"82",
          1995 => x"90",
          1996 => x"05",
          1997 => x"08",
          1998 => x"82",
          1999 => x"90",
          2000 => x"2e",
          2001 => x"d5",
          2002 => x"05",
          2003 => x"33",
          2004 => x"08",
          2005 => x"81",
          2006 => x"84",
          2007 => x"0c",
          2008 => x"08",
          2009 => x"52",
          2010 => x"34",
          2011 => x"08",
          2012 => x"81",
          2013 => x"84",
          2014 => x"0c",
          2015 => x"82",
          2016 => x"88",
          2017 => x"82",
          2018 => x"51",
          2019 => x"82",
          2020 => x"04",
          2021 => x"08",
          2022 => x"84",
          2023 => x"0d",
          2024 => x"08",
          2025 => x"80",
          2026 => x"38",
          2027 => x"08",
          2028 => x"52",
          2029 => x"d5",
          2030 => x"05",
          2031 => x"82",
          2032 => x"8c",
          2033 => x"d5",
          2034 => x"05",
          2035 => x"72",
          2036 => x"53",
          2037 => x"71",
          2038 => x"38",
          2039 => x"82",
          2040 => x"88",
          2041 => x"71",
          2042 => x"84",
          2043 => x"08",
          2044 => x"d5",
          2045 => x"05",
          2046 => x"ff",
          2047 => x"70",
          2048 => x"0b",
          2049 => x"08",
          2050 => x"81",
          2051 => x"d5",
          2052 => x"05",
          2053 => x"82",
          2054 => x"90",
          2055 => x"d5",
          2056 => x"05",
          2057 => x"84",
          2058 => x"39",
          2059 => x"08",
          2060 => x"80",
          2061 => x"38",
          2062 => x"08",
          2063 => x"70",
          2064 => x"70",
          2065 => x"0b",
          2066 => x"08",
          2067 => x"80",
          2068 => x"d5",
          2069 => x"05",
          2070 => x"82",
          2071 => x"8c",
          2072 => x"d5",
          2073 => x"05",
          2074 => x"52",
          2075 => x"38",
          2076 => x"d5",
          2077 => x"05",
          2078 => x"82",
          2079 => x"88",
          2080 => x"33",
          2081 => x"08",
          2082 => x"70",
          2083 => x"31",
          2084 => x"84",
          2085 => x"0c",
          2086 => x"52",
          2087 => x"80",
          2088 => x"84",
          2089 => x"0c",
          2090 => x"08",
          2091 => x"82",
          2092 => x"85",
          2093 => x"d5",
          2094 => x"82",
          2095 => x"02",
          2096 => x"0c",
          2097 => x"82",
          2098 => x"8c",
          2099 => x"82",
          2100 => x"88",
          2101 => x"81",
          2102 => x"d4",
          2103 => x"82",
          2104 => x"f8",
          2105 => x"d5",
          2106 => x"05",
          2107 => x"70",
          2108 => x"80",
          2109 => x"82",
          2110 => x"70",
          2111 => x"08",
          2112 => x"54",
          2113 => x"08",
          2114 => x"8c",
          2115 => x"82",
          2116 => x"f4",
          2117 => x"39",
          2118 => x"08",
          2119 => x"82",
          2120 => x"f8",
          2121 => x"54",
          2122 => x"82",
          2123 => x"f8",
          2124 => x"82",
          2125 => x"88",
          2126 => x"82",
          2127 => x"fc",
          2128 => x"fb",
          2129 => x"d4",
          2130 => x"82",
          2131 => x"f4",
          2132 => x"82",
          2133 => x"f4",
          2134 => x"d4",
          2135 => x"3d",
          2136 => x"84",
          2137 => x"d5",
          2138 => x"82",
          2139 => x"fd",
          2140 => x"d5",
          2141 => x"05",
          2142 => x"84",
          2143 => x"0c",
          2144 => x"08",
          2145 => x"8d",
          2146 => x"82",
          2147 => x"fc",
          2148 => x"ec",
          2149 => x"84",
          2150 => x"08",
          2151 => x"82",
          2152 => x"f8",
          2153 => x"05",
          2154 => x"08",
          2155 => x"70",
          2156 => x"51",
          2157 => x"2e",
          2158 => x"d5",
          2159 => x"05",
          2160 => x"82",
          2161 => x"8c",
          2162 => x"d5",
          2163 => x"05",
          2164 => x"84",
          2165 => x"39",
          2166 => x"08",
          2167 => x"ff",
          2168 => x"84",
          2169 => x"0c",
          2170 => x"08",
          2171 => x"82",
          2172 => x"88",
          2173 => x"70",
          2174 => x"08",
          2175 => x"51",
          2176 => x"08",
          2177 => x"82",
          2178 => x"85",
          2179 => x"d5",
          2180 => x"82",
          2181 => x"02",
          2182 => x"0c",
          2183 => x"82",
          2184 => x"88",
          2185 => x"d5",
          2186 => x"05",
          2187 => x"84",
          2188 => x"08",
          2189 => x"d4",
          2190 => x"84",
          2191 => x"08",
          2192 => x"d5",
          2193 => x"05",
          2194 => x"84",
          2195 => x"08",
          2196 => x"d5",
          2197 => x"05",
          2198 => x"84",
          2199 => x"08",
          2200 => x"38",
          2201 => x"08",
          2202 => x"51",
          2203 => x"84",
          2204 => x"08",
          2205 => x"71",
          2206 => x"84",
          2207 => x"08",
          2208 => x"d5",
          2209 => x"05",
          2210 => x"39",
          2211 => x"08",
          2212 => x"70",
          2213 => x"0c",
          2214 => x"0d",
          2215 => x"0c",
          2216 => x"84",
          2217 => x"d5",
          2218 => x"3d",
          2219 => x"82",
          2220 => x"fc",
          2221 => x"d5",
          2222 => x"05",
          2223 => x"b9",
          2224 => x"84",
          2225 => x"08",
          2226 => x"84",
          2227 => x"0c",
          2228 => x"d5",
          2229 => x"05",
          2230 => x"84",
          2231 => x"08",
          2232 => x"0b",
          2233 => x"08",
          2234 => x"82",
          2235 => x"f4",
          2236 => x"d5",
          2237 => x"05",
          2238 => x"84",
          2239 => x"08",
          2240 => x"38",
          2241 => x"08",
          2242 => x"30",
          2243 => x"08",
          2244 => x"80",
          2245 => x"84",
          2246 => x"0c",
          2247 => x"08",
          2248 => x"8a",
          2249 => x"82",
          2250 => x"f0",
          2251 => x"d5",
          2252 => x"05",
          2253 => x"84",
          2254 => x"0c",
          2255 => x"d5",
          2256 => x"05",
          2257 => x"d5",
          2258 => x"05",
          2259 => x"c5",
          2260 => x"f8",
          2261 => x"d5",
          2262 => x"05",
          2263 => x"d5",
          2264 => x"05",
          2265 => x"90",
          2266 => x"84",
          2267 => x"08",
          2268 => x"84",
          2269 => x"0c",
          2270 => x"08",
          2271 => x"70",
          2272 => x"0c",
          2273 => x"0d",
          2274 => x"0c",
          2275 => x"84",
          2276 => x"d5",
          2277 => x"3d",
          2278 => x"82",
          2279 => x"fc",
          2280 => x"d5",
          2281 => x"05",
          2282 => x"99",
          2283 => x"84",
          2284 => x"08",
          2285 => x"84",
          2286 => x"0c",
          2287 => x"d5",
          2288 => x"05",
          2289 => x"84",
          2290 => x"08",
          2291 => x"38",
          2292 => x"08",
          2293 => x"30",
          2294 => x"08",
          2295 => x"81",
          2296 => x"84",
          2297 => x"08",
          2298 => x"84",
          2299 => x"08",
          2300 => x"3f",
          2301 => x"08",
          2302 => x"84",
          2303 => x"0c",
          2304 => x"84",
          2305 => x"08",
          2306 => x"38",
          2307 => x"08",
          2308 => x"30",
          2309 => x"08",
          2310 => x"82",
          2311 => x"f8",
          2312 => x"82",
          2313 => x"54",
          2314 => x"82",
          2315 => x"04",
          2316 => x"08",
          2317 => x"84",
          2318 => x"0d",
          2319 => x"d5",
          2320 => x"05",
          2321 => x"d5",
          2322 => x"05",
          2323 => x"c5",
          2324 => x"f8",
          2325 => x"d4",
          2326 => x"85",
          2327 => x"d5",
          2328 => x"82",
          2329 => x"02",
          2330 => x"0c",
          2331 => x"81",
          2332 => x"84",
          2333 => x"08",
          2334 => x"84",
          2335 => x"08",
          2336 => x"82",
          2337 => x"70",
          2338 => x"0c",
          2339 => x"0d",
          2340 => x"0c",
          2341 => x"84",
          2342 => x"d5",
          2343 => x"3d",
          2344 => x"82",
          2345 => x"fc",
          2346 => x"0b",
          2347 => x"08",
          2348 => x"82",
          2349 => x"8c",
          2350 => x"d5",
          2351 => x"05",
          2352 => x"38",
          2353 => x"08",
          2354 => x"80",
          2355 => x"80",
          2356 => x"84",
          2357 => x"08",
          2358 => x"82",
          2359 => x"8c",
          2360 => x"82",
          2361 => x"8c",
          2362 => x"d5",
          2363 => x"05",
          2364 => x"d5",
          2365 => x"05",
          2366 => x"39",
          2367 => x"08",
          2368 => x"80",
          2369 => x"38",
          2370 => x"08",
          2371 => x"82",
          2372 => x"88",
          2373 => x"ad",
          2374 => x"84",
          2375 => x"08",
          2376 => x"08",
          2377 => x"31",
          2378 => x"08",
          2379 => x"82",
          2380 => x"f8",
          2381 => x"d5",
          2382 => x"05",
          2383 => x"d5",
          2384 => x"05",
          2385 => x"84",
          2386 => x"08",
          2387 => x"d5",
          2388 => x"05",
          2389 => x"84",
          2390 => x"08",
          2391 => x"d5",
          2392 => x"05",
          2393 => x"39",
          2394 => x"08",
          2395 => x"80",
          2396 => x"82",
          2397 => x"88",
          2398 => x"82",
          2399 => x"f4",
          2400 => x"91",
          2401 => x"84",
          2402 => x"08",
          2403 => x"84",
          2404 => x"0c",
          2405 => x"84",
          2406 => x"08",
          2407 => x"0c",
          2408 => x"82",
          2409 => x"04",
          2410 => x"08",
          2411 => x"84",
          2412 => x"0d",
          2413 => x"d5",
          2414 => x"05",
          2415 => x"84",
          2416 => x"08",
          2417 => x"0c",
          2418 => x"08",
          2419 => x"70",
          2420 => x"72",
          2421 => x"82",
          2422 => x"f8",
          2423 => x"81",
          2424 => x"72",
          2425 => x"81",
          2426 => x"82",
          2427 => x"88",
          2428 => x"08",
          2429 => x"0c",
          2430 => x"82",
          2431 => x"f8",
          2432 => x"72",
          2433 => x"81",
          2434 => x"81",
          2435 => x"84",
          2436 => x"34",
          2437 => x"08",
          2438 => x"70",
          2439 => x"71",
          2440 => x"51",
          2441 => x"82",
          2442 => x"f8",
          2443 => x"d5",
          2444 => x"05",
          2445 => x"b0",
          2446 => x"06",
          2447 => x"82",
          2448 => x"88",
          2449 => x"08",
          2450 => x"0c",
          2451 => x"53",
          2452 => x"d5",
          2453 => x"05",
          2454 => x"84",
          2455 => x"33",
          2456 => x"08",
          2457 => x"82",
          2458 => x"e8",
          2459 => x"e2",
          2460 => x"82",
          2461 => x"e8",
          2462 => x"f8",
          2463 => x"80",
          2464 => x"0b",
          2465 => x"08",
          2466 => x"82",
          2467 => x"88",
          2468 => x"08",
          2469 => x"0c",
          2470 => x"53",
          2471 => x"d5",
          2472 => x"05",
          2473 => x"39",
          2474 => x"d5",
          2475 => x"05",
          2476 => x"84",
          2477 => x"08",
          2478 => x"05",
          2479 => x"08",
          2480 => x"33",
          2481 => x"08",
          2482 => x"80",
          2483 => x"d5",
          2484 => x"05",
          2485 => x"a0",
          2486 => x"81",
          2487 => x"84",
          2488 => x"0c",
          2489 => x"82",
          2490 => x"f8",
          2491 => x"af",
          2492 => x"38",
          2493 => x"08",
          2494 => x"53",
          2495 => x"83",
          2496 => x"80",
          2497 => x"84",
          2498 => x"0c",
          2499 => x"88",
          2500 => x"84",
          2501 => x"34",
          2502 => x"d5",
          2503 => x"05",
          2504 => x"73",
          2505 => x"82",
          2506 => x"f8",
          2507 => x"72",
          2508 => x"38",
          2509 => x"0b",
          2510 => x"08",
          2511 => x"82",
          2512 => x"0b",
          2513 => x"08",
          2514 => x"80",
          2515 => x"84",
          2516 => x"0c",
          2517 => x"08",
          2518 => x"53",
          2519 => x"81",
          2520 => x"d5",
          2521 => x"05",
          2522 => x"e0",
          2523 => x"38",
          2524 => x"08",
          2525 => x"e0",
          2526 => x"72",
          2527 => x"08",
          2528 => x"82",
          2529 => x"f8",
          2530 => x"11",
          2531 => x"82",
          2532 => x"f8",
          2533 => x"d5",
          2534 => x"05",
          2535 => x"73",
          2536 => x"82",
          2537 => x"f8",
          2538 => x"11",
          2539 => x"82",
          2540 => x"f8",
          2541 => x"d5",
          2542 => x"05",
          2543 => x"89",
          2544 => x"80",
          2545 => x"84",
          2546 => x"0c",
          2547 => x"82",
          2548 => x"f8",
          2549 => x"d5",
          2550 => x"05",
          2551 => x"72",
          2552 => x"38",
          2553 => x"d5",
          2554 => x"05",
          2555 => x"39",
          2556 => x"08",
          2557 => x"70",
          2558 => x"08",
          2559 => x"29",
          2560 => x"08",
          2561 => x"70",
          2562 => x"84",
          2563 => x"0c",
          2564 => x"08",
          2565 => x"70",
          2566 => x"71",
          2567 => x"51",
          2568 => x"53",
          2569 => x"d5",
          2570 => x"05",
          2571 => x"39",
          2572 => x"08",
          2573 => x"53",
          2574 => x"90",
          2575 => x"84",
          2576 => x"08",
          2577 => x"84",
          2578 => x"0c",
          2579 => x"08",
          2580 => x"82",
          2581 => x"fc",
          2582 => x"0c",
          2583 => x"82",
          2584 => x"ec",
          2585 => x"d5",
          2586 => x"05",
          2587 => x"f8",
          2588 => x"0d",
          2589 => x"0c",
          2590 => x"84",
          2591 => x"d5",
          2592 => x"3d",
          2593 => x"82",
          2594 => x"f0",
          2595 => x"d5",
          2596 => x"05",
          2597 => x"73",
          2598 => x"84",
          2599 => x"08",
          2600 => x"53",
          2601 => x"72",
          2602 => x"08",
          2603 => x"72",
          2604 => x"53",
          2605 => x"09",
          2606 => x"38",
          2607 => x"08",
          2608 => x"70",
          2609 => x"71",
          2610 => x"39",
          2611 => x"08",
          2612 => x"53",
          2613 => x"09",
          2614 => x"38",
          2615 => x"d5",
          2616 => x"05",
          2617 => x"84",
          2618 => x"08",
          2619 => x"05",
          2620 => x"08",
          2621 => x"33",
          2622 => x"08",
          2623 => x"82",
          2624 => x"f8",
          2625 => x"72",
          2626 => x"81",
          2627 => x"38",
          2628 => x"08",
          2629 => x"70",
          2630 => x"71",
          2631 => x"51",
          2632 => x"82",
          2633 => x"f8",
          2634 => x"d5",
          2635 => x"05",
          2636 => x"84",
          2637 => x"0c",
          2638 => x"08",
          2639 => x"80",
          2640 => x"38",
          2641 => x"08",
          2642 => x"80",
          2643 => x"38",
          2644 => x"90",
          2645 => x"84",
          2646 => x"34",
          2647 => x"08",
          2648 => x"70",
          2649 => x"71",
          2650 => x"51",
          2651 => x"82",
          2652 => x"f8",
          2653 => x"a4",
          2654 => x"82",
          2655 => x"f4",
          2656 => x"d5",
          2657 => x"05",
          2658 => x"81",
          2659 => x"70",
          2660 => x"72",
          2661 => x"84",
          2662 => x"34",
          2663 => x"82",
          2664 => x"f8",
          2665 => x"72",
          2666 => x"38",
          2667 => x"d5",
          2668 => x"05",
          2669 => x"39",
          2670 => x"08",
          2671 => x"53",
          2672 => x"90",
          2673 => x"84",
          2674 => x"33",
          2675 => x"26",
          2676 => x"39",
          2677 => x"d5",
          2678 => x"05",
          2679 => x"39",
          2680 => x"d5",
          2681 => x"05",
          2682 => x"82",
          2683 => x"f8",
          2684 => x"af",
          2685 => x"38",
          2686 => x"08",
          2687 => x"53",
          2688 => x"83",
          2689 => x"80",
          2690 => x"84",
          2691 => x"0c",
          2692 => x"8a",
          2693 => x"84",
          2694 => x"34",
          2695 => x"d5",
          2696 => x"05",
          2697 => x"84",
          2698 => x"33",
          2699 => x"27",
          2700 => x"82",
          2701 => x"f8",
          2702 => x"80",
          2703 => x"94",
          2704 => x"84",
          2705 => x"33",
          2706 => x"53",
          2707 => x"84",
          2708 => x"34",
          2709 => x"08",
          2710 => x"d0",
          2711 => x"72",
          2712 => x"08",
          2713 => x"82",
          2714 => x"f8",
          2715 => x"90",
          2716 => x"38",
          2717 => x"08",
          2718 => x"f9",
          2719 => x"72",
          2720 => x"08",
          2721 => x"82",
          2722 => x"f8",
          2723 => x"72",
          2724 => x"38",
          2725 => x"d5",
          2726 => x"05",
          2727 => x"39",
          2728 => x"08",
          2729 => x"82",
          2730 => x"f4",
          2731 => x"54",
          2732 => x"8d",
          2733 => x"82",
          2734 => x"ec",
          2735 => x"f7",
          2736 => x"84",
          2737 => x"33",
          2738 => x"84",
          2739 => x"08",
          2740 => x"84",
          2741 => x"33",
          2742 => x"d5",
          2743 => x"05",
          2744 => x"84",
          2745 => x"08",
          2746 => x"05",
          2747 => x"08",
          2748 => x"55",
          2749 => x"82",
          2750 => x"f8",
          2751 => x"a5",
          2752 => x"84",
          2753 => x"33",
          2754 => x"2e",
          2755 => x"d5",
          2756 => x"05",
          2757 => x"d5",
          2758 => x"05",
          2759 => x"84",
          2760 => x"08",
          2761 => x"08",
          2762 => x"71",
          2763 => x"0b",
          2764 => x"08",
          2765 => x"82",
          2766 => x"ec",
          2767 => x"d4",
          2768 => x"3d",
          2769 => x"84",
          2770 => x"3d",
          2771 => x"08",
          2772 => x"59",
          2773 => x"80",
          2774 => x"39",
          2775 => x"0c",
          2776 => x"54",
          2777 => x"74",
          2778 => x"a0",
          2779 => x"06",
          2780 => x"15",
          2781 => x"80",
          2782 => x"29",
          2783 => x"05",
          2784 => x"56",
          2785 => x"82",
          2786 => x"82",
          2787 => x"54",
          2788 => x"08",
          2789 => x"fc",
          2790 => x"f8",
          2791 => x"84",
          2792 => x"73",
          2793 => x"b4",
          2794 => x"70",
          2795 => x"58",
          2796 => x"27",
          2797 => x"54",
          2798 => x"f8",
          2799 => x"0d",
          2800 => x"0d",
          2801 => x"93",
          2802 => x"38",
          2803 => x"82",
          2804 => x"52",
          2805 => x"82",
          2806 => x"81",
          2807 => x"b2",
          2808 => x"f9",
          2809 => x"a4",
          2810 => x"39",
          2811 => x"51",
          2812 => x"82",
          2813 => x"80",
          2814 => x"b2",
          2815 => x"dd",
          2816 => x"e8",
          2817 => x"39",
          2818 => x"51",
          2819 => x"82",
          2820 => x"80",
          2821 => x"b3",
          2822 => x"c1",
          2823 => x"c0",
          2824 => x"82",
          2825 => x"b5",
          2826 => x"f0",
          2827 => x"82",
          2828 => x"a9",
          2829 => x"a8",
          2830 => x"82",
          2831 => x"9d",
          2832 => x"d8",
          2833 => x"82",
          2834 => x"91",
          2835 => x"88",
          2836 => x"82",
          2837 => x"85",
          2838 => x"ac",
          2839 => x"3f",
          2840 => x"04",
          2841 => x"77",
          2842 => x"74",
          2843 => x"8a",
          2844 => x"75",
          2845 => x"51",
          2846 => x"e8",
          2847 => x"ef",
          2848 => x"d4",
          2849 => x"75",
          2850 => x"3f",
          2851 => x"08",
          2852 => x"75",
          2853 => x"bc",
          2854 => x"be",
          2855 => x"0d",
          2856 => x"0d",
          2857 => x"05",
          2858 => x"33",
          2859 => x"68",
          2860 => x"7a",
          2861 => x"51",
          2862 => x"78",
          2863 => x"ff",
          2864 => x"81",
          2865 => x"07",
          2866 => x"06",
          2867 => x"56",
          2868 => x"38",
          2869 => x"52",
          2870 => x"52",
          2871 => x"8d",
          2872 => x"f8",
          2873 => x"d4",
          2874 => x"38",
          2875 => x"08",
          2876 => x"88",
          2877 => x"f8",
          2878 => x"3d",
          2879 => x"84",
          2880 => x"52",
          2881 => x"96",
          2882 => x"d4",
          2883 => x"82",
          2884 => x"90",
          2885 => x"74",
          2886 => x"38",
          2887 => x"19",
          2888 => x"39",
          2889 => x"05",
          2890 => x"c0",
          2891 => x"70",
          2892 => x"25",
          2893 => x"9f",
          2894 => x"51",
          2895 => x"74",
          2896 => x"38",
          2897 => x"53",
          2898 => x"88",
          2899 => x"51",
          2900 => x"76",
          2901 => x"d4",
          2902 => x"3d",
          2903 => x"3d",
          2904 => x"84",
          2905 => x"33",
          2906 => x"59",
          2907 => x"52",
          2908 => x"ad",
          2909 => x"f8",
          2910 => x"38",
          2911 => x"88",
          2912 => x"2e",
          2913 => x"39",
          2914 => x"57",
          2915 => x"56",
          2916 => x"55",
          2917 => x"08",
          2918 => x"dc",
          2919 => x"f0",
          2920 => x"82",
          2921 => x"ff",
          2922 => x"82",
          2923 => x"62",
          2924 => x"82",
          2925 => x"60",
          2926 => x"79",
          2927 => x"f8",
          2928 => x"39",
          2929 => x"82",
          2930 => x"8b",
          2931 => x"f3",
          2932 => x"61",
          2933 => x"05",
          2934 => x"33",
          2935 => x"68",
          2936 => x"5c",
          2937 => x"7a",
          2938 => x"9c",
          2939 => x"ea",
          2940 => x"a4",
          2941 => x"e2",
          2942 => x"74",
          2943 => x"80",
          2944 => x"2e",
          2945 => x"a0",
          2946 => x"80",
          2947 => x"18",
          2948 => x"27",
          2949 => x"22",
          2950 => x"a8",
          2951 => x"ba",
          2952 => x"82",
          2953 => x"ff",
          2954 => x"82",
          2955 => x"c3",
          2956 => x"53",
          2957 => x"8e",
          2958 => x"52",
          2959 => x"51",
          2960 => x"3f",
          2961 => x"b6",
          2962 => x"b7",
          2963 => x"15",
          2964 => x"74",
          2965 => x"7a",
          2966 => x"72",
          2967 => x"b6",
          2968 => x"b6",
          2969 => x"39",
          2970 => x"51",
          2971 => x"3f",
          2972 => x"82",
          2973 => x"52",
          2974 => x"b8",
          2975 => x"39",
          2976 => x"51",
          2977 => x"3f",
          2978 => x"79",
          2979 => x"38",
          2980 => x"33",
          2981 => x"56",
          2982 => x"83",
          2983 => x"80",
          2984 => x"27",
          2985 => x"53",
          2986 => x"70",
          2987 => x"51",
          2988 => x"2e",
          2989 => x"80",
          2990 => x"38",
          2991 => x"08",
          2992 => x"88",
          2993 => x"dc",
          2994 => x"51",
          2995 => x"81",
          2996 => x"b6",
          2997 => x"cc",
          2998 => x"3f",
          2999 => x"1c",
          3000 => x"bd",
          3001 => x"f8",
          3002 => x"70",
          3003 => x"57",
          3004 => x"09",
          3005 => x"38",
          3006 => x"82",
          3007 => x"98",
          3008 => x"2c",
          3009 => x"70",
          3010 => x"32",
          3011 => x"72",
          3012 => x"07",
          3013 => x"58",
          3014 => x"57",
          3015 => x"d8",
          3016 => x"2e",
          3017 => x"85",
          3018 => x"8c",
          3019 => x"53",
          3020 => x"fd",
          3021 => x"53",
          3022 => x"f8",
          3023 => x"0d",
          3024 => x"0d",
          3025 => x"33",
          3026 => x"53",
          3027 => x"52",
          3028 => x"86",
          3029 => x"d0",
          3030 => x"96",
          3031 => x"e0",
          3032 => x"ec",
          3033 => x"d1",
          3034 => x"b6",
          3035 => x"b4",
          3036 => x"80",
          3037 => x"a1",
          3038 => x"3d",
          3039 => x"3d",
          3040 => x"96",
          3041 => x"a6",
          3042 => x"51",
          3043 => x"82",
          3044 => x"9a",
          3045 => x"51",
          3046 => x"72",
          3047 => x"81",
          3048 => x"71",
          3049 => x"38",
          3050 => x"e2",
          3051 => x"a8",
          3052 => x"3f",
          3053 => x"d6",
          3054 => x"2a",
          3055 => x"51",
          3056 => x"2e",
          3057 => x"51",
          3058 => x"82",
          3059 => x"99",
          3060 => x"51",
          3061 => x"72",
          3062 => x"81",
          3063 => x"71",
          3064 => x"38",
          3065 => x"a6",
          3066 => x"c8",
          3067 => x"3f",
          3068 => x"9a",
          3069 => x"2a",
          3070 => x"51",
          3071 => x"2e",
          3072 => x"51",
          3073 => x"82",
          3074 => x"99",
          3075 => x"51",
          3076 => x"72",
          3077 => x"81",
          3078 => x"71",
          3079 => x"38",
          3080 => x"ea",
          3081 => x"f0",
          3082 => x"3f",
          3083 => x"de",
          3084 => x"2a",
          3085 => x"51",
          3086 => x"2e",
          3087 => x"51",
          3088 => x"82",
          3089 => x"98",
          3090 => x"51",
          3091 => x"72",
          3092 => x"81",
          3093 => x"71",
          3094 => x"38",
          3095 => x"ae",
          3096 => x"98",
          3097 => x"3f",
          3098 => x"a2",
          3099 => x"2a",
          3100 => x"51",
          3101 => x"2e",
          3102 => x"51",
          3103 => x"82",
          3104 => x"98",
          3105 => x"51",
          3106 => x"a4",
          3107 => x"3d",
          3108 => x"3d",
          3109 => x"84",
          3110 => x"33",
          3111 => x"56",
          3112 => x"51",
          3113 => x"0b",
          3114 => x"f4",
          3115 => x"a9",
          3116 => x"82",
          3117 => x"82",
          3118 => x"81",
          3119 => x"82",
          3120 => x"30",
          3121 => x"f8",
          3122 => x"25",
          3123 => x"51",
          3124 => x"0b",
          3125 => x"f4",
          3126 => x"82",
          3127 => x"54",
          3128 => x"09",
          3129 => x"38",
          3130 => x"53",
          3131 => x"51",
          3132 => x"3f",
          3133 => x"08",
          3134 => x"38",
          3135 => x"08",
          3136 => x"3f",
          3137 => x"ec",
          3138 => x"96",
          3139 => x"0b",
          3140 => x"cf",
          3141 => x"0b",
          3142 => x"33",
          3143 => x"2e",
          3144 => x"8c",
          3145 => x"f8",
          3146 => x"75",
          3147 => x"3f",
          3148 => x"d4",
          3149 => x"3d",
          3150 => x"3d",
          3151 => x"41",
          3152 => x"82",
          3153 => x"5f",
          3154 => x"51",
          3155 => x"3f",
          3156 => x"08",
          3157 => x"59",
          3158 => x"09",
          3159 => x"38",
          3160 => x"83",
          3161 => x"80",
          3162 => x"da",
          3163 => x"53",
          3164 => x"d6",
          3165 => x"88",
          3166 => x"d4",
          3167 => x"2e",
          3168 => x"b9",
          3169 => x"df",
          3170 => x"41",
          3171 => x"bc",
          3172 => x"c6",
          3173 => x"70",
          3174 => x"f8",
          3175 => x"fd",
          3176 => x"3d",
          3177 => x"51",
          3178 => x"82",
          3179 => x"90",
          3180 => x"2c",
          3181 => x"80",
          3182 => x"a3",
          3183 => x"c2",
          3184 => x"78",
          3185 => x"d2",
          3186 => x"24",
          3187 => x"80",
          3188 => x"38",
          3189 => x"80",
          3190 => x"d6",
          3191 => x"c0",
          3192 => x"38",
          3193 => x"24",
          3194 => x"78",
          3195 => x"8c",
          3196 => x"39",
          3197 => x"2e",
          3198 => x"78",
          3199 => x"92",
          3200 => x"c3",
          3201 => x"38",
          3202 => x"2e",
          3203 => x"8a",
          3204 => x"81",
          3205 => x"88",
          3206 => x"83",
          3207 => x"78",
          3208 => x"89",
          3209 => x"8a",
          3210 => x"85",
          3211 => x"38",
          3212 => x"b5",
          3213 => x"11",
          3214 => x"05",
          3215 => x"3f",
          3216 => x"08",
          3217 => x"c5",
          3218 => x"fe",
          3219 => x"ff",
          3220 => x"ec",
          3221 => x"d4",
          3222 => x"2e",
          3223 => x"b5",
          3224 => x"11",
          3225 => x"05",
          3226 => x"3f",
          3227 => x"08",
          3228 => x"d4",
          3229 => x"82",
          3230 => x"ff",
          3231 => x"64",
          3232 => x"79",
          3233 => x"ec",
          3234 => x"78",
          3235 => x"05",
          3236 => x"7a",
          3237 => x"81",
          3238 => x"3d",
          3239 => x"53",
          3240 => x"51",
          3241 => x"82",
          3242 => x"80",
          3243 => x"38",
          3244 => x"fc",
          3245 => x"84",
          3246 => x"bd",
          3247 => x"f8",
          3248 => x"fd",
          3249 => x"3d",
          3250 => x"53",
          3251 => x"51",
          3252 => x"82",
          3253 => x"80",
          3254 => x"38",
          3255 => x"51",
          3256 => x"3f",
          3257 => x"64",
          3258 => x"38",
          3259 => x"70",
          3260 => x"33",
          3261 => x"81",
          3262 => x"39",
          3263 => x"80",
          3264 => x"84",
          3265 => x"f1",
          3266 => x"f8",
          3267 => x"fc",
          3268 => x"3d",
          3269 => x"53",
          3270 => x"51",
          3271 => x"82",
          3272 => x"80",
          3273 => x"38",
          3274 => x"f8",
          3275 => x"84",
          3276 => x"c5",
          3277 => x"f8",
          3278 => x"fc",
          3279 => x"b9",
          3280 => x"ad",
          3281 => x"5a",
          3282 => x"a8",
          3283 => x"33",
          3284 => x"5a",
          3285 => x"2e",
          3286 => x"55",
          3287 => x"33",
          3288 => x"82",
          3289 => x"ff",
          3290 => x"81",
          3291 => x"05",
          3292 => x"39",
          3293 => x"8f",
          3294 => x"39",
          3295 => x"80",
          3296 => x"84",
          3297 => x"f1",
          3298 => x"f8",
          3299 => x"38",
          3300 => x"33",
          3301 => x"2e",
          3302 => x"d3",
          3303 => x"80",
          3304 => x"d3",
          3305 => x"78",
          3306 => x"38",
          3307 => x"08",
          3308 => x"82",
          3309 => x"59",
          3310 => x"88",
          3311 => x"ac",
          3312 => x"39",
          3313 => x"33",
          3314 => x"2e",
          3315 => x"d3",
          3316 => x"9a",
          3317 => x"e2",
          3318 => x"80",
          3319 => x"82",
          3320 => x"45",
          3321 => x"d3",
          3322 => x"80",
          3323 => x"3d",
          3324 => x"53",
          3325 => x"51",
          3326 => x"82",
          3327 => x"80",
          3328 => x"d3",
          3329 => x"78",
          3330 => x"38",
          3331 => x"08",
          3332 => x"39",
          3333 => x"33",
          3334 => x"2e",
          3335 => x"d3",
          3336 => x"bb",
          3337 => x"e6",
          3338 => x"80",
          3339 => x"82",
          3340 => x"44",
          3341 => x"d3",
          3342 => x"78",
          3343 => x"38",
          3344 => x"08",
          3345 => x"82",
          3346 => x"59",
          3347 => x"88",
          3348 => x"c0",
          3349 => x"39",
          3350 => x"08",
          3351 => x"b5",
          3352 => x"11",
          3353 => x"05",
          3354 => x"3f",
          3355 => x"08",
          3356 => x"38",
          3357 => x"5c",
          3358 => x"83",
          3359 => x"7a",
          3360 => x"30",
          3361 => x"9f",
          3362 => x"06",
          3363 => x"5a",
          3364 => x"88",
          3365 => x"2e",
          3366 => x"43",
          3367 => x"51",
          3368 => x"a0",
          3369 => x"62",
          3370 => x"64",
          3371 => x"3f",
          3372 => x"51",
          3373 => x"b5",
          3374 => x"11",
          3375 => x"05",
          3376 => x"3f",
          3377 => x"08",
          3378 => x"c1",
          3379 => x"fe",
          3380 => x"ff",
          3381 => x"e7",
          3382 => x"d4",
          3383 => x"2e",
          3384 => x"59",
          3385 => x"05",
          3386 => x"64",
          3387 => x"b5",
          3388 => x"11",
          3389 => x"05",
          3390 => x"3f",
          3391 => x"08",
          3392 => x"89",
          3393 => x"33",
          3394 => x"ba",
          3395 => x"a9",
          3396 => x"f0",
          3397 => x"80",
          3398 => x"51",
          3399 => x"3f",
          3400 => x"33",
          3401 => x"2e",
          3402 => x"9f",
          3403 => x"38",
          3404 => x"fc",
          3405 => x"84",
          3406 => x"bd",
          3407 => x"f8",
          3408 => x"91",
          3409 => x"02",
          3410 => x"33",
          3411 => x"81",
          3412 => x"b1",
          3413 => x"ac",
          3414 => x"3f",
          3415 => x"b5",
          3416 => x"11",
          3417 => x"05",
          3418 => x"3f",
          3419 => x"08",
          3420 => x"99",
          3421 => x"fe",
          3422 => x"ff",
          3423 => x"e0",
          3424 => x"d4",
          3425 => x"2e",
          3426 => x"59",
          3427 => x"05",
          3428 => x"82",
          3429 => x"78",
          3430 => x"fe",
          3431 => x"ff",
          3432 => x"e0",
          3433 => x"d4",
          3434 => x"38",
          3435 => x"61",
          3436 => x"52",
          3437 => x"51",
          3438 => x"3f",
          3439 => x"08",
          3440 => x"52",
          3441 => x"a8",
          3442 => x"46",
          3443 => x"78",
          3444 => x"b9",
          3445 => x"26",
          3446 => x"82",
          3447 => x"39",
          3448 => x"f0",
          3449 => x"84",
          3450 => x"bc",
          3451 => x"f8",
          3452 => x"93",
          3453 => x"02",
          3454 => x"22",
          3455 => x"05",
          3456 => x"42",
          3457 => x"82",
          3458 => x"c3",
          3459 => x"9f",
          3460 => x"fe",
          3461 => x"ff",
          3462 => x"df",
          3463 => x"d4",
          3464 => x"2e",
          3465 => x"b5",
          3466 => x"11",
          3467 => x"05",
          3468 => x"3f",
          3469 => x"08",
          3470 => x"38",
          3471 => x"0c",
          3472 => x"05",
          3473 => x"fe",
          3474 => x"ff",
          3475 => x"de",
          3476 => x"d4",
          3477 => x"38",
          3478 => x"61",
          3479 => x"52",
          3480 => x"51",
          3481 => x"3f",
          3482 => x"08",
          3483 => x"52",
          3484 => x"a7",
          3485 => x"46",
          3486 => x"78",
          3487 => x"8d",
          3488 => x"27",
          3489 => x"3d",
          3490 => x"53",
          3491 => x"51",
          3492 => x"82",
          3493 => x"80",
          3494 => x"61",
          3495 => x"59",
          3496 => x"42",
          3497 => x"82",
          3498 => x"c2",
          3499 => x"ab",
          3500 => x"ff",
          3501 => x"ff",
          3502 => x"e3",
          3503 => x"d4",
          3504 => x"2e",
          3505 => x"64",
          3506 => x"cc",
          3507 => x"8a",
          3508 => x"78",
          3509 => x"ff",
          3510 => x"ff",
          3511 => x"e3",
          3512 => x"d4",
          3513 => x"2e",
          3514 => x"64",
          3515 => x"e8",
          3516 => x"e6",
          3517 => x"78",
          3518 => x"f8",
          3519 => x"f5",
          3520 => x"d4",
          3521 => x"82",
          3522 => x"ff",
          3523 => x"f4",
          3524 => x"bb",
          3525 => x"cd",
          3526 => x"9f",
          3527 => x"39",
          3528 => x"51",
          3529 => x"80",
          3530 => x"39",
          3531 => x"f4",
          3532 => x"3d",
          3533 => x"80",
          3534 => x"38",
          3535 => x"79",
          3536 => x"3f",
          3537 => x"08",
          3538 => x"f8",
          3539 => x"82",
          3540 => x"d4",
          3541 => x"b5",
          3542 => x"05",
          3543 => x"3f",
          3544 => x"08",
          3545 => x"5a",
          3546 => x"2e",
          3547 => x"82",
          3548 => x"51",
          3549 => x"82",
          3550 => x"8f",
          3551 => x"38",
          3552 => x"82",
          3553 => x"7a",
          3554 => x"38",
          3555 => x"8c",
          3556 => x"39",
          3557 => x"ad",
          3558 => x"39",
          3559 => x"56",
          3560 => x"bb",
          3561 => x"53",
          3562 => x"52",
          3563 => x"b0",
          3564 => x"a7",
          3565 => x"39",
          3566 => x"3d",
          3567 => x"51",
          3568 => x"ab",
          3569 => x"82",
          3570 => x"80",
          3571 => x"e8",
          3572 => x"ff",
          3573 => x"ff",
          3574 => x"93",
          3575 => x"80",
          3576 => x"f4",
          3577 => x"ff",
          3578 => x"ff",
          3579 => x"82",
          3580 => x"82",
          3581 => x"7c",
          3582 => x"80",
          3583 => x"80",
          3584 => x"80",
          3585 => x"ff",
          3586 => x"ea",
          3587 => x"d4",
          3588 => x"d4",
          3589 => x"70",
          3590 => x"07",
          3591 => x"5b",
          3592 => x"5a",
          3593 => x"83",
          3594 => x"78",
          3595 => x"78",
          3596 => x"38",
          3597 => x"81",
          3598 => x"59",
          3599 => x"38",
          3600 => x"7e",
          3601 => x"59",
          3602 => x"7e",
          3603 => x"81",
          3604 => x"82",
          3605 => x"ff",
          3606 => x"7c",
          3607 => x"3f",
          3608 => x"82",
          3609 => x"ff",
          3610 => x"f2",
          3611 => x"3d",
          3612 => x"82",
          3613 => x"87",
          3614 => x"08",
          3615 => x"80",
          3616 => x"d7",
          3617 => x"d4",
          3618 => x"2b",
          3619 => x"8c",
          3620 => x"87",
          3621 => x"73",
          3622 => x"3f",
          3623 => x"f8",
          3624 => x"c0",
          3625 => x"87",
          3626 => x"08",
          3627 => x"80",
          3628 => x"d6",
          3629 => x"d4",
          3630 => x"2b",
          3631 => x"9c",
          3632 => x"87",
          3633 => x"73",
          3634 => x"3f",
          3635 => x"f8",
          3636 => x"c0",
          3637 => x"8c",
          3638 => x"87",
          3639 => x"0c",
          3640 => x"0b",
          3641 => x"94",
          3642 => x"0a",
          3643 => x"86",
          3644 => x"84",
          3645 => x"87",
          3646 => x"73",
          3647 => x"8e",
          3648 => x"fa",
          3649 => x"f6",
          3650 => x"05",
          3651 => x"9f",
          3652 => x"27",
          3653 => x"f8",
          3654 => x"fb",
          3655 => x"02",
          3656 => x"05",
          3657 => x"85",
          3658 => x"f0",
          3659 => x"82",
          3660 => x"82",
          3661 => x"89",
          3662 => x"ff",
          3663 => x"b8",
          3664 => x"a1",
          3665 => x"c4",
          3666 => x"99",
          3667 => x"fc",
          3668 => x"3f",
          3669 => x"e9",
          3670 => x"3f",
          3671 => x"3d",
          3672 => x"83",
          3673 => x"2b",
          3674 => x"3f",
          3675 => x"08",
          3676 => x"72",
          3677 => x"54",
          3678 => x"25",
          3679 => x"82",
          3680 => x"84",
          3681 => x"fc",
          3682 => x"70",
          3683 => x"80",
          3684 => x"72",
          3685 => x"8a",
          3686 => x"51",
          3687 => x"09",
          3688 => x"38",
          3689 => x"f1",
          3690 => x"51",
          3691 => x"09",
          3692 => x"38",
          3693 => x"81",
          3694 => x"73",
          3695 => x"81",
          3696 => x"84",
          3697 => x"52",
          3698 => x"52",
          3699 => x"2e",
          3700 => x"54",
          3701 => x"9d",
          3702 => x"38",
          3703 => x"12",
          3704 => x"33",
          3705 => x"a0",
          3706 => x"81",
          3707 => x"2e",
          3708 => x"ea",
          3709 => x"33",
          3710 => x"a0",
          3711 => x"06",
          3712 => x"54",
          3713 => x"70",
          3714 => x"25",
          3715 => x"51",
          3716 => x"2e",
          3717 => x"72",
          3718 => x"54",
          3719 => x"0c",
          3720 => x"82",
          3721 => x"86",
          3722 => x"fc",
          3723 => x"53",
          3724 => x"2e",
          3725 => x"3d",
          3726 => x"72",
          3727 => x"3f",
          3728 => x"08",
          3729 => x"53",
          3730 => x"53",
          3731 => x"f8",
          3732 => x"0d",
          3733 => x"0d",
          3734 => x"33",
          3735 => x"53",
          3736 => x"8b",
          3737 => x"38",
          3738 => x"ff",
          3739 => x"52",
          3740 => x"81",
          3741 => x"13",
          3742 => x"52",
          3743 => x"80",
          3744 => x"13",
          3745 => x"52",
          3746 => x"80",
          3747 => x"13",
          3748 => x"52",
          3749 => x"80",
          3750 => x"13",
          3751 => x"52",
          3752 => x"26",
          3753 => x"8a",
          3754 => x"87",
          3755 => x"e7",
          3756 => x"38",
          3757 => x"c0",
          3758 => x"72",
          3759 => x"98",
          3760 => x"13",
          3761 => x"98",
          3762 => x"13",
          3763 => x"98",
          3764 => x"13",
          3765 => x"98",
          3766 => x"13",
          3767 => x"98",
          3768 => x"13",
          3769 => x"98",
          3770 => x"87",
          3771 => x"0c",
          3772 => x"98",
          3773 => x"0b",
          3774 => x"9c",
          3775 => x"71",
          3776 => x"0c",
          3777 => x"04",
          3778 => x"7f",
          3779 => x"98",
          3780 => x"7d",
          3781 => x"98",
          3782 => x"7d",
          3783 => x"c0",
          3784 => x"5a",
          3785 => x"34",
          3786 => x"b4",
          3787 => x"83",
          3788 => x"c0",
          3789 => x"5a",
          3790 => x"34",
          3791 => x"ac",
          3792 => x"85",
          3793 => x"c0",
          3794 => x"5a",
          3795 => x"34",
          3796 => x"a4",
          3797 => x"88",
          3798 => x"c0",
          3799 => x"5a",
          3800 => x"23",
          3801 => x"79",
          3802 => x"06",
          3803 => x"ff",
          3804 => x"86",
          3805 => x"85",
          3806 => x"84",
          3807 => x"83",
          3808 => x"82",
          3809 => x"7d",
          3810 => x"06",
          3811 => x"dc",
          3812 => x"c6",
          3813 => x"0d",
          3814 => x"0d",
          3815 => x"33",
          3816 => x"33",
          3817 => x"06",
          3818 => x"87",
          3819 => x"51",
          3820 => x"86",
          3821 => x"94",
          3822 => x"08",
          3823 => x"70",
          3824 => x"54",
          3825 => x"2e",
          3826 => x"91",
          3827 => x"06",
          3828 => x"d7",
          3829 => x"32",
          3830 => x"51",
          3831 => x"2e",
          3832 => x"93",
          3833 => x"06",
          3834 => x"ff",
          3835 => x"81",
          3836 => x"87",
          3837 => x"52",
          3838 => x"86",
          3839 => x"94",
          3840 => x"72",
          3841 => x"d4",
          3842 => x"3d",
          3843 => x"3d",
          3844 => x"05",
          3845 => x"70",
          3846 => x"52",
          3847 => x"d3",
          3848 => x"3d",
          3849 => x"3d",
          3850 => x"05",
          3851 => x"8a",
          3852 => x"06",
          3853 => x"52",
          3854 => x"3f",
          3855 => x"33",
          3856 => x"06",
          3857 => x"c0",
          3858 => x"76",
          3859 => x"38",
          3860 => x"94",
          3861 => x"70",
          3862 => x"81",
          3863 => x"54",
          3864 => x"8c",
          3865 => x"2a",
          3866 => x"51",
          3867 => x"38",
          3868 => x"70",
          3869 => x"53",
          3870 => x"8d",
          3871 => x"2a",
          3872 => x"51",
          3873 => x"be",
          3874 => x"ff",
          3875 => x"c0",
          3876 => x"72",
          3877 => x"38",
          3878 => x"90",
          3879 => x"0c",
          3880 => x"d4",
          3881 => x"3d",
          3882 => x"3d",
          3883 => x"80",
          3884 => x"81",
          3885 => x"53",
          3886 => x"2e",
          3887 => x"71",
          3888 => x"81",
          3889 => x"98",
          3890 => x"ff",
          3891 => x"55",
          3892 => x"94",
          3893 => x"80",
          3894 => x"87",
          3895 => x"51",
          3896 => x"96",
          3897 => x"06",
          3898 => x"70",
          3899 => x"38",
          3900 => x"70",
          3901 => x"51",
          3902 => x"72",
          3903 => x"81",
          3904 => x"70",
          3905 => x"38",
          3906 => x"70",
          3907 => x"51",
          3908 => x"38",
          3909 => x"06",
          3910 => x"94",
          3911 => x"80",
          3912 => x"87",
          3913 => x"52",
          3914 => x"81",
          3915 => x"70",
          3916 => x"53",
          3917 => x"ff",
          3918 => x"82",
          3919 => x"89",
          3920 => x"fe",
          3921 => x"d3",
          3922 => x"81",
          3923 => x"52",
          3924 => x"84",
          3925 => x"2e",
          3926 => x"c0",
          3927 => x"70",
          3928 => x"2a",
          3929 => x"51",
          3930 => x"80",
          3931 => x"71",
          3932 => x"51",
          3933 => x"80",
          3934 => x"2e",
          3935 => x"c0",
          3936 => x"71",
          3937 => x"ff",
          3938 => x"f8",
          3939 => x"3d",
          3940 => x"af",
          3941 => x"f8",
          3942 => x"06",
          3943 => x"0c",
          3944 => x"0d",
          3945 => x"33",
          3946 => x"06",
          3947 => x"c0",
          3948 => x"70",
          3949 => x"38",
          3950 => x"94",
          3951 => x"70",
          3952 => x"81",
          3953 => x"51",
          3954 => x"80",
          3955 => x"72",
          3956 => x"51",
          3957 => x"80",
          3958 => x"2e",
          3959 => x"c0",
          3960 => x"71",
          3961 => x"2b",
          3962 => x"51",
          3963 => x"82",
          3964 => x"84",
          3965 => x"ff",
          3966 => x"c0",
          3967 => x"70",
          3968 => x"06",
          3969 => x"80",
          3970 => x"38",
          3971 => x"a4",
          3972 => x"9c",
          3973 => x"9e",
          3974 => x"d3",
          3975 => x"c0",
          3976 => x"82",
          3977 => x"87",
          3978 => x"08",
          3979 => x"0c",
          3980 => x"9c",
          3981 => x"ac",
          3982 => x"9e",
          3983 => x"d3",
          3984 => x"c0",
          3985 => x"82",
          3986 => x"87",
          3987 => x"08",
          3988 => x"0c",
          3989 => x"b4",
          3990 => x"bc",
          3991 => x"9e",
          3992 => x"d3",
          3993 => x"c0",
          3994 => x"82",
          3995 => x"87",
          3996 => x"08",
          3997 => x"0c",
          3998 => x"c4",
          3999 => x"cc",
          4000 => x"9e",
          4001 => x"70",
          4002 => x"23",
          4003 => x"84",
          4004 => x"d4",
          4005 => x"9e",
          4006 => x"d3",
          4007 => x"c0",
          4008 => x"82",
          4009 => x"81",
          4010 => x"e0",
          4011 => x"87",
          4012 => x"08",
          4013 => x"0a",
          4014 => x"52",
          4015 => x"83",
          4016 => x"71",
          4017 => x"34",
          4018 => x"c0",
          4019 => x"70",
          4020 => x"06",
          4021 => x"70",
          4022 => x"38",
          4023 => x"82",
          4024 => x"80",
          4025 => x"9e",
          4026 => x"90",
          4027 => x"51",
          4028 => x"80",
          4029 => x"81",
          4030 => x"d3",
          4031 => x"0b",
          4032 => x"90",
          4033 => x"80",
          4034 => x"52",
          4035 => x"2e",
          4036 => x"52",
          4037 => x"e4",
          4038 => x"87",
          4039 => x"08",
          4040 => x"80",
          4041 => x"52",
          4042 => x"83",
          4043 => x"71",
          4044 => x"34",
          4045 => x"c0",
          4046 => x"70",
          4047 => x"06",
          4048 => x"70",
          4049 => x"38",
          4050 => x"82",
          4051 => x"80",
          4052 => x"9e",
          4053 => x"84",
          4054 => x"51",
          4055 => x"80",
          4056 => x"81",
          4057 => x"d3",
          4058 => x"0b",
          4059 => x"90",
          4060 => x"80",
          4061 => x"52",
          4062 => x"2e",
          4063 => x"52",
          4064 => x"e8",
          4065 => x"87",
          4066 => x"08",
          4067 => x"80",
          4068 => x"52",
          4069 => x"83",
          4070 => x"71",
          4071 => x"34",
          4072 => x"c0",
          4073 => x"70",
          4074 => x"06",
          4075 => x"70",
          4076 => x"38",
          4077 => x"82",
          4078 => x"80",
          4079 => x"9e",
          4080 => x"a0",
          4081 => x"52",
          4082 => x"2e",
          4083 => x"52",
          4084 => x"eb",
          4085 => x"9e",
          4086 => x"98",
          4087 => x"8a",
          4088 => x"51",
          4089 => x"ec",
          4090 => x"87",
          4091 => x"08",
          4092 => x"06",
          4093 => x"70",
          4094 => x"38",
          4095 => x"82",
          4096 => x"87",
          4097 => x"08",
          4098 => x"06",
          4099 => x"51",
          4100 => x"82",
          4101 => x"80",
          4102 => x"9e",
          4103 => x"88",
          4104 => x"52",
          4105 => x"83",
          4106 => x"71",
          4107 => x"34",
          4108 => x"90",
          4109 => x"06",
          4110 => x"82",
          4111 => x"83",
          4112 => x"fb",
          4113 => x"bc",
          4114 => x"93",
          4115 => x"d3",
          4116 => x"73",
          4117 => x"38",
          4118 => x"51",
          4119 => x"3f",
          4120 => x"51",
          4121 => x"3f",
          4122 => x"33",
          4123 => x"2e",
          4124 => x"d3",
          4125 => x"d3",
          4126 => x"54",
          4127 => x"b4",
          4128 => x"d6",
          4129 => x"e7",
          4130 => x"80",
          4131 => x"82",
          4132 => x"82",
          4133 => x"11",
          4134 => x"bd",
          4135 => x"92",
          4136 => x"d3",
          4137 => x"73",
          4138 => x"38",
          4139 => x"08",
          4140 => x"08",
          4141 => x"82",
          4142 => x"ff",
          4143 => x"82",
          4144 => x"54",
          4145 => x"94",
          4146 => x"a4",
          4147 => x"a8",
          4148 => x"52",
          4149 => x"51",
          4150 => x"3f",
          4151 => x"33",
          4152 => x"2e",
          4153 => x"d3",
          4154 => x"d3",
          4155 => x"54",
          4156 => x"a4",
          4157 => x"e2",
          4158 => x"eb",
          4159 => x"80",
          4160 => x"82",
          4161 => x"52",
          4162 => x"51",
          4163 => x"3f",
          4164 => x"33",
          4165 => x"2e",
          4166 => x"d3",
          4167 => x"82",
          4168 => x"ff",
          4169 => x"82",
          4170 => x"54",
          4171 => x"8e",
          4172 => x"ee",
          4173 => x"bf",
          4174 => x"91",
          4175 => x"d3",
          4176 => x"73",
          4177 => x"38",
          4178 => x"51",
          4179 => x"3f",
          4180 => x"33",
          4181 => x"2e",
          4182 => x"bf",
          4183 => x"ad",
          4184 => x"d3",
          4185 => x"73",
          4186 => x"38",
          4187 => x"51",
          4188 => x"3f",
          4189 => x"33",
          4190 => x"2e",
          4191 => x"bf",
          4192 => x"ac",
          4193 => x"d3",
          4194 => x"73",
          4195 => x"38",
          4196 => x"51",
          4197 => x"3f",
          4198 => x"51",
          4199 => x"3f",
          4200 => x"08",
          4201 => x"e8",
          4202 => x"ae",
          4203 => x"c8",
          4204 => x"c0",
          4205 => x"90",
          4206 => x"d3",
          4207 => x"82",
          4208 => x"ff",
          4209 => x"82",
          4210 => x"ff",
          4211 => x"82",
          4212 => x"52",
          4213 => x"51",
          4214 => x"3f",
          4215 => x"08",
          4216 => x"c0",
          4217 => x"c4",
          4218 => x"d4",
          4219 => x"84",
          4220 => x"71",
          4221 => x"82",
          4222 => x"52",
          4223 => x"51",
          4224 => x"3f",
          4225 => x"33",
          4226 => x"2e",
          4227 => x"d3",
          4228 => x"bd",
          4229 => x"75",
          4230 => x"3f",
          4231 => x"08",
          4232 => x"29",
          4233 => x"54",
          4234 => x"f8",
          4235 => x"c1",
          4236 => x"8f",
          4237 => x"d3",
          4238 => x"73",
          4239 => x"38",
          4240 => x"08",
          4241 => x"c0",
          4242 => x"c3",
          4243 => x"d4",
          4244 => x"84",
          4245 => x"71",
          4246 => x"82",
          4247 => x"52",
          4248 => x"51",
          4249 => x"3f",
          4250 => x"ae",
          4251 => x"3d",
          4252 => x"3d",
          4253 => x"05",
          4254 => x"52",
          4255 => x"aa",
          4256 => x"29",
          4257 => x"05",
          4258 => x"04",
          4259 => x"51",
          4260 => x"c2",
          4261 => x"39",
          4262 => x"51",
          4263 => x"c2",
          4264 => x"39",
          4265 => x"51",
          4266 => x"c2",
          4267 => x"8e",
          4268 => x"3d",
          4269 => x"88",
          4270 => x"80",
          4271 => x"96",
          4272 => x"82",
          4273 => x"87",
          4274 => x"0c",
          4275 => x"0d",
          4276 => x"70",
          4277 => x"98",
          4278 => x"2c",
          4279 => x"70",
          4280 => x"53",
          4281 => x"51",
          4282 => x"c2",
          4283 => x"55",
          4284 => x"25",
          4285 => x"c2",
          4286 => x"12",
          4287 => x"97",
          4288 => x"33",
          4289 => x"70",
          4290 => x"81",
          4291 => x"81",
          4292 => x"d4",
          4293 => x"3d",
          4294 => x"3d",
          4295 => x"84",
          4296 => x"33",
          4297 => x"56",
          4298 => x"2e",
          4299 => x"f0",
          4300 => x"88",
          4301 => x"fc",
          4302 => x"dc",
          4303 => x"51",
          4304 => x"3f",
          4305 => x"08",
          4306 => x"ff",
          4307 => x"73",
          4308 => x"53",
          4309 => x"72",
          4310 => x"53",
          4311 => x"51",
          4312 => x"3f",
          4313 => x"87",
          4314 => x"f6",
          4315 => x"02",
          4316 => x"05",
          4317 => x"05",
          4318 => x"82",
          4319 => x"70",
          4320 => x"d3",
          4321 => x"08",
          4322 => x"5a",
          4323 => x"80",
          4324 => x"74",
          4325 => x"3f",
          4326 => x"33",
          4327 => x"82",
          4328 => x"81",
          4329 => x"58",
          4330 => x"fc",
          4331 => x"f8",
          4332 => x"82",
          4333 => x"70",
          4334 => x"d3",
          4335 => x"08",
          4336 => x"74",
          4337 => x"38",
          4338 => x"52",
          4339 => x"b6",
          4340 => x"d4",
          4341 => x"05",
          4342 => x"d4",
          4343 => x"81",
          4344 => x"93",
          4345 => x"38",
          4346 => x"d4",
          4347 => x"80",
          4348 => x"82",
          4349 => x"56",
          4350 => x"ac",
          4351 => x"c8",
          4352 => x"a4",
          4353 => x"fc",
          4354 => x"53",
          4355 => x"51",
          4356 => x"3f",
          4357 => x"08",
          4358 => x"81",
          4359 => x"82",
          4360 => x"51",
          4361 => x"3f",
          4362 => x"04",
          4363 => x"82",
          4364 => x"93",
          4365 => x"52",
          4366 => x"89",
          4367 => x"99",
          4368 => x"73",
          4369 => x"84",
          4370 => x"73",
          4371 => x"38",
          4372 => x"d4",
          4373 => x"d4",
          4374 => x"71",
          4375 => x"38",
          4376 => x"f0",
          4377 => x"d4",
          4378 => x"99",
          4379 => x"0b",
          4380 => x"0c",
          4381 => x"04",
          4382 => x"81",
          4383 => x"82",
          4384 => x"51",
          4385 => x"3f",
          4386 => x"08",
          4387 => x"82",
          4388 => x"53",
          4389 => x"88",
          4390 => x"56",
          4391 => x"3f",
          4392 => x"08",
          4393 => x"38",
          4394 => x"b2",
          4395 => x"d4",
          4396 => x"80",
          4397 => x"f8",
          4398 => x"38",
          4399 => x"08",
          4400 => x"17",
          4401 => x"74",
          4402 => x"76",
          4403 => x"82",
          4404 => x"57",
          4405 => x"3f",
          4406 => x"09",
          4407 => x"af",
          4408 => x"0d",
          4409 => x"0d",
          4410 => x"ad",
          4411 => x"5a",
          4412 => x"58",
          4413 => x"d4",
          4414 => x"80",
          4415 => x"82",
          4416 => x"81",
          4417 => x"0b",
          4418 => x"08",
          4419 => x"f8",
          4420 => x"70",
          4421 => x"9c",
          4422 => x"d4",
          4423 => x"2e",
          4424 => x"51",
          4425 => x"3f",
          4426 => x"08",
          4427 => x"55",
          4428 => x"d4",
          4429 => x"8e",
          4430 => x"f8",
          4431 => x"70",
          4432 => x"80",
          4433 => x"09",
          4434 => x"72",
          4435 => x"51",
          4436 => x"77",
          4437 => x"73",
          4438 => x"82",
          4439 => x"8c",
          4440 => x"51",
          4441 => x"3f",
          4442 => x"08",
          4443 => x"38",
          4444 => x"51",
          4445 => x"3f",
          4446 => x"09",
          4447 => x"38",
          4448 => x"51",
          4449 => x"3f",
          4450 => x"b0",
          4451 => x"3d",
          4452 => x"d4",
          4453 => x"34",
          4454 => x"82",
          4455 => x"a9",
          4456 => x"f6",
          4457 => x"7e",
          4458 => x"72",
          4459 => x"5a",
          4460 => x"2e",
          4461 => x"a2",
          4462 => x"78",
          4463 => x"76",
          4464 => x"81",
          4465 => x"70",
          4466 => x"58",
          4467 => x"2e",
          4468 => x"86",
          4469 => x"26",
          4470 => x"54",
          4471 => x"82",
          4472 => x"70",
          4473 => x"ff",
          4474 => x"82",
          4475 => x"53",
          4476 => x"08",
          4477 => x"9c",
          4478 => x"f8",
          4479 => x"38",
          4480 => x"55",
          4481 => x"88",
          4482 => x"2e",
          4483 => x"39",
          4484 => x"ac",
          4485 => x"5a",
          4486 => x"11",
          4487 => x"51",
          4488 => x"82",
          4489 => x"80",
          4490 => x"ff",
          4491 => x"52",
          4492 => x"b1",
          4493 => x"f8",
          4494 => x"06",
          4495 => x"38",
          4496 => x"39",
          4497 => x"81",
          4498 => x"54",
          4499 => x"ff",
          4500 => x"54",
          4501 => x"f8",
          4502 => x"0d",
          4503 => x"0d",
          4504 => x"b2",
          4505 => x"3d",
          4506 => x"5a",
          4507 => x"3d",
          4508 => x"d0",
          4509 => x"cc",
          4510 => x"73",
          4511 => x"73",
          4512 => x"33",
          4513 => x"83",
          4514 => x"76",
          4515 => x"bc",
          4516 => x"76",
          4517 => x"73",
          4518 => x"ad",
          4519 => x"98",
          4520 => x"d4",
          4521 => x"d4",
          4522 => x"d4",
          4523 => x"2e",
          4524 => x"93",
          4525 => x"82",
          4526 => x"51",
          4527 => x"3f",
          4528 => x"08",
          4529 => x"38",
          4530 => x"51",
          4531 => x"3f",
          4532 => x"82",
          4533 => x"5b",
          4534 => x"08",
          4535 => x"52",
          4536 => x"52",
          4537 => x"8a",
          4538 => x"f8",
          4539 => x"d4",
          4540 => x"2e",
          4541 => x"80",
          4542 => x"d4",
          4543 => x"ff",
          4544 => x"82",
          4545 => x"55",
          4546 => x"d4",
          4547 => x"a9",
          4548 => x"f8",
          4549 => x"70",
          4550 => x"80",
          4551 => x"53",
          4552 => x"06",
          4553 => x"f8",
          4554 => x"1b",
          4555 => x"06",
          4556 => x"7b",
          4557 => x"80",
          4558 => x"2e",
          4559 => x"ff",
          4560 => x"39",
          4561 => x"c8",
          4562 => x"38",
          4563 => x"08",
          4564 => x"38",
          4565 => x"8f",
          4566 => x"c5",
          4567 => x"f8",
          4568 => x"70",
          4569 => x"59",
          4570 => x"ee",
          4571 => x"ff",
          4572 => x"b4",
          4573 => x"2b",
          4574 => x"82",
          4575 => x"70",
          4576 => x"97",
          4577 => x"2c",
          4578 => x"29",
          4579 => x"05",
          4580 => x"70",
          4581 => x"51",
          4582 => x"51",
          4583 => x"81",
          4584 => x"2e",
          4585 => x"77",
          4586 => x"38",
          4587 => x"0a",
          4588 => x"0a",
          4589 => x"2c",
          4590 => x"75",
          4591 => x"38",
          4592 => x"52",
          4593 => x"85",
          4594 => x"f8",
          4595 => x"06",
          4596 => x"2e",
          4597 => x"82",
          4598 => x"81",
          4599 => x"74",
          4600 => x"29",
          4601 => x"05",
          4602 => x"70",
          4603 => x"56",
          4604 => x"95",
          4605 => x"76",
          4606 => x"77",
          4607 => x"3f",
          4608 => x"08",
          4609 => x"54",
          4610 => x"d3",
          4611 => x"75",
          4612 => x"ca",
          4613 => x"55",
          4614 => x"b4",
          4615 => x"2b",
          4616 => x"82",
          4617 => x"70",
          4618 => x"98",
          4619 => x"11",
          4620 => x"82",
          4621 => x"33",
          4622 => x"51",
          4623 => x"55",
          4624 => x"09",
          4625 => x"92",
          4626 => x"c8",
          4627 => x"0c",
          4628 => x"ec",
          4629 => x"0b",
          4630 => x"34",
          4631 => x"82",
          4632 => x"75",
          4633 => x"34",
          4634 => x"34",
          4635 => x"7e",
          4636 => x"26",
          4637 => x"73",
          4638 => x"ac",
          4639 => x"73",
          4640 => x"ec",
          4641 => x"73",
          4642 => x"cb",
          4643 => x"b8",
          4644 => x"75",
          4645 => x"74",
          4646 => x"98",
          4647 => x"73",
          4648 => x"38",
          4649 => x"73",
          4650 => x"34",
          4651 => x"0a",
          4652 => x"0a",
          4653 => x"2c",
          4654 => x"33",
          4655 => x"df",
          4656 => x"bc",
          4657 => x"56",
          4658 => x"ec",
          4659 => x"1a",
          4660 => x"33",
          4661 => x"ec",
          4662 => x"73",
          4663 => x"38",
          4664 => x"73",
          4665 => x"34",
          4666 => x"33",
          4667 => x"0a",
          4668 => x"0a",
          4669 => x"2c",
          4670 => x"33",
          4671 => x"56",
          4672 => x"a8",
          4673 => x"dc",
          4674 => x"1a",
          4675 => x"54",
          4676 => x"3f",
          4677 => x"0a",
          4678 => x"0a",
          4679 => x"2c",
          4680 => x"33",
          4681 => x"73",
          4682 => x"38",
          4683 => x"33",
          4684 => x"70",
          4685 => x"ec",
          4686 => x"51",
          4687 => x"77",
          4688 => x"38",
          4689 => x"08",
          4690 => x"ff",
          4691 => x"74",
          4692 => x"29",
          4693 => x"05",
          4694 => x"82",
          4695 => x"56",
          4696 => x"75",
          4697 => x"fb",
          4698 => x"7a",
          4699 => x"81",
          4700 => x"ec",
          4701 => x"52",
          4702 => x"51",
          4703 => x"81",
          4704 => x"ec",
          4705 => x"81",
          4706 => x"55",
          4707 => x"fb",
          4708 => x"ec",
          4709 => x"05",
          4710 => x"ec",
          4711 => x"15",
          4712 => x"ec",
          4713 => x"f0",
          4714 => x"88",
          4715 => x"84",
          4716 => x"bc",
          4717 => x"2b",
          4718 => x"82",
          4719 => x"57",
          4720 => x"74",
          4721 => x"38",
          4722 => x"81",
          4723 => x"34",
          4724 => x"08",
          4725 => x"51",
          4726 => x"3f",
          4727 => x"0a",
          4728 => x"0a",
          4729 => x"2c",
          4730 => x"33",
          4731 => x"75",
          4732 => x"38",
          4733 => x"08",
          4734 => x"ff",
          4735 => x"82",
          4736 => x"70",
          4737 => x"98",
          4738 => x"b8",
          4739 => x"56",
          4740 => x"24",
          4741 => x"82",
          4742 => x"52",
          4743 => x"9f",
          4744 => x"81",
          4745 => x"81",
          4746 => x"70",
          4747 => x"ec",
          4748 => x"51",
          4749 => x"25",
          4750 => x"9b",
          4751 => x"b8",
          4752 => x"54",
          4753 => x"82",
          4754 => x"52",
          4755 => x"9e",
          4756 => x"ec",
          4757 => x"51",
          4758 => x"82",
          4759 => x"81",
          4760 => x"73",
          4761 => x"ec",
          4762 => x"73",
          4763 => x"38",
          4764 => x"52",
          4765 => x"f3",
          4766 => x"80",
          4767 => x"0b",
          4768 => x"34",
          4769 => x"ec",
          4770 => x"82",
          4771 => x"af",
          4772 => x"82",
          4773 => x"54",
          4774 => x"f9",
          4775 => x"f0",
          4776 => x"88",
          4777 => x"8c",
          4778 => x"bc",
          4779 => x"54",
          4780 => x"bc",
          4781 => x"ff",
          4782 => x"39",
          4783 => x"33",
          4784 => x"33",
          4785 => x"75",
          4786 => x"38",
          4787 => x"73",
          4788 => x"34",
          4789 => x"70",
          4790 => x"81",
          4791 => x"51",
          4792 => x"25",
          4793 => x"1a",
          4794 => x"33",
          4795 => x"f0",
          4796 => x"73",
          4797 => x"9d",
          4798 => x"81",
          4799 => x"81",
          4800 => x"70",
          4801 => x"ec",
          4802 => x"51",
          4803 => x"24",
          4804 => x"f0",
          4805 => x"a0",
          4806 => x"98",
          4807 => x"bc",
          4808 => x"2b",
          4809 => x"82",
          4810 => x"57",
          4811 => x"74",
          4812 => x"a3",
          4813 => x"dc",
          4814 => x"51",
          4815 => x"3f",
          4816 => x"0a",
          4817 => x"0a",
          4818 => x"2c",
          4819 => x"33",
          4820 => x"75",
          4821 => x"38",
          4822 => x"82",
          4823 => x"70",
          4824 => x"82",
          4825 => x"59",
          4826 => x"77",
          4827 => x"38",
          4828 => x"08",
          4829 => x"54",
          4830 => x"bc",
          4831 => x"70",
          4832 => x"ff",
          4833 => x"82",
          4834 => x"70",
          4835 => x"82",
          4836 => x"58",
          4837 => x"75",
          4838 => x"f7",
          4839 => x"ec",
          4840 => x"52",
          4841 => x"51",
          4842 => x"80",
          4843 => x"bc",
          4844 => x"82",
          4845 => x"f7",
          4846 => x"b0",
          4847 => x"c4",
          4848 => x"80",
          4849 => x"74",
          4850 => x"bb",
          4851 => x"f8",
          4852 => x"b8",
          4853 => x"f8",
          4854 => x"06",
          4855 => x"74",
          4856 => x"ff",
          4857 => x"93",
          4858 => x"39",
          4859 => x"82",
          4860 => x"fc",
          4861 => x"54",
          4862 => x"a7",
          4863 => x"ff",
          4864 => x"82",
          4865 => x"82",
          4866 => x"82",
          4867 => x"81",
          4868 => x"05",
          4869 => x"79",
          4870 => x"cb",
          4871 => x"54",
          4872 => x"73",
          4873 => x"80",
          4874 => x"38",
          4875 => x"a3",
          4876 => x"39",
          4877 => x"09",
          4878 => x"38",
          4879 => x"08",
          4880 => x"2e",
          4881 => x"51",
          4882 => x"3f",
          4883 => x"08",
          4884 => x"34",
          4885 => x"08",
          4886 => x"81",
          4887 => x"52",
          4888 => x"a5",
          4889 => x"c3",
          4890 => x"29",
          4891 => x"05",
          4892 => x"54",
          4893 => x"ab",
          4894 => x"ff",
          4895 => x"82",
          4896 => x"82",
          4897 => x"82",
          4898 => x"81",
          4899 => x"05",
          4900 => x"79",
          4901 => x"cf",
          4902 => x"54",
          4903 => x"06",
          4904 => x"74",
          4905 => x"34",
          4906 => x"82",
          4907 => x"82",
          4908 => x"52",
          4909 => x"e2",
          4910 => x"39",
          4911 => x"33",
          4912 => x"06",
          4913 => x"33",
          4914 => x"74",
          4915 => x"87",
          4916 => x"dc",
          4917 => x"14",
          4918 => x"ec",
          4919 => x"1a",
          4920 => x"54",
          4921 => x"3f",
          4922 => x"82",
          4923 => x"54",
          4924 => x"f4",
          4925 => x"f0",
          4926 => x"88",
          4927 => x"b4",
          4928 => x"bc",
          4929 => x"54",
          4930 => x"bc",
          4931 => x"39",
          4932 => x"86",
          4933 => x"82",
          4934 => x"8c",
          4935 => x"d4",
          4936 => x"e0",
          4937 => x"52",
          4938 => x"51",
          4939 => x"3f",
          4940 => x"08",
          4941 => x"77",
          4942 => x"57",
          4943 => x"34",
          4944 => x"08",
          4945 => x"15",
          4946 => x"15",
          4947 => x"f0",
          4948 => x"86",
          4949 => x"87",
          4950 => x"d4",
          4951 => x"d4",
          4952 => x"05",
          4953 => x"07",
          4954 => x"ff",
          4955 => x"2a",
          4956 => x"56",
          4957 => x"34",
          4958 => x"34",
          4959 => x"22",
          4960 => x"82",
          4961 => x"05",
          4962 => x"55",
          4963 => x"15",
          4964 => x"15",
          4965 => x"0d",
          4966 => x"0d",
          4967 => x"51",
          4968 => x"8f",
          4969 => x"83",
          4970 => x"70",
          4971 => x"06",
          4972 => x"70",
          4973 => x"0c",
          4974 => x"04",
          4975 => x"02",
          4976 => x"02",
          4977 => x"05",
          4978 => x"82",
          4979 => x"71",
          4980 => x"11",
          4981 => x"73",
          4982 => x"81",
          4983 => x"88",
          4984 => x"a4",
          4985 => x"22",
          4986 => x"ff",
          4987 => x"88",
          4988 => x"52",
          4989 => x"5b",
          4990 => x"55",
          4991 => x"70",
          4992 => x"82",
          4993 => x"14",
          4994 => x"52",
          4995 => x"15",
          4996 => x"15",
          4997 => x"f0",
          4998 => x"70",
          4999 => x"33",
          5000 => x"07",
          5001 => x"8f",
          5002 => x"51",
          5003 => x"71",
          5004 => x"ff",
          5005 => x"88",
          5006 => x"51",
          5007 => x"34",
          5008 => x"06",
          5009 => x"12",
          5010 => x"f0",
          5011 => x"71",
          5012 => x"81",
          5013 => x"3d",
          5014 => x"3d",
          5015 => x"f0",
          5016 => x"05",
          5017 => x"70",
          5018 => x"11",
          5019 => x"87",
          5020 => x"8b",
          5021 => x"2b",
          5022 => x"59",
          5023 => x"72",
          5024 => x"33",
          5025 => x"71",
          5026 => x"70",
          5027 => x"56",
          5028 => x"84",
          5029 => x"85",
          5030 => x"d4",
          5031 => x"14",
          5032 => x"85",
          5033 => x"8b",
          5034 => x"2b",
          5035 => x"57",
          5036 => x"86",
          5037 => x"13",
          5038 => x"2b",
          5039 => x"2a",
          5040 => x"52",
          5041 => x"34",
          5042 => x"34",
          5043 => x"08",
          5044 => x"81",
          5045 => x"88",
          5046 => x"81",
          5047 => x"70",
          5048 => x"51",
          5049 => x"71",
          5050 => x"81",
          5051 => x"3d",
          5052 => x"3d",
          5053 => x"05",
          5054 => x"f0",
          5055 => x"2b",
          5056 => x"33",
          5057 => x"71",
          5058 => x"70",
          5059 => x"70",
          5060 => x"33",
          5061 => x"71",
          5062 => x"53",
          5063 => x"52",
          5064 => x"53",
          5065 => x"25",
          5066 => x"72",
          5067 => x"3f",
          5068 => x"08",
          5069 => x"33",
          5070 => x"71",
          5071 => x"83",
          5072 => x"11",
          5073 => x"12",
          5074 => x"2b",
          5075 => x"2b",
          5076 => x"06",
          5077 => x"51",
          5078 => x"53",
          5079 => x"88",
          5080 => x"72",
          5081 => x"73",
          5082 => x"82",
          5083 => x"70",
          5084 => x"81",
          5085 => x"8b",
          5086 => x"2b",
          5087 => x"57",
          5088 => x"70",
          5089 => x"33",
          5090 => x"07",
          5091 => x"ff",
          5092 => x"2a",
          5093 => x"58",
          5094 => x"34",
          5095 => x"34",
          5096 => x"04",
          5097 => x"82",
          5098 => x"02",
          5099 => x"05",
          5100 => x"2b",
          5101 => x"11",
          5102 => x"33",
          5103 => x"71",
          5104 => x"59",
          5105 => x"56",
          5106 => x"71",
          5107 => x"33",
          5108 => x"07",
          5109 => x"a2",
          5110 => x"07",
          5111 => x"53",
          5112 => x"53",
          5113 => x"70",
          5114 => x"82",
          5115 => x"70",
          5116 => x"81",
          5117 => x"8b",
          5118 => x"2b",
          5119 => x"57",
          5120 => x"82",
          5121 => x"13",
          5122 => x"2b",
          5123 => x"2a",
          5124 => x"52",
          5125 => x"34",
          5126 => x"34",
          5127 => x"08",
          5128 => x"33",
          5129 => x"71",
          5130 => x"82",
          5131 => x"52",
          5132 => x"0d",
          5133 => x"0d",
          5134 => x"f0",
          5135 => x"2a",
          5136 => x"ff",
          5137 => x"57",
          5138 => x"3f",
          5139 => x"08",
          5140 => x"71",
          5141 => x"33",
          5142 => x"71",
          5143 => x"83",
          5144 => x"11",
          5145 => x"12",
          5146 => x"2b",
          5147 => x"07",
          5148 => x"51",
          5149 => x"55",
          5150 => x"80",
          5151 => x"82",
          5152 => x"75",
          5153 => x"3f",
          5154 => x"84",
          5155 => x"15",
          5156 => x"2b",
          5157 => x"07",
          5158 => x"88",
          5159 => x"55",
          5160 => x"86",
          5161 => x"81",
          5162 => x"75",
          5163 => x"82",
          5164 => x"70",
          5165 => x"33",
          5166 => x"71",
          5167 => x"70",
          5168 => x"57",
          5169 => x"72",
          5170 => x"73",
          5171 => x"82",
          5172 => x"18",
          5173 => x"86",
          5174 => x"0b",
          5175 => x"82",
          5176 => x"53",
          5177 => x"34",
          5178 => x"34",
          5179 => x"08",
          5180 => x"81",
          5181 => x"88",
          5182 => x"82",
          5183 => x"70",
          5184 => x"51",
          5185 => x"74",
          5186 => x"81",
          5187 => x"3d",
          5188 => x"3d",
          5189 => x"82",
          5190 => x"84",
          5191 => x"3f",
          5192 => x"86",
          5193 => x"fe",
          5194 => x"3d",
          5195 => x"3d",
          5196 => x"52",
          5197 => x"3f",
          5198 => x"08",
          5199 => x"06",
          5200 => x"08",
          5201 => x"85",
          5202 => x"88",
          5203 => x"5f",
          5204 => x"5a",
          5205 => x"59",
          5206 => x"80",
          5207 => x"88",
          5208 => x"33",
          5209 => x"71",
          5210 => x"70",
          5211 => x"06",
          5212 => x"83",
          5213 => x"70",
          5214 => x"53",
          5215 => x"55",
          5216 => x"8a",
          5217 => x"2e",
          5218 => x"78",
          5219 => x"15",
          5220 => x"33",
          5221 => x"07",
          5222 => x"c2",
          5223 => x"ff",
          5224 => x"38",
          5225 => x"56",
          5226 => x"2b",
          5227 => x"08",
          5228 => x"81",
          5229 => x"88",
          5230 => x"81",
          5231 => x"51",
          5232 => x"5c",
          5233 => x"2e",
          5234 => x"55",
          5235 => x"78",
          5236 => x"38",
          5237 => x"80",
          5238 => x"38",
          5239 => x"09",
          5240 => x"38",
          5241 => x"f2",
          5242 => x"39",
          5243 => x"53",
          5244 => x"51",
          5245 => x"82",
          5246 => x"70",
          5247 => x"33",
          5248 => x"71",
          5249 => x"83",
          5250 => x"5a",
          5251 => x"05",
          5252 => x"83",
          5253 => x"70",
          5254 => x"59",
          5255 => x"84",
          5256 => x"81",
          5257 => x"76",
          5258 => x"82",
          5259 => x"75",
          5260 => x"11",
          5261 => x"11",
          5262 => x"33",
          5263 => x"07",
          5264 => x"53",
          5265 => x"5a",
          5266 => x"86",
          5267 => x"87",
          5268 => x"d4",
          5269 => x"1c",
          5270 => x"85",
          5271 => x"8b",
          5272 => x"2b",
          5273 => x"5a",
          5274 => x"54",
          5275 => x"34",
          5276 => x"34",
          5277 => x"08",
          5278 => x"1d",
          5279 => x"85",
          5280 => x"88",
          5281 => x"88",
          5282 => x"5f",
          5283 => x"73",
          5284 => x"75",
          5285 => x"82",
          5286 => x"1b",
          5287 => x"73",
          5288 => x"0c",
          5289 => x"04",
          5290 => x"74",
          5291 => x"f0",
          5292 => x"f4",
          5293 => x"53",
          5294 => x"8b",
          5295 => x"fc",
          5296 => x"d4",
          5297 => x"72",
          5298 => x"0c",
          5299 => x"04",
          5300 => x"64",
          5301 => x"80",
          5302 => x"82",
          5303 => x"60",
          5304 => x"06",
          5305 => x"a8",
          5306 => x"38",
          5307 => x"b8",
          5308 => x"f8",
          5309 => x"c7",
          5310 => x"38",
          5311 => x"92",
          5312 => x"83",
          5313 => x"51",
          5314 => x"82",
          5315 => x"83",
          5316 => x"82",
          5317 => x"7d",
          5318 => x"2a",
          5319 => x"ff",
          5320 => x"2b",
          5321 => x"33",
          5322 => x"71",
          5323 => x"70",
          5324 => x"83",
          5325 => x"70",
          5326 => x"05",
          5327 => x"1a",
          5328 => x"12",
          5329 => x"2b",
          5330 => x"2b",
          5331 => x"53",
          5332 => x"5c",
          5333 => x"5c",
          5334 => x"73",
          5335 => x"38",
          5336 => x"ff",
          5337 => x"70",
          5338 => x"06",
          5339 => x"16",
          5340 => x"33",
          5341 => x"07",
          5342 => x"1c",
          5343 => x"12",
          5344 => x"2b",
          5345 => x"07",
          5346 => x"52",
          5347 => x"80",
          5348 => x"78",
          5349 => x"83",
          5350 => x"41",
          5351 => x"27",
          5352 => x"60",
          5353 => x"7b",
          5354 => x"06",
          5355 => x"51",
          5356 => x"7a",
          5357 => x"06",
          5358 => x"39",
          5359 => x"7a",
          5360 => x"38",
          5361 => x"aa",
          5362 => x"39",
          5363 => x"7a",
          5364 => x"c8",
          5365 => x"82",
          5366 => x"12",
          5367 => x"2b",
          5368 => x"54",
          5369 => x"80",
          5370 => x"f7",
          5371 => x"d4",
          5372 => x"ff",
          5373 => x"54",
          5374 => x"83",
          5375 => x"f0",
          5376 => x"05",
          5377 => x"ff",
          5378 => x"82",
          5379 => x"14",
          5380 => x"83",
          5381 => x"59",
          5382 => x"39",
          5383 => x"7a",
          5384 => x"d4",
          5385 => x"f5",
          5386 => x"d4",
          5387 => x"82",
          5388 => x"12",
          5389 => x"2b",
          5390 => x"54",
          5391 => x"80",
          5392 => x"f6",
          5393 => x"d4",
          5394 => x"ff",
          5395 => x"54",
          5396 => x"83",
          5397 => x"f0",
          5398 => x"05",
          5399 => x"ff",
          5400 => x"82",
          5401 => x"14",
          5402 => x"62",
          5403 => x"5c",
          5404 => x"ff",
          5405 => x"39",
          5406 => x"54",
          5407 => x"82",
          5408 => x"5c",
          5409 => x"08",
          5410 => x"38",
          5411 => x"52",
          5412 => x"08",
          5413 => x"cf",
          5414 => x"f7",
          5415 => x"58",
          5416 => x"99",
          5417 => x"7a",
          5418 => x"f2",
          5419 => x"19",
          5420 => x"d4",
          5421 => x"84",
          5422 => x"f9",
          5423 => x"73",
          5424 => x"0c",
          5425 => x"04",
          5426 => x"77",
          5427 => x"52",
          5428 => x"3f",
          5429 => x"08",
          5430 => x"f8",
          5431 => x"8e",
          5432 => x"80",
          5433 => x"f8",
          5434 => x"9a",
          5435 => x"82",
          5436 => x"86",
          5437 => x"ff",
          5438 => x"8f",
          5439 => x"81",
          5440 => x"26",
          5441 => x"d4",
          5442 => x"52",
          5443 => x"f8",
          5444 => x"0d",
          5445 => x"0d",
          5446 => x"33",
          5447 => x"9f",
          5448 => x"53",
          5449 => x"81",
          5450 => x"38",
          5451 => x"87",
          5452 => x"11",
          5453 => x"54",
          5454 => x"84",
          5455 => x"54",
          5456 => x"87",
          5457 => x"11",
          5458 => x"0c",
          5459 => x"c0",
          5460 => x"70",
          5461 => x"70",
          5462 => x"51",
          5463 => x"8a",
          5464 => x"98",
          5465 => x"70",
          5466 => x"08",
          5467 => x"06",
          5468 => x"38",
          5469 => x"8c",
          5470 => x"80",
          5471 => x"71",
          5472 => x"14",
          5473 => x"f4",
          5474 => x"70",
          5475 => x"0c",
          5476 => x"04",
          5477 => x"60",
          5478 => x"8c",
          5479 => x"33",
          5480 => x"5b",
          5481 => x"5a",
          5482 => x"82",
          5483 => x"81",
          5484 => x"52",
          5485 => x"38",
          5486 => x"84",
          5487 => x"92",
          5488 => x"c0",
          5489 => x"87",
          5490 => x"13",
          5491 => x"57",
          5492 => x"0b",
          5493 => x"8c",
          5494 => x"0c",
          5495 => x"75",
          5496 => x"2a",
          5497 => x"51",
          5498 => x"80",
          5499 => x"7b",
          5500 => x"7b",
          5501 => x"5d",
          5502 => x"59",
          5503 => x"06",
          5504 => x"73",
          5505 => x"81",
          5506 => x"ff",
          5507 => x"72",
          5508 => x"38",
          5509 => x"8c",
          5510 => x"c3",
          5511 => x"98",
          5512 => x"71",
          5513 => x"38",
          5514 => x"2e",
          5515 => x"76",
          5516 => x"92",
          5517 => x"72",
          5518 => x"06",
          5519 => x"f7",
          5520 => x"5a",
          5521 => x"80",
          5522 => x"70",
          5523 => x"5a",
          5524 => x"80",
          5525 => x"73",
          5526 => x"06",
          5527 => x"38",
          5528 => x"fe",
          5529 => x"fc",
          5530 => x"52",
          5531 => x"83",
          5532 => x"71",
          5533 => x"d4",
          5534 => x"3d",
          5535 => x"3d",
          5536 => x"64",
          5537 => x"bf",
          5538 => x"40",
          5539 => x"59",
          5540 => x"58",
          5541 => x"82",
          5542 => x"81",
          5543 => x"52",
          5544 => x"09",
          5545 => x"b1",
          5546 => x"84",
          5547 => x"92",
          5548 => x"c0",
          5549 => x"87",
          5550 => x"13",
          5551 => x"56",
          5552 => x"87",
          5553 => x"0c",
          5554 => x"82",
          5555 => x"58",
          5556 => x"84",
          5557 => x"06",
          5558 => x"71",
          5559 => x"38",
          5560 => x"05",
          5561 => x"0c",
          5562 => x"73",
          5563 => x"81",
          5564 => x"71",
          5565 => x"38",
          5566 => x"8c",
          5567 => x"d0",
          5568 => x"98",
          5569 => x"71",
          5570 => x"38",
          5571 => x"2e",
          5572 => x"76",
          5573 => x"92",
          5574 => x"72",
          5575 => x"06",
          5576 => x"f7",
          5577 => x"59",
          5578 => x"1a",
          5579 => x"06",
          5580 => x"59",
          5581 => x"80",
          5582 => x"73",
          5583 => x"06",
          5584 => x"38",
          5585 => x"fe",
          5586 => x"fc",
          5587 => x"52",
          5588 => x"83",
          5589 => x"71",
          5590 => x"d4",
          5591 => x"3d",
          5592 => x"3d",
          5593 => x"84",
          5594 => x"33",
          5595 => x"a7",
          5596 => x"54",
          5597 => x"fa",
          5598 => x"d4",
          5599 => x"06",
          5600 => x"72",
          5601 => x"85",
          5602 => x"98",
          5603 => x"56",
          5604 => x"80",
          5605 => x"76",
          5606 => x"74",
          5607 => x"c0",
          5608 => x"54",
          5609 => x"2e",
          5610 => x"d4",
          5611 => x"2e",
          5612 => x"80",
          5613 => x"08",
          5614 => x"70",
          5615 => x"51",
          5616 => x"2e",
          5617 => x"c0",
          5618 => x"52",
          5619 => x"87",
          5620 => x"08",
          5621 => x"38",
          5622 => x"87",
          5623 => x"14",
          5624 => x"70",
          5625 => x"52",
          5626 => x"96",
          5627 => x"92",
          5628 => x"0a",
          5629 => x"39",
          5630 => x"0c",
          5631 => x"39",
          5632 => x"54",
          5633 => x"f8",
          5634 => x"0d",
          5635 => x"0d",
          5636 => x"33",
          5637 => x"88",
          5638 => x"d4",
          5639 => x"51",
          5640 => x"04",
          5641 => x"75",
          5642 => x"82",
          5643 => x"90",
          5644 => x"2b",
          5645 => x"33",
          5646 => x"88",
          5647 => x"71",
          5648 => x"f8",
          5649 => x"54",
          5650 => x"85",
          5651 => x"ff",
          5652 => x"02",
          5653 => x"05",
          5654 => x"70",
          5655 => x"05",
          5656 => x"88",
          5657 => x"72",
          5658 => x"0d",
          5659 => x"0d",
          5660 => x"52",
          5661 => x"81",
          5662 => x"70",
          5663 => x"70",
          5664 => x"05",
          5665 => x"88",
          5666 => x"72",
          5667 => x"54",
          5668 => x"2a",
          5669 => x"34",
          5670 => x"04",
          5671 => x"76",
          5672 => x"54",
          5673 => x"2e",
          5674 => x"70",
          5675 => x"33",
          5676 => x"05",
          5677 => x"11",
          5678 => x"84",
          5679 => x"fe",
          5680 => x"77",
          5681 => x"53",
          5682 => x"81",
          5683 => x"ff",
          5684 => x"f4",
          5685 => x"0d",
          5686 => x"0d",
          5687 => x"56",
          5688 => x"70",
          5689 => x"33",
          5690 => x"05",
          5691 => x"71",
          5692 => x"56",
          5693 => x"72",
          5694 => x"38",
          5695 => x"e2",
          5696 => x"d4",
          5697 => x"3d",
          5698 => x"3d",
          5699 => x"54",
          5700 => x"71",
          5701 => x"38",
          5702 => x"70",
          5703 => x"f3",
          5704 => x"82",
          5705 => x"84",
          5706 => x"80",
          5707 => x"f8",
          5708 => x"3d",
          5709 => x"08",
          5710 => x"05",
          5711 => x"54",
          5712 => x"e7",
          5713 => x"82",
          5714 => x"a2",
          5715 => x"2e",
          5716 => x"b5",
          5717 => x"80",
          5718 => x"82",
          5719 => x"83",
          5720 => x"53",
          5721 => x"86",
          5722 => x"0c",
          5723 => x"82",
          5724 => x"87",
          5725 => x"f7",
          5726 => x"56",
          5727 => x"17",
          5728 => x"74",
          5729 => x"d6",
          5730 => x"b4",
          5731 => x"b8",
          5732 => x"81",
          5733 => x"59",
          5734 => x"82",
          5735 => x"7a",
          5736 => x"06",
          5737 => x"d4",
          5738 => x"17",
          5739 => x"08",
          5740 => x"08",
          5741 => x"08",
          5742 => x"74",
          5743 => x"38",
          5744 => x"55",
          5745 => x"09",
          5746 => x"38",
          5747 => x"18",
          5748 => x"81",
          5749 => x"f9",
          5750 => x"39",
          5751 => x"82",
          5752 => x"8b",
          5753 => x"fa",
          5754 => x"7a",
          5755 => x"57",
          5756 => x"08",
          5757 => x"75",
          5758 => x"3f",
          5759 => x"08",
          5760 => x"f8",
          5761 => x"81",
          5762 => x"b8",
          5763 => x"16",
          5764 => x"80",
          5765 => x"f8",
          5766 => x"85",
          5767 => x"81",
          5768 => x"17",
          5769 => x"d4",
          5770 => x"3d",
          5771 => x"3d",
          5772 => x"52",
          5773 => x"3f",
          5774 => x"08",
          5775 => x"f8",
          5776 => x"38",
          5777 => x"74",
          5778 => x"81",
          5779 => x"38",
          5780 => x"59",
          5781 => x"09",
          5782 => x"e3",
          5783 => x"53",
          5784 => x"08",
          5785 => x"70",
          5786 => x"d3",
          5787 => x"d5",
          5788 => x"17",
          5789 => x"3f",
          5790 => x"a4",
          5791 => x"51",
          5792 => x"86",
          5793 => x"f2",
          5794 => x"17",
          5795 => x"3f",
          5796 => x"52",
          5797 => x"51",
          5798 => x"90",
          5799 => x"84",
          5800 => x"fb",
          5801 => x"17",
          5802 => x"70",
          5803 => x"79",
          5804 => x"52",
          5805 => x"51",
          5806 => x"77",
          5807 => x"80",
          5808 => x"81",
          5809 => x"f9",
          5810 => x"d4",
          5811 => x"2e",
          5812 => x"58",
          5813 => x"f8",
          5814 => x"0d",
          5815 => x"0d",
          5816 => x"9c",
          5817 => x"05",
          5818 => x"80",
          5819 => x"27",
          5820 => x"14",
          5821 => x"29",
          5822 => x"05",
          5823 => x"82",
          5824 => x"87",
          5825 => x"f9",
          5826 => x"7a",
          5827 => x"54",
          5828 => x"27",
          5829 => x"76",
          5830 => x"27",
          5831 => x"ff",
          5832 => x"58",
          5833 => x"80",
          5834 => x"82",
          5835 => x"72",
          5836 => x"38",
          5837 => x"72",
          5838 => x"8e",
          5839 => x"39",
          5840 => x"17",
          5841 => x"a8",
          5842 => x"53",
          5843 => x"fd",
          5844 => x"d4",
          5845 => x"9f",
          5846 => x"ff",
          5847 => x"11",
          5848 => x"70",
          5849 => x"18",
          5850 => x"76",
          5851 => x"53",
          5852 => x"82",
          5853 => x"80",
          5854 => x"83",
          5855 => x"b8",
          5856 => x"88",
          5857 => x"79",
          5858 => x"84",
          5859 => x"58",
          5860 => x"80",
          5861 => x"9f",
          5862 => x"80",
          5863 => x"88",
          5864 => x"08",
          5865 => x"51",
          5866 => x"82",
          5867 => x"80",
          5868 => x"10",
          5869 => x"74",
          5870 => x"51",
          5871 => x"82",
          5872 => x"83",
          5873 => x"58",
          5874 => x"87",
          5875 => x"08",
          5876 => x"51",
          5877 => x"82",
          5878 => x"9b",
          5879 => x"2b",
          5880 => x"74",
          5881 => x"51",
          5882 => x"82",
          5883 => x"f0",
          5884 => x"83",
          5885 => x"77",
          5886 => x"0c",
          5887 => x"04",
          5888 => x"7a",
          5889 => x"58",
          5890 => x"81",
          5891 => x"9e",
          5892 => x"17",
          5893 => x"96",
          5894 => x"53",
          5895 => x"81",
          5896 => x"79",
          5897 => x"72",
          5898 => x"38",
          5899 => x"72",
          5900 => x"b8",
          5901 => x"39",
          5902 => x"17",
          5903 => x"a8",
          5904 => x"53",
          5905 => x"fb",
          5906 => x"d4",
          5907 => x"82",
          5908 => x"81",
          5909 => x"83",
          5910 => x"b8",
          5911 => x"78",
          5912 => x"56",
          5913 => x"76",
          5914 => x"38",
          5915 => x"9f",
          5916 => x"33",
          5917 => x"07",
          5918 => x"74",
          5919 => x"83",
          5920 => x"89",
          5921 => x"08",
          5922 => x"51",
          5923 => x"82",
          5924 => x"59",
          5925 => x"08",
          5926 => x"74",
          5927 => x"16",
          5928 => x"84",
          5929 => x"76",
          5930 => x"88",
          5931 => x"81",
          5932 => x"8f",
          5933 => x"53",
          5934 => x"80",
          5935 => x"88",
          5936 => x"08",
          5937 => x"51",
          5938 => x"82",
          5939 => x"59",
          5940 => x"08",
          5941 => x"77",
          5942 => x"06",
          5943 => x"83",
          5944 => x"05",
          5945 => x"f6",
          5946 => x"39",
          5947 => x"a8",
          5948 => x"52",
          5949 => x"ef",
          5950 => x"f8",
          5951 => x"d4",
          5952 => x"38",
          5953 => x"06",
          5954 => x"83",
          5955 => x"18",
          5956 => x"54",
          5957 => x"f6",
          5958 => x"d4",
          5959 => x"0a",
          5960 => x"52",
          5961 => x"c5",
          5962 => x"83",
          5963 => x"82",
          5964 => x"8a",
          5965 => x"f8",
          5966 => x"7c",
          5967 => x"59",
          5968 => x"81",
          5969 => x"38",
          5970 => x"08",
          5971 => x"73",
          5972 => x"38",
          5973 => x"52",
          5974 => x"a4",
          5975 => x"f8",
          5976 => x"d4",
          5977 => x"f2",
          5978 => x"82",
          5979 => x"39",
          5980 => x"e6",
          5981 => x"f8",
          5982 => x"de",
          5983 => x"78",
          5984 => x"3f",
          5985 => x"08",
          5986 => x"f8",
          5987 => x"80",
          5988 => x"d4",
          5989 => x"2e",
          5990 => x"d4",
          5991 => x"2e",
          5992 => x"53",
          5993 => x"51",
          5994 => x"82",
          5995 => x"c5",
          5996 => x"08",
          5997 => x"18",
          5998 => x"57",
          5999 => x"90",
          6000 => x"94",
          6001 => x"16",
          6002 => x"54",
          6003 => x"34",
          6004 => x"78",
          6005 => x"38",
          6006 => x"82",
          6007 => x"8a",
          6008 => x"f6",
          6009 => x"7e",
          6010 => x"5b",
          6011 => x"38",
          6012 => x"58",
          6013 => x"88",
          6014 => x"08",
          6015 => x"38",
          6016 => x"39",
          6017 => x"51",
          6018 => x"81",
          6019 => x"d4",
          6020 => x"82",
          6021 => x"d4",
          6022 => x"82",
          6023 => x"ff",
          6024 => x"38",
          6025 => x"82",
          6026 => x"26",
          6027 => x"79",
          6028 => x"08",
          6029 => x"73",
          6030 => x"b9",
          6031 => x"2e",
          6032 => x"80",
          6033 => x"1a",
          6034 => x"08",
          6035 => x"38",
          6036 => x"52",
          6037 => x"af",
          6038 => x"82",
          6039 => x"81",
          6040 => x"06",
          6041 => x"d4",
          6042 => x"82",
          6043 => x"09",
          6044 => x"72",
          6045 => x"70",
          6046 => x"d4",
          6047 => x"51",
          6048 => x"73",
          6049 => x"82",
          6050 => x"80",
          6051 => x"90",
          6052 => x"81",
          6053 => x"38",
          6054 => x"08",
          6055 => x"73",
          6056 => x"75",
          6057 => x"77",
          6058 => x"56",
          6059 => x"76",
          6060 => x"82",
          6061 => x"26",
          6062 => x"75",
          6063 => x"f8",
          6064 => x"d4",
          6065 => x"2e",
          6066 => x"59",
          6067 => x"08",
          6068 => x"81",
          6069 => x"82",
          6070 => x"59",
          6071 => x"08",
          6072 => x"70",
          6073 => x"25",
          6074 => x"51",
          6075 => x"73",
          6076 => x"75",
          6077 => x"81",
          6078 => x"38",
          6079 => x"f5",
          6080 => x"75",
          6081 => x"f9",
          6082 => x"d4",
          6083 => x"d4",
          6084 => x"70",
          6085 => x"08",
          6086 => x"51",
          6087 => x"80",
          6088 => x"73",
          6089 => x"38",
          6090 => x"52",
          6091 => x"d0",
          6092 => x"f8",
          6093 => x"a5",
          6094 => x"18",
          6095 => x"08",
          6096 => x"18",
          6097 => x"74",
          6098 => x"38",
          6099 => x"18",
          6100 => x"33",
          6101 => x"73",
          6102 => x"97",
          6103 => x"74",
          6104 => x"38",
          6105 => x"55",
          6106 => x"d4",
          6107 => x"85",
          6108 => x"75",
          6109 => x"d4",
          6110 => x"3d",
          6111 => x"3d",
          6112 => x"52",
          6113 => x"3f",
          6114 => x"08",
          6115 => x"82",
          6116 => x"80",
          6117 => x"52",
          6118 => x"c1",
          6119 => x"f8",
          6120 => x"f8",
          6121 => x"0c",
          6122 => x"53",
          6123 => x"15",
          6124 => x"f2",
          6125 => x"56",
          6126 => x"16",
          6127 => x"22",
          6128 => x"27",
          6129 => x"54",
          6130 => x"76",
          6131 => x"33",
          6132 => x"3f",
          6133 => x"08",
          6134 => x"38",
          6135 => x"76",
          6136 => x"70",
          6137 => x"9f",
          6138 => x"56",
          6139 => x"d4",
          6140 => x"3d",
          6141 => x"3d",
          6142 => x"71",
          6143 => x"57",
          6144 => x"0a",
          6145 => x"38",
          6146 => x"53",
          6147 => x"38",
          6148 => x"0c",
          6149 => x"54",
          6150 => x"75",
          6151 => x"73",
          6152 => x"ac",
          6153 => x"73",
          6154 => x"85",
          6155 => x"0b",
          6156 => x"5a",
          6157 => x"27",
          6158 => x"ac",
          6159 => x"18",
          6160 => x"39",
          6161 => x"70",
          6162 => x"58",
          6163 => x"b2",
          6164 => x"76",
          6165 => x"3f",
          6166 => x"08",
          6167 => x"f8",
          6168 => x"bd",
          6169 => x"82",
          6170 => x"27",
          6171 => x"16",
          6172 => x"f8",
          6173 => x"38",
          6174 => x"39",
          6175 => x"55",
          6176 => x"52",
          6177 => x"d5",
          6178 => x"f8",
          6179 => x"0c",
          6180 => x"0c",
          6181 => x"53",
          6182 => x"80",
          6183 => x"85",
          6184 => x"94",
          6185 => x"2a",
          6186 => x"0c",
          6187 => x"06",
          6188 => x"9c",
          6189 => x"58",
          6190 => x"f8",
          6191 => x"0d",
          6192 => x"0d",
          6193 => x"90",
          6194 => x"05",
          6195 => x"f0",
          6196 => x"27",
          6197 => x"0b",
          6198 => x"98",
          6199 => x"84",
          6200 => x"2e",
          6201 => x"76",
          6202 => x"58",
          6203 => x"38",
          6204 => x"15",
          6205 => x"08",
          6206 => x"38",
          6207 => x"88",
          6208 => x"53",
          6209 => x"81",
          6210 => x"c0",
          6211 => x"22",
          6212 => x"89",
          6213 => x"72",
          6214 => x"74",
          6215 => x"f3",
          6216 => x"d4",
          6217 => x"82",
          6218 => x"82",
          6219 => x"27",
          6220 => x"81",
          6221 => x"f8",
          6222 => x"80",
          6223 => x"16",
          6224 => x"f8",
          6225 => x"ca",
          6226 => x"38",
          6227 => x"0c",
          6228 => x"dd",
          6229 => x"08",
          6230 => x"f9",
          6231 => x"d4",
          6232 => x"87",
          6233 => x"f8",
          6234 => x"80",
          6235 => x"55",
          6236 => x"08",
          6237 => x"38",
          6238 => x"d4",
          6239 => x"2e",
          6240 => x"d4",
          6241 => x"75",
          6242 => x"3f",
          6243 => x"08",
          6244 => x"94",
          6245 => x"52",
          6246 => x"c1",
          6247 => x"f8",
          6248 => x"0c",
          6249 => x"0c",
          6250 => x"05",
          6251 => x"80",
          6252 => x"d4",
          6253 => x"3d",
          6254 => x"3d",
          6255 => x"71",
          6256 => x"57",
          6257 => x"51",
          6258 => x"82",
          6259 => x"54",
          6260 => x"08",
          6261 => x"82",
          6262 => x"56",
          6263 => x"52",
          6264 => x"83",
          6265 => x"f8",
          6266 => x"d4",
          6267 => x"d2",
          6268 => x"f8",
          6269 => x"08",
          6270 => x"54",
          6271 => x"e5",
          6272 => x"06",
          6273 => x"58",
          6274 => x"08",
          6275 => x"38",
          6276 => x"75",
          6277 => x"80",
          6278 => x"81",
          6279 => x"7a",
          6280 => x"06",
          6281 => x"39",
          6282 => x"08",
          6283 => x"76",
          6284 => x"3f",
          6285 => x"08",
          6286 => x"f8",
          6287 => x"ff",
          6288 => x"84",
          6289 => x"06",
          6290 => x"54",
          6291 => x"f8",
          6292 => x"0d",
          6293 => x"0d",
          6294 => x"52",
          6295 => x"3f",
          6296 => x"08",
          6297 => x"06",
          6298 => x"51",
          6299 => x"83",
          6300 => x"06",
          6301 => x"14",
          6302 => x"3f",
          6303 => x"08",
          6304 => x"07",
          6305 => x"d4",
          6306 => x"3d",
          6307 => x"3d",
          6308 => x"70",
          6309 => x"06",
          6310 => x"53",
          6311 => x"af",
          6312 => x"33",
          6313 => x"83",
          6314 => x"06",
          6315 => x"90",
          6316 => x"15",
          6317 => x"3f",
          6318 => x"04",
          6319 => x"75",
          6320 => x"8b",
          6321 => x"2a",
          6322 => x"29",
          6323 => x"81",
          6324 => x"71",
          6325 => x"ff",
          6326 => x"56",
          6327 => x"72",
          6328 => x"82",
          6329 => x"85",
          6330 => x"f2",
          6331 => x"62",
          6332 => x"79",
          6333 => x"81",
          6334 => x"5d",
          6335 => x"80",
          6336 => x"38",
          6337 => x"52",
          6338 => x"db",
          6339 => x"f8",
          6340 => x"d4",
          6341 => x"eb",
          6342 => x"08",
          6343 => x"55",
          6344 => x"84",
          6345 => x"39",
          6346 => x"bf",
          6347 => x"ff",
          6348 => x"72",
          6349 => x"82",
          6350 => x"56",
          6351 => x"2e",
          6352 => x"83",
          6353 => x"82",
          6354 => x"53",
          6355 => x"09",
          6356 => x"38",
          6357 => x"73",
          6358 => x"99",
          6359 => x"f8",
          6360 => x"06",
          6361 => x"88",
          6362 => x"06",
          6363 => x"56",
          6364 => x"87",
          6365 => x"5c",
          6366 => x"76",
          6367 => x"81",
          6368 => x"38",
          6369 => x"70",
          6370 => x"53",
          6371 => x"92",
          6372 => x"33",
          6373 => x"06",
          6374 => x"08",
          6375 => x"56",
          6376 => x"7c",
          6377 => x"06",
          6378 => x"8d",
          6379 => x"7c",
          6380 => x"81",
          6381 => x"38",
          6382 => x"9a",
          6383 => x"e8",
          6384 => x"d4",
          6385 => x"ff",
          6386 => x"72",
          6387 => x"74",
          6388 => x"bf",
          6389 => x"f3",
          6390 => x"81",
          6391 => x"82",
          6392 => x"33",
          6393 => x"e8",
          6394 => x"d4",
          6395 => x"ff",
          6396 => x"77",
          6397 => x"38",
          6398 => x"26",
          6399 => x"73",
          6400 => x"59",
          6401 => x"23",
          6402 => x"8b",
          6403 => x"ff",
          6404 => x"81",
          6405 => x"81",
          6406 => x"77",
          6407 => x"74",
          6408 => x"2a",
          6409 => x"51",
          6410 => x"80",
          6411 => x"73",
          6412 => x"92",
          6413 => x"1a",
          6414 => x"23",
          6415 => x"81",
          6416 => x"53",
          6417 => x"ff",
          6418 => x"9d",
          6419 => x"38",
          6420 => x"e8",
          6421 => x"f8",
          6422 => x"06",
          6423 => x"2e",
          6424 => x"0b",
          6425 => x"a0",
          6426 => x"78",
          6427 => x"3f",
          6428 => x"08",
          6429 => x"f8",
          6430 => x"98",
          6431 => x"84",
          6432 => x"80",
          6433 => x"0c",
          6434 => x"f8",
          6435 => x"0d",
          6436 => x"0d",
          6437 => x"40",
          6438 => x"78",
          6439 => x"3f",
          6440 => x"08",
          6441 => x"f8",
          6442 => x"38",
          6443 => x"5f",
          6444 => x"ac",
          6445 => x"19",
          6446 => x"51",
          6447 => x"82",
          6448 => x"58",
          6449 => x"08",
          6450 => x"9c",
          6451 => x"33",
          6452 => x"86",
          6453 => x"82",
          6454 => x"17",
          6455 => x"70",
          6456 => x"56",
          6457 => x"1a",
          6458 => x"e5",
          6459 => x"38",
          6460 => x"70",
          6461 => x"54",
          6462 => x"8e",
          6463 => x"b2",
          6464 => x"2e",
          6465 => x"81",
          6466 => x"19",
          6467 => x"2a",
          6468 => x"51",
          6469 => x"82",
          6470 => x"86",
          6471 => x"06",
          6472 => x"80",
          6473 => x"8d",
          6474 => x"81",
          6475 => x"90",
          6476 => x"1d",
          6477 => x"5e",
          6478 => x"09",
          6479 => x"b9",
          6480 => x"33",
          6481 => x"2e",
          6482 => x"81",
          6483 => x"1f",
          6484 => x"52",
          6485 => x"3f",
          6486 => x"08",
          6487 => x"06",
          6488 => x"95",
          6489 => x"70",
          6490 => x"29",
          6491 => x"56",
          6492 => x"5a",
          6493 => x"1b",
          6494 => x"51",
          6495 => x"82",
          6496 => x"83",
          6497 => x"56",
          6498 => x"b1",
          6499 => x"fe",
          6500 => x"38",
          6501 => x"df",
          6502 => x"d4",
          6503 => x"10",
          6504 => x"53",
          6505 => x"59",
          6506 => x"a1",
          6507 => x"d4",
          6508 => x"09",
          6509 => x"c1",
          6510 => x"8b",
          6511 => x"ff",
          6512 => x"81",
          6513 => x"81",
          6514 => x"7b",
          6515 => x"38",
          6516 => x"86",
          6517 => x"06",
          6518 => x"79",
          6519 => x"38",
          6520 => x"8b",
          6521 => x"1d",
          6522 => x"54",
          6523 => x"ff",
          6524 => x"ff",
          6525 => x"84",
          6526 => x"54",
          6527 => x"39",
          6528 => x"76",
          6529 => x"3f",
          6530 => x"08",
          6531 => x"54",
          6532 => x"bb",
          6533 => x"33",
          6534 => x"73",
          6535 => x"53",
          6536 => x"9c",
          6537 => x"e5",
          6538 => x"d4",
          6539 => x"2e",
          6540 => x"ff",
          6541 => x"ac",
          6542 => x"52",
          6543 => x"81",
          6544 => x"f8",
          6545 => x"d4",
          6546 => x"2e",
          6547 => x"77",
          6548 => x"0c",
          6549 => x"04",
          6550 => x"64",
          6551 => x"12",
          6552 => x"06",
          6553 => x"86",
          6554 => x"b5",
          6555 => x"1d",
          6556 => x"56",
          6557 => x"80",
          6558 => x"81",
          6559 => x"16",
          6560 => x"55",
          6561 => x"8c",
          6562 => x"70",
          6563 => x"70",
          6564 => x"e4",
          6565 => x"80",
          6566 => x"81",
          6567 => x"80",
          6568 => x"38",
          6569 => x"ab",
          6570 => x"5b",
          6571 => x"7b",
          6572 => x"53",
          6573 => x"51",
          6574 => x"85",
          6575 => x"c6",
          6576 => x"77",
          6577 => x"ff",
          6578 => x"55",
          6579 => x"b4",
          6580 => x"ff",
          6581 => x"19",
          6582 => x"57",
          6583 => x"76",
          6584 => x"81",
          6585 => x"2a",
          6586 => x"51",
          6587 => x"73",
          6588 => x"38",
          6589 => x"a1",
          6590 => x"17",
          6591 => x"25",
          6592 => x"39",
          6593 => x"02",
          6594 => x"05",
          6595 => x"b0",
          6596 => x"54",
          6597 => x"84",
          6598 => x"54",
          6599 => x"ff",
          6600 => x"76",
          6601 => x"58",
          6602 => x"38",
          6603 => x"05",
          6604 => x"fe",
          6605 => x"77",
          6606 => x"78",
          6607 => x"a0",
          6608 => x"74",
          6609 => x"52",
          6610 => x"3f",
          6611 => x"08",
          6612 => x"38",
          6613 => x"74",
          6614 => x"38",
          6615 => x"81",
          6616 => x"77",
          6617 => x"74",
          6618 => x"51",
          6619 => x"94",
          6620 => x"eb",
          6621 => x"15",
          6622 => x"58",
          6623 => x"87",
          6624 => x"81",
          6625 => x"70",
          6626 => x"57",
          6627 => x"87",
          6628 => x"38",
          6629 => x"f9",
          6630 => x"f8",
          6631 => x"81",
          6632 => x"e3",
          6633 => x"84",
          6634 => x"7a",
          6635 => x"82",
          6636 => x"d4",
          6637 => x"82",
          6638 => x"84",
          6639 => x"06",
          6640 => x"02",
          6641 => x"33",
          6642 => x"02",
          6643 => x"33",
          6644 => x"70",
          6645 => x"55",
          6646 => x"73",
          6647 => x"38",
          6648 => x"1d",
          6649 => x"c8",
          6650 => x"f8",
          6651 => x"78",
          6652 => x"f3",
          6653 => x"d4",
          6654 => x"82",
          6655 => x"82",
          6656 => x"19",
          6657 => x"2e",
          6658 => x"78",
          6659 => x"1b",
          6660 => x"53",
          6661 => x"ef",
          6662 => x"d4",
          6663 => x"82",
          6664 => x"81",
          6665 => x"1a",
          6666 => x"3f",
          6667 => x"08",
          6668 => x"5d",
          6669 => x"52",
          6670 => x"ab",
          6671 => x"f8",
          6672 => x"d4",
          6673 => x"d7",
          6674 => x"08",
          6675 => x"7a",
          6676 => x"5a",
          6677 => x"8d",
          6678 => x"0b",
          6679 => x"82",
          6680 => x"8c",
          6681 => x"d4",
          6682 => x"9a",
          6683 => x"df",
          6684 => x"29",
          6685 => x"55",
          6686 => x"ff",
          6687 => x"38",
          6688 => x"70",
          6689 => x"57",
          6690 => x"52",
          6691 => x"17",
          6692 => x"51",
          6693 => x"73",
          6694 => x"ff",
          6695 => x"17",
          6696 => x"27",
          6697 => x"83",
          6698 => x"8b",
          6699 => x"1b",
          6700 => x"54",
          6701 => x"77",
          6702 => x"58",
          6703 => x"81",
          6704 => x"34",
          6705 => x"51",
          6706 => x"82",
          6707 => x"57",
          6708 => x"08",
          6709 => x"ff",
          6710 => x"fe",
          6711 => x"1a",
          6712 => x"51",
          6713 => x"82",
          6714 => x"57",
          6715 => x"08",
          6716 => x"53",
          6717 => x"08",
          6718 => x"08",
          6719 => x"3f",
          6720 => x"1a",
          6721 => x"08",
          6722 => x"3f",
          6723 => x"ab",
          6724 => x"06",
          6725 => x"8c",
          6726 => x"0b",
          6727 => x"76",
          6728 => x"d4",
          6729 => x"3d",
          6730 => x"3d",
          6731 => x"08",
          6732 => x"ac",
          6733 => x"59",
          6734 => x"ff",
          6735 => x"72",
          6736 => x"ed",
          6737 => x"d4",
          6738 => x"82",
          6739 => x"80",
          6740 => x"15",
          6741 => x"51",
          6742 => x"82",
          6743 => x"54",
          6744 => x"08",
          6745 => x"15",
          6746 => x"73",
          6747 => x"83",
          6748 => x"15",
          6749 => x"a2",
          6750 => x"f8",
          6751 => x"51",
          6752 => x"82",
          6753 => x"54",
          6754 => x"08",
          6755 => x"38",
          6756 => x"09",
          6757 => x"38",
          6758 => x"82",
          6759 => x"88",
          6760 => x"f4",
          6761 => x"60",
          6762 => x"59",
          6763 => x"96",
          6764 => x"1c",
          6765 => x"83",
          6766 => x"1c",
          6767 => x"81",
          6768 => x"70",
          6769 => x"05",
          6770 => x"57",
          6771 => x"57",
          6772 => x"81",
          6773 => x"10",
          6774 => x"81",
          6775 => x"53",
          6776 => x"80",
          6777 => x"70",
          6778 => x"06",
          6779 => x"8f",
          6780 => x"38",
          6781 => x"df",
          6782 => x"96",
          6783 => x"79",
          6784 => x"54",
          6785 => x"7a",
          6786 => x"07",
          6787 => x"98",
          6788 => x"f8",
          6789 => x"ff",
          6790 => x"ff",
          6791 => x"38",
          6792 => x"a5",
          6793 => x"2a",
          6794 => x"34",
          6795 => x"34",
          6796 => x"39",
          6797 => x"30",
          6798 => x"80",
          6799 => x"25",
          6800 => x"54",
          6801 => x"85",
          6802 => x"9a",
          6803 => x"34",
          6804 => x"17",
          6805 => x"8c",
          6806 => x"10",
          6807 => x"51",
          6808 => x"fe",
          6809 => x"30",
          6810 => x"70",
          6811 => x"59",
          6812 => x"17",
          6813 => x"80",
          6814 => x"34",
          6815 => x"1a",
          6816 => x"9c",
          6817 => x"70",
          6818 => x"5b",
          6819 => x"a0",
          6820 => x"74",
          6821 => x"81",
          6822 => x"81",
          6823 => x"89",
          6824 => x"70",
          6825 => x"25",
          6826 => x"76",
          6827 => x"38",
          6828 => x"8b",
          6829 => x"70",
          6830 => x"34",
          6831 => x"74",
          6832 => x"05",
          6833 => x"17",
          6834 => x"27",
          6835 => x"77",
          6836 => x"53",
          6837 => x"14",
          6838 => x"33",
          6839 => x"87",
          6840 => x"38",
          6841 => x"19",
          6842 => x"80",
          6843 => x"73",
          6844 => x"55",
          6845 => x"80",
          6846 => x"38",
          6847 => x"19",
          6848 => x"33",
          6849 => x"54",
          6850 => x"26",
          6851 => x"1c",
          6852 => x"33",
          6853 => x"79",
          6854 => x"72",
          6855 => x"85",
          6856 => x"2a",
          6857 => x"06",
          6858 => x"2e",
          6859 => x"15",
          6860 => x"ff",
          6861 => x"74",
          6862 => x"05",
          6863 => x"19",
          6864 => x"19",
          6865 => x"59",
          6866 => x"ff",
          6867 => x"17",
          6868 => x"80",
          6869 => x"34",
          6870 => x"8c",
          6871 => x"53",
          6872 => x"72",
          6873 => x"9c",
          6874 => x"8b",
          6875 => x"19",
          6876 => x"08",
          6877 => x"53",
          6878 => x"82",
          6879 => x"78",
          6880 => x"51",
          6881 => x"82",
          6882 => x"86",
          6883 => x"13",
          6884 => x"3f",
          6885 => x"08",
          6886 => x"8e",
          6887 => x"f0",
          6888 => x"70",
          6889 => x"80",
          6890 => x"51",
          6891 => x"af",
          6892 => x"81",
          6893 => x"dc",
          6894 => x"74",
          6895 => x"38",
          6896 => x"08",
          6897 => x"aa",
          6898 => x"44",
          6899 => x"33",
          6900 => x"73",
          6901 => x"81",
          6902 => x"81",
          6903 => x"dc",
          6904 => x"70",
          6905 => x"07",
          6906 => x"73",
          6907 => x"88",
          6908 => x"70",
          6909 => x"73",
          6910 => x"38",
          6911 => x"ab",
          6912 => x"52",
          6913 => x"ee",
          6914 => x"f8",
          6915 => x"e1",
          6916 => x"7d",
          6917 => x"08",
          6918 => x"59",
          6919 => x"05",
          6920 => x"3f",
          6921 => x"08",
          6922 => x"b1",
          6923 => x"ff",
          6924 => x"f8",
          6925 => x"38",
          6926 => x"82",
          6927 => x"90",
          6928 => x"73",
          6929 => x"19",
          6930 => x"f8",
          6931 => x"ff",
          6932 => x"32",
          6933 => x"73",
          6934 => x"25",
          6935 => x"55",
          6936 => x"38",
          6937 => x"2e",
          6938 => x"80",
          6939 => x"38",
          6940 => x"c6",
          6941 => x"92",
          6942 => x"f8",
          6943 => x"38",
          6944 => x"26",
          6945 => x"78",
          6946 => x"75",
          6947 => x"19",
          6948 => x"39",
          6949 => x"80",
          6950 => x"56",
          6951 => x"af",
          6952 => x"06",
          6953 => x"57",
          6954 => x"32",
          6955 => x"80",
          6956 => x"51",
          6957 => x"dc",
          6958 => x"9f",
          6959 => x"2b",
          6960 => x"2e",
          6961 => x"8c",
          6962 => x"54",
          6963 => x"a5",
          6964 => x"39",
          6965 => x"09",
          6966 => x"c9",
          6967 => x"22",
          6968 => x"2e",
          6969 => x"80",
          6970 => x"22",
          6971 => x"2e",
          6972 => x"b6",
          6973 => x"1a",
          6974 => x"23",
          6975 => x"1f",
          6976 => x"54",
          6977 => x"83",
          6978 => x"73",
          6979 => x"05",
          6980 => x"18",
          6981 => x"27",
          6982 => x"a0",
          6983 => x"ab",
          6984 => x"c4",
          6985 => x"2e",
          6986 => x"10",
          6987 => x"55",
          6988 => x"16",
          6989 => x"32",
          6990 => x"9f",
          6991 => x"53",
          6992 => x"75",
          6993 => x"38",
          6994 => x"ff",
          6995 => x"e0",
          6996 => x"7a",
          6997 => x"80",
          6998 => x"8d",
          6999 => x"85",
          7000 => x"83",
          7001 => x"99",
          7002 => x"22",
          7003 => x"ff",
          7004 => x"5d",
          7005 => x"09",
          7006 => x"38",
          7007 => x"10",
          7008 => x"51",
          7009 => x"a0",
          7010 => x"7c",
          7011 => x"83",
          7012 => x"54",
          7013 => x"09",
          7014 => x"38",
          7015 => x"57",
          7016 => x"aa",
          7017 => x"fe",
          7018 => x"51",
          7019 => x"2e",
          7020 => x"10",
          7021 => x"55",
          7022 => x"78",
          7023 => x"38",
          7024 => x"22",
          7025 => x"ae",
          7026 => x"06",
          7027 => x"53",
          7028 => x"1e",
          7029 => x"3f",
          7030 => x"5c",
          7031 => x"10",
          7032 => x"81",
          7033 => x"54",
          7034 => x"82",
          7035 => x"a0",
          7036 => x"75",
          7037 => x"30",
          7038 => x"51",
          7039 => x"79",
          7040 => x"73",
          7041 => x"38",
          7042 => x"57",
          7043 => x"54",
          7044 => x"78",
          7045 => x"81",
          7046 => x"32",
          7047 => x"72",
          7048 => x"70",
          7049 => x"51",
          7050 => x"80",
          7051 => x"7e",
          7052 => x"ae",
          7053 => x"2e",
          7054 => x"83",
          7055 => x"79",
          7056 => x"38",
          7057 => x"58",
          7058 => x"2b",
          7059 => x"5d",
          7060 => x"39",
          7061 => x"27",
          7062 => x"82",
          7063 => x"b5",
          7064 => x"80",
          7065 => x"82",
          7066 => x"83",
          7067 => x"70",
          7068 => x"81",
          7069 => x"56",
          7070 => x"8c",
          7071 => x"ff",
          7072 => x"90",
          7073 => x"54",
          7074 => x"27",
          7075 => x"1f",
          7076 => x"26",
          7077 => x"83",
          7078 => x"57",
          7079 => x"7d",
          7080 => x"76",
          7081 => x"55",
          7082 => x"81",
          7083 => x"c3",
          7084 => x"2e",
          7085 => x"52",
          7086 => x"51",
          7087 => x"82",
          7088 => x"80",
          7089 => x"80",
          7090 => x"07",
          7091 => x"39",
          7092 => x"54",
          7093 => x"85",
          7094 => x"07",
          7095 => x"16",
          7096 => x"26",
          7097 => x"81",
          7098 => x"70",
          7099 => x"06",
          7100 => x"7d",
          7101 => x"54",
          7102 => x"81",
          7103 => x"de",
          7104 => x"33",
          7105 => x"e5",
          7106 => x"06",
          7107 => x"0b",
          7108 => x"7e",
          7109 => x"81",
          7110 => x"7b",
          7111 => x"fc",
          7112 => x"8c",
          7113 => x"8c",
          7114 => x"7b",
          7115 => x"73",
          7116 => x"81",
          7117 => x"76",
          7118 => x"76",
          7119 => x"81",
          7120 => x"73",
          7121 => x"81",
          7122 => x"80",
          7123 => x"76",
          7124 => x"7b",
          7125 => x"81",
          7126 => x"73",
          7127 => x"38",
          7128 => x"57",
          7129 => x"34",
          7130 => x"a5",
          7131 => x"f8",
          7132 => x"33",
          7133 => x"d4",
          7134 => x"2e",
          7135 => x"d4",
          7136 => x"2e",
          7137 => x"80",
          7138 => x"85",
          7139 => x"06",
          7140 => x"57",
          7141 => x"80",
          7142 => x"74",
          7143 => x"73",
          7144 => x"ed",
          7145 => x"0b",
          7146 => x"80",
          7147 => x"39",
          7148 => x"54",
          7149 => x"85",
          7150 => x"74",
          7151 => x"81",
          7152 => x"73",
          7153 => x"1e",
          7154 => x"2a",
          7155 => x"51",
          7156 => x"80",
          7157 => x"90",
          7158 => x"ff",
          7159 => x"b8",
          7160 => x"51",
          7161 => x"82",
          7162 => x"88",
          7163 => x"a1",
          7164 => x"d4",
          7165 => x"3d",
          7166 => x"3d",
          7167 => x"ff",
          7168 => x"71",
          7169 => x"5c",
          7170 => x"80",
          7171 => x"38",
          7172 => x"05",
          7173 => x"9f",
          7174 => x"71",
          7175 => x"38",
          7176 => x"71",
          7177 => x"81",
          7178 => x"38",
          7179 => x"11",
          7180 => x"06",
          7181 => x"70",
          7182 => x"38",
          7183 => x"81",
          7184 => x"05",
          7185 => x"76",
          7186 => x"38",
          7187 => x"c6",
          7188 => x"77",
          7189 => x"57",
          7190 => x"05",
          7191 => x"70",
          7192 => x"33",
          7193 => x"53",
          7194 => x"99",
          7195 => x"e0",
          7196 => x"ff",
          7197 => x"ff",
          7198 => x"70",
          7199 => x"38",
          7200 => x"81",
          7201 => x"51",
          7202 => x"9f",
          7203 => x"72",
          7204 => x"81",
          7205 => x"70",
          7206 => x"72",
          7207 => x"32",
          7208 => x"72",
          7209 => x"73",
          7210 => x"53",
          7211 => x"70",
          7212 => x"38",
          7213 => x"19",
          7214 => x"75",
          7215 => x"38",
          7216 => x"83",
          7217 => x"74",
          7218 => x"59",
          7219 => x"39",
          7220 => x"33",
          7221 => x"d4",
          7222 => x"3d",
          7223 => x"3d",
          7224 => x"80",
          7225 => x"34",
          7226 => x"17",
          7227 => x"75",
          7228 => x"3f",
          7229 => x"d4",
          7230 => x"80",
          7231 => x"16",
          7232 => x"3f",
          7233 => x"08",
          7234 => x"06",
          7235 => x"73",
          7236 => x"2e",
          7237 => x"80",
          7238 => x"0b",
          7239 => x"56",
          7240 => x"e9",
          7241 => x"06",
          7242 => x"57",
          7243 => x"32",
          7244 => x"80",
          7245 => x"51",
          7246 => x"8a",
          7247 => x"e8",
          7248 => x"06",
          7249 => x"53",
          7250 => x"52",
          7251 => x"51",
          7252 => x"82",
          7253 => x"55",
          7254 => x"08",
          7255 => x"38",
          7256 => x"c6",
          7257 => x"8a",
          7258 => x"ed",
          7259 => x"f8",
          7260 => x"d4",
          7261 => x"2e",
          7262 => x"55",
          7263 => x"f8",
          7264 => x"0d",
          7265 => x"0d",
          7266 => x"05",
          7267 => x"33",
          7268 => x"75",
          7269 => x"fc",
          7270 => x"d4",
          7271 => x"8b",
          7272 => x"82",
          7273 => x"24",
          7274 => x"82",
          7275 => x"84",
          7276 => x"c0",
          7277 => x"55",
          7278 => x"73",
          7279 => x"ee",
          7280 => x"0c",
          7281 => x"06",
          7282 => x"57",
          7283 => x"ae",
          7284 => x"33",
          7285 => x"3f",
          7286 => x"08",
          7287 => x"70",
          7288 => x"55",
          7289 => x"76",
          7290 => x"c0",
          7291 => x"2a",
          7292 => x"51",
          7293 => x"72",
          7294 => x"86",
          7295 => x"74",
          7296 => x"15",
          7297 => x"81",
          7298 => x"c6",
          7299 => x"d4",
          7300 => x"ff",
          7301 => x"06",
          7302 => x"56",
          7303 => x"38",
          7304 => x"8f",
          7305 => x"2a",
          7306 => x"51",
          7307 => x"72",
          7308 => x"80",
          7309 => x"52",
          7310 => x"3f",
          7311 => x"08",
          7312 => x"57",
          7313 => x"09",
          7314 => x"e2",
          7315 => x"74",
          7316 => x"56",
          7317 => x"33",
          7318 => x"72",
          7319 => x"38",
          7320 => x"51",
          7321 => x"82",
          7322 => x"57",
          7323 => x"84",
          7324 => x"ff",
          7325 => x"56",
          7326 => x"25",
          7327 => x"0b",
          7328 => x"56",
          7329 => x"05",
          7330 => x"83",
          7331 => x"2e",
          7332 => x"52",
          7333 => x"c6",
          7334 => x"f8",
          7335 => x"06",
          7336 => x"27",
          7337 => x"16",
          7338 => x"27",
          7339 => x"56",
          7340 => x"84",
          7341 => x"56",
          7342 => x"84",
          7343 => x"c3",
          7344 => x"c9",
          7345 => x"f8",
          7346 => x"ff",
          7347 => x"84",
          7348 => x"81",
          7349 => x"38",
          7350 => x"51",
          7351 => x"82",
          7352 => x"83",
          7353 => x"58",
          7354 => x"80",
          7355 => x"ca",
          7356 => x"d4",
          7357 => x"77",
          7358 => x"80",
          7359 => x"82",
          7360 => x"c8",
          7361 => x"11",
          7362 => x"06",
          7363 => x"8d",
          7364 => x"26",
          7365 => x"74",
          7366 => x"78",
          7367 => x"c5",
          7368 => x"59",
          7369 => x"15",
          7370 => x"2e",
          7371 => x"13",
          7372 => x"72",
          7373 => x"38",
          7374 => x"f2",
          7375 => x"14",
          7376 => x"3f",
          7377 => x"08",
          7378 => x"f8",
          7379 => x"23",
          7380 => x"57",
          7381 => x"83",
          7382 => x"cb",
          7383 => x"ad",
          7384 => x"f8",
          7385 => x"ff",
          7386 => x"8d",
          7387 => x"14",
          7388 => x"3f",
          7389 => x"08",
          7390 => x"14",
          7391 => x"3f",
          7392 => x"08",
          7393 => x"06",
          7394 => x"72",
          7395 => x"9e",
          7396 => x"22",
          7397 => x"84",
          7398 => x"5a",
          7399 => x"83",
          7400 => x"14",
          7401 => x"79",
          7402 => x"e1",
          7403 => x"d4",
          7404 => x"82",
          7405 => x"80",
          7406 => x"38",
          7407 => x"08",
          7408 => x"ff",
          7409 => x"38",
          7410 => x"83",
          7411 => x"83",
          7412 => x"74",
          7413 => x"85",
          7414 => x"89",
          7415 => x"76",
          7416 => x"ca",
          7417 => x"70",
          7418 => x"7b",
          7419 => x"73",
          7420 => x"17",
          7421 => x"b0",
          7422 => x"55",
          7423 => x"09",
          7424 => x"38",
          7425 => x"51",
          7426 => x"82",
          7427 => x"83",
          7428 => x"53",
          7429 => x"82",
          7430 => x"82",
          7431 => x"e4",
          7432 => x"80",
          7433 => x"f8",
          7434 => x"0c",
          7435 => x"53",
          7436 => x"56",
          7437 => x"81",
          7438 => x"13",
          7439 => x"74",
          7440 => x"82",
          7441 => x"74",
          7442 => x"81",
          7443 => x"06",
          7444 => x"83",
          7445 => x"2a",
          7446 => x"72",
          7447 => x"26",
          7448 => x"ff",
          7449 => x"0c",
          7450 => x"15",
          7451 => x"0b",
          7452 => x"76",
          7453 => x"81",
          7454 => x"38",
          7455 => x"51",
          7456 => x"82",
          7457 => x"83",
          7458 => x"53",
          7459 => x"09",
          7460 => x"f9",
          7461 => x"52",
          7462 => x"cb",
          7463 => x"f8",
          7464 => x"38",
          7465 => x"08",
          7466 => x"84",
          7467 => x"c6",
          7468 => x"d4",
          7469 => x"ff",
          7470 => x"72",
          7471 => x"2e",
          7472 => x"80",
          7473 => x"14",
          7474 => x"3f",
          7475 => x"08",
          7476 => x"a4",
          7477 => x"81",
          7478 => x"84",
          7479 => x"c6",
          7480 => x"d4",
          7481 => x"8a",
          7482 => x"2e",
          7483 => x"9d",
          7484 => x"14",
          7485 => x"3f",
          7486 => x"08",
          7487 => x"84",
          7488 => x"c6",
          7489 => x"d4",
          7490 => x"15",
          7491 => x"34",
          7492 => x"22",
          7493 => x"72",
          7494 => x"23",
          7495 => x"23",
          7496 => x"0b",
          7497 => x"80",
          7498 => x"0c",
          7499 => x"82",
          7500 => x"90",
          7501 => x"fb",
          7502 => x"54",
          7503 => x"80",
          7504 => x"73",
          7505 => x"80",
          7506 => x"72",
          7507 => x"80",
          7508 => x"86",
          7509 => x"15",
          7510 => x"71",
          7511 => x"81",
          7512 => x"81",
          7513 => x"ff",
          7514 => x"82",
          7515 => x"81",
          7516 => x"88",
          7517 => x"08",
          7518 => x"39",
          7519 => x"73",
          7520 => x"74",
          7521 => x"0c",
          7522 => x"04",
          7523 => x"02",
          7524 => x"7a",
          7525 => x"fc",
          7526 => x"f4",
          7527 => x"54",
          7528 => x"d4",
          7529 => x"bc",
          7530 => x"f8",
          7531 => x"82",
          7532 => x"70",
          7533 => x"73",
          7534 => x"38",
          7535 => x"78",
          7536 => x"2e",
          7537 => x"74",
          7538 => x"0c",
          7539 => x"80",
          7540 => x"80",
          7541 => x"70",
          7542 => x"51",
          7543 => x"82",
          7544 => x"54",
          7545 => x"f8",
          7546 => x"0d",
          7547 => x"0d",
          7548 => x"05",
          7549 => x"33",
          7550 => x"54",
          7551 => x"84",
          7552 => x"bf",
          7553 => x"99",
          7554 => x"53",
          7555 => x"05",
          7556 => x"f1",
          7557 => x"f8",
          7558 => x"d4",
          7559 => x"a4",
          7560 => x"69",
          7561 => x"70",
          7562 => x"f3",
          7563 => x"f8",
          7564 => x"d4",
          7565 => x"38",
          7566 => x"05",
          7567 => x"2b",
          7568 => x"80",
          7569 => x"86",
          7570 => x"06",
          7571 => x"2e",
          7572 => x"74",
          7573 => x"38",
          7574 => x"09",
          7575 => x"38",
          7576 => x"f4",
          7577 => x"f8",
          7578 => x"39",
          7579 => x"33",
          7580 => x"73",
          7581 => x"77",
          7582 => x"81",
          7583 => x"73",
          7584 => x"38",
          7585 => x"bc",
          7586 => x"07",
          7587 => x"b4",
          7588 => x"2a",
          7589 => x"51",
          7590 => x"2e",
          7591 => x"62",
          7592 => x"d7",
          7593 => x"d4",
          7594 => x"82",
          7595 => x"52",
          7596 => x"51",
          7597 => x"62",
          7598 => x"8b",
          7599 => x"53",
          7600 => x"51",
          7601 => x"80",
          7602 => x"05",
          7603 => x"3f",
          7604 => x"0b",
          7605 => x"75",
          7606 => x"f1",
          7607 => x"11",
          7608 => x"80",
          7609 => x"98",
          7610 => x"51",
          7611 => x"82",
          7612 => x"55",
          7613 => x"08",
          7614 => x"b7",
          7615 => x"c4",
          7616 => x"05",
          7617 => x"2a",
          7618 => x"51",
          7619 => x"80",
          7620 => x"84",
          7621 => x"39",
          7622 => x"70",
          7623 => x"54",
          7624 => x"a9",
          7625 => x"06",
          7626 => x"2e",
          7627 => x"55",
          7628 => x"73",
          7629 => x"c5",
          7630 => x"d4",
          7631 => x"ff",
          7632 => x"0c",
          7633 => x"d4",
          7634 => x"f8",
          7635 => x"2a",
          7636 => x"51",
          7637 => x"2e",
          7638 => x"80",
          7639 => x"7a",
          7640 => x"a0",
          7641 => x"a4",
          7642 => x"53",
          7643 => x"d5",
          7644 => x"d4",
          7645 => x"d4",
          7646 => x"1b",
          7647 => x"05",
          7648 => x"a0",
          7649 => x"f8",
          7650 => x"f8",
          7651 => x"0c",
          7652 => x"56",
          7653 => x"84",
          7654 => x"90",
          7655 => x"0b",
          7656 => x"80",
          7657 => x"0c",
          7658 => x"1a",
          7659 => x"2a",
          7660 => x"51",
          7661 => x"2e",
          7662 => x"82",
          7663 => x"80",
          7664 => x"38",
          7665 => x"08",
          7666 => x"8a",
          7667 => x"89",
          7668 => x"59",
          7669 => x"76",
          7670 => x"c6",
          7671 => x"d4",
          7672 => x"82",
          7673 => x"81",
          7674 => x"82",
          7675 => x"f8",
          7676 => x"09",
          7677 => x"38",
          7678 => x"78",
          7679 => x"30",
          7680 => x"80",
          7681 => x"77",
          7682 => x"38",
          7683 => x"06",
          7684 => x"c3",
          7685 => x"1a",
          7686 => x"38",
          7687 => x"06",
          7688 => x"2e",
          7689 => x"52",
          7690 => x"b1",
          7691 => x"f8",
          7692 => x"82",
          7693 => x"75",
          7694 => x"d4",
          7695 => x"9c",
          7696 => x"39",
          7697 => x"74",
          7698 => x"d4",
          7699 => x"3d",
          7700 => x"3d",
          7701 => x"65",
          7702 => x"5d",
          7703 => x"0c",
          7704 => x"05",
          7705 => x"f9",
          7706 => x"d4",
          7707 => x"82",
          7708 => x"8a",
          7709 => x"33",
          7710 => x"2e",
          7711 => x"56",
          7712 => x"90",
          7713 => x"06",
          7714 => x"74",
          7715 => x"b9",
          7716 => x"82",
          7717 => x"34",
          7718 => x"ad",
          7719 => x"91",
          7720 => x"56",
          7721 => x"8c",
          7722 => x"1a",
          7723 => x"74",
          7724 => x"38",
          7725 => x"80",
          7726 => x"38",
          7727 => x"70",
          7728 => x"56",
          7729 => x"b4",
          7730 => x"11",
          7731 => x"77",
          7732 => x"5b",
          7733 => x"38",
          7734 => x"88",
          7735 => x"8f",
          7736 => x"08",
          7737 => x"c4",
          7738 => x"d4",
          7739 => x"81",
          7740 => x"9f",
          7741 => x"2e",
          7742 => x"74",
          7743 => x"98",
          7744 => x"7e",
          7745 => x"3f",
          7746 => x"08",
          7747 => x"83",
          7748 => x"f8",
          7749 => x"89",
          7750 => x"77",
          7751 => x"d8",
          7752 => x"7f",
          7753 => x"58",
          7754 => x"75",
          7755 => x"75",
          7756 => x"77",
          7757 => x"7c",
          7758 => x"33",
          7759 => x"d4",
          7760 => x"f8",
          7761 => x"38",
          7762 => x"33",
          7763 => x"80",
          7764 => x"b4",
          7765 => x"31",
          7766 => x"27",
          7767 => x"80",
          7768 => x"52",
          7769 => x"77",
          7770 => x"7d",
          7771 => x"be",
          7772 => x"89",
          7773 => x"39",
          7774 => x"0c",
          7775 => x"83",
          7776 => x"80",
          7777 => x"55",
          7778 => x"83",
          7779 => x"9c",
          7780 => x"7e",
          7781 => x"3f",
          7782 => x"08",
          7783 => x"75",
          7784 => x"08",
          7785 => x"1f",
          7786 => x"7c",
          7787 => x"ec",
          7788 => x"31",
          7789 => x"7f",
          7790 => x"94",
          7791 => x"94",
          7792 => x"5c",
          7793 => x"80",
          7794 => x"d4",
          7795 => x"3d",
          7796 => x"3d",
          7797 => x"65",
          7798 => x"5d",
          7799 => x"0c",
          7800 => x"05",
          7801 => x"f6",
          7802 => x"d4",
          7803 => x"82",
          7804 => x"8a",
          7805 => x"33",
          7806 => x"2e",
          7807 => x"56",
          7808 => x"90",
          7809 => x"81",
          7810 => x"06",
          7811 => x"87",
          7812 => x"2e",
          7813 => x"95",
          7814 => x"91",
          7815 => x"56",
          7816 => x"81",
          7817 => x"34",
          7818 => x"94",
          7819 => x"08",
          7820 => x"56",
          7821 => x"84",
          7822 => x"5c",
          7823 => x"82",
          7824 => x"18",
          7825 => x"ff",
          7826 => x"74",
          7827 => x"7e",
          7828 => x"ff",
          7829 => x"2a",
          7830 => x"7a",
          7831 => x"8c",
          7832 => x"08",
          7833 => x"38",
          7834 => x"39",
          7835 => x"52",
          7836 => x"ef",
          7837 => x"f8",
          7838 => x"d4",
          7839 => x"2e",
          7840 => x"74",
          7841 => x"91",
          7842 => x"2e",
          7843 => x"74",
          7844 => x"88",
          7845 => x"38",
          7846 => x"0c",
          7847 => x"15",
          7848 => x"08",
          7849 => x"06",
          7850 => x"51",
          7851 => x"3f",
          7852 => x"08",
          7853 => x"98",
          7854 => x"7e",
          7855 => x"3f",
          7856 => x"08",
          7857 => x"d1",
          7858 => x"f8",
          7859 => x"89",
          7860 => x"78",
          7861 => x"d7",
          7862 => x"7f",
          7863 => x"58",
          7864 => x"75",
          7865 => x"75",
          7866 => x"78",
          7867 => x"7c",
          7868 => x"33",
          7869 => x"86",
          7870 => x"f8",
          7871 => x"38",
          7872 => x"08",
          7873 => x"56",
          7874 => x"9c",
          7875 => x"53",
          7876 => x"77",
          7877 => x"7d",
          7878 => x"16",
          7879 => x"fc",
          7880 => x"80",
          7881 => x"34",
          7882 => x"56",
          7883 => x"8c",
          7884 => x"19",
          7885 => x"38",
          7886 => x"bc",
          7887 => x"d4",
          7888 => x"df",
          7889 => x"b4",
          7890 => x"76",
          7891 => x"94",
          7892 => x"ff",
          7893 => x"71",
          7894 => x"7b",
          7895 => x"38",
          7896 => x"18",
          7897 => x"51",
          7898 => x"3f",
          7899 => x"08",
          7900 => x"75",
          7901 => x"94",
          7902 => x"ff",
          7903 => x"05",
          7904 => x"98",
          7905 => x"81",
          7906 => x"34",
          7907 => x"7e",
          7908 => x"0c",
          7909 => x"1a",
          7910 => x"94",
          7911 => x"1b",
          7912 => x"5e",
          7913 => x"27",
          7914 => x"55",
          7915 => x"0c",
          7916 => x"90",
          7917 => x"c0",
          7918 => x"90",
          7919 => x"56",
          7920 => x"f8",
          7921 => x"0d",
          7922 => x"0d",
          7923 => x"fc",
          7924 => x"52",
          7925 => x"3f",
          7926 => x"08",
          7927 => x"f8",
          7928 => x"38",
          7929 => x"70",
          7930 => x"81",
          7931 => x"55",
          7932 => x"80",
          7933 => x"16",
          7934 => x"51",
          7935 => x"3f",
          7936 => x"08",
          7937 => x"f8",
          7938 => x"38",
          7939 => x"8b",
          7940 => x"07",
          7941 => x"8b",
          7942 => x"16",
          7943 => x"52",
          7944 => x"cc",
          7945 => x"16",
          7946 => x"15",
          7947 => x"bd",
          7948 => x"b2",
          7949 => x"15",
          7950 => x"b1",
          7951 => x"92",
          7952 => x"b8",
          7953 => x"54",
          7954 => x"15",
          7955 => x"ff",
          7956 => x"82",
          7957 => x"90",
          7958 => x"bf",
          7959 => x"73",
          7960 => x"76",
          7961 => x"0c",
          7962 => x"04",
          7963 => x"76",
          7964 => x"fe",
          7965 => x"d4",
          7966 => x"82",
          7967 => x"9c",
          7968 => x"fc",
          7969 => x"51",
          7970 => x"82",
          7971 => x"53",
          7972 => x"08",
          7973 => x"d4",
          7974 => x"0c",
          7975 => x"f8",
          7976 => x"0d",
          7977 => x"0d",
          7978 => x"e6",
          7979 => x"52",
          7980 => x"d4",
          7981 => x"8b",
          7982 => x"f8",
          7983 => x"d4",
          7984 => x"71",
          7985 => x"0c",
          7986 => x"04",
          7987 => x"80",
          7988 => x"cc",
          7989 => x"3d",
          7990 => x"3f",
          7991 => x"08",
          7992 => x"f8",
          7993 => x"38",
          7994 => x"52",
          7995 => x"05",
          7996 => x"3f",
          7997 => x"08",
          7998 => x"f8",
          7999 => x"02",
          8000 => x"33",
          8001 => x"55",
          8002 => x"25",
          8003 => x"7a",
          8004 => x"54",
          8005 => x"a2",
          8006 => x"84",
          8007 => x"06",
          8008 => x"73",
          8009 => x"38",
          8010 => x"70",
          8011 => x"a5",
          8012 => x"f8",
          8013 => x"0c",
          8014 => x"d4",
          8015 => x"2e",
          8016 => x"83",
          8017 => x"74",
          8018 => x"0c",
          8019 => x"04",
          8020 => x"0d",
          8021 => x"08",
          8022 => x"08",
          8023 => x"7a",
          8024 => x"80",
          8025 => x"b4",
          8026 => x"e0",
          8027 => x"95",
          8028 => x"f8",
          8029 => x"d4",
          8030 => x"a1",
          8031 => x"d4",
          8032 => x"7c",
          8033 => x"80",
          8034 => x"55",
          8035 => x"3d",
          8036 => x"80",
          8037 => x"38",
          8038 => x"d3",
          8039 => x"55",
          8040 => x"82",
          8041 => x"57",
          8042 => x"08",
          8043 => x"80",
          8044 => x"52",
          8045 => x"b8",
          8046 => x"d4",
          8047 => x"82",
          8048 => x"82",
          8049 => x"da",
          8050 => x"7b",
          8051 => x"3f",
          8052 => x"08",
          8053 => x"0c",
          8054 => x"51",
          8055 => x"82",
          8056 => x"57",
          8057 => x"08",
          8058 => x"80",
          8059 => x"c9",
          8060 => x"d4",
          8061 => x"82",
          8062 => x"a7",
          8063 => x"3d",
          8064 => x"51",
          8065 => x"73",
          8066 => x"08",
          8067 => x"76",
          8068 => x"c5",
          8069 => x"d4",
          8070 => x"82",
          8071 => x"80",
          8072 => x"76",
          8073 => x"81",
          8074 => x"82",
          8075 => x"39",
          8076 => x"38",
          8077 => x"fd",
          8078 => x"74",
          8079 => x"3f",
          8080 => x"78",
          8081 => x"33",
          8082 => x"56",
          8083 => x"92",
          8084 => x"c6",
          8085 => x"16",
          8086 => x"33",
          8087 => x"73",
          8088 => x"16",
          8089 => x"26",
          8090 => x"75",
          8091 => x"38",
          8092 => x"05",
          8093 => x"80",
          8094 => x"11",
          8095 => x"18",
          8096 => x"58",
          8097 => x"34",
          8098 => x"ff",
          8099 => x"3d",
          8100 => x"58",
          8101 => x"fd",
          8102 => x"7b",
          8103 => x"06",
          8104 => x"18",
          8105 => x"08",
          8106 => x"af",
          8107 => x"0b",
          8108 => x"33",
          8109 => x"82",
          8110 => x"70",
          8111 => x"52",
          8112 => x"56",
          8113 => x"8d",
          8114 => x"70",
          8115 => x"51",
          8116 => x"f5",
          8117 => x"54",
          8118 => x"a7",
          8119 => x"74",
          8120 => x"38",
          8121 => x"73",
          8122 => x"81",
          8123 => x"81",
          8124 => x"39",
          8125 => x"81",
          8126 => x"74",
          8127 => x"81",
          8128 => x"91",
          8129 => x"80",
          8130 => x"18",
          8131 => x"54",
          8132 => x"70",
          8133 => x"34",
          8134 => x"eb",
          8135 => x"34",
          8136 => x"f8",
          8137 => x"3d",
          8138 => x"3d",
          8139 => x"8d",
          8140 => x"54",
          8141 => x"55",
          8142 => x"82",
          8143 => x"53",
          8144 => x"08",
          8145 => x"91",
          8146 => x"72",
          8147 => x"8c",
          8148 => x"73",
          8149 => x"38",
          8150 => x"70",
          8151 => x"81",
          8152 => x"57",
          8153 => x"73",
          8154 => x"08",
          8155 => x"94",
          8156 => x"75",
          8157 => x"9b",
          8158 => x"11",
          8159 => x"2b",
          8160 => x"73",
          8161 => x"38",
          8162 => x"16",
          8163 => x"a0",
          8164 => x"f8",
          8165 => x"78",
          8166 => x"55",
          8167 => x"90",
          8168 => x"f8",
          8169 => x"96",
          8170 => x"70",
          8171 => x"94",
          8172 => x"71",
          8173 => x"08",
          8174 => x"53",
          8175 => x"15",
          8176 => x"a7",
          8177 => x"74",
          8178 => x"97",
          8179 => x"f8",
          8180 => x"d4",
          8181 => x"2e",
          8182 => x"82",
          8183 => x"ff",
          8184 => x"38",
          8185 => x"08",
          8186 => x"73",
          8187 => x"73",
          8188 => x"9f",
          8189 => x"27",
          8190 => x"75",
          8191 => x"16",
          8192 => x"17",
          8193 => x"33",
          8194 => x"70",
          8195 => x"55",
          8196 => x"80",
          8197 => x"73",
          8198 => x"ff",
          8199 => x"82",
          8200 => x"54",
          8201 => x"08",
          8202 => x"d4",
          8203 => x"a8",
          8204 => x"74",
          8205 => x"cf",
          8206 => x"f8",
          8207 => x"ff",
          8208 => x"81",
          8209 => x"38",
          8210 => x"9c",
          8211 => x"a7",
          8212 => x"16",
          8213 => x"39",
          8214 => x"16",
          8215 => x"75",
          8216 => x"53",
          8217 => x"ab",
          8218 => x"79",
          8219 => x"ed",
          8220 => x"f8",
          8221 => x"82",
          8222 => x"34",
          8223 => x"c4",
          8224 => x"91",
          8225 => x"53",
          8226 => x"89",
          8227 => x"f8",
          8228 => x"94",
          8229 => x"8c",
          8230 => x"27",
          8231 => x"8c",
          8232 => x"15",
          8233 => x"07",
          8234 => x"16",
          8235 => x"ff",
          8236 => x"80",
          8237 => x"77",
          8238 => x"2e",
          8239 => x"9c",
          8240 => x"53",
          8241 => x"f8",
          8242 => x"0d",
          8243 => x"0d",
          8244 => x"54",
          8245 => x"81",
          8246 => x"53",
          8247 => x"05",
          8248 => x"84",
          8249 => x"9d",
          8250 => x"f8",
          8251 => x"d4",
          8252 => x"eb",
          8253 => x"0c",
          8254 => x"51",
          8255 => x"82",
          8256 => x"55",
          8257 => x"08",
          8258 => x"ab",
          8259 => x"98",
          8260 => x"80",
          8261 => x"38",
          8262 => x"70",
          8263 => x"81",
          8264 => x"57",
          8265 => x"ae",
          8266 => x"08",
          8267 => x"c2",
          8268 => x"d4",
          8269 => x"17",
          8270 => x"86",
          8271 => x"17",
          8272 => x"75",
          8273 => x"ae",
          8274 => x"f8",
          8275 => x"84",
          8276 => x"06",
          8277 => x"55",
          8278 => x"80",
          8279 => x"80",
          8280 => x"54",
          8281 => x"f8",
          8282 => x"0d",
          8283 => x"0d",
          8284 => x"fc",
          8285 => x"52",
          8286 => x"3f",
          8287 => x"08",
          8288 => x"d4",
          8289 => x"0c",
          8290 => x"04",
          8291 => x"77",
          8292 => x"fc",
          8293 => x"53",
          8294 => x"9b",
          8295 => x"f8",
          8296 => x"d4",
          8297 => x"e1",
          8298 => x"38",
          8299 => x"08",
          8300 => x"ff",
          8301 => x"82",
          8302 => x"53",
          8303 => x"82",
          8304 => x"52",
          8305 => x"a3",
          8306 => x"f8",
          8307 => x"d4",
          8308 => x"2e",
          8309 => x"85",
          8310 => x"87",
          8311 => x"f8",
          8312 => x"74",
          8313 => x"cf",
          8314 => x"52",
          8315 => x"bd",
          8316 => x"d4",
          8317 => x"32",
          8318 => x"72",
          8319 => x"70",
          8320 => x"08",
          8321 => x"54",
          8322 => x"d4",
          8323 => x"3d",
          8324 => x"3d",
          8325 => x"80",
          8326 => x"70",
          8327 => x"52",
          8328 => x"3f",
          8329 => x"08",
          8330 => x"f8",
          8331 => x"65",
          8332 => x"d2",
          8333 => x"d4",
          8334 => x"82",
          8335 => x"a0",
          8336 => x"cb",
          8337 => x"98",
          8338 => x"73",
          8339 => x"38",
          8340 => x"39",
          8341 => x"88",
          8342 => x"75",
          8343 => x"3f",
          8344 => x"f8",
          8345 => x"0d",
          8346 => x"0d",
          8347 => x"5c",
          8348 => x"3d",
          8349 => x"93",
          8350 => x"89",
          8351 => x"f8",
          8352 => x"d4",
          8353 => x"82",
          8354 => x"0c",
          8355 => x"11",
          8356 => x"94",
          8357 => x"56",
          8358 => x"74",
          8359 => x"75",
          8360 => x"e6",
          8361 => x"81",
          8362 => x"5b",
          8363 => x"82",
          8364 => x"75",
          8365 => x"73",
          8366 => x"81",
          8367 => x"38",
          8368 => x"57",
          8369 => x"3d",
          8370 => x"ff",
          8371 => x"82",
          8372 => x"ff",
          8373 => x"82",
          8374 => x"81",
          8375 => x"82",
          8376 => x"30",
          8377 => x"f8",
          8378 => x"25",
          8379 => x"19",
          8380 => x"5a",
          8381 => x"08",
          8382 => x"38",
          8383 => x"a8",
          8384 => x"d4",
          8385 => x"58",
          8386 => x"77",
          8387 => x"7d",
          8388 => x"ad",
          8389 => x"d4",
          8390 => x"82",
          8391 => x"80",
          8392 => x"70",
          8393 => x"ff",
          8394 => x"56",
          8395 => x"2e",
          8396 => x"9e",
          8397 => x"51",
          8398 => x"3f",
          8399 => x"08",
          8400 => x"06",
          8401 => x"80",
          8402 => x"19",
          8403 => x"54",
          8404 => x"14",
          8405 => x"cc",
          8406 => x"f8",
          8407 => x"06",
          8408 => x"80",
          8409 => x"19",
          8410 => x"54",
          8411 => x"06",
          8412 => x"79",
          8413 => x"78",
          8414 => x"79",
          8415 => x"84",
          8416 => x"07",
          8417 => x"84",
          8418 => x"82",
          8419 => x"92",
          8420 => x"f9",
          8421 => x"8a",
          8422 => x"53",
          8423 => x"e3",
          8424 => x"d4",
          8425 => x"82",
          8426 => x"81",
          8427 => x"17",
          8428 => x"81",
          8429 => x"17",
          8430 => x"2a",
          8431 => x"51",
          8432 => x"55",
          8433 => x"81",
          8434 => x"17",
          8435 => x"8c",
          8436 => x"81",
          8437 => x"9c",
          8438 => x"f8",
          8439 => x"17",
          8440 => x"51",
          8441 => x"3f",
          8442 => x"08",
          8443 => x"0c",
          8444 => x"39",
          8445 => x"52",
          8446 => x"ae",
          8447 => x"d4",
          8448 => x"2e",
          8449 => x"83",
          8450 => x"82",
          8451 => x"81",
          8452 => x"06",
          8453 => x"56",
          8454 => x"a1",
          8455 => x"82",
          8456 => x"9c",
          8457 => x"95",
          8458 => x"08",
          8459 => x"f8",
          8460 => x"51",
          8461 => x"3f",
          8462 => x"08",
          8463 => x"08",
          8464 => x"90",
          8465 => x"c0",
          8466 => x"90",
          8467 => x"80",
          8468 => x"75",
          8469 => x"75",
          8470 => x"d4",
          8471 => x"3d",
          8472 => x"3d",
          8473 => x"a2",
          8474 => x"05",
          8475 => x"51",
          8476 => x"82",
          8477 => x"55",
          8478 => x"08",
          8479 => x"78",
          8480 => x"08",
          8481 => x"70",
          8482 => x"93",
          8483 => x"f8",
          8484 => x"d4",
          8485 => x"df",
          8486 => x"ff",
          8487 => x"85",
          8488 => x"06",
          8489 => x"86",
          8490 => x"cb",
          8491 => x"2b",
          8492 => x"24",
          8493 => x"02",
          8494 => x"33",
          8495 => x"58",
          8496 => x"76",
          8497 => x"6c",
          8498 => x"ff",
          8499 => x"82",
          8500 => x"74",
          8501 => x"81",
          8502 => x"56",
          8503 => x"80",
          8504 => x"54",
          8505 => x"08",
          8506 => x"2e",
          8507 => x"73",
          8508 => x"f8",
          8509 => x"52",
          8510 => x"52",
          8511 => x"f6",
          8512 => x"f8",
          8513 => x"d4",
          8514 => x"eb",
          8515 => x"f8",
          8516 => x"51",
          8517 => x"3f",
          8518 => x"08",
          8519 => x"f8",
          8520 => x"87",
          8521 => x"39",
          8522 => x"08",
          8523 => x"38",
          8524 => x"08",
          8525 => x"77",
          8526 => x"3f",
          8527 => x"08",
          8528 => x"08",
          8529 => x"d4",
          8530 => x"80",
          8531 => x"55",
          8532 => x"95",
          8533 => x"2e",
          8534 => x"53",
          8535 => x"51",
          8536 => x"3f",
          8537 => x"08",
          8538 => x"38",
          8539 => x"a9",
          8540 => x"d4",
          8541 => x"74",
          8542 => x"0c",
          8543 => x"04",
          8544 => x"82",
          8545 => x"ff",
          8546 => x"9b",
          8547 => x"f5",
          8548 => x"f8",
          8549 => x"d4",
          8550 => x"b7",
          8551 => x"6a",
          8552 => x"70",
          8553 => x"f7",
          8554 => x"f8",
          8555 => x"d4",
          8556 => x"38",
          8557 => x"9b",
          8558 => x"f8",
          8559 => x"09",
          8560 => x"8f",
          8561 => x"df",
          8562 => x"85",
          8563 => x"51",
          8564 => x"74",
          8565 => x"78",
          8566 => x"8a",
          8567 => x"57",
          8568 => x"3f",
          8569 => x"08",
          8570 => x"82",
          8571 => x"83",
          8572 => x"82",
          8573 => x"81",
          8574 => x"06",
          8575 => x"54",
          8576 => x"08",
          8577 => x"81",
          8578 => x"81",
          8579 => x"39",
          8580 => x"38",
          8581 => x"08",
          8582 => x"ff",
          8583 => x"82",
          8584 => x"54",
          8585 => x"08",
          8586 => x"8b",
          8587 => x"b8",
          8588 => x"a5",
          8589 => x"54",
          8590 => x"15",
          8591 => x"90",
          8592 => x"15",
          8593 => x"b2",
          8594 => x"ce",
          8595 => x"a4",
          8596 => x"53",
          8597 => x"53",
          8598 => x"b2",
          8599 => x"78",
          8600 => x"80",
          8601 => x"ff",
          8602 => x"78",
          8603 => x"80",
          8604 => x"7f",
          8605 => x"d8",
          8606 => x"ff",
          8607 => x"78",
          8608 => x"83",
          8609 => x"51",
          8610 => x"3f",
          8611 => x"08",
          8612 => x"f8",
          8613 => x"82",
          8614 => x"52",
          8615 => x"51",
          8616 => x"3f",
          8617 => x"52",
          8618 => x"b7",
          8619 => x"54",
          8620 => x"15",
          8621 => x"81",
          8622 => x"34",
          8623 => x"a6",
          8624 => x"d4",
          8625 => x"8b",
          8626 => x"75",
          8627 => x"ff",
          8628 => x"73",
          8629 => x"0c",
          8630 => x"04",
          8631 => x"ab",
          8632 => x"51",
          8633 => x"82",
          8634 => x"fe",
          8635 => x"ab",
          8636 => x"91",
          8637 => x"f8",
          8638 => x"d4",
          8639 => x"d8",
          8640 => x"ab",
          8641 => x"9e",
          8642 => x"58",
          8643 => x"82",
          8644 => x"55",
          8645 => x"08",
          8646 => x"02",
          8647 => x"33",
          8648 => x"54",
          8649 => x"82",
          8650 => x"53",
          8651 => x"52",
          8652 => x"80",
          8653 => x"a2",
          8654 => x"53",
          8655 => x"3d",
          8656 => x"ff",
          8657 => x"ac",
          8658 => x"73",
          8659 => x"3f",
          8660 => x"08",
          8661 => x"f8",
          8662 => x"63",
          8663 => x"2e",
          8664 => x"88",
          8665 => x"3d",
          8666 => x"38",
          8667 => x"e8",
          8668 => x"f8",
          8669 => x"09",
          8670 => x"bb",
          8671 => x"ff",
          8672 => x"82",
          8673 => x"55",
          8674 => x"08",
          8675 => x"68",
          8676 => x"aa",
          8677 => x"05",
          8678 => x"51",
          8679 => x"3f",
          8680 => x"33",
          8681 => x"8b",
          8682 => x"84",
          8683 => x"06",
          8684 => x"73",
          8685 => x"a0",
          8686 => x"8b",
          8687 => x"54",
          8688 => x"15",
          8689 => x"33",
          8690 => x"70",
          8691 => x"55",
          8692 => x"2e",
          8693 => x"6f",
          8694 => x"e1",
          8695 => x"78",
          8696 => x"f1",
          8697 => x"f8",
          8698 => x"51",
          8699 => x"3f",
          8700 => x"d4",
          8701 => x"2e",
          8702 => x"82",
          8703 => x"52",
          8704 => x"a3",
          8705 => x"d4",
          8706 => x"80",
          8707 => x"58",
          8708 => x"f8",
          8709 => x"38",
          8710 => x"54",
          8711 => x"09",
          8712 => x"38",
          8713 => x"52",
          8714 => x"b4",
          8715 => x"54",
          8716 => x"15",
          8717 => x"82",
          8718 => x"9c",
          8719 => x"c1",
          8720 => x"d4",
          8721 => x"82",
          8722 => x"8c",
          8723 => x"ff",
          8724 => x"82",
          8725 => x"55",
          8726 => x"f8",
          8727 => x"0d",
          8728 => x"0d",
          8729 => x"05",
          8730 => x"05",
          8731 => x"33",
          8732 => x"53",
          8733 => x"05",
          8734 => x"51",
          8735 => x"82",
          8736 => x"55",
          8737 => x"08",
          8738 => x"78",
          8739 => x"96",
          8740 => x"51",
          8741 => x"82",
          8742 => x"55",
          8743 => x"08",
          8744 => x"80",
          8745 => x"81",
          8746 => x"86",
          8747 => x"38",
          8748 => x"61",
          8749 => x"12",
          8750 => x"7a",
          8751 => x"51",
          8752 => x"74",
          8753 => x"78",
          8754 => x"83",
          8755 => x"51",
          8756 => x"3f",
          8757 => x"08",
          8758 => x"d4",
          8759 => x"3d",
          8760 => x"3d",
          8761 => x"82",
          8762 => x"cc",
          8763 => x"3d",
          8764 => x"3f",
          8765 => x"08",
          8766 => x"f8",
          8767 => x"38",
          8768 => x"52",
          8769 => x"05",
          8770 => x"3f",
          8771 => x"08",
          8772 => x"f8",
          8773 => x"02",
          8774 => x"33",
          8775 => x"54",
          8776 => x"a6",
          8777 => x"22",
          8778 => x"71",
          8779 => x"53",
          8780 => x"51",
          8781 => x"3f",
          8782 => x"0b",
          8783 => x"76",
          8784 => x"ea",
          8785 => x"f8",
          8786 => x"82",
          8787 => x"94",
          8788 => x"e9",
          8789 => x"6c",
          8790 => x"53",
          8791 => x"05",
          8792 => x"51",
          8793 => x"82",
          8794 => x"82",
          8795 => x"30",
          8796 => x"f8",
          8797 => x"25",
          8798 => x"79",
          8799 => x"86",
          8800 => x"75",
          8801 => x"73",
          8802 => x"fa",
          8803 => x"80",
          8804 => x"8d",
          8805 => x"54",
          8806 => x"3f",
          8807 => x"08",
          8808 => x"f8",
          8809 => x"38",
          8810 => x"51",
          8811 => x"3f",
          8812 => x"08",
          8813 => x"f8",
          8814 => x"82",
          8815 => x"82",
          8816 => x"65",
          8817 => x"78",
          8818 => x"7b",
          8819 => x"55",
          8820 => x"34",
          8821 => x"8a",
          8822 => x"38",
          8823 => x"1a",
          8824 => x"34",
          8825 => x"9e",
          8826 => x"70",
          8827 => x"51",
          8828 => x"a0",
          8829 => x"8e",
          8830 => x"2e",
          8831 => x"86",
          8832 => x"34",
          8833 => x"30",
          8834 => x"80",
          8835 => x"7a",
          8836 => x"c1",
          8837 => x"2e",
          8838 => x"a4",
          8839 => x"51",
          8840 => x"3f",
          8841 => x"08",
          8842 => x"f8",
          8843 => x"7b",
          8844 => x"55",
          8845 => x"73",
          8846 => x"38",
          8847 => x"73",
          8848 => x"38",
          8849 => x"15",
          8850 => x"ff",
          8851 => x"82",
          8852 => x"7b",
          8853 => x"d4",
          8854 => x"3d",
          8855 => x"3d",
          8856 => x"9c",
          8857 => x"05",
          8858 => x"51",
          8859 => x"82",
          8860 => x"82",
          8861 => x"56",
          8862 => x"f8",
          8863 => x"38",
          8864 => x"52",
          8865 => x"52",
          8866 => x"b3",
          8867 => x"70",
          8868 => x"56",
          8869 => x"81",
          8870 => x"57",
          8871 => x"ff",
          8872 => x"82",
          8873 => x"83",
          8874 => x"80",
          8875 => x"d4",
          8876 => x"95",
          8877 => x"b5",
          8878 => x"f8",
          8879 => x"e8",
          8880 => x"f8",
          8881 => x"ff",
          8882 => x"80",
          8883 => x"74",
          8884 => x"90",
          8885 => x"b2",
          8886 => x"f8",
          8887 => x"81",
          8888 => x"88",
          8889 => x"26",
          8890 => x"39",
          8891 => x"86",
          8892 => x"81",
          8893 => x"ff",
          8894 => x"38",
          8895 => x"54",
          8896 => x"81",
          8897 => x"81",
          8898 => x"77",
          8899 => x"59",
          8900 => x"6d",
          8901 => x"55",
          8902 => x"26",
          8903 => x"8a",
          8904 => x"86",
          8905 => x"e5",
          8906 => x"38",
          8907 => x"99",
          8908 => x"05",
          8909 => x"70",
          8910 => x"73",
          8911 => x"81",
          8912 => x"ff",
          8913 => x"ed",
          8914 => x"80",
          8915 => x"90",
          8916 => x"55",
          8917 => x"3f",
          8918 => x"08",
          8919 => x"f8",
          8920 => x"38",
          8921 => x"51",
          8922 => x"3f",
          8923 => x"08",
          8924 => x"f8",
          8925 => x"75",
          8926 => x"66",
          8927 => x"34",
          8928 => x"82",
          8929 => x"84",
          8930 => x"06",
          8931 => x"80",
          8932 => x"2e",
          8933 => x"81",
          8934 => x"ff",
          8935 => x"82",
          8936 => x"54",
          8937 => x"08",
          8938 => x"53",
          8939 => x"08",
          8940 => x"ff",
          8941 => x"66",
          8942 => x"8b",
          8943 => x"53",
          8944 => x"51",
          8945 => x"3f",
          8946 => x"0b",
          8947 => x"78",
          8948 => x"da",
          8949 => x"f8",
          8950 => x"55",
          8951 => x"f8",
          8952 => x"0d",
          8953 => x"0d",
          8954 => x"88",
          8955 => x"05",
          8956 => x"fc",
          8957 => x"54",
          8958 => x"d2",
          8959 => x"d4",
          8960 => x"82",
          8961 => x"82",
          8962 => x"1a",
          8963 => x"82",
          8964 => x"80",
          8965 => x"8c",
          8966 => x"78",
          8967 => x"1a",
          8968 => x"2a",
          8969 => x"51",
          8970 => x"90",
          8971 => x"82",
          8972 => x"58",
          8973 => x"81",
          8974 => x"39",
          8975 => x"22",
          8976 => x"70",
          8977 => x"56",
          8978 => x"af",
          8979 => x"14",
          8980 => x"30",
          8981 => x"9f",
          8982 => x"f8",
          8983 => x"19",
          8984 => x"5a",
          8985 => x"81",
          8986 => x"38",
          8987 => x"77",
          8988 => x"82",
          8989 => x"56",
          8990 => x"74",
          8991 => x"ff",
          8992 => x"81",
          8993 => x"55",
          8994 => x"75",
          8995 => x"82",
          8996 => x"f8",
          8997 => x"ff",
          8998 => x"d4",
          8999 => x"2e",
          9000 => x"82",
          9001 => x"8e",
          9002 => x"56",
          9003 => x"09",
          9004 => x"38",
          9005 => x"59",
          9006 => x"77",
          9007 => x"06",
          9008 => x"87",
          9009 => x"39",
          9010 => x"ba",
          9011 => x"55",
          9012 => x"2e",
          9013 => x"15",
          9014 => x"2e",
          9015 => x"83",
          9016 => x"75",
          9017 => x"7e",
          9018 => x"94",
          9019 => x"f8",
          9020 => x"d4",
          9021 => x"ce",
          9022 => x"16",
          9023 => x"56",
          9024 => x"38",
          9025 => x"19",
          9026 => x"90",
          9027 => x"7d",
          9028 => x"38",
          9029 => x"0c",
          9030 => x"0c",
          9031 => x"80",
          9032 => x"73",
          9033 => x"9c",
          9034 => x"05",
          9035 => x"57",
          9036 => x"26",
          9037 => x"7b",
          9038 => x"0c",
          9039 => x"81",
          9040 => x"84",
          9041 => x"54",
          9042 => x"f8",
          9043 => x"0d",
          9044 => x"0d",
          9045 => x"88",
          9046 => x"05",
          9047 => x"54",
          9048 => x"c5",
          9049 => x"56",
          9050 => x"d4",
          9051 => x"8b",
          9052 => x"d4",
          9053 => x"29",
          9054 => x"05",
          9055 => x"55",
          9056 => x"84",
          9057 => x"34",
          9058 => x"08",
          9059 => x"5f",
          9060 => x"51",
          9061 => x"3f",
          9062 => x"08",
          9063 => x"70",
          9064 => x"57",
          9065 => x"8b",
          9066 => x"82",
          9067 => x"06",
          9068 => x"56",
          9069 => x"38",
          9070 => x"05",
          9071 => x"7e",
          9072 => x"9e",
          9073 => x"f8",
          9074 => x"67",
          9075 => x"2e",
          9076 => x"82",
          9077 => x"8b",
          9078 => x"75",
          9079 => x"80",
          9080 => x"81",
          9081 => x"2e",
          9082 => x"80",
          9083 => x"38",
          9084 => x"0a",
          9085 => x"ff",
          9086 => x"55",
          9087 => x"86",
          9088 => x"8a",
          9089 => x"89",
          9090 => x"2a",
          9091 => x"77",
          9092 => x"59",
          9093 => x"81",
          9094 => x"70",
          9095 => x"07",
          9096 => x"56",
          9097 => x"38",
          9098 => x"05",
          9099 => x"7e",
          9100 => x"ae",
          9101 => x"82",
          9102 => x"8a",
          9103 => x"83",
          9104 => x"06",
          9105 => x"08",
          9106 => x"74",
          9107 => x"41",
          9108 => x"56",
          9109 => x"8a",
          9110 => x"61",
          9111 => x"55",
          9112 => x"27",
          9113 => x"93",
          9114 => x"80",
          9115 => x"38",
          9116 => x"70",
          9117 => x"43",
          9118 => x"95",
          9119 => x"06",
          9120 => x"2e",
          9121 => x"77",
          9122 => x"74",
          9123 => x"83",
          9124 => x"06",
          9125 => x"82",
          9126 => x"2e",
          9127 => x"78",
          9128 => x"2e",
          9129 => x"80",
          9130 => x"ae",
          9131 => x"2a",
          9132 => x"82",
          9133 => x"56",
          9134 => x"2e",
          9135 => x"77",
          9136 => x"82",
          9137 => x"79",
          9138 => x"70",
          9139 => x"5a",
          9140 => x"86",
          9141 => x"27",
          9142 => x"52",
          9143 => x"aa",
          9144 => x"d4",
          9145 => x"29",
          9146 => x"70",
          9147 => x"55",
          9148 => x"0b",
          9149 => x"08",
          9150 => x"05",
          9151 => x"ff",
          9152 => x"27",
          9153 => x"88",
          9154 => x"ae",
          9155 => x"2a",
          9156 => x"82",
          9157 => x"56",
          9158 => x"2e",
          9159 => x"77",
          9160 => x"82",
          9161 => x"79",
          9162 => x"70",
          9163 => x"5a",
          9164 => x"86",
          9165 => x"27",
          9166 => x"52",
          9167 => x"a9",
          9168 => x"d4",
          9169 => x"84",
          9170 => x"d4",
          9171 => x"f5",
          9172 => x"81",
          9173 => x"f8",
          9174 => x"d4",
          9175 => x"71",
          9176 => x"83",
          9177 => x"5e",
          9178 => x"89",
          9179 => x"5c",
          9180 => x"1c",
          9181 => x"05",
          9182 => x"ff",
          9183 => x"70",
          9184 => x"31",
          9185 => x"57",
          9186 => x"83",
          9187 => x"06",
          9188 => x"1c",
          9189 => x"5c",
          9190 => x"1d",
          9191 => x"29",
          9192 => x"31",
          9193 => x"55",
          9194 => x"87",
          9195 => x"7c",
          9196 => x"7a",
          9197 => x"31",
          9198 => x"a8",
          9199 => x"d4",
          9200 => x"7d",
          9201 => x"81",
          9202 => x"82",
          9203 => x"83",
          9204 => x"80",
          9205 => x"87",
          9206 => x"81",
          9207 => x"fd",
          9208 => x"f8",
          9209 => x"2e",
          9210 => x"80",
          9211 => x"ff",
          9212 => x"d4",
          9213 => x"a0",
          9214 => x"38",
          9215 => x"74",
          9216 => x"86",
          9217 => x"fd",
          9218 => x"81",
          9219 => x"80",
          9220 => x"83",
          9221 => x"39",
          9222 => x"08",
          9223 => x"92",
          9224 => x"b8",
          9225 => x"59",
          9226 => x"27",
          9227 => x"86",
          9228 => x"55",
          9229 => x"09",
          9230 => x"38",
          9231 => x"f5",
          9232 => x"38",
          9233 => x"55",
          9234 => x"86",
          9235 => x"80",
          9236 => x"7a",
          9237 => x"e7",
          9238 => x"82",
          9239 => x"7a",
          9240 => x"b8",
          9241 => x"52",
          9242 => x"ff",
          9243 => x"79",
          9244 => x"7b",
          9245 => x"06",
          9246 => x"51",
          9247 => x"3f",
          9248 => x"1c",
          9249 => x"32",
          9250 => x"96",
          9251 => x"06",
          9252 => x"91",
          9253 => x"8f",
          9254 => x"55",
          9255 => x"ff",
          9256 => x"74",
          9257 => x"06",
          9258 => x"51",
          9259 => x"3f",
          9260 => x"52",
          9261 => x"ff",
          9262 => x"f8",
          9263 => x"34",
          9264 => x"1b",
          9265 => x"87",
          9266 => x"52",
          9267 => x"ff",
          9268 => x"60",
          9269 => x"51",
          9270 => x"3f",
          9271 => x"09",
          9272 => x"cb",
          9273 => x"b2",
          9274 => x"c3",
          9275 => x"8e",
          9276 => x"52",
          9277 => x"ff",
          9278 => x"82",
          9279 => x"51",
          9280 => x"3f",
          9281 => x"1b",
          9282 => x"c3",
          9283 => x"b2",
          9284 => x"8e",
          9285 => x"80",
          9286 => x"1c",
          9287 => x"80",
          9288 => x"93",
          9289 => x"c8",
          9290 => x"1b",
          9291 => x"82",
          9292 => x"52",
          9293 => x"ff",
          9294 => x"7c",
          9295 => x"06",
          9296 => x"51",
          9297 => x"3f",
          9298 => x"a4",
          9299 => x"0b",
          9300 => x"93",
          9301 => x"dc",
          9302 => x"51",
          9303 => x"3f",
          9304 => x"52",
          9305 => x"70",
          9306 => x"8d",
          9307 => x"54",
          9308 => x"52",
          9309 => x"8a",
          9310 => x"56",
          9311 => x"08",
          9312 => x"7d",
          9313 => x"81",
          9314 => x"38",
          9315 => x"86",
          9316 => x"52",
          9317 => x"89",
          9318 => x"80",
          9319 => x"7a",
          9320 => x"9b",
          9321 => x"85",
          9322 => x"7a",
          9323 => x"bd",
          9324 => x"85",
          9325 => x"83",
          9326 => x"ff",
          9327 => x"ff",
          9328 => x"e8",
          9329 => x"8d",
          9330 => x"52",
          9331 => x"51",
          9332 => x"3f",
          9333 => x"52",
          9334 => x"8c",
          9335 => x"54",
          9336 => x"53",
          9337 => x"51",
          9338 => x"3f",
          9339 => x"16",
          9340 => x"7e",
          9341 => x"86",
          9342 => x"80",
          9343 => x"ff",
          9344 => x"7f",
          9345 => x"7d",
          9346 => x"81",
          9347 => x"f8",
          9348 => x"ff",
          9349 => x"ff",
          9350 => x"51",
          9351 => x"3f",
          9352 => x"88",
          9353 => x"39",
          9354 => x"f8",
          9355 => x"2e",
          9356 => x"55",
          9357 => x"51",
          9358 => x"3f",
          9359 => x"57",
          9360 => x"83",
          9361 => x"76",
          9362 => x"7a",
          9363 => x"ff",
          9364 => x"82",
          9365 => x"82",
          9366 => x"80",
          9367 => x"f8",
          9368 => x"51",
          9369 => x"3f",
          9370 => x"78",
          9371 => x"74",
          9372 => x"18",
          9373 => x"2e",
          9374 => x"79",
          9375 => x"2e",
          9376 => x"55",
          9377 => x"62",
          9378 => x"74",
          9379 => x"75",
          9380 => x"7e",
          9381 => x"e6",
          9382 => x"f8",
          9383 => x"38",
          9384 => x"78",
          9385 => x"74",
          9386 => x"56",
          9387 => x"93",
          9388 => x"66",
          9389 => x"26",
          9390 => x"56",
          9391 => x"83",
          9392 => x"64",
          9393 => x"77",
          9394 => x"84",
          9395 => x"52",
          9396 => x"8b",
          9397 => x"d4",
          9398 => x"51",
          9399 => x"3f",
          9400 => x"55",
          9401 => x"81",
          9402 => x"34",
          9403 => x"16",
          9404 => x"16",
          9405 => x"16",
          9406 => x"05",
          9407 => x"c1",
          9408 => x"fe",
          9409 => x"fe",
          9410 => x"34",
          9411 => x"08",
          9412 => x"07",
          9413 => x"16",
          9414 => x"f8",
          9415 => x"34",
          9416 => x"c6",
          9417 => x"8a",
          9418 => x"52",
          9419 => x"51",
          9420 => x"3f",
          9421 => x"53",
          9422 => x"51",
          9423 => x"3f",
          9424 => x"d4",
          9425 => x"38",
          9426 => x"52",
          9427 => x"88",
          9428 => x"56",
          9429 => x"08",
          9430 => x"39",
          9431 => x"39",
          9432 => x"39",
          9433 => x"08",
          9434 => x"d4",
          9435 => x"3d",
          9436 => x"3d",
          9437 => x"5b",
          9438 => x"60",
          9439 => x"57",
          9440 => x"25",
          9441 => x"3d",
          9442 => x"55",
          9443 => x"15",
          9444 => x"c9",
          9445 => x"81",
          9446 => x"06",
          9447 => x"3d",
          9448 => x"8d",
          9449 => x"74",
          9450 => x"05",
          9451 => x"17",
          9452 => x"2e",
          9453 => x"c9",
          9454 => x"34",
          9455 => x"83",
          9456 => x"74",
          9457 => x"0c",
          9458 => x"04",
          9459 => x"7b",
          9460 => x"b3",
          9461 => x"57",
          9462 => x"09",
          9463 => x"38",
          9464 => x"51",
          9465 => x"17",
          9466 => x"76",
          9467 => x"88",
          9468 => x"17",
          9469 => x"59",
          9470 => x"81",
          9471 => x"76",
          9472 => x"8b",
          9473 => x"54",
          9474 => x"17",
          9475 => x"51",
          9476 => x"79",
          9477 => x"30",
          9478 => x"9f",
          9479 => x"53",
          9480 => x"75",
          9481 => x"81",
          9482 => x"0c",
          9483 => x"04",
          9484 => x"79",
          9485 => x"56",
          9486 => x"24",
          9487 => x"3d",
          9488 => x"74",
          9489 => x"52",
          9490 => x"cb",
          9491 => x"d4",
          9492 => x"38",
          9493 => x"78",
          9494 => x"06",
          9495 => x"16",
          9496 => x"39",
          9497 => x"82",
          9498 => x"89",
          9499 => x"fd",
          9500 => x"54",
          9501 => x"80",
          9502 => x"ff",
          9503 => x"76",
          9504 => x"3d",
          9505 => x"3d",
          9506 => x"e3",
          9507 => x"53",
          9508 => x"53",
          9509 => x"3f",
          9510 => x"51",
          9511 => x"72",
          9512 => x"3f",
          9513 => x"04",
          9514 => x"75",
          9515 => x"9a",
          9516 => x"53",
          9517 => x"80",
          9518 => x"38",
          9519 => x"ff",
          9520 => x"c3",
          9521 => x"ff",
          9522 => x"73",
          9523 => x"09",
          9524 => x"38",
          9525 => x"af",
          9526 => x"c4",
          9527 => x"71",
          9528 => x"81",
          9529 => x"ff",
          9530 => x"51",
          9531 => x"26",
          9532 => x"10",
          9533 => x"05",
          9534 => x"51",
          9535 => x"80",
          9536 => x"ff",
          9537 => x"71",
          9538 => x"0c",
          9539 => x"04",
          9540 => x"02",
          9541 => x"02",
          9542 => x"05",
          9543 => x"80",
          9544 => x"ff",
          9545 => x"70",
          9546 => x"71",
          9547 => x"09",
          9548 => x"38",
          9549 => x"26",
          9550 => x"10",
          9551 => x"05",
          9552 => x"51",
          9553 => x"f8",
          9554 => x"0d",
          9555 => x"0d",
          9556 => x"83",
          9557 => x"81",
          9558 => x"83",
          9559 => x"82",
          9560 => x"52",
          9561 => x"27",
          9562 => x"ce",
          9563 => x"70",
          9564 => x"22",
          9565 => x"80",
          9566 => x"26",
          9567 => x"55",
          9568 => x"38",
          9569 => x"05",
          9570 => x"88",
          9571 => x"ff",
          9572 => x"54",
          9573 => x"71",
          9574 => x"d7",
          9575 => x"26",
          9576 => x"73",
          9577 => x"ad",
          9578 => x"70",
          9579 => x"75",
          9580 => x"11",
          9581 => x"51",
          9582 => x"39",
          9583 => x"81",
          9584 => x"31",
          9585 => x"39",
          9586 => x"9f",
          9587 => x"51",
          9588 => x"12",
          9589 => x"e6",
          9590 => x"39",
          9591 => x"8b",
          9592 => x"12",
          9593 => x"c7",
          9594 => x"70",
          9595 => x"06",
          9596 => x"73",
          9597 => x"72",
          9598 => x"fe",
          9599 => x"51",
          9600 => x"f8",
          9601 => x"0d",
          9602 => x"ff",
          9603 => x"00",
          9604 => x"ff",
          9605 => x"ff",
          9606 => x"00",
          9607 => x"00",
          9608 => x"00",
          9609 => x"00",
          9610 => x"00",
          9611 => x"00",
          9612 => x"00",
          9613 => x"00",
          9614 => x"00",
          9615 => x"00",
          9616 => x"00",
          9617 => x"00",
          9618 => x"00",
          9619 => x"00",
          9620 => x"00",
          9621 => x"00",
          9622 => x"00",
          9623 => x"00",
          9624 => x"00",
          9625 => x"00",
          9626 => x"00",
          9627 => x"00",
          9628 => x"00",
          9629 => x"00",
          9630 => x"00",
          9631 => x"00",
          9632 => x"00",
          9633 => x"00",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"00",
          9638 => x"00",
          9639 => x"00",
          9640 => x"00",
          9641 => x"00",
          9642 => x"00",
          9643 => x"00",
          9644 => x"00",
          9645 => x"00",
          9646 => x"00",
          9647 => x"00",
          9648 => x"00",
          9649 => x"00",
          9650 => x"00",
          9651 => x"00",
          9652 => x"00",
          9653 => x"00",
          9654 => x"00",
          9655 => x"00",
          9656 => x"00",
          9657 => x"00",
          9658 => x"00",
          9659 => x"00",
          9660 => x"00",
          9661 => x"00",
          9662 => x"00",
          9663 => x"00",
          9664 => x"00",
          9665 => x"00",
          9666 => x"00",
          9667 => x"00",
          9668 => x"00",
          9669 => x"00",
          9670 => x"00",
          9671 => x"00",
          9672 => x"00",
          9673 => x"00",
          9674 => x"00",
          9675 => x"00",
          9676 => x"00",
          9677 => x"00",
          9678 => x"00",
          9679 => x"00",
          9680 => x"00",
          9681 => x"00",
          9682 => x"00",
          9683 => x"00",
          9684 => x"00",
          9685 => x"00",
          9686 => x"00",
          9687 => x"00",
          9688 => x"00",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"00",
          9693 => x"00",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"00",
          9721 => x"00",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"00",
          9726 => x"00",
          9727 => x"00",
          9728 => x"00",
          9729 => x"00",
          9730 => x"00",
          9731 => x"00",
          9732 => x"00",
          9733 => x"00",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"69",
          9752 => x"00",
          9753 => x"69",
          9754 => x"6c",
          9755 => x"69",
          9756 => x"00",
          9757 => x"6c",
          9758 => x"00",
          9759 => x"65",
          9760 => x"00",
          9761 => x"63",
          9762 => x"72",
          9763 => x"63",
          9764 => x"00",
          9765 => x"64",
          9766 => x"00",
          9767 => x"64",
          9768 => x"00",
          9769 => x"65",
          9770 => x"65",
          9771 => x"65",
          9772 => x"69",
          9773 => x"69",
          9774 => x"66",
          9775 => x"66",
          9776 => x"61",
          9777 => x"00",
          9778 => x"6d",
          9779 => x"65",
          9780 => x"72",
          9781 => x"65",
          9782 => x"00",
          9783 => x"6e",
          9784 => x"00",
          9785 => x"65",
          9786 => x"00",
          9787 => x"62",
          9788 => x"63",
          9789 => x"62",
          9790 => x"63",
          9791 => x"69",
          9792 => x"00",
          9793 => x"64",
          9794 => x"69",
          9795 => x"45",
          9796 => x"72",
          9797 => x"6e",
          9798 => x"6e",
          9799 => x"65",
          9800 => x"72",
          9801 => x"69",
          9802 => x"6e",
          9803 => x"72",
          9804 => x"79",
          9805 => x"6f",
          9806 => x"6c",
          9807 => x"6f",
          9808 => x"2e",
          9809 => x"6f",
          9810 => x"74",
          9811 => x"6f",
          9812 => x"2e",
          9813 => x"6e",
          9814 => x"69",
          9815 => x"69",
          9816 => x"61",
          9817 => x"00",
          9818 => x"63",
          9819 => x"73",
          9820 => x"6e",
          9821 => x"2e",
          9822 => x"69",
          9823 => x"61",
          9824 => x"61",
          9825 => x"65",
          9826 => x"74",
          9827 => x"00",
          9828 => x"69",
          9829 => x"68",
          9830 => x"6c",
          9831 => x"6e",
          9832 => x"69",
          9833 => x"00",
          9834 => x"44",
          9835 => x"20",
          9836 => x"74",
          9837 => x"72",
          9838 => x"63",
          9839 => x"2e",
          9840 => x"72",
          9841 => x"20",
          9842 => x"62",
          9843 => x"69",
          9844 => x"6e",
          9845 => x"69",
          9846 => x"00",
          9847 => x"69",
          9848 => x"6e",
          9849 => x"65",
          9850 => x"6c",
          9851 => x"00",
          9852 => x"6f",
          9853 => x"6d",
          9854 => x"69",
          9855 => x"20",
          9856 => x"65",
          9857 => x"74",
          9858 => x"66",
          9859 => x"64",
          9860 => x"20",
          9861 => x"6b",
          9862 => x"6f",
          9863 => x"74",
          9864 => x"6f",
          9865 => x"64",
          9866 => x"69",
          9867 => x"75",
          9868 => x"6f",
          9869 => x"61",
          9870 => x"6e",
          9871 => x"6e",
          9872 => x"6c",
          9873 => x"00",
          9874 => x"69",
          9875 => x"69",
          9876 => x"6f",
          9877 => x"64",
          9878 => x"6e",
          9879 => x"66",
          9880 => x"65",
          9881 => x"6d",
          9882 => x"72",
          9883 => x"00",
          9884 => x"6f",
          9885 => x"61",
          9886 => x"6f",
          9887 => x"20",
          9888 => x"65",
          9889 => x"00",
          9890 => x"61",
          9891 => x"65",
          9892 => x"73",
          9893 => x"63",
          9894 => x"65",
          9895 => x"00",
          9896 => x"75",
          9897 => x"73",
          9898 => x"00",
          9899 => x"6e",
          9900 => x"77",
          9901 => x"72",
          9902 => x"2e",
          9903 => x"25",
          9904 => x"62",
          9905 => x"73",
          9906 => x"20",
          9907 => x"25",
          9908 => x"62",
          9909 => x"73",
          9910 => x"63",
          9911 => x"00",
          9912 => x"65",
          9913 => x"00",
          9914 => x"3d",
          9915 => x"6c",
          9916 => x"31",
          9917 => x"38",
          9918 => x"20",
          9919 => x"30",
          9920 => x"2c",
          9921 => x"4f",
          9922 => x"30",
          9923 => x"20",
          9924 => x"6c",
          9925 => x"30",
          9926 => x"0a",
          9927 => x"30",
          9928 => x"00",
          9929 => x"20",
          9930 => x"30",
          9931 => x"00",
          9932 => x"20",
          9933 => x"20",
          9934 => x"00",
          9935 => x"30",
          9936 => x"00",
          9937 => x"20",
          9938 => x"7c",
          9939 => x"00",
          9940 => x"4f",
          9941 => x"2a",
          9942 => x"73",
          9943 => x"00",
          9944 => x"35",
          9945 => x"2f",
          9946 => x"30",
          9947 => x"31",
          9948 => x"65",
          9949 => x"5a",
          9950 => x"20",
          9951 => x"20",
          9952 => x"78",
          9953 => x"73",
          9954 => x"20",
          9955 => x"0a",
          9956 => x"50",
          9957 => x"6e",
          9958 => x"72",
          9959 => x"20",
          9960 => x"64",
          9961 => x"00",
          9962 => x"69",
          9963 => x"20",
          9964 => x"65",
          9965 => x"70",
          9966 => x"53",
          9967 => x"6e",
          9968 => x"72",
          9969 => x"00",
          9970 => x"4f",
          9971 => x"20",
          9972 => x"69",
          9973 => x"72",
          9974 => x"74",
          9975 => x"4f",
          9976 => x"20",
          9977 => x"69",
          9978 => x"72",
          9979 => x"74",
          9980 => x"41",
          9981 => x"20",
          9982 => x"69",
          9983 => x"72",
          9984 => x"74",
          9985 => x"41",
          9986 => x"20",
          9987 => x"69",
          9988 => x"72",
          9989 => x"74",
          9990 => x"41",
          9991 => x"20",
          9992 => x"69",
          9993 => x"72",
          9994 => x"74",
          9995 => x"41",
          9996 => x"20",
          9997 => x"69",
          9998 => x"72",
          9999 => x"74",
         10000 => x"65",
         10001 => x"6e",
         10002 => x"70",
         10003 => x"6d",
         10004 => x"2e",
         10005 => x"6e",
         10006 => x"69",
         10007 => x"74",
         10008 => x"72",
         10009 => x"00",
         10010 => x"75",
         10011 => x"78",
         10012 => x"62",
         10013 => x"00",
         10014 => x"4f",
         10015 => x"73",
         10016 => x"3a",
         10017 => x"61",
         10018 => x"64",
         10019 => x"20",
         10020 => x"74",
         10021 => x"69",
         10022 => x"73",
         10023 => x"61",
         10024 => x"30",
         10025 => x"6c",
         10026 => x"65",
         10027 => x"69",
         10028 => x"61",
         10029 => x"6c",
         10030 => x"00",
         10031 => x"20",
         10032 => x"6c",
         10033 => x"69",
         10034 => x"2e",
         10035 => x"00",
         10036 => x"6f",
         10037 => x"6e",
         10038 => x"2e",
         10039 => x"6f",
         10040 => x"72",
         10041 => x"2e",
         10042 => x"00",
         10043 => x"30",
         10044 => x"28",
         10045 => x"78",
         10046 => x"25",
         10047 => x"78",
         10048 => x"38",
         10049 => x"00",
         10050 => x"75",
         10051 => x"4d",
         10052 => x"72",
         10053 => x"43",
         10054 => x"6c",
         10055 => x"2e",
         10056 => x"30",
         10057 => x"20",
         10058 => x"58",
         10059 => x"3f",
         10060 => x"30",
         10061 => x"20",
         10062 => x"58",
         10063 => x"30",
         10064 => x"20",
         10065 => x"6c",
         10066 => x"00",
         10067 => x"78",
         10068 => x"74",
         10069 => x"20",
         10070 => x"65",
         10071 => x"25",
         10072 => x"78",
         10073 => x"2e",
         10074 => x"61",
         10075 => x"6e",
         10076 => x"6f",
         10077 => x"40",
         10078 => x"38",
         10079 => x"2e",
         10080 => x"00",
         10081 => x"61",
         10082 => x"72",
         10083 => x"72",
         10084 => x"20",
         10085 => x"65",
         10086 => x"64",
         10087 => x"00",
         10088 => x"65",
         10089 => x"72",
         10090 => x"67",
         10091 => x"70",
         10092 => x"61",
         10093 => x"6e",
         10094 => x"00",
         10095 => x"6f",
         10096 => x"72",
         10097 => x"6f",
         10098 => x"67",
         10099 => x"00",
         10100 => x"50",
         10101 => x"69",
         10102 => x"64",
         10103 => x"73",
         10104 => x"2e",
         10105 => x"00",
         10106 => x"64",
         10107 => x"73",
         10108 => x"00",
         10109 => x"64",
         10110 => x"73",
         10111 => x"61",
         10112 => x"6f",
         10113 => x"6e",
         10114 => x"00",
         10115 => x"65",
         10116 => x"79",
         10117 => x"68",
         10118 => x"74",
         10119 => x"20",
         10120 => x"6e",
         10121 => x"70",
         10122 => x"65",
         10123 => x"63",
         10124 => x"61",
         10125 => x"00",
         10126 => x"75",
         10127 => x"6e",
         10128 => x"2e",
         10129 => x"6e",
         10130 => x"69",
         10131 => x"69",
         10132 => x"72",
         10133 => x"74",
         10134 => x"2e",
         10135 => x"64",
         10136 => x"2f",
         10137 => x"25",
         10138 => x"64",
         10139 => x"2e",
         10140 => x"64",
         10141 => x"6f",
         10142 => x"6f",
         10143 => x"67",
         10144 => x"74",
         10145 => x"00",
         10146 => x"28",
         10147 => x"6d",
         10148 => x"43",
         10149 => x"6e",
         10150 => x"29",
         10151 => x"0a",
         10152 => x"69",
         10153 => x"20",
         10154 => x"6c",
         10155 => x"6e",
         10156 => x"3a",
         10157 => x"20",
         10158 => x"42",
         10159 => x"52",
         10160 => x"20",
         10161 => x"38",
         10162 => x"30",
         10163 => x"2e",
         10164 => x"20",
         10165 => x"44",
         10166 => x"20",
         10167 => x"20",
         10168 => x"38",
         10169 => x"30",
         10170 => x"2e",
         10171 => x"20",
         10172 => x"4e",
         10173 => x"42",
         10174 => x"20",
         10175 => x"38",
         10176 => x"30",
         10177 => x"2e",
         10178 => x"20",
         10179 => x"52",
         10180 => x"20",
         10181 => x"20",
         10182 => x"38",
         10183 => x"30",
         10184 => x"2e",
         10185 => x"20",
         10186 => x"41",
         10187 => x"20",
         10188 => x"20",
         10189 => x"38",
         10190 => x"30",
         10191 => x"2e",
         10192 => x"20",
         10193 => x"44",
         10194 => x"52",
         10195 => x"20",
         10196 => x"76",
         10197 => x"73",
         10198 => x"30",
         10199 => x"2e",
         10200 => x"20",
         10201 => x"49",
         10202 => x"31",
         10203 => x"20",
         10204 => x"6d",
         10205 => x"20",
         10206 => x"30",
         10207 => x"2e",
         10208 => x"20",
         10209 => x"4e",
         10210 => x"43",
         10211 => x"20",
         10212 => x"61",
         10213 => x"6c",
         10214 => x"30",
         10215 => x"2e",
         10216 => x"20",
         10217 => x"49",
         10218 => x"4f",
         10219 => x"42",
         10220 => x"00",
         10221 => x"20",
         10222 => x"42",
         10223 => x"43",
         10224 => x"20",
         10225 => x"4f",
         10226 => x"00",
         10227 => x"20",
         10228 => x"53",
         10229 => x"20",
         10230 => x"50",
         10231 => x"64",
         10232 => x"73",
         10233 => x"3a",
         10234 => x"20",
         10235 => x"50",
         10236 => x"65",
         10237 => x"20",
         10238 => x"74",
         10239 => x"41",
         10240 => x"65",
         10241 => x"3d",
         10242 => x"38",
         10243 => x"00",
         10244 => x"20",
         10245 => x"50",
         10246 => x"65",
         10247 => x"79",
         10248 => x"61",
         10249 => x"41",
         10250 => x"65",
         10251 => x"3d",
         10252 => x"38",
         10253 => x"00",
         10254 => x"20",
         10255 => x"74",
         10256 => x"20",
         10257 => x"72",
         10258 => x"64",
         10259 => x"73",
         10260 => x"20",
         10261 => x"3d",
         10262 => x"38",
         10263 => x"00",
         10264 => x"69",
         10265 => x"00",
         10266 => x"20",
         10267 => x"50",
         10268 => x"64",
         10269 => x"20",
         10270 => x"20",
         10271 => x"20",
         10272 => x"20",
         10273 => x"3d",
         10274 => x"34",
         10275 => x"00",
         10276 => x"20",
         10277 => x"79",
         10278 => x"6d",
         10279 => x"6f",
         10280 => x"46",
         10281 => x"20",
         10282 => x"20",
         10283 => x"3d",
         10284 => x"2e",
         10285 => x"64",
         10286 => x"0a",
         10287 => x"20",
         10288 => x"44",
         10289 => x"20",
         10290 => x"63",
         10291 => x"72",
         10292 => x"20",
         10293 => x"20",
         10294 => x"3d",
         10295 => x"2e",
         10296 => x"64",
         10297 => x"0a",
         10298 => x"20",
         10299 => x"69",
         10300 => x"6f",
         10301 => x"53",
         10302 => x"4d",
         10303 => x"6f",
         10304 => x"46",
         10305 => x"3d",
         10306 => x"2e",
         10307 => x"64",
         10308 => x"0a",
         10309 => x"6d",
         10310 => x"00",
         10311 => x"65",
         10312 => x"6d",
         10313 => x"6c",
         10314 => x"00",
         10315 => x"56",
         10316 => x"56",
         10317 => x"00",
         10318 => x"6e",
         10319 => x"77",
         10320 => x"00",
         10321 => x"00",
         10322 => x"00",
         10323 => x"00",
         10324 => x"00",
         10325 => x"00",
         10326 => x"00",
         10327 => x"00",
         10328 => x"00",
         10329 => x"00",
         10330 => x"00",
         10331 => x"00",
         10332 => x"00",
         10333 => x"00",
         10334 => x"00",
         10335 => x"00",
         10336 => x"00",
         10337 => x"00",
         10338 => x"00",
         10339 => x"00",
         10340 => x"00",
         10341 => x"00",
         10342 => x"00",
         10343 => x"00",
         10344 => x"00",
         10345 => x"00",
         10346 => x"00",
         10347 => x"00",
         10348 => x"00",
         10349 => x"00",
         10350 => x"00",
         10351 => x"00",
         10352 => x"00",
         10353 => x"00",
         10354 => x"00",
         10355 => x"00",
         10356 => x"00",
         10357 => x"00",
         10358 => x"00",
         10359 => x"00",
         10360 => x"00",
         10361 => x"00",
         10362 => x"00",
         10363 => x"00",
         10364 => x"00",
         10365 => x"00",
         10366 => x"00",
         10367 => x"00",
         10368 => x"00",
         10369 => x"00",
         10370 => x"00",
         10371 => x"00",
         10372 => x"00",
         10373 => x"00",
         10374 => x"00",
         10375 => x"00",
         10376 => x"00",
         10377 => x"00",
         10378 => x"00",
         10379 => x"00",
         10380 => x"00",
         10381 => x"00",
         10382 => x"00",
         10383 => x"00",
         10384 => x"00",
         10385 => x"00",
         10386 => x"5b",
         10387 => x"5b",
         10388 => x"5b",
         10389 => x"5b",
         10390 => x"5b",
         10391 => x"5b",
         10392 => x"5b",
         10393 => x"30",
         10394 => x"5b",
         10395 => x"5b",
         10396 => x"5b",
         10397 => x"00",
         10398 => x"00",
         10399 => x"00",
         10400 => x"00",
         10401 => x"00",
         10402 => x"00",
         10403 => x"00",
         10404 => x"00",
         10405 => x"00",
         10406 => x"00",
         10407 => x"00",
         10408 => x"69",
         10409 => x"72",
         10410 => x"69",
         10411 => x"00",
         10412 => x"00",
         10413 => x"30",
         10414 => x"20",
         10415 => x"0a",
         10416 => x"61",
         10417 => x"64",
         10418 => x"20",
         10419 => x"65",
         10420 => x"68",
         10421 => x"69",
         10422 => x"72",
         10423 => x"69",
         10424 => x"74",
         10425 => x"4f",
         10426 => x"00",
         10427 => x"61",
         10428 => x"74",
         10429 => x"65",
         10430 => x"72",
         10431 => x"65",
         10432 => x"73",
         10433 => x"79",
         10434 => x"6c",
         10435 => x"64",
         10436 => x"62",
         10437 => x"67",
         10438 => x"44",
         10439 => x"2a",
         10440 => x"3f",
         10441 => x"00",
         10442 => x"2c",
         10443 => x"5d",
         10444 => x"41",
         10445 => x"41",
         10446 => x"00",
         10447 => x"fe",
         10448 => x"44",
         10449 => x"2e",
         10450 => x"4f",
         10451 => x"4d",
         10452 => x"20",
         10453 => x"54",
         10454 => x"20",
         10455 => x"4f",
         10456 => x"4d",
         10457 => x"20",
         10458 => x"54",
         10459 => x"20",
         10460 => x"00",
         10461 => x"00",
         10462 => x"00",
         10463 => x"00",
         10464 => x"03",
         10465 => x"0e",
         10466 => x"16",
         10467 => x"00",
         10468 => x"9a",
         10469 => x"41",
         10470 => x"45",
         10471 => x"49",
         10472 => x"92",
         10473 => x"4f",
         10474 => x"99",
         10475 => x"9d",
         10476 => x"49",
         10477 => x"a5",
         10478 => x"a9",
         10479 => x"ad",
         10480 => x"b1",
         10481 => x"b5",
         10482 => x"b9",
         10483 => x"bd",
         10484 => x"c1",
         10485 => x"c5",
         10486 => x"c9",
         10487 => x"cd",
         10488 => x"d1",
         10489 => x"d5",
         10490 => x"d9",
         10491 => x"dd",
         10492 => x"e1",
         10493 => x"e5",
         10494 => x"e9",
         10495 => x"ed",
         10496 => x"f1",
         10497 => x"f5",
         10498 => x"f9",
         10499 => x"fd",
         10500 => x"2e",
         10501 => x"5b",
         10502 => x"22",
         10503 => x"3e",
         10504 => x"00",
         10505 => x"01",
         10506 => x"10",
         10507 => x"00",
         10508 => x"00",
         10509 => x"01",
         10510 => x"04",
         10511 => x"10",
         10512 => x"00",
         10513 => x"c7",
         10514 => x"e9",
         10515 => x"e4",
         10516 => x"e5",
         10517 => x"ea",
         10518 => x"e8",
         10519 => x"ee",
         10520 => x"c4",
         10521 => x"c9",
         10522 => x"c6",
         10523 => x"f6",
         10524 => x"fb",
         10525 => x"ff",
         10526 => x"dc",
         10527 => x"a3",
         10528 => x"a7",
         10529 => x"e1",
         10530 => x"f3",
         10531 => x"f1",
         10532 => x"aa",
         10533 => x"bf",
         10534 => x"ac",
         10535 => x"bc",
         10536 => x"ab",
         10537 => x"91",
         10538 => x"93",
         10539 => x"24",
         10540 => x"62",
         10541 => x"55",
         10542 => x"51",
         10543 => x"5d",
         10544 => x"5b",
         10545 => x"14",
         10546 => x"2c",
         10547 => x"00",
         10548 => x"5e",
         10549 => x"5a",
         10550 => x"69",
         10551 => x"60",
         10552 => x"6c",
         10553 => x"68",
         10554 => x"65",
         10555 => x"58",
         10556 => x"53",
         10557 => x"6a",
         10558 => x"0c",
         10559 => x"84",
         10560 => x"90",
         10561 => x"b1",
         10562 => x"93",
         10563 => x"a3",
         10564 => x"b5",
         10565 => x"a6",
         10566 => x"a9",
         10567 => x"1e",
         10568 => x"b5",
         10569 => x"61",
         10570 => x"65",
         10571 => x"20",
         10572 => x"f7",
         10573 => x"b0",
         10574 => x"b7",
         10575 => x"7f",
         10576 => x"a0",
         10577 => x"61",
         10578 => x"e0",
         10579 => x"f8",
         10580 => x"ff",
         10581 => x"78",
         10582 => x"30",
         10583 => x"06",
         10584 => x"10",
         10585 => x"2e",
         10586 => x"06",
         10587 => x"4d",
         10588 => x"81",
         10589 => x"82",
         10590 => x"84",
         10591 => x"87",
         10592 => x"89",
         10593 => x"8b",
         10594 => x"8d",
         10595 => x"8f",
         10596 => x"91",
         10597 => x"93",
         10598 => x"f6",
         10599 => x"97",
         10600 => x"98",
         10601 => x"9b",
         10602 => x"9d",
         10603 => x"9f",
         10604 => x"a0",
         10605 => x"a2",
         10606 => x"a4",
         10607 => x"a7",
         10608 => x"a9",
         10609 => x"ab",
         10610 => x"ac",
         10611 => x"af",
         10612 => x"b1",
         10613 => x"b3",
         10614 => x"b5",
         10615 => x"b7",
         10616 => x"b8",
         10617 => x"bb",
         10618 => x"bc",
         10619 => x"f7",
         10620 => x"c1",
         10621 => x"c3",
         10622 => x"c5",
         10623 => x"c7",
         10624 => x"c7",
         10625 => x"cb",
         10626 => x"cd",
         10627 => x"dd",
         10628 => x"8e",
         10629 => x"12",
         10630 => x"03",
         10631 => x"f4",
         10632 => x"f8",
         10633 => x"22",
         10634 => x"3a",
         10635 => x"65",
         10636 => x"3b",
         10637 => x"66",
         10638 => x"40",
         10639 => x"41",
         10640 => x"0a",
         10641 => x"40",
         10642 => x"86",
         10643 => x"89",
         10644 => x"58",
         10645 => x"5a",
         10646 => x"5c",
         10647 => x"5e",
         10648 => x"93",
         10649 => x"62",
         10650 => x"64",
         10651 => x"66",
         10652 => x"97",
         10653 => x"6a",
         10654 => x"6c",
         10655 => x"6e",
         10656 => x"70",
         10657 => x"9d",
         10658 => x"74",
         10659 => x"76",
         10660 => x"78",
         10661 => x"7a",
         10662 => x"7c",
         10663 => x"7e",
         10664 => x"a6",
         10665 => x"82",
         10666 => x"84",
         10667 => x"86",
         10668 => x"ae",
         10669 => x"b1",
         10670 => x"45",
         10671 => x"8e",
         10672 => x"90",
         10673 => x"b7",
         10674 => x"03",
         10675 => x"fe",
         10676 => x"ac",
         10677 => x"86",
         10678 => x"89",
         10679 => x"b1",
         10680 => x"c2",
         10681 => x"a3",
         10682 => x"c4",
         10683 => x"cc",
         10684 => x"8c",
         10685 => x"8f",
         10686 => x"18",
         10687 => x"0a",
         10688 => x"f3",
         10689 => x"f5",
         10690 => x"f7",
         10691 => x"f9",
         10692 => x"fa",
         10693 => x"20",
         10694 => x"10",
         10695 => x"22",
         10696 => x"36",
         10697 => x"0e",
         10698 => x"01",
         10699 => x"d0",
         10700 => x"61",
         10701 => x"00",
         10702 => x"7d",
         10703 => x"63",
         10704 => x"96",
         10705 => x"5a",
         10706 => x"08",
         10707 => x"06",
         10708 => x"08",
         10709 => x"08",
         10710 => x"06",
         10711 => x"07",
         10712 => x"52",
         10713 => x"54",
         10714 => x"56",
         10715 => x"60",
         10716 => x"70",
         10717 => x"ba",
         10718 => x"c8",
         10719 => x"ca",
         10720 => x"da",
         10721 => x"f8",
         10722 => x"ea",
         10723 => x"fa",
         10724 => x"80",
         10725 => x"90",
         10726 => x"a0",
         10727 => x"b0",
         10728 => x"b8",
         10729 => x"b2",
         10730 => x"cc",
         10731 => x"c3",
         10732 => x"02",
         10733 => x"02",
         10734 => x"01",
         10735 => x"f3",
         10736 => x"fc",
         10737 => x"01",
         10738 => x"70",
         10739 => x"84",
         10740 => x"83",
         10741 => x"1a",
         10742 => x"2f",
         10743 => x"02",
         10744 => x"06",
         10745 => x"02",
         10746 => x"64",
         10747 => x"26",
         10748 => x"1a",
         10749 => x"00",
         10750 => x"00",
         10751 => x"02",
         10752 => x"00",
         10753 => x"00",
         10754 => x"00",
         10755 => x"04",
         10756 => x"00",
         10757 => x"00",
         10758 => x"00",
         10759 => x"14",
         10760 => x"00",
         10761 => x"00",
         10762 => x"00",
         10763 => x"2b",
         10764 => x"00",
         10765 => x"00",
         10766 => x"00",
         10767 => x"30",
         10768 => x"00",
         10769 => x"00",
         10770 => x"00",
         10771 => x"3c",
         10772 => x"00",
         10773 => x"00",
         10774 => x"00",
         10775 => x"3d",
         10776 => x"00",
         10777 => x"00",
         10778 => x"00",
         10779 => x"3f",
         10780 => x"00",
         10781 => x"00",
         10782 => x"00",
         10783 => x"40",
         10784 => x"00",
         10785 => x"00",
         10786 => x"00",
         10787 => x"41",
         10788 => x"00",
         10789 => x"00",
         10790 => x"00",
         10791 => x"42",
         10792 => x"00",
         10793 => x"00",
         10794 => x"00",
         10795 => x"43",
         10796 => x"00",
         10797 => x"00",
         10798 => x"00",
         10799 => x"50",
         10800 => x"00",
         10801 => x"00",
         10802 => x"00",
         10803 => x"51",
         10804 => x"00",
         10805 => x"00",
         10806 => x"00",
         10807 => x"54",
         10808 => x"00",
         10809 => x"00",
         10810 => x"00",
         10811 => x"55",
         10812 => x"00",
         10813 => x"00",
         10814 => x"00",
         10815 => x"79",
         10816 => x"00",
         10817 => x"00",
         10818 => x"00",
         10819 => x"78",
         10820 => x"00",
         10821 => x"00",
         10822 => x"00",
         10823 => x"82",
         10824 => x"00",
         10825 => x"00",
         10826 => x"00",
         10827 => x"83",
         10828 => x"00",
         10829 => x"00",
         10830 => x"00",
         10831 => x"85",
         10832 => x"00",
         10833 => x"00",
         10834 => x"00",
         10835 => x"87",
         10836 => x"00",
         10837 => x"00",
         10838 => x"00",
         10839 => x"8c",
         10840 => x"00",
         10841 => x"00",
         10842 => x"00",
         10843 => x"8d",
         10844 => x"00",
         10845 => x"00",
         10846 => x"00",
         10847 => x"8e",
         10848 => x"00",
         10849 => x"00",
         10850 => x"00",
         10851 => x"8f",
         10852 => x"00",
         10853 => x"00",
         10854 => x"00",
         10855 => x"00",
         10856 => x"00",
         10857 => x"00",
         10858 => x"00",
         10859 => x"01",
         10860 => x"00",
         10861 => x"01",
         10862 => x"81",
         10863 => x"00",
         10864 => x"7f",
         10865 => x"00",
         10866 => x"00",
         10867 => x"00",
         10868 => x"00",
         10869 => x"f5",
         10870 => x"f5",
         10871 => x"f5",
         10872 => x"00",
         10873 => x"01",
         10874 => x"01",
         10875 => x"01",
         10876 => x"00",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"00",
         10884 => x"00",
         10885 => x"00",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"00",
         10890 => x"00",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"00",
         10895 => x"00",
         10896 => x"00",
         10897 => x"00",
         10898 => x"00",
         10899 => x"00",
         10900 => x"00",
         10901 => x"00",
         10902 => x"00",
         10903 => x"00",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"9d",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"88",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"9f",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"8b",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"95",
           269 => x"0b",
           270 => x"0b",
           271 => x"b3",
           272 => x"0b",
           273 => x"0b",
           274 => x"d1",
           275 => x"0b",
           276 => x"0b",
           277 => x"f0",
           278 => x"0b",
           279 => x"0b",
           280 => x"8f",
           281 => x"0b",
           282 => x"0b",
           283 => x"ad",
           284 => x"0b",
           285 => x"0b",
           286 => x"cd",
           287 => x"0b",
           288 => x"0b",
           289 => x"ed",
           290 => x"0b",
           291 => x"0b",
           292 => x"8d",
           293 => x"0b",
           294 => x"0b",
           295 => x"ad",
           296 => x"0b",
           297 => x"0b",
           298 => x"cd",
           299 => x"0b",
           300 => x"0b",
           301 => x"ed",
           302 => x"0b",
           303 => x"0b",
           304 => x"8d",
           305 => x"0b",
           306 => x"0b",
           307 => x"ad",
           308 => x"0b",
           309 => x"0b",
           310 => x"cd",
           311 => x"0b",
           312 => x"0b",
           313 => x"ed",
           314 => x"0b",
           315 => x"0b",
           316 => x"8d",
           317 => x"0b",
           318 => x"0b",
           319 => x"ad",
           320 => x"0b",
           321 => x"0b",
           322 => x"cd",
           323 => x"0b",
           324 => x"0b",
           325 => x"ed",
           326 => x"0b",
           327 => x"0b",
           328 => x"8d",
           329 => x"0b",
           330 => x"0b",
           331 => x"ad",
           332 => x"0b",
           333 => x"0b",
           334 => x"cd",
           335 => x"0b",
           336 => x"0b",
           337 => x"ed",
           338 => x"0b",
           339 => x"0b",
           340 => x"8d",
           341 => x"0b",
           342 => x"0b",
           343 => x"ad",
           344 => x"0b",
           345 => x"0b",
           346 => x"cd",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"04",
           390 => x"0c",
           391 => x"82",
           392 => x"84",
           393 => x"82",
           394 => x"af",
           395 => x"d5",
           396 => x"80",
           397 => x"d5",
           398 => x"ad",
           399 => x"84",
           400 => x"90",
           401 => x"84",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"82",
           407 => x"84",
           408 => x"82",
           409 => x"80",
           410 => x"82",
           411 => x"84",
           412 => x"82",
           413 => x"80",
           414 => x"82",
           415 => x"84",
           416 => x"82",
           417 => x"93",
           418 => x"d5",
           419 => x"80",
           420 => x"d5",
           421 => x"c0",
           422 => x"84",
           423 => x"90",
           424 => x"84",
           425 => x"2d",
           426 => x"08",
           427 => x"04",
           428 => x"0c",
           429 => x"2d",
           430 => x"08",
           431 => x"04",
           432 => x"0c",
           433 => x"2d",
           434 => x"08",
           435 => x"04",
           436 => x"0c",
           437 => x"2d",
           438 => x"08",
           439 => x"04",
           440 => x"0c",
           441 => x"2d",
           442 => x"08",
           443 => x"04",
           444 => x"0c",
           445 => x"2d",
           446 => x"08",
           447 => x"04",
           448 => x"0c",
           449 => x"2d",
           450 => x"08",
           451 => x"04",
           452 => x"0c",
           453 => x"2d",
           454 => x"08",
           455 => x"04",
           456 => x"0c",
           457 => x"2d",
           458 => x"08",
           459 => x"04",
           460 => x"0c",
           461 => x"2d",
           462 => x"08",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"04",
           480 => x"0c",
           481 => x"2d",
           482 => x"08",
           483 => x"04",
           484 => x"0c",
           485 => x"2d",
           486 => x"08",
           487 => x"04",
           488 => x"0c",
           489 => x"2d",
           490 => x"08",
           491 => x"04",
           492 => x"0c",
           493 => x"2d",
           494 => x"08",
           495 => x"04",
           496 => x"0c",
           497 => x"2d",
           498 => x"08",
           499 => x"04",
           500 => x"0c",
           501 => x"2d",
           502 => x"08",
           503 => x"04",
           504 => x"0c",
           505 => x"2d",
           506 => x"08",
           507 => x"04",
           508 => x"0c",
           509 => x"2d",
           510 => x"08",
           511 => x"04",
           512 => x"0c",
           513 => x"2d",
           514 => x"08",
           515 => x"04",
           516 => x"0c",
           517 => x"2d",
           518 => x"08",
           519 => x"04",
           520 => x"0c",
           521 => x"2d",
           522 => x"08",
           523 => x"04",
           524 => x"0c",
           525 => x"2d",
           526 => x"08",
           527 => x"04",
           528 => x"0c",
           529 => x"2d",
           530 => x"08",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"04",
           548 => x"0c",
           549 => x"2d",
           550 => x"08",
           551 => x"04",
           552 => x"0c",
           553 => x"2d",
           554 => x"08",
           555 => x"04",
           556 => x"0c",
           557 => x"2d",
           558 => x"08",
           559 => x"04",
           560 => x"0c",
           561 => x"2d",
           562 => x"08",
           563 => x"04",
           564 => x"0c",
           565 => x"2d",
           566 => x"08",
           567 => x"04",
           568 => x"0c",
           569 => x"2d",
           570 => x"08",
           571 => x"04",
           572 => x"0c",
           573 => x"2d",
           574 => x"08",
           575 => x"04",
           576 => x"0c",
           577 => x"2d",
           578 => x"08",
           579 => x"04",
           580 => x"0c",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"0c",
           589 => x"2d",
           590 => x"08",
           591 => x"04",
           592 => x"0c",
           593 => x"2d",
           594 => x"08",
           595 => x"04",
           596 => x"0c",
           597 => x"2d",
           598 => x"08",
           599 => x"04",
           600 => x"00",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"53",
           609 => x"00",
           610 => x"06",
           611 => x"09",
           612 => x"05",
           613 => x"2b",
           614 => x"06",
           615 => x"04",
           616 => x"72",
           617 => x"05",
           618 => x"05",
           619 => x"72",
           620 => x"53",
           621 => x"51",
           622 => x"04",
           623 => x"70",
           624 => x"27",
           625 => x"71",
           626 => x"53",
           627 => x"0b",
           628 => x"8c",
           629 => x"f0",
           630 => x"82",
           631 => x"02",
           632 => x"0c",
           633 => x"82",
           634 => x"8c",
           635 => x"d5",
           636 => x"05",
           637 => x"84",
           638 => x"08",
           639 => x"84",
           640 => x"08",
           641 => x"dc",
           642 => x"84",
           643 => x"d4",
           644 => x"82",
           645 => x"f8",
           646 => x"d5",
           647 => x"05",
           648 => x"d4",
           649 => x"54",
           650 => x"82",
           651 => x"04",
           652 => x"08",
           653 => x"84",
           654 => x"0d",
           655 => x"08",
           656 => x"85",
           657 => x"81",
           658 => x"06",
           659 => x"52",
           660 => x"80",
           661 => x"84",
           662 => x"08",
           663 => x"8d",
           664 => x"82",
           665 => x"f4",
           666 => x"c4",
           667 => x"84",
           668 => x"08",
           669 => x"d5",
           670 => x"05",
           671 => x"82",
           672 => x"f8",
           673 => x"d5",
           674 => x"05",
           675 => x"84",
           676 => x"0c",
           677 => x"08",
           678 => x"8a",
           679 => x"38",
           680 => x"d5",
           681 => x"05",
           682 => x"e9",
           683 => x"84",
           684 => x"08",
           685 => x"3f",
           686 => x"08",
           687 => x"84",
           688 => x"0c",
           689 => x"84",
           690 => x"08",
           691 => x"81",
           692 => x"80",
           693 => x"84",
           694 => x"0c",
           695 => x"82",
           696 => x"fc",
           697 => x"d5",
           698 => x"05",
           699 => x"71",
           700 => x"d5",
           701 => x"05",
           702 => x"82",
           703 => x"8c",
           704 => x"d5",
           705 => x"05",
           706 => x"82",
           707 => x"fc",
           708 => x"80",
           709 => x"84",
           710 => x"08",
           711 => x"34",
           712 => x"08",
           713 => x"70",
           714 => x"08",
           715 => x"52",
           716 => x"08",
           717 => x"82",
           718 => x"87",
           719 => x"d5",
           720 => x"82",
           721 => x"02",
           722 => x"0c",
           723 => x"86",
           724 => x"84",
           725 => x"34",
           726 => x"08",
           727 => x"82",
           728 => x"e0",
           729 => x"0a",
           730 => x"84",
           731 => x"0c",
           732 => x"08",
           733 => x"82",
           734 => x"fc",
           735 => x"d5",
           736 => x"05",
           737 => x"d5",
           738 => x"05",
           739 => x"d5",
           740 => x"05",
           741 => x"54",
           742 => x"82",
           743 => x"70",
           744 => x"08",
           745 => x"82",
           746 => x"ec",
           747 => x"d5",
           748 => x"05",
           749 => x"54",
           750 => x"82",
           751 => x"dc",
           752 => x"82",
           753 => x"54",
           754 => x"82",
           755 => x"04",
           756 => x"08",
           757 => x"84",
           758 => x"0d",
           759 => x"08",
           760 => x"82",
           761 => x"fc",
           762 => x"d5",
           763 => x"05",
           764 => x"d5",
           765 => x"05",
           766 => x"d5",
           767 => x"05",
           768 => x"a3",
           769 => x"f8",
           770 => x"d5",
           771 => x"05",
           772 => x"84",
           773 => x"08",
           774 => x"f8",
           775 => x"87",
           776 => x"d5",
           777 => x"82",
           778 => x"02",
           779 => x"0c",
           780 => x"80",
           781 => x"84",
           782 => x"23",
           783 => x"08",
           784 => x"53",
           785 => x"14",
           786 => x"84",
           787 => x"08",
           788 => x"70",
           789 => x"81",
           790 => x"06",
           791 => x"51",
           792 => x"2e",
           793 => x"0b",
           794 => x"08",
           795 => x"96",
           796 => x"d5",
           797 => x"05",
           798 => x"33",
           799 => x"d5",
           800 => x"05",
           801 => x"ff",
           802 => x"80",
           803 => x"38",
           804 => x"08",
           805 => x"81",
           806 => x"84",
           807 => x"0c",
           808 => x"08",
           809 => x"70",
           810 => x"53",
           811 => x"95",
           812 => x"d5",
           813 => x"05",
           814 => x"73",
           815 => x"38",
           816 => x"08",
           817 => x"53",
           818 => x"81",
           819 => x"d5",
           820 => x"05",
           821 => x"b0",
           822 => x"06",
           823 => x"82",
           824 => x"e8",
           825 => x"98",
           826 => x"2c",
           827 => x"72",
           828 => x"d5",
           829 => x"05",
           830 => x"2a",
           831 => x"70",
           832 => x"51",
           833 => x"80",
           834 => x"82",
           835 => x"e4",
           836 => x"82",
           837 => x"53",
           838 => x"84",
           839 => x"23",
           840 => x"82",
           841 => x"e8",
           842 => x"98",
           843 => x"2c",
           844 => x"2b",
           845 => x"11",
           846 => x"53",
           847 => x"72",
           848 => x"08",
           849 => x"82",
           850 => x"e8",
           851 => x"82",
           852 => x"f8",
           853 => x"15",
           854 => x"51",
           855 => x"d5",
           856 => x"05",
           857 => x"84",
           858 => x"33",
           859 => x"70",
           860 => x"51",
           861 => x"25",
           862 => x"ff",
           863 => x"84",
           864 => x"34",
           865 => x"08",
           866 => x"70",
           867 => x"81",
           868 => x"53",
           869 => x"38",
           870 => x"08",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"53",
           876 => x"84",
           877 => x"23",
           878 => x"82",
           879 => x"e4",
           880 => x"83",
           881 => x"06",
           882 => x"72",
           883 => x"38",
           884 => x"08",
           885 => x"70",
           886 => x"98",
           887 => x"53",
           888 => x"81",
           889 => x"84",
           890 => x"34",
           891 => x"08",
           892 => x"e0",
           893 => x"84",
           894 => x"0c",
           895 => x"84",
           896 => x"08",
           897 => x"92",
           898 => x"d5",
           899 => x"05",
           900 => x"2b",
           901 => x"11",
           902 => x"51",
           903 => x"04",
           904 => x"08",
           905 => x"70",
           906 => x"53",
           907 => x"84",
           908 => x"23",
           909 => x"08",
           910 => x"70",
           911 => x"53",
           912 => x"84",
           913 => x"23",
           914 => x"82",
           915 => x"e4",
           916 => x"81",
           917 => x"53",
           918 => x"84",
           919 => x"23",
           920 => x"82",
           921 => x"e4",
           922 => x"80",
           923 => x"53",
           924 => x"84",
           925 => x"23",
           926 => x"82",
           927 => x"e4",
           928 => x"88",
           929 => x"72",
           930 => x"08",
           931 => x"80",
           932 => x"84",
           933 => x"34",
           934 => x"82",
           935 => x"e4",
           936 => x"84",
           937 => x"72",
           938 => x"08",
           939 => x"fb",
           940 => x"0b",
           941 => x"08",
           942 => x"82",
           943 => x"ec",
           944 => x"11",
           945 => x"82",
           946 => x"ec",
           947 => x"e3",
           948 => x"84",
           949 => x"34",
           950 => x"82",
           951 => x"90",
           952 => x"d5",
           953 => x"05",
           954 => x"82",
           955 => x"90",
           956 => x"08",
           957 => x"82",
           958 => x"fc",
           959 => x"d5",
           960 => x"05",
           961 => x"51",
           962 => x"d5",
           963 => x"05",
           964 => x"39",
           965 => x"08",
           966 => x"82",
           967 => x"90",
           968 => x"05",
           969 => x"08",
           970 => x"70",
           971 => x"84",
           972 => x"0c",
           973 => x"08",
           974 => x"70",
           975 => x"81",
           976 => x"51",
           977 => x"2e",
           978 => x"d5",
           979 => x"05",
           980 => x"2b",
           981 => x"2c",
           982 => x"84",
           983 => x"08",
           984 => x"83",
           985 => x"f8",
           986 => x"82",
           987 => x"f4",
           988 => x"39",
           989 => x"08",
           990 => x"51",
           991 => x"82",
           992 => x"53",
           993 => x"84",
           994 => x"23",
           995 => x"08",
           996 => x"53",
           997 => x"08",
           998 => x"73",
           999 => x"54",
          1000 => x"84",
          1001 => x"23",
          1002 => x"82",
          1003 => x"90",
          1004 => x"d5",
          1005 => x"05",
          1006 => x"82",
          1007 => x"90",
          1008 => x"08",
          1009 => x"08",
          1010 => x"82",
          1011 => x"e4",
          1012 => x"83",
          1013 => x"06",
          1014 => x"53",
          1015 => x"ab",
          1016 => x"84",
          1017 => x"33",
          1018 => x"53",
          1019 => x"53",
          1020 => x"08",
          1021 => x"52",
          1022 => x"3f",
          1023 => x"08",
          1024 => x"d5",
          1025 => x"05",
          1026 => x"82",
          1027 => x"fc",
          1028 => x"9b",
          1029 => x"d4",
          1030 => x"72",
          1031 => x"08",
          1032 => x"82",
          1033 => x"ec",
          1034 => x"82",
          1035 => x"f4",
          1036 => x"71",
          1037 => x"72",
          1038 => x"08",
          1039 => x"8a",
          1040 => x"d5",
          1041 => x"05",
          1042 => x"2a",
          1043 => x"51",
          1044 => x"80",
          1045 => x"82",
          1046 => x"90",
          1047 => x"d5",
          1048 => x"05",
          1049 => x"82",
          1050 => x"90",
          1051 => x"08",
          1052 => x"08",
          1053 => x"53",
          1054 => x"d5",
          1055 => x"05",
          1056 => x"84",
          1057 => x"08",
          1058 => x"d5",
          1059 => x"05",
          1060 => x"82",
          1061 => x"dc",
          1062 => x"82",
          1063 => x"dc",
          1064 => x"d5",
          1065 => x"05",
          1066 => x"84",
          1067 => x"08",
          1068 => x"38",
          1069 => x"08",
          1070 => x"70",
          1071 => x"53",
          1072 => x"84",
          1073 => x"23",
          1074 => x"08",
          1075 => x"30",
          1076 => x"08",
          1077 => x"82",
          1078 => x"e4",
          1079 => x"ff",
          1080 => x"53",
          1081 => x"84",
          1082 => x"23",
          1083 => x"88",
          1084 => x"84",
          1085 => x"23",
          1086 => x"d5",
          1087 => x"05",
          1088 => x"c0",
          1089 => x"72",
          1090 => x"08",
          1091 => x"80",
          1092 => x"d5",
          1093 => x"05",
          1094 => x"82",
          1095 => x"f4",
          1096 => x"d5",
          1097 => x"05",
          1098 => x"2a",
          1099 => x"51",
          1100 => x"80",
          1101 => x"82",
          1102 => x"90",
          1103 => x"d5",
          1104 => x"05",
          1105 => x"82",
          1106 => x"90",
          1107 => x"08",
          1108 => x"08",
          1109 => x"53",
          1110 => x"d5",
          1111 => x"05",
          1112 => x"84",
          1113 => x"08",
          1114 => x"d5",
          1115 => x"05",
          1116 => x"82",
          1117 => x"d8",
          1118 => x"82",
          1119 => x"d8",
          1120 => x"d5",
          1121 => x"05",
          1122 => x"84",
          1123 => x"22",
          1124 => x"51",
          1125 => x"d5",
          1126 => x"05",
          1127 => x"88",
          1128 => x"84",
          1129 => x"0c",
          1130 => x"08",
          1131 => x"82",
          1132 => x"f4",
          1133 => x"d5",
          1134 => x"05",
          1135 => x"70",
          1136 => x"55",
          1137 => x"82",
          1138 => x"53",
          1139 => x"82",
          1140 => x"f0",
          1141 => x"d5",
          1142 => x"05",
          1143 => x"84",
          1144 => x"08",
          1145 => x"53",
          1146 => x"a4",
          1147 => x"84",
          1148 => x"08",
          1149 => x"54",
          1150 => x"08",
          1151 => x"70",
          1152 => x"51",
          1153 => x"82",
          1154 => x"d0",
          1155 => x"39",
          1156 => x"08",
          1157 => x"53",
          1158 => x"11",
          1159 => x"82",
          1160 => x"d0",
          1161 => x"d5",
          1162 => x"05",
          1163 => x"d5",
          1164 => x"05",
          1165 => x"82",
          1166 => x"f0",
          1167 => x"05",
          1168 => x"08",
          1169 => x"82",
          1170 => x"f4",
          1171 => x"53",
          1172 => x"08",
          1173 => x"52",
          1174 => x"3f",
          1175 => x"08",
          1176 => x"84",
          1177 => x"0c",
          1178 => x"84",
          1179 => x"08",
          1180 => x"38",
          1181 => x"82",
          1182 => x"f0",
          1183 => x"d5",
          1184 => x"72",
          1185 => x"75",
          1186 => x"72",
          1187 => x"08",
          1188 => x"82",
          1189 => x"e4",
          1190 => x"b2",
          1191 => x"72",
          1192 => x"38",
          1193 => x"08",
          1194 => x"ff",
          1195 => x"72",
          1196 => x"08",
          1197 => x"82",
          1198 => x"e4",
          1199 => x"86",
          1200 => x"06",
          1201 => x"72",
          1202 => x"e7",
          1203 => x"84",
          1204 => x"22",
          1205 => x"82",
          1206 => x"cc",
          1207 => x"d5",
          1208 => x"05",
          1209 => x"82",
          1210 => x"cc",
          1211 => x"d5",
          1212 => x"05",
          1213 => x"72",
          1214 => x"81",
          1215 => x"82",
          1216 => x"cc",
          1217 => x"05",
          1218 => x"d5",
          1219 => x"05",
          1220 => x"82",
          1221 => x"cc",
          1222 => x"05",
          1223 => x"d5",
          1224 => x"05",
          1225 => x"84",
          1226 => x"22",
          1227 => x"08",
          1228 => x"82",
          1229 => x"e4",
          1230 => x"83",
          1231 => x"06",
          1232 => x"72",
          1233 => x"d0",
          1234 => x"84",
          1235 => x"33",
          1236 => x"70",
          1237 => x"d5",
          1238 => x"05",
          1239 => x"51",
          1240 => x"24",
          1241 => x"d5",
          1242 => x"05",
          1243 => x"06",
          1244 => x"82",
          1245 => x"e4",
          1246 => x"39",
          1247 => x"08",
          1248 => x"53",
          1249 => x"08",
          1250 => x"73",
          1251 => x"54",
          1252 => x"84",
          1253 => x"34",
          1254 => x"08",
          1255 => x"70",
          1256 => x"81",
          1257 => x"53",
          1258 => x"b1",
          1259 => x"84",
          1260 => x"33",
          1261 => x"70",
          1262 => x"90",
          1263 => x"2c",
          1264 => x"51",
          1265 => x"82",
          1266 => x"ec",
          1267 => x"75",
          1268 => x"72",
          1269 => x"08",
          1270 => x"af",
          1271 => x"84",
          1272 => x"33",
          1273 => x"70",
          1274 => x"90",
          1275 => x"2c",
          1276 => x"51",
          1277 => x"82",
          1278 => x"ec",
          1279 => x"75",
          1280 => x"72",
          1281 => x"08",
          1282 => x"82",
          1283 => x"e4",
          1284 => x"83",
          1285 => x"53",
          1286 => x"82",
          1287 => x"ec",
          1288 => x"11",
          1289 => x"82",
          1290 => x"ec",
          1291 => x"90",
          1292 => x"2c",
          1293 => x"73",
          1294 => x"82",
          1295 => x"88",
          1296 => x"a0",
          1297 => x"3f",
          1298 => x"d5",
          1299 => x"05",
          1300 => x"2a",
          1301 => x"51",
          1302 => x"80",
          1303 => x"82",
          1304 => x"88",
          1305 => x"ad",
          1306 => x"3f",
          1307 => x"82",
          1308 => x"e4",
          1309 => x"84",
          1310 => x"06",
          1311 => x"72",
          1312 => x"38",
          1313 => x"08",
          1314 => x"52",
          1315 => x"a5",
          1316 => x"82",
          1317 => x"e4",
          1318 => x"85",
          1319 => x"06",
          1320 => x"72",
          1321 => x"38",
          1322 => x"08",
          1323 => x"52",
          1324 => x"81",
          1325 => x"84",
          1326 => x"22",
          1327 => x"70",
          1328 => x"51",
          1329 => x"2e",
          1330 => x"d5",
          1331 => x"05",
          1332 => x"51",
          1333 => x"82",
          1334 => x"f4",
          1335 => x"72",
          1336 => x"81",
          1337 => x"82",
          1338 => x"88",
          1339 => x"82",
          1340 => x"f8",
          1341 => x"89",
          1342 => x"d5",
          1343 => x"05",
          1344 => x"2a",
          1345 => x"51",
          1346 => x"80",
          1347 => x"82",
          1348 => x"ec",
          1349 => x"11",
          1350 => x"82",
          1351 => x"ec",
          1352 => x"90",
          1353 => x"2c",
          1354 => x"73",
          1355 => x"82",
          1356 => x"88",
          1357 => x"b0",
          1358 => x"3f",
          1359 => x"d5",
          1360 => x"05",
          1361 => x"2a",
          1362 => x"51",
          1363 => x"80",
          1364 => x"82",
          1365 => x"e8",
          1366 => x"11",
          1367 => x"82",
          1368 => x"e8",
          1369 => x"98",
          1370 => x"2c",
          1371 => x"73",
          1372 => x"82",
          1373 => x"88",
          1374 => x"b0",
          1375 => x"3f",
          1376 => x"d5",
          1377 => x"05",
          1378 => x"2a",
          1379 => x"51",
          1380 => x"b0",
          1381 => x"84",
          1382 => x"22",
          1383 => x"54",
          1384 => x"84",
          1385 => x"23",
          1386 => x"70",
          1387 => x"53",
          1388 => x"90",
          1389 => x"84",
          1390 => x"08",
          1391 => x"87",
          1392 => x"39",
          1393 => x"08",
          1394 => x"53",
          1395 => x"2e",
          1396 => x"97",
          1397 => x"84",
          1398 => x"08",
          1399 => x"84",
          1400 => x"33",
          1401 => x"3f",
          1402 => x"82",
          1403 => x"f8",
          1404 => x"72",
          1405 => x"09",
          1406 => x"cb",
          1407 => x"84",
          1408 => x"22",
          1409 => x"53",
          1410 => x"84",
          1411 => x"23",
          1412 => x"ff",
          1413 => x"83",
          1414 => x"81",
          1415 => x"d5",
          1416 => x"05",
          1417 => x"d5",
          1418 => x"05",
          1419 => x"52",
          1420 => x"08",
          1421 => x"81",
          1422 => x"84",
          1423 => x"0c",
          1424 => x"3f",
          1425 => x"82",
          1426 => x"f8",
          1427 => x"72",
          1428 => x"09",
          1429 => x"cb",
          1430 => x"84",
          1431 => x"22",
          1432 => x"53",
          1433 => x"84",
          1434 => x"23",
          1435 => x"ff",
          1436 => x"83",
          1437 => x"80",
          1438 => x"d5",
          1439 => x"05",
          1440 => x"d5",
          1441 => x"05",
          1442 => x"52",
          1443 => x"3f",
          1444 => x"08",
          1445 => x"81",
          1446 => x"84",
          1447 => x"0c",
          1448 => x"82",
          1449 => x"f0",
          1450 => x"d5",
          1451 => x"38",
          1452 => x"08",
          1453 => x"52",
          1454 => x"08",
          1455 => x"ff",
          1456 => x"84",
          1457 => x"0c",
          1458 => x"08",
          1459 => x"70",
          1460 => x"85",
          1461 => x"39",
          1462 => x"08",
          1463 => x"70",
          1464 => x"81",
          1465 => x"53",
          1466 => x"80",
          1467 => x"d5",
          1468 => x"05",
          1469 => x"54",
          1470 => x"d5",
          1471 => x"05",
          1472 => x"2b",
          1473 => x"51",
          1474 => x"25",
          1475 => x"d5",
          1476 => x"05",
          1477 => x"51",
          1478 => x"d2",
          1479 => x"84",
          1480 => x"08",
          1481 => x"84",
          1482 => x"33",
          1483 => x"3f",
          1484 => x"d5",
          1485 => x"05",
          1486 => x"39",
          1487 => x"08",
          1488 => x"53",
          1489 => x"09",
          1490 => x"38",
          1491 => x"d5",
          1492 => x"05",
          1493 => x"82",
          1494 => x"ec",
          1495 => x"0b",
          1496 => x"08",
          1497 => x"8a",
          1498 => x"84",
          1499 => x"23",
          1500 => x"82",
          1501 => x"88",
          1502 => x"82",
          1503 => x"f8",
          1504 => x"84",
          1505 => x"ea",
          1506 => x"84",
          1507 => x"08",
          1508 => x"70",
          1509 => x"08",
          1510 => x"51",
          1511 => x"84",
          1512 => x"08",
          1513 => x"0c",
          1514 => x"82",
          1515 => x"04",
          1516 => x"08",
          1517 => x"84",
          1518 => x"0d",
          1519 => x"08",
          1520 => x"84",
          1521 => x"08",
          1522 => x"84",
          1523 => x"08",
          1524 => x"3f",
          1525 => x"08",
          1526 => x"f8",
          1527 => x"3d",
          1528 => x"84",
          1529 => x"d5",
          1530 => x"82",
          1531 => x"fb",
          1532 => x"0b",
          1533 => x"08",
          1534 => x"82",
          1535 => x"85",
          1536 => x"81",
          1537 => x"32",
          1538 => x"51",
          1539 => x"53",
          1540 => x"8d",
          1541 => x"82",
          1542 => x"f4",
          1543 => x"92",
          1544 => x"84",
          1545 => x"08",
          1546 => x"82",
          1547 => x"88",
          1548 => x"05",
          1549 => x"08",
          1550 => x"53",
          1551 => x"84",
          1552 => x"34",
          1553 => x"06",
          1554 => x"2e",
          1555 => x"f0",
          1556 => x"f0",
          1557 => x"82",
          1558 => x"fc",
          1559 => x"90",
          1560 => x"53",
          1561 => x"d4",
          1562 => x"72",
          1563 => x"b1",
          1564 => x"82",
          1565 => x"f8",
          1566 => x"a5",
          1567 => x"dc",
          1568 => x"dc",
          1569 => x"8a",
          1570 => x"08",
          1571 => x"82",
          1572 => x"53",
          1573 => x"8a",
          1574 => x"82",
          1575 => x"f8",
          1576 => x"d5",
          1577 => x"05",
          1578 => x"d5",
          1579 => x"05",
          1580 => x"d5",
          1581 => x"05",
          1582 => x"f8",
          1583 => x"0d",
          1584 => x"0c",
          1585 => x"84",
          1586 => x"d5",
          1587 => x"3d",
          1588 => x"82",
          1589 => x"f8",
          1590 => x"d5",
          1591 => x"05",
          1592 => x"33",
          1593 => x"70",
          1594 => x"81",
          1595 => x"51",
          1596 => x"80",
          1597 => x"ff",
          1598 => x"84",
          1599 => x"0c",
          1600 => x"82",
          1601 => x"88",
          1602 => x"72",
          1603 => x"84",
          1604 => x"08",
          1605 => x"d5",
          1606 => x"05",
          1607 => x"82",
          1608 => x"fc",
          1609 => x"81",
          1610 => x"72",
          1611 => x"38",
          1612 => x"08",
          1613 => x"82",
          1614 => x"8c",
          1615 => x"82",
          1616 => x"fc",
          1617 => x"90",
          1618 => x"53",
          1619 => x"d4",
          1620 => x"72",
          1621 => x"ab",
          1622 => x"82",
          1623 => x"f8",
          1624 => x"9f",
          1625 => x"84",
          1626 => x"08",
          1627 => x"84",
          1628 => x"0c",
          1629 => x"84",
          1630 => x"08",
          1631 => x"0c",
          1632 => x"82",
          1633 => x"04",
          1634 => x"08",
          1635 => x"84",
          1636 => x"0d",
          1637 => x"08",
          1638 => x"84",
          1639 => x"08",
          1640 => x"82",
          1641 => x"70",
          1642 => x"0c",
          1643 => x"0d",
          1644 => x"0c",
          1645 => x"84",
          1646 => x"d5",
          1647 => x"3d",
          1648 => x"84",
          1649 => x"08",
          1650 => x"70",
          1651 => x"81",
          1652 => x"06",
          1653 => x"51",
          1654 => x"2e",
          1655 => x"0b",
          1656 => x"08",
          1657 => x"81",
          1658 => x"d5",
          1659 => x"05",
          1660 => x"33",
          1661 => x"70",
          1662 => x"51",
          1663 => x"80",
          1664 => x"38",
          1665 => x"08",
          1666 => x"82",
          1667 => x"8c",
          1668 => x"54",
          1669 => x"88",
          1670 => x"9f",
          1671 => x"84",
          1672 => x"08",
          1673 => x"82",
          1674 => x"88",
          1675 => x"57",
          1676 => x"75",
          1677 => x"81",
          1678 => x"82",
          1679 => x"8c",
          1680 => x"11",
          1681 => x"8c",
          1682 => x"d5",
          1683 => x"05",
          1684 => x"d5",
          1685 => x"05",
          1686 => x"80",
          1687 => x"d5",
          1688 => x"05",
          1689 => x"84",
          1690 => x"08",
          1691 => x"84",
          1692 => x"08",
          1693 => x"06",
          1694 => x"08",
          1695 => x"72",
          1696 => x"f8",
          1697 => x"a3",
          1698 => x"84",
          1699 => x"08",
          1700 => x"81",
          1701 => x"0c",
          1702 => x"08",
          1703 => x"70",
          1704 => x"08",
          1705 => x"51",
          1706 => x"ff",
          1707 => x"84",
          1708 => x"0c",
          1709 => x"08",
          1710 => x"82",
          1711 => x"87",
          1712 => x"d5",
          1713 => x"82",
          1714 => x"02",
          1715 => x"0c",
          1716 => x"82",
          1717 => x"88",
          1718 => x"11",
          1719 => x"32",
          1720 => x"51",
          1721 => x"71",
          1722 => x"38",
          1723 => x"d5",
          1724 => x"05",
          1725 => x"39",
          1726 => x"08",
          1727 => x"85",
          1728 => x"86",
          1729 => x"06",
          1730 => x"52",
          1731 => x"80",
          1732 => x"d5",
          1733 => x"05",
          1734 => x"84",
          1735 => x"08",
          1736 => x"12",
          1737 => x"bf",
          1738 => x"71",
          1739 => x"82",
          1740 => x"88",
          1741 => x"11",
          1742 => x"8c",
          1743 => x"d5",
          1744 => x"05",
          1745 => x"33",
          1746 => x"84",
          1747 => x"0c",
          1748 => x"82",
          1749 => x"d5",
          1750 => x"05",
          1751 => x"33",
          1752 => x"70",
          1753 => x"51",
          1754 => x"80",
          1755 => x"38",
          1756 => x"08",
          1757 => x"70",
          1758 => x"82",
          1759 => x"fc",
          1760 => x"52",
          1761 => x"08",
          1762 => x"a9",
          1763 => x"84",
          1764 => x"08",
          1765 => x"08",
          1766 => x"53",
          1767 => x"33",
          1768 => x"51",
          1769 => x"14",
          1770 => x"82",
          1771 => x"f8",
          1772 => x"d7",
          1773 => x"84",
          1774 => x"08",
          1775 => x"05",
          1776 => x"81",
          1777 => x"d5",
          1778 => x"05",
          1779 => x"84",
          1780 => x"08",
          1781 => x"08",
          1782 => x"2d",
          1783 => x"08",
          1784 => x"84",
          1785 => x"0c",
          1786 => x"84",
          1787 => x"08",
          1788 => x"f2",
          1789 => x"84",
          1790 => x"08",
          1791 => x"08",
          1792 => x"82",
          1793 => x"88",
          1794 => x"11",
          1795 => x"84",
          1796 => x"0c",
          1797 => x"84",
          1798 => x"08",
          1799 => x"81",
          1800 => x"82",
          1801 => x"f0",
          1802 => x"07",
          1803 => x"d5",
          1804 => x"05",
          1805 => x"82",
          1806 => x"f0",
          1807 => x"07",
          1808 => x"d5",
          1809 => x"05",
          1810 => x"84",
          1811 => x"08",
          1812 => x"84",
          1813 => x"33",
          1814 => x"ff",
          1815 => x"84",
          1816 => x"0c",
          1817 => x"d5",
          1818 => x"05",
          1819 => x"08",
          1820 => x"12",
          1821 => x"84",
          1822 => x"08",
          1823 => x"06",
          1824 => x"84",
          1825 => x"0c",
          1826 => x"82",
          1827 => x"f8",
          1828 => x"d4",
          1829 => x"3d",
          1830 => x"84",
          1831 => x"d5",
          1832 => x"82",
          1833 => x"fd",
          1834 => x"d5",
          1835 => x"05",
          1836 => x"84",
          1837 => x"0c",
          1838 => x"08",
          1839 => x"82",
          1840 => x"f8",
          1841 => x"d5",
          1842 => x"05",
          1843 => x"82",
          1844 => x"d5",
          1845 => x"05",
          1846 => x"84",
          1847 => x"08",
          1848 => x"38",
          1849 => x"08",
          1850 => x"82",
          1851 => x"90",
          1852 => x"51",
          1853 => x"08",
          1854 => x"71",
          1855 => x"38",
          1856 => x"08",
          1857 => x"82",
          1858 => x"90",
          1859 => x"82",
          1860 => x"fc",
          1861 => x"d5",
          1862 => x"05",
          1863 => x"84",
          1864 => x"08",
          1865 => x"84",
          1866 => x"0c",
          1867 => x"08",
          1868 => x"81",
          1869 => x"84",
          1870 => x"0c",
          1871 => x"08",
          1872 => x"ff",
          1873 => x"84",
          1874 => x"0c",
          1875 => x"08",
          1876 => x"80",
          1877 => x"38",
          1878 => x"08",
          1879 => x"ff",
          1880 => x"84",
          1881 => x"0c",
          1882 => x"08",
          1883 => x"ff",
          1884 => x"84",
          1885 => x"0c",
          1886 => x"08",
          1887 => x"82",
          1888 => x"f8",
          1889 => x"51",
          1890 => x"34",
          1891 => x"82",
          1892 => x"90",
          1893 => x"05",
          1894 => x"08",
          1895 => x"82",
          1896 => x"90",
          1897 => x"05",
          1898 => x"08",
          1899 => x"82",
          1900 => x"90",
          1901 => x"2e",
          1902 => x"d5",
          1903 => x"05",
          1904 => x"33",
          1905 => x"08",
          1906 => x"81",
          1907 => x"84",
          1908 => x"0c",
          1909 => x"08",
          1910 => x"52",
          1911 => x"34",
          1912 => x"08",
          1913 => x"81",
          1914 => x"84",
          1915 => x"0c",
          1916 => x"82",
          1917 => x"88",
          1918 => x"82",
          1919 => x"51",
          1920 => x"82",
          1921 => x"04",
          1922 => x"08",
          1923 => x"84",
          1924 => x"0d",
          1925 => x"08",
          1926 => x"82",
          1927 => x"fc",
          1928 => x"d5",
          1929 => x"05",
          1930 => x"33",
          1931 => x"08",
          1932 => x"81",
          1933 => x"84",
          1934 => x"0c",
          1935 => x"06",
          1936 => x"80",
          1937 => x"da",
          1938 => x"84",
          1939 => x"08",
          1940 => x"d5",
          1941 => x"05",
          1942 => x"84",
          1943 => x"08",
          1944 => x"08",
          1945 => x"31",
          1946 => x"f8",
          1947 => x"3d",
          1948 => x"84",
          1949 => x"d5",
          1950 => x"82",
          1951 => x"fe",
          1952 => x"d5",
          1953 => x"05",
          1954 => x"84",
          1955 => x"0c",
          1956 => x"08",
          1957 => x"52",
          1958 => x"d5",
          1959 => x"05",
          1960 => x"82",
          1961 => x"8c",
          1962 => x"d5",
          1963 => x"05",
          1964 => x"70",
          1965 => x"d5",
          1966 => x"05",
          1967 => x"82",
          1968 => x"fc",
          1969 => x"81",
          1970 => x"70",
          1971 => x"38",
          1972 => x"82",
          1973 => x"88",
          1974 => x"82",
          1975 => x"51",
          1976 => x"82",
          1977 => x"04",
          1978 => x"08",
          1979 => x"84",
          1980 => x"0d",
          1981 => x"08",
          1982 => x"82",
          1983 => x"fc",
          1984 => x"d5",
          1985 => x"05",
          1986 => x"84",
          1987 => x"0c",
          1988 => x"08",
          1989 => x"80",
          1990 => x"38",
          1991 => x"08",
          1992 => x"81",
          1993 => x"84",
          1994 => x"0c",
          1995 => x"08",
          1996 => x"ff",
          1997 => x"84",
          1998 => x"0c",
          1999 => x"08",
          2000 => x"80",
          2001 => x"82",
          2002 => x"f8",
          2003 => x"70",
          2004 => x"84",
          2005 => x"08",
          2006 => x"d5",
          2007 => x"05",
          2008 => x"84",
          2009 => x"08",
          2010 => x"71",
          2011 => x"84",
          2012 => x"08",
          2013 => x"d5",
          2014 => x"05",
          2015 => x"39",
          2016 => x"08",
          2017 => x"70",
          2018 => x"0c",
          2019 => x"0d",
          2020 => x"0c",
          2021 => x"84",
          2022 => x"d5",
          2023 => x"3d",
          2024 => x"84",
          2025 => x"08",
          2026 => x"f4",
          2027 => x"84",
          2028 => x"08",
          2029 => x"82",
          2030 => x"8c",
          2031 => x"05",
          2032 => x"08",
          2033 => x"82",
          2034 => x"88",
          2035 => x"33",
          2036 => x"06",
          2037 => x"51",
          2038 => x"84",
          2039 => x"39",
          2040 => x"08",
          2041 => x"52",
          2042 => x"d5",
          2043 => x"05",
          2044 => x"82",
          2045 => x"88",
          2046 => x"81",
          2047 => x"51",
          2048 => x"80",
          2049 => x"84",
          2050 => x"0c",
          2051 => x"82",
          2052 => x"90",
          2053 => x"05",
          2054 => x"08",
          2055 => x"82",
          2056 => x"90",
          2057 => x"2e",
          2058 => x"81",
          2059 => x"84",
          2060 => x"08",
          2061 => x"e8",
          2062 => x"84",
          2063 => x"08",
          2064 => x"53",
          2065 => x"ff",
          2066 => x"84",
          2067 => x"0c",
          2068 => x"82",
          2069 => x"8c",
          2070 => x"05",
          2071 => x"08",
          2072 => x"82",
          2073 => x"8c",
          2074 => x"33",
          2075 => x"8c",
          2076 => x"82",
          2077 => x"fc",
          2078 => x"39",
          2079 => x"08",
          2080 => x"70",
          2081 => x"84",
          2082 => x"08",
          2083 => x"71",
          2084 => x"d5",
          2085 => x"05",
          2086 => x"52",
          2087 => x"39",
          2088 => x"d5",
          2089 => x"05",
          2090 => x"84",
          2091 => x"08",
          2092 => x"0c",
          2093 => x"82",
          2094 => x"04",
          2095 => x"08",
          2096 => x"84",
          2097 => x"0d",
          2098 => x"08",
          2099 => x"52",
          2100 => x"08",
          2101 => x"51",
          2102 => x"82",
          2103 => x"70",
          2104 => x"08",
          2105 => x"82",
          2106 => x"f8",
          2107 => x"05",
          2108 => x"54",
          2109 => x"3f",
          2110 => x"08",
          2111 => x"84",
          2112 => x"0c",
          2113 => x"84",
          2114 => x"08",
          2115 => x"0b",
          2116 => x"08",
          2117 => x"bc",
          2118 => x"84",
          2119 => x"08",
          2120 => x"08",
          2121 => x"05",
          2122 => x"34",
          2123 => x"08",
          2124 => x"53",
          2125 => x"08",
          2126 => x"52",
          2127 => x"08",
          2128 => x"51",
          2129 => x"82",
          2130 => x"70",
          2131 => x"08",
          2132 => x"54",
          2133 => x"08",
          2134 => x"82",
          2135 => x"88",
          2136 => x"d5",
          2137 => x"82",
          2138 => x"02",
          2139 => x"0c",
          2140 => x"82",
          2141 => x"88",
          2142 => x"d5",
          2143 => x"05",
          2144 => x"84",
          2145 => x"08",
          2146 => x"0b",
          2147 => x"08",
          2148 => x"80",
          2149 => x"d5",
          2150 => x"05",
          2151 => x"33",
          2152 => x"08",
          2153 => x"81",
          2154 => x"84",
          2155 => x"0c",
          2156 => x"06",
          2157 => x"80",
          2158 => x"82",
          2159 => x"8c",
          2160 => x"05",
          2161 => x"08",
          2162 => x"82",
          2163 => x"8c",
          2164 => x"2e",
          2165 => x"be",
          2166 => x"84",
          2167 => x"08",
          2168 => x"d5",
          2169 => x"05",
          2170 => x"84",
          2171 => x"08",
          2172 => x"08",
          2173 => x"31",
          2174 => x"84",
          2175 => x"0c",
          2176 => x"84",
          2177 => x"08",
          2178 => x"0c",
          2179 => x"82",
          2180 => x"04",
          2181 => x"08",
          2182 => x"84",
          2183 => x"0d",
          2184 => x"08",
          2185 => x"82",
          2186 => x"fc",
          2187 => x"d5",
          2188 => x"05",
          2189 => x"80",
          2190 => x"d5",
          2191 => x"05",
          2192 => x"82",
          2193 => x"90",
          2194 => x"d5",
          2195 => x"05",
          2196 => x"82",
          2197 => x"90",
          2198 => x"d5",
          2199 => x"05",
          2200 => x"a9",
          2201 => x"84",
          2202 => x"08",
          2203 => x"d5",
          2204 => x"05",
          2205 => x"71",
          2206 => x"d5",
          2207 => x"05",
          2208 => x"82",
          2209 => x"fc",
          2210 => x"be",
          2211 => x"84",
          2212 => x"08",
          2213 => x"f8",
          2214 => x"3d",
          2215 => x"84",
          2216 => x"d5",
          2217 => x"82",
          2218 => x"f9",
          2219 => x"0b",
          2220 => x"08",
          2221 => x"82",
          2222 => x"88",
          2223 => x"25",
          2224 => x"d5",
          2225 => x"05",
          2226 => x"d5",
          2227 => x"05",
          2228 => x"82",
          2229 => x"f4",
          2230 => x"d5",
          2231 => x"05",
          2232 => x"81",
          2233 => x"84",
          2234 => x"0c",
          2235 => x"08",
          2236 => x"82",
          2237 => x"fc",
          2238 => x"d5",
          2239 => x"05",
          2240 => x"b9",
          2241 => x"84",
          2242 => x"08",
          2243 => x"84",
          2244 => x"0c",
          2245 => x"d5",
          2246 => x"05",
          2247 => x"84",
          2248 => x"08",
          2249 => x"0b",
          2250 => x"08",
          2251 => x"82",
          2252 => x"f0",
          2253 => x"d5",
          2254 => x"05",
          2255 => x"82",
          2256 => x"8c",
          2257 => x"82",
          2258 => x"88",
          2259 => x"82",
          2260 => x"d4",
          2261 => x"82",
          2262 => x"f8",
          2263 => x"82",
          2264 => x"fc",
          2265 => x"2e",
          2266 => x"d5",
          2267 => x"05",
          2268 => x"d5",
          2269 => x"05",
          2270 => x"84",
          2271 => x"08",
          2272 => x"f8",
          2273 => x"3d",
          2274 => x"84",
          2275 => x"d5",
          2276 => x"82",
          2277 => x"fb",
          2278 => x"0b",
          2279 => x"08",
          2280 => x"82",
          2281 => x"88",
          2282 => x"25",
          2283 => x"d5",
          2284 => x"05",
          2285 => x"d5",
          2286 => x"05",
          2287 => x"82",
          2288 => x"fc",
          2289 => x"d5",
          2290 => x"05",
          2291 => x"90",
          2292 => x"84",
          2293 => x"08",
          2294 => x"84",
          2295 => x"0c",
          2296 => x"d5",
          2297 => x"05",
          2298 => x"d5",
          2299 => x"05",
          2300 => x"a2",
          2301 => x"f8",
          2302 => x"d5",
          2303 => x"05",
          2304 => x"d5",
          2305 => x"05",
          2306 => x"90",
          2307 => x"84",
          2308 => x"08",
          2309 => x"84",
          2310 => x"0c",
          2311 => x"08",
          2312 => x"70",
          2313 => x"0c",
          2314 => x"0d",
          2315 => x"0c",
          2316 => x"84",
          2317 => x"d5",
          2318 => x"3d",
          2319 => x"82",
          2320 => x"8c",
          2321 => x"82",
          2322 => x"88",
          2323 => x"80",
          2324 => x"d4",
          2325 => x"82",
          2326 => x"54",
          2327 => x"82",
          2328 => x"04",
          2329 => x"08",
          2330 => x"84",
          2331 => x"0d",
          2332 => x"d5",
          2333 => x"05",
          2334 => x"d5",
          2335 => x"05",
          2336 => x"3f",
          2337 => x"08",
          2338 => x"f8",
          2339 => x"3d",
          2340 => x"84",
          2341 => x"d5",
          2342 => x"82",
          2343 => x"fd",
          2344 => x"0b",
          2345 => x"08",
          2346 => x"80",
          2347 => x"84",
          2348 => x"0c",
          2349 => x"08",
          2350 => x"82",
          2351 => x"88",
          2352 => x"b9",
          2353 => x"84",
          2354 => x"08",
          2355 => x"38",
          2356 => x"d5",
          2357 => x"05",
          2358 => x"38",
          2359 => x"08",
          2360 => x"10",
          2361 => x"08",
          2362 => x"82",
          2363 => x"fc",
          2364 => x"82",
          2365 => x"fc",
          2366 => x"b8",
          2367 => x"84",
          2368 => x"08",
          2369 => x"e1",
          2370 => x"84",
          2371 => x"08",
          2372 => x"08",
          2373 => x"26",
          2374 => x"d5",
          2375 => x"05",
          2376 => x"84",
          2377 => x"08",
          2378 => x"84",
          2379 => x"0c",
          2380 => x"08",
          2381 => x"82",
          2382 => x"fc",
          2383 => x"82",
          2384 => x"f8",
          2385 => x"d5",
          2386 => x"05",
          2387 => x"82",
          2388 => x"fc",
          2389 => x"d5",
          2390 => x"05",
          2391 => x"82",
          2392 => x"8c",
          2393 => x"95",
          2394 => x"84",
          2395 => x"08",
          2396 => x"38",
          2397 => x"08",
          2398 => x"70",
          2399 => x"08",
          2400 => x"51",
          2401 => x"d5",
          2402 => x"05",
          2403 => x"d5",
          2404 => x"05",
          2405 => x"d5",
          2406 => x"05",
          2407 => x"f8",
          2408 => x"0d",
          2409 => x"0c",
          2410 => x"84",
          2411 => x"d5",
          2412 => x"3d",
          2413 => x"82",
          2414 => x"f0",
          2415 => x"d5",
          2416 => x"05",
          2417 => x"73",
          2418 => x"84",
          2419 => x"08",
          2420 => x"53",
          2421 => x"72",
          2422 => x"08",
          2423 => x"72",
          2424 => x"53",
          2425 => x"09",
          2426 => x"38",
          2427 => x"08",
          2428 => x"70",
          2429 => x"71",
          2430 => x"39",
          2431 => x"08",
          2432 => x"53",
          2433 => x"09",
          2434 => x"38",
          2435 => x"d5",
          2436 => x"05",
          2437 => x"84",
          2438 => x"08",
          2439 => x"05",
          2440 => x"08",
          2441 => x"33",
          2442 => x"08",
          2443 => x"82",
          2444 => x"f8",
          2445 => x"72",
          2446 => x"81",
          2447 => x"38",
          2448 => x"08",
          2449 => x"70",
          2450 => x"71",
          2451 => x"51",
          2452 => x"82",
          2453 => x"f8",
          2454 => x"d5",
          2455 => x"05",
          2456 => x"84",
          2457 => x"0c",
          2458 => x"08",
          2459 => x"80",
          2460 => x"38",
          2461 => x"08",
          2462 => x"80",
          2463 => x"38",
          2464 => x"90",
          2465 => x"84",
          2466 => x"34",
          2467 => x"08",
          2468 => x"70",
          2469 => x"71",
          2470 => x"51",
          2471 => x"82",
          2472 => x"f8",
          2473 => x"a4",
          2474 => x"82",
          2475 => x"f4",
          2476 => x"d5",
          2477 => x"05",
          2478 => x"81",
          2479 => x"70",
          2480 => x"72",
          2481 => x"84",
          2482 => x"34",
          2483 => x"82",
          2484 => x"f8",
          2485 => x"72",
          2486 => x"38",
          2487 => x"d5",
          2488 => x"05",
          2489 => x"39",
          2490 => x"08",
          2491 => x"53",
          2492 => x"90",
          2493 => x"84",
          2494 => x"33",
          2495 => x"26",
          2496 => x"39",
          2497 => x"d5",
          2498 => x"05",
          2499 => x"39",
          2500 => x"d5",
          2501 => x"05",
          2502 => x"82",
          2503 => x"f8",
          2504 => x"af",
          2505 => x"38",
          2506 => x"08",
          2507 => x"53",
          2508 => x"83",
          2509 => x"80",
          2510 => x"84",
          2511 => x"0c",
          2512 => x"8a",
          2513 => x"84",
          2514 => x"34",
          2515 => x"d5",
          2516 => x"05",
          2517 => x"84",
          2518 => x"33",
          2519 => x"27",
          2520 => x"82",
          2521 => x"f8",
          2522 => x"80",
          2523 => x"94",
          2524 => x"84",
          2525 => x"33",
          2526 => x"53",
          2527 => x"84",
          2528 => x"34",
          2529 => x"08",
          2530 => x"d0",
          2531 => x"72",
          2532 => x"08",
          2533 => x"82",
          2534 => x"f8",
          2535 => x"90",
          2536 => x"38",
          2537 => x"08",
          2538 => x"f9",
          2539 => x"72",
          2540 => x"08",
          2541 => x"82",
          2542 => x"f8",
          2543 => x"72",
          2544 => x"38",
          2545 => x"d5",
          2546 => x"05",
          2547 => x"39",
          2548 => x"08",
          2549 => x"82",
          2550 => x"f4",
          2551 => x"54",
          2552 => x"8d",
          2553 => x"82",
          2554 => x"ec",
          2555 => x"f7",
          2556 => x"84",
          2557 => x"33",
          2558 => x"84",
          2559 => x"08",
          2560 => x"84",
          2561 => x"33",
          2562 => x"d5",
          2563 => x"05",
          2564 => x"84",
          2565 => x"08",
          2566 => x"05",
          2567 => x"08",
          2568 => x"55",
          2569 => x"82",
          2570 => x"f8",
          2571 => x"a5",
          2572 => x"84",
          2573 => x"33",
          2574 => x"2e",
          2575 => x"d5",
          2576 => x"05",
          2577 => x"d5",
          2578 => x"05",
          2579 => x"84",
          2580 => x"08",
          2581 => x"08",
          2582 => x"71",
          2583 => x"0b",
          2584 => x"08",
          2585 => x"82",
          2586 => x"ec",
          2587 => x"d4",
          2588 => x"3d",
          2589 => x"84",
          2590 => x"d5",
          2591 => x"82",
          2592 => x"f7",
          2593 => x"0b",
          2594 => x"08",
          2595 => x"82",
          2596 => x"8c",
          2597 => x"80",
          2598 => x"d5",
          2599 => x"05",
          2600 => x"51",
          2601 => x"53",
          2602 => x"84",
          2603 => x"34",
          2604 => x"06",
          2605 => x"2e",
          2606 => x"91",
          2607 => x"84",
          2608 => x"08",
          2609 => x"05",
          2610 => x"ce",
          2611 => x"84",
          2612 => x"33",
          2613 => x"2e",
          2614 => x"a4",
          2615 => x"82",
          2616 => x"f0",
          2617 => x"d5",
          2618 => x"05",
          2619 => x"81",
          2620 => x"70",
          2621 => x"72",
          2622 => x"84",
          2623 => x"34",
          2624 => x"08",
          2625 => x"53",
          2626 => x"09",
          2627 => x"dc",
          2628 => x"84",
          2629 => x"08",
          2630 => x"05",
          2631 => x"08",
          2632 => x"33",
          2633 => x"08",
          2634 => x"82",
          2635 => x"f8",
          2636 => x"d5",
          2637 => x"05",
          2638 => x"84",
          2639 => x"08",
          2640 => x"b6",
          2641 => x"84",
          2642 => x"08",
          2643 => x"84",
          2644 => x"39",
          2645 => x"d5",
          2646 => x"05",
          2647 => x"84",
          2648 => x"08",
          2649 => x"05",
          2650 => x"08",
          2651 => x"33",
          2652 => x"08",
          2653 => x"81",
          2654 => x"0b",
          2655 => x"08",
          2656 => x"82",
          2657 => x"88",
          2658 => x"08",
          2659 => x"0c",
          2660 => x"53",
          2661 => x"d5",
          2662 => x"05",
          2663 => x"39",
          2664 => x"08",
          2665 => x"53",
          2666 => x"8d",
          2667 => x"82",
          2668 => x"ec",
          2669 => x"80",
          2670 => x"84",
          2671 => x"33",
          2672 => x"27",
          2673 => x"d5",
          2674 => x"05",
          2675 => x"b9",
          2676 => x"8d",
          2677 => x"82",
          2678 => x"ec",
          2679 => x"d8",
          2680 => x"82",
          2681 => x"f4",
          2682 => x"39",
          2683 => x"08",
          2684 => x"53",
          2685 => x"90",
          2686 => x"84",
          2687 => x"33",
          2688 => x"26",
          2689 => x"39",
          2690 => x"d5",
          2691 => x"05",
          2692 => x"39",
          2693 => x"d5",
          2694 => x"05",
          2695 => x"82",
          2696 => x"fc",
          2697 => x"d5",
          2698 => x"05",
          2699 => x"73",
          2700 => x"38",
          2701 => x"08",
          2702 => x"53",
          2703 => x"27",
          2704 => x"d5",
          2705 => x"05",
          2706 => x"51",
          2707 => x"d5",
          2708 => x"05",
          2709 => x"84",
          2710 => x"33",
          2711 => x"53",
          2712 => x"84",
          2713 => x"34",
          2714 => x"08",
          2715 => x"53",
          2716 => x"ad",
          2717 => x"84",
          2718 => x"33",
          2719 => x"53",
          2720 => x"84",
          2721 => x"34",
          2722 => x"08",
          2723 => x"53",
          2724 => x"8d",
          2725 => x"82",
          2726 => x"ec",
          2727 => x"98",
          2728 => x"84",
          2729 => x"33",
          2730 => x"08",
          2731 => x"54",
          2732 => x"26",
          2733 => x"0b",
          2734 => x"08",
          2735 => x"80",
          2736 => x"d5",
          2737 => x"05",
          2738 => x"d5",
          2739 => x"05",
          2740 => x"d5",
          2741 => x"05",
          2742 => x"82",
          2743 => x"fc",
          2744 => x"d5",
          2745 => x"05",
          2746 => x"81",
          2747 => x"70",
          2748 => x"52",
          2749 => x"33",
          2750 => x"08",
          2751 => x"fe",
          2752 => x"d5",
          2753 => x"05",
          2754 => x"80",
          2755 => x"82",
          2756 => x"fc",
          2757 => x"82",
          2758 => x"fc",
          2759 => x"d5",
          2760 => x"05",
          2761 => x"84",
          2762 => x"08",
          2763 => x"81",
          2764 => x"84",
          2765 => x"0c",
          2766 => x"08",
          2767 => x"82",
          2768 => x"8b",
          2769 => x"d5",
          2770 => x"f8",
          2771 => x"70",
          2772 => x"56",
          2773 => x"2e",
          2774 => x"8c",
          2775 => x"79",
          2776 => x"33",
          2777 => x"39",
          2778 => x"73",
          2779 => x"81",
          2780 => x"81",
          2781 => x"39",
          2782 => x"90",
          2783 => x"f8",
          2784 => x"52",
          2785 => x"3f",
          2786 => x"08",
          2787 => x"08",
          2788 => x"76",
          2789 => x"e7",
          2790 => x"d4",
          2791 => x"38",
          2792 => x"54",
          2793 => x"ff",
          2794 => x"17",
          2795 => x"06",
          2796 => x"77",
          2797 => x"ff",
          2798 => x"d4",
          2799 => x"3d",
          2800 => x"3d",
          2801 => x"71",
          2802 => x"8e",
          2803 => x"29",
          2804 => x"05",
          2805 => x"04",
          2806 => x"51",
          2807 => x"82",
          2808 => x"80",
          2809 => x"b2",
          2810 => x"f2",
          2811 => x"b4",
          2812 => x"39",
          2813 => x"51",
          2814 => x"82",
          2815 => x"80",
          2816 => x"b2",
          2817 => x"d6",
          2818 => x"f8",
          2819 => x"39",
          2820 => x"51",
          2821 => x"82",
          2822 => x"80",
          2823 => x"b3",
          2824 => x"39",
          2825 => x"51",
          2826 => x"b3",
          2827 => x"39",
          2828 => x"51",
          2829 => x"b4",
          2830 => x"39",
          2831 => x"51",
          2832 => x"b4",
          2833 => x"39",
          2834 => x"51",
          2835 => x"b5",
          2836 => x"39",
          2837 => x"51",
          2838 => x"b5",
          2839 => x"86",
          2840 => x"0d",
          2841 => x"0d",
          2842 => x"56",
          2843 => x"26",
          2844 => x"52",
          2845 => x"29",
          2846 => x"87",
          2847 => x"51",
          2848 => x"82",
          2849 => x"52",
          2850 => x"a5",
          2851 => x"f8",
          2852 => x"53",
          2853 => x"b5",
          2854 => x"ba",
          2855 => x"3d",
          2856 => x"3d",
          2857 => x"84",
          2858 => x"05",
          2859 => x"80",
          2860 => x"70",
          2861 => x"25",
          2862 => x"59",
          2863 => x"87",
          2864 => x"38",
          2865 => x"76",
          2866 => x"ff",
          2867 => x"93",
          2868 => x"82",
          2869 => x"76",
          2870 => x"70",
          2871 => x"92",
          2872 => x"d4",
          2873 => x"82",
          2874 => x"b9",
          2875 => x"f8",
          2876 => x"98",
          2877 => x"d4",
          2878 => x"96",
          2879 => x"54",
          2880 => x"77",
          2881 => x"81",
          2882 => x"82",
          2883 => x"57",
          2884 => x"08",
          2885 => x"55",
          2886 => x"89",
          2887 => x"75",
          2888 => x"d7",
          2889 => x"d8",
          2890 => x"9e",
          2891 => x"30",
          2892 => x"80",
          2893 => x"70",
          2894 => x"06",
          2895 => x"56",
          2896 => x"90",
          2897 => x"e0",
          2898 => x"98",
          2899 => x"78",
          2900 => x"3f",
          2901 => x"82",
          2902 => x"96",
          2903 => x"f7",
          2904 => x"02",
          2905 => x"05",
          2906 => x"ff",
          2907 => x"7c",
          2908 => x"fe",
          2909 => x"d4",
          2910 => x"cb",
          2911 => x"2e",
          2912 => x"81",
          2913 => x"bf",
          2914 => x"d8",
          2915 => x"d8",
          2916 => x"d8",
          2917 => x"e0",
          2918 => x"f0",
          2919 => x"82",
          2920 => x"52",
          2921 => x"51",
          2922 => x"3f",
          2923 => x"56",
          2924 => x"54",
          2925 => x"53",
          2926 => x"51",
          2927 => x"d4",
          2928 => x"83",
          2929 => x"78",
          2930 => x"0c",
          2931 => x"04",
          2932 => x"7f",
          2933 => x"8c",
          2934 => x"05",
          2935 => x"15",
          2936 => x"5c",
          2937 => x"5e",
          2938 => x"b6",
          2939 => x"b7",
          2940 => x"b6",
          2941 => x"b7",
          2942 => x"55",
          2943 => x"81",
          2944 => x"90",
          2945 => x"7b",
          2946 => x"38",
          2947 => x"74",
          2948 => x"7a",
          2949 => x"72",
          2950 => x"b6",
          2951 => x"b7",
          2952 => x"39",
          2953 => x"51",
          2954 => x"3f",
          2955 => x"80",
          2956 => x"18",
          2957 => x"27",
          2958 => x"08",
          2959 => x"9c",
          2960 => x"97",
          2961 => x"82",
          2962 => x"ff",
          2963 => x"84",
          2964 => x"39",
          2965 => x"72",
          2966 => x"38",
          2967 => x"82",
          2968 => x"ff",
          2969 => x"89",
          2970 => x"c4",
          2971 => x"eb",
          2972 => x"55",
          2973 => x"08",
          2974 => x"d6",
          2975 => x"fc",
          2976 => x"c8",
          2977 => x"d3",
          2978 => x"74",
          2979 => x"c6",
          2980 => x"70",
          2981 => x"80",
          2982 => x"27",
          2983 => x"56",
          2984 => x"74",
          2985 => x"81",
          2986 => x"06",
          2987 => x"06",
          2988 => x"80",
          2989 => x"73",
          2990 => x"8a",
          2991 => x"dc",
          2992 => x"51",
          2993 => x"f0",
          2994 => x"a0",
          2995 => x"3f",
          2996 => x"ff",
          2997 => x"b6",
          2998 => x"8a",
          2999 => x"79",
          3000 => x"9d",
          3001 => x"d4",
          3002 => x"2b",
          3003 => x"51",
          3004 => x"2e",
          3005 => x"aa",
          3006 => x"3f",
          3007 => x"08",
          3008 => x"98",
          3009 => x"32",
          3010 => x"9b",
          3011 => x"70",
          3012 => x"75",
          3013 => x"58",
          3014 => x"51",
          3015 => x"24",
          3016 => x"9b",
          3017 => x"06",
          3018 => x"53",
          3019 => x"1e",
          3020 => x"26",
          3021 => x"ff",
          3022 => x"d4",
          3023 => x"3d",
          3024 => x"3d",
          3025 => x"05",
          3026 => x"d0",
          3027 => x"d4",
          3028 => x"b5",
          3029 => x"d3",
          3030 => x"a6",
          3031 => x"b6",
          3032 => x"b6",
          3033 => x"d3",
          3034 => x"82",
          3035 => x"ff",
          3036 => x"74",
          3037 => x"38",
          3038 => x"86",
          3039 => x"fe",
          3040 => x"c0",
          3041 => x"53",
          3042 => x"81",
          3043 => x"3f",
          3044 => x"51",
          3045 => x"80",
          3046 => x"3f",
          3047 => x"70",
          3048 => x"52",
          3049 => x"92",
          3050 => x"98",
          3051 => x"b7",
          3052 => x"f7",
          3053 => x"98",
          3054 => x"82",
          3055 => x"06",
          3056 => x"80",
          3057 => x"81",
          3058 => x"3f",
          3059 => x"51",
          3060 => x"80",
          3061 => x"3f",
          3062 => x"70",
          3063 => x"52",
          3064 => x"92",
          3065 => x"98",
          3066 => x"b7",
          3067 => x"bb",
          3068 => x"98",
          3069 => x"84",
          3070 => x"06",
          3071 => x"80",
          3072 => x"81",
          3073 => x"3f",
          3074 => x"51",
          3075 => x"80",
          3076 => x"3f",
          3077 => x"70",
          3078 => x"52",
          3079 => x"92",
          3080 => x"97",
          3081 => x"b7",
          3082 => x"ff",
          3083 => x"97",
          3084 => x"86",
          3085 => x"06",
          3086 => x"80",
          3087 => x"81",
          3088 => x"3f",
          3089 => x"51",
          3090 => x"80",
          3091 => x"3f",
          3092 => x"70",
          3093 => x"52",
          3094 => x"92",
          3095 => x"97",
          3096 => x"b8",
          3097 => x"c3",
          3098 => x"97",
          3099 => x"88",
          3100 => x"06",
          3101 => x"80",
          3102 => x"81",
          3103 => x"3f",
          3104 => x"51",
          3105 => x"80",
          3106 => x"3f",
          3107 => x"84",
          3108 => x"fb",
          3109 => x"02",
          3110 => x"05",
          3111 => x"56",
          3112 => x"75",
          3113 => x"3f",
          3114 => x"cf",
          3115 => x"73",
          3116 => x"53",
          3117 => x"52",
          3118 => x"51",
          3119 => x"3f",
          3120 => x"08",
          3121 => x"d4",
          3122 => x"80",
          3123 => x"31",
          3124 => x"73",
          3125 => x"cf",
          3126 => x"0b",
          3127 => x"33",
          3128 => x"2e",
          3129 => x"af",
          3130 => x"88",
          3131 => x"75",
          3132 => x"ff",
          3133 => x"f8",
          3134 => x"8b",
          3135 => x"f8",
          3136 => x"e2",
          3137 => x"82",
          3138 => x"81",
          3139 => x"82",
          3140 => x"82",
          3141 => x"0b",
          3142 => x"f4",
          3143 => x"82",
          3144 => x"06",
          3145 => x"b8",
          3146 => x"52",
          3147 => x"ae",
          3148 => x"82",
          3149 => x"87",
          3150 => x"cd",
          3151 => x"70",
          3152 => x"7e",
          3153 => x"0c",
          3154 => x"7d",
          3155 => x"c6",
          3156 => x"f8",
          3157 => x"06",
          3158 => x"2e",
          3159 => x"a3",
          3160 => x"59",
          3161 => x"b9",
          3162 => x"51",
          3163 => x"7d",
          3164 => x"82",
          3165 => x"81",
          3166 => x"82",
          3167 => x"7e",
          3168 => x"82",
          3169 => x"8d",
          3170 => x"70",
          3171 => x"b9",
          3172 => x"b0",
          3173 => x"3d",
          3174 => x"80",
          3175 => x"51",
          3176 => x"b5",
          3177 => x"05",
          3178 => x"3f",
          3179 => x"08",
          3180 => x"90",
          3181 => x"78",
          3182 => x"87",
          3183 => x"80",
          3184 => x"38",
          3185 => x"81",
          3186 => x"bd",
          3187 => x"78",
          3188 => x"ba",
          3189 => x"2e",
          3190 => x"8a",
          3191 => x"80",
          3192 => x"99",
          3193 => x"c0",
          3194 => x"38",
          3195 => x"82",
          3196 => x"bf",
          3197 => x"f9",
          3198 => x"38",
          3199 => x"24",
          3200 => x"80",
          3201 => x"8a",
          3202 => x"f8",
          3203 => x"38",
          3204 => x"78",
          3205 => x"8a",
          3206 => x"81",
          3207 => x"38",
          3208 => x"2e",
          3209 => x"8a",
          3210 => x"81",
          3211 => x"fd",
          3212 => x"39",
          3213 => x"80",
          3214 => x"84",
          3215 => x"ba",
          3216 => x"f8",
          3217 => x"fe",
          3218 => x"3d",
          3219 => x"53",
          3220 => x"51",
          3221 => x"82",
          3222 => x"80",
          3223 => x"38",
          3224 => x"f8",
          3225 => x"84",
          3226 => x"8e",
          3227 => x"f8",
          3228 => x"82",
          3229 => x"43",
          3230 => x"51",
          3231 => x"3f",
          3232 => x"5a",
          3233 => x"81",
          3234 => x"59",
          3235 => x"84",
          3236 => x"7a",
          3237 => x"38",
          3238 => x"b5",
          3239 => x"11",
          3240 => x"05",
          3241 => x"3f",
          3242 => x"08",
          3243 => x"de",
          3244 => x"fe",
          3245 => x"ff",
          3246 => x"eb",
          3247 => x"d4",
          3248 => x"2e",
          3249 => x"b5",
          3250 => x"11",
          3251 => x"05",
          3252 => x"3f",
          3253 => x"08",
          3254 => x"b2",
          3255 => x"d0",
          3256 => x"f7",
          3257 => x"79",
          3258 => x"89",
          3259 => x"79",
          3260 => x"5b",
          3261 => x"62",
          3262 => x"eb",
          3263 => x"ff",
          3264 => x"ff",
          3265 => x"ea",
          3266 => x"d4",
          3267 => x"2e",
          3268 => x"b5",
          3269 => x"11",
          3270 => x"05",
          3271 => x"3f",
          3272 => x"08",
          3273 => x"e6",
          3274 => x"fe",
          3275 => x"ff",
          3276 => x"ea",
          3277 => x"d4",
          3278 => x"2e",
          3279 => x"82",
          3280 => x"ff",
          3281 => x"64",
          3282 => x"27",
          3283 => x"70",
          3284 => x"5e",
          3285 => x"7c",
          3286 => x"78",
          3287 => x"79",
          3288 => x"52",
          3289 => x"51",
          3290 => x"3f",
          3291 => x"81",
          3292 => x"d5",
          3293 => x"cc",
          3294 => x"92",
          3295 => x"ff",
          3296 => x"ff",
          3297 => x"e9",
          3298 => x"d4",
          3299 => x"df",
          3300 => x"e4",
          3301 => x"80",
          3302 => x"82",
          3303 => x"45",
          3304 => x"82",
          3305 => x"59",
          3306 => x"88",
          3307 => x"a4",
          3308 => x"39",
          3309 => x"33",
          3310 => x"2e",
          3311 => x"d3",
          3312 => x"ab",
          3313 => x"e7",
          3314 => x"80",
          3315 => x"82",
          3316 => x"45",
          3317 => x"d3",
          3318 => x"78",
          3319 => x"38",
          3320 => x"08",
          3321 => x"82",
          3322 => x"fc",
          3323 => x"b5",
          3324 => x"11",
          3325 => x"05",
          3326 => x"3f",
          3327 => x"08",
          3328 => x"82",
          3329 => x"59",
          3330 => x"89",
          3331 => x"a0",
          3332 => x"cc",
          3333 => x"e5",
          3334 => x"80",
          3335 => x"82",
          3336 => x"44",
          3337 => x"d3",
          3338 => x"78",
          3339 => x"38",
          3340 => x"08",
          3341 => x"82",
          3342 => x"59",
          3343 => x"88",
          3344 => x"b8",
          3345 => x"39",
          3346 => x"33",
          3347 => x"2e",
          3348 => x"d3",
          3349 => x"88",
          3350 => x"cc",
          3351 => x"44",
          3352 => x"f8",
          3353 => x"84",
          3354 => x"8e",
          3355 => x"f8",
          3356 => x"a7",
          3357 => x"5c",
          3358 => x"2e",
          3359 => x"5c",
          3360 => x"70",
          3361 => x"07",
          3362 => x"7f",
          3363 => x"5a",
          3364 => x"2e",
          3365 => x"a0",
          3366 => x"88",
          3367 => x"88",
          3368 => x"3f",
          3369 => x"54",
          3370 => x"52",
          3371 => x"a0",
          3372 => x"94",
          3373 => x"39",
          3374 => x"80",
          3375 => x"84",
          3376 => x"b6",
          3377 => x"f8",
          3378 => x"f9",
          3379 => x"3d",
          3380 => x"53",
          3381 => x"51",
          3382 => x"82",
          3383 => x"80",
          3384 => x"64",
          3385 => x"cf",
          3386 => x"34",
          3387 => x"45",
          3388 => x"fc",
          3389 => x"84",
          3390 => x"fe",
          3391 => x"f8",
          3392 => x"f9",
          3393 => x"70",
          3394 => x"82",
          3395 => x"ff",
          3396 => x"82",
          3397 => x"53",
          3398 => x"79",
          3399 => x"90",
          3400 => x"79",
          3401 => x"ae",
          3402 => x"38",
          3403 => x"9f",
          3404 => x"fe",
          3405 => x"ff",
          3406 => x"e6",
          3407 => x"d4",
          3408 => x"2e",
          3409 => x"59",
          3410 => x"05",
          3411 => x"64",
          3412 => x"ff",
          3413 => x"ba",
          3414 => x"8a",
          3415 => x"39",
          3416 => x"f4",
          3417 => x"84",
          3418 => x"bd",
          3419 => x"f8",
          3420 => x"f8",
          3421 => x"3d",
          3422 => x"53",
          3423 => x"51",
          3424 => x"82",
          3425 => x"80",
          3426 => x"61",
          3427 => x"c2",
          3428 => x"70",
          3429 => x"23",
          3430 => x"3d",
          3431 => x"53",
          3432 => x"51",
          3433 => x"82",
          3434 => x"df",
          3435 => x"39",
          3436 => x"54",
          3437 => x"b0",
          3438 => x"9f",
          3439 => x"d8",
          3440 => x"f8",
          3441 => x"ff",
          3442 => x"79",
          3443 => x"59",
          3444 => x"f7",
          3445 => x"9f",
          3446 => x"61",
          3447 => x"d0",
          3448 => x"fe",
          3449 => x"ff",
          3450 => x"df",
          3451 => x"d4",
          3452 => x"2e",
          3453 => x"59",
          3454 => x"05",
          3455 => x"82",
          3456 => x"78",
          3457 => x"39",
          3458 => x"51",
          3459 => x"ff",
          3460 => x"3d",
          3461 => x"53",
          3462 => x"51",
          3463 => x"82",
          3464 => x"80",
          3465 => x"38",
          3466 => x"f0",
          3467 => x"84",
          3468 => x"f5",
          3469 => x"f8",
          3470 => x"a0",
          3471 => x"71",
          3472 => x"84",
          3473 => x"3d",
          3474 => x"53",
          3475 => x"51",
          3476 => x"82",
          3477 => x"e5",
          3478 => x"39",
          3479 => x"54",
          3480 => x"bc",
          3481 => x"f3",
          3482 => x"d8",
          3483 => x"f8",
          3484 => x"ff",
          3485 => x"79",
          3486 => x"59",
          3487 => x"f6",
          3488 => x"79",
          3489 => x"b5",
          3490 => x"11",
          3491 => x"05",
          3492 => x"3f",
          3493 => x"08",
          3494 => x"38",
          3495 => x"0c",
          3496 => x"05",
          3497 => x"39",
          3498 => x"51",
          3499 => x"ff",
          3500 => x"3d",
          3501 => x"53",
          3502 => x"51",
          3503 => x"82",
          3504 => x"80",
          3505 => x"38",
          3506 => x"ba",
          3507 => x"a6",
          3508 => x"59",
          3509 => x"3d",
          3510 => x"53",
          3511 => x"51",
          3512 => x"82",
          3513 => x"80",
          3514 => x"38",
          3515 => x"ba",
          3516 => x"a5",
          3517 => x"59",
          3518 => x"d4",
          3519 => x"2e",
          3520 => x"82",
          3521 => x"52",
          3522 => x"51",
          3523 => x"3f",
          3524 => x"82",
          3525 => x"c1",
          3526 => x"a5",
          3527 => x"ee",
          3528 => x"bc",
          3529 => x"3f",
          3530 => x"a8",
          3531 => x"3f",
          3532 => x"97",
          3533 => x"78",
          3534 => x"d2",
          3535 => x"52",
          3536 => x"f8",
          3537 => x"f8",
          3538 => x"d4",
          3539 => x"2e",
          3540 => x"82",
          3541 => x"46",
          3542 => x"84",
          3543 => x"a8",
          3544 => x"f8",
          3545 => x"06",
          3546 => x"80",
          3547 => x"38",
          3548 => x"08",
          3549 => x"3f",
          3550 => x"08",
          3551 => x"c1",
          3552 => x"7a",
          3553 => x"38",
          3554 => x"89",
          3555 => x"2e",
          3556 => x"ca",
          3557 => x"2e",
          3558 => x"c2",
          3559 => x"d0",
          3560 => x"82",
          3561 => x"80",
          3562 => x"d8",
          3563 => x"ff",
          3564 => x"ff",
          3565 => x"b8",
          3566 => x"b5",
          3567 => x"05",
          3568 => x"3f",
          3569 => x"55",
          3570 => x"54",
          3571 => x"bb",
          3572 => x"3d",
          3573 => x"51",
          3574 => x"3f",
          3575 => x"54",
          3576 => x"bb",
          3577 => x"3d",
          3578 => x"51",
          3579 => x"3f",
          3580 => x"58",
          3581 => x"57",
          3582 => x"55",
          3583 => x"80",
          3584 => x"80",
          3585 => x"3d",
          3586 => x"51",
          3587 => x"82",
          3588 => x"82",
          3589 => x"09",
          3590 => x"72",
          3591 => x"51",
          3592 => x"80",
          3593 => x"26",
          3594 => x"5a",
          3595 => x"59",
          3596 => x"8d",
          3597 => x"70",
          3598 => x"5c",
          3599 => x"c3",
          3600 => x"32",
          3601 => x"07",
          3602 => x"38",
          3603 => x"09",
          3604 => x"38",
          3605 => x"51",
          3606 => x"3f",
          3607 => x"b3",
          3608 => x"39",
          3609 => x"51",
          3610 => x"3f",
          3611 => x"f6",
          3612 => x"0b",
          3613 => x"34",
          3614 => x"8c",
          3615 => x"84",
          3616 => x"51",
          3617 => x"82",
          3618 => x"90",
          3619 => x"94",
          3620 => x"53",
          3621 => x"52",
          3622 => x"95",
          3623 => x"d4",
          3624 => x"87",
          3625 => x"0c",
          3626 => x"9c",
          3627 => x"84",
          3628 => x"51",
          3629 => x"82",
          3630 => x"90",
          3631 => x"94",
          3632 => x"53",
          3633 => x"52",
          3634 => x"e5",
          3635 => x"d4",
          3636 => x"87",
          3637 => x"0c",
          3638 => x"0b",
          3639 => x"84",
          3640 => x"83",
          3641 => x"94",
          3642 => x"80",
          3643 => x"88",
          3644 => x"70",
          3645 => x"0c",
          3646 => x"fe",
          3647 => x"38",
          3648 => x"53",
          3649 => x"b0",
          3650 => x"84",
          3651 => x"87",
          3652 => x"73",
          3653 => x"80",
          3654 => x"80",
          3655 => x"83",
          3656 => x"95",
          3657 => x"5b",
          3658 => x"82",
          3659 => x"70",
          3660 => x"0c",
          3661 => x"0c",
          3662 => x"92",
          3663 => x"bc",
          3664 => x"bd",
          3665 => x"bc",
          3666 => x"bd",
          3667 => x"de",
          3668 => x"e3",
          3669 => x"eb",
          3670 => x"df",
          3671 => x"fe",
          3672 => x"52",
          3673 => x"88",
          3674 => x"d8",
          3675 => x"f8",
          3676 => x"06",
          3677 => x"14",
          3678 => x"80",
          3679 => x"71",
          3680 => x"0c",
          3681 => x"04",
          3682 => x"76",
          3683 => x"55",
          3684 => x"54",
          3685 => x"81",
          3686 => x"33",
          3687 => x"2e",
          3688 => x"86",
          3689 => x"53",
          3690 => x"33",
          3691 => x"2e",
          3692 => x"86",
          3693 => x"53",
          3694 => x"52",
          3695 => x"09",
          3696 => x"38",
          3697 => x"12",
          3698 => x"33",
          3699 => x"a2",
          3700 => x"81",
          3701 => x"2e",
          3702 => x"ea",
          3703 => x"81",
          3704 => x"72",
          3705 => x"70",
          3706 => x"38",
          3707 => x"80",
          3708 => x"73",
          3709 => x"72",
          3710 => x"70",
          3711 => x"81",
          3712 => x"81",
          3713 => x"32",
          3714 => x"80",
          3715 => x"51",
          3716 => x"80",
          3717 => x"80",
          3718 => x"05",
          3719 => x"75",
          3720 => x"70",
          3721 => x"0c",
          3722 => x"04",
          3723 => x"76",
          3724 => x"80",
          3725 => x"86",
          3726 => x"52",
          3727 => x"e9",
          3728 => x"f8",
          3729 => x"80",
          3730 => x"74",
          3731 => x"d4",
          3732 => x"3d",
          3733 => x"3d",
          3734 => x"11",
          3735 => x"52",
          3736 => x"70",
          3737 => x"98",
          3738 => x"33",
          3739 => x"82",
          3740 => x"26",
          3741 => x"84",
          3742 => x"83",
          3743 => x"26",
          3744 => x"85",
          3745 => x"84",
          3746 => x"26",
          3747 => x"86",
          3748 => x"85",
          3749 => x"26",
          3750 => x"88",
          3751 => x"86",
          3752 => x"e7",
          3753 => x"38",
          3754 => x"54",
          3755 => x"87",
          3756 => x"cc",
          3757 => x"87",
          3758 => x"0c",
          3759 => x"c0",
          3760 => x"82",
          3761 => x"c0",
          3762 => x"83",
          3763 => x"c0",
          3764 => x"84",
          3765 => x"c0",
          3766 => x"85",
          3767 => x"c0",
          3768 => x"86",
          3769 => x"c0",
          3770 => x"74",
          3771 => x"a4",
          3772 => x"c0",
          3773 => x"80",
          3774 => x"98",
          3775 => x"52",
          3776 => x"f8",
          3777 => x"0d",
          3778 => x"0d",
          3779 => x"c0",
          3780 => x"81",
          3781 => x"c0",
          3782 => x"5e",
          3783 => x"87",
          3784 => x"08",
          3785 => x"1c",
          3786 => x"98",
          3787 => x"79",
          3788 => x"87",
          3789 => x"08",
          3790 => x"1c",
          3791 => x"98",
          3792 => x"79",
          3793 => x"87",
          3794 => x"08",
          3795 => x"1c",
          3796 => x"98",
          3797 => x"7b",
          3798 => x"87",
          3799 => x"08",
          3800 => x"1c",
          3801 => x"0c",
          3802 => x"ff",
          3803 => x"83",
          3804 => x"58",
          3805 => x"57",
          3806 => x"56",
          3807 => x"55",
          3808 => x"54",
          3809 => x"53",
          3810 => x"ff",
          3811 => x"bc",
          3812 => x"9c",
          3813 => x"3d",
          3814 => x"3d",
          3815 => x"05",
          3816 => x"98",
          3817 => x"ff",
          3818 => x"55",
          3819 => x"84",
          3820 => x"2e",
          3821 => x"c0",
          3822 => x"70",
          3823 => x"2a",
          3824 => x"53",
          3825 => x"80",
          3826 => x"71",
          3827 => x"81",
          3828 => x"70",
          3829 => x"81",
          3830 => x"06",
          3831 => x"80",
          3832 => x"71",
          3833 => x"81",
          3834 => x"70",
          3835 => x"73",
          3836 => x"51",
          3837 => x"80",
          3838 => x"2e",
          3839 => x"c0",
          3840 => x"74",
          3841 => x"82",
          3842 => x"87",
          3843 => x"ff",
          3844 => x"8f",
          3845 => x"30",
          3846 => x"51",
          3847 => x"82",
          3848 => x"83",
          3849 => x"f9",
          3850 => x"a7",
          3851 => x"77",
          3852 => x"81",
          3853 => x"7a",
          3854 => x"eb",
          3855 => x"98",
          3856 => x"ff",
          3857 => x"87",
          3858 => x"53",
          3859 => x"86",
          3860 => x"94",
          3861 => x"08",
          3862 => x"70",
          3863 => x"56",
          3864 => x"2e",
          3865 => x"91",
          3866 => x"06",
          3867 => x"d7",
          3868 => x"32",
          3869 => x"51",
          3870 => x"2e",
          3871 => x"93",
          3872 => x"06",
          3873 => x"ff",
          3874 => x"81",
          3875 => x"87",
          3876 => x"54",
          3877 => x"86",
          3878 => x"94",
          3879 => x"74",
          3880 => x"82",
          3881 => x"89",
          3882 => x"f9",
          3883 => x"54",
          3884 => x"70",
          3885 => x"53",
          3886 => x"77",
          3887 => x"38",
          3888 => x"06",
          3889 => x"d3",
          3890 => x"81",
          3891 => x"57",
          3892 => x"c0",
          3893 => x"75",
          3894 => x"38",
          3895 => x"94",
          3896 => x"70",
          3897 => x"81",
          3898 => x"52",
          3899 => x"8c",
          3900 => x"2a",
          3901 => x"51",
          3902 => x"38",
          3903 => x"70",
          3904 => x"51",
          3905 => x"8d",
          3906 => x"2a",
          3907 => x"51",
          3908 => x"be",
          3909 => x"ff",
          3910 => x"c0",
          3911 => x"70",
          3912 => x"38",
          3913 => x"90",
          3914 => x"0c",
          3915 => x"33",
          3916 => x"06",
          3917 => x"70",
          3918 => x"76",
          3919 => x"0c",
          3920 => x"04",
          3921 => x"82",
          3922 => x"70",
          3923 => x"54",
          3924 => x"94",
          3925 => x"80",
          3926 => x"87",
          3927 => x"51",
          3928 => x"82",
          3929 => x"06",
          3930 => x"70",
          3931 => x"38",
          3932 => x"06",
          3933 => x"94",
          3934 => x"80",
          3935 => x"87",
          3936 => x"52",
          3937 => x"81",
          3938 => x"d4",
          3939 => x"84",
          3940 => x"ff",
          3941 => x"d4",
          3942 => x"ff",
          3943 => x"f8",
          3944 => x"3d",
          3945 => x"98",
          3946 => x"ff",
          3947 => x"87",
          3948 => x"52",
          3949 => x"86",
          3950 => x"94",
          3951 => x"08",
          3952 => x"70",
          3953 => x"51",
          3954 => x"70",
          3955 => x"38",
          3956 => x"06",
          3957 => x"94",
          3958 => x"80",
          3959 => x"87",
          3960 => x"52",
          3961 => x"98",
          3962 => x"2c",
          3963 => x"71",
          3964 => x"0c",
          3965 => x"04",
          3966 => x"87",
          3967 => x"08",
          3968 => x"8a",
          3969 => x"70",
          3970 => x"b4",
          3971 => x"9e",
          3972 => x"d3",
          3973 => x"c0",
          3974 => x"82",
          3975 => x"87",
          3976 => x"08",
          3977 => x"0c",
          3978 => x"98",
          3979 => x"a8",
          3980 => x"9e",
          3981 => x"d3",
          3982 => x"c0",
          3983 => x"82",
          3984 => x"87",
          3985 => x"08",
          3986 => x"0c",
          3987 => x"b0",
          3988 => x"b8",
          3989 => x"9e",
          3990 => x"d3",
          3991 => x"c0",
          3992 => x"82",
          3993 => x"87",
          3994 => x"08",
          3995 => x"0c",
          3996 => x"c0",
          3997 => x"c8",
          3998 => x"9e",
          3999 => x"d3",
          4000 => x"c0",
          4001 => x"51",
          4002 => x"d0",
          4003 => x"9e",
          4004 => x"d3",
          4005 => x"c0",
          4006 => x"82",
          4007 => x"87",
          4008 => x"08",
          4009 => x"0c",
          4010 => x"d3",
          4011 => x"0b",
          4012 => x"90",
          4013 => x"80",
          4014 => x"52",
          4015 => x"2e",
          4016 => x"52",
          4017 => x"e1",
          4018 => x"87",
          4019 => x"08",
          4020 => x"0a",
          4021 => x"52",
          4022 => x"83",
          4023 => x"71",
          4024 => x"34",
          4025 => x"c0",
          4026 => x"70",
          4027 => x"06",
          4028 => x"70",
          4029 => x"38",
          4030 => x"82",
          4031 => x"80",
          4032 => x"9e",
          4033 => x"88",
          4034 => x"51",
          4035 => x"80",
          4036 => x"81",
          4037 => x"d3",
          4038 => x"0b",
          4039 => x"90",
          4040 => x"80",
          4041 => x"52",
          4042 => x"2e",
          4043 => x"52",
          4044 => x"e5",
          4045 => x"87",
          4046 => x"08",
          4047 => x"80",
          4048 => x"52",
          4049 => x"83",
          4050 => x"71",
          4051 => x"34",
          4052 => x"c0",
          4053 => x"70",
          4054 => x"06",
          4055 => x"70",
          4056 => x"38",
          4057 => x"82",
          4058 => x"80",
          4059 => x"9e",
          4060 => x"82",
          4061 => x"51",
          4062 => x"80",
          4063 => x"81",
          4064 => x"d3",
          4065 => x"0b",
          4066 => x"90",
          4067 => x"80",
          4068 => x"52",
          4069 => x"2e",
          4070 => x"52",
          4071 => x"e9",
          4072 => x"87",
          4073 => x"08",
          4074 => x"80",
          4075 => x"52",
          4076 => x"83",
          4077 => x"71",
          4078 => x"34",
          4079 => x"c0",
          4080 => x"70",
          4081 => x"51",
          4082 => x"80",
          4083 => x"81",
          4084 => x"d3",
          4085 => x"c0",
          4086 => x"70",
          4087 => x"70",
          4088 => x"51",
          4089 => x"d3",
          4090 => x"0b",
          4091 => x"90",
          4092 => x"80",
          4093 => x"52",
          4094 => x"83",
          4095 => x"71",
          4096 => x"34",
          4097 => x"90",
          4098 => x"f0",
          4099 => x"2a",
          4100 => x"70",
          4101 => x"34",
          4102 => x"c0",
          4103 => x"70",
          4104 => x"52",
          4105 => x"2e",
          4106 => x"52",
          4107 => x"ef",
          4108 => x"9e",
          4109 => x"87",
          4110 => x"70",
          4111 => x"34",
          4112 => x"04",
          4113 => x"82",
          4114 => x"ff",
          4115 => x"82",
          4116 => x"54",
          4117 => x"89",
          4118 => x"88",
          4119 => x"fb",
          4120 => x"9c",
          4121 => x"fe",
          4122 => x"e2",
          4123 => x"80",
          4124 => x"82",
          4125 => x"82",
          4126 => x"11",
          4127 => x"bd",
          4128 => x"92",
          4129 => x"d3",
          4130 => x"73",
          4131 => x"38",
          4132 => x"08",
          4133 => x"08",
          4134 => x"82",
          4135 => x"ff",
          4136 => x"82",
          4137 => x"54",
          4138 => x"94",
          4139 => x"9c",
          4140 => x"a0",
          4141 => x"52",
          4142 => x"51",
          4143 => x"3f",
          4144 => x"33",
          4145 => x"2e",
          4146 => x"d3",
          4147 => x"d3",
          4148 => x"54",
          4149 => x"88",
          4150 => x"ff",
          4151 => x"e6",
          4152 => x"80",
          4153 => x"82",
          4154 => x"82",
          4155 => x"11",
          4156 => x"be",
          4157 => x"91",
          4158 => x"d3",
          4159 => x"73",
          4160 => x"38",
          4161 => x"33",
          4162 => x"c0",
          4163 => x"cb",
          4164 => x"ef",
          4165 => x"80",
          4166 => x"82",
          4167 => x"52",
          4168 => x"51",
          4169 => x"3f",
          4170 => x"33",
          4171 => x"2e",
          4172 => x"d3",
          4173 => x"82",
          4174 => x"ff",
          4175 => x"82",
          4176 => x"54",
          4177 => x"89",
          4178 => x"a0",
          4179 => x"96",
          4180 => x"e3",
          4181 => x"80",
          4182 => x"82",
          4183 => x"ff",
          4184 => x"82",
          4185 => x"54",
          4186 => x"89",
          4187 => x"c0",
          4188 => x"f2",
          4189 => x"e9",
          4190 => x"80",
          4191 => x"82",
          4192 => x"ff",
          4193 => x"82",
          4194 => x"54",
          4195 => x"89",
          4196 => x"d4",
          4197 => x"ce",
          4198 => x"dc",
          4199 => x"c6",
          4200 => x"c4",
          4201 => x"bf",
          4202 => x"90",
          4203 => x"d3",
          4204 => x"82",
          4205 => x"ff",
          4206 => x"82",
          4207 => x"52",
          4208 => x"51",
          4209 => x"3f",
          4210 => x"51",
          4211 => x"3f",
          4212 => x"22",
          4213 => x"e8",
          4214 => x"ff",
          4215 => x"d4",
          4216 => x"84",
          4217 => x"51",
          4218 => x"82",
          4219 => x"bd",
          4220 => x"76",
          4221 => x"54",
          4222 => x"08",
          4223 => x"90",
          4224 => x"d7",
          4225 => x"e7",
          4226 => x"80",
          4227 => x"82",
          4228 => x"56",
          4229 => x"52",
          4230 => x"95",
          4231 => x"f8",
          4232 => x"c0",
          4233 => x"31",
          4234 => x"d4",
          4235 => x"82",
          4236 => x"ff",
          4237 => x"82",
          4238 => x"54",
          4239 => x"a9",
          4240 => x"dc",
          4241 => x"84",
          4242 => x"51",
          4243 => x"82",
          4244 => x"bd",
          4245 => x"76",
          4246 => x"54",
          4247 => x"08",
          4248 => x"e8",
          4249 => x"f3",
          4250 => x"ff",
          4251 => x"87",
          4252 => x"fe",
          4253 => x"92",
          4254 => x"05",
          4255 => x"26",
          4256 => x"84",
          4257 => x"e8",
          4258 => x"08",
          4259 => x"94",
          4260 => x"82",
          4261 => x"97",
          4262 => x"a4",
          4263 => x"82",
          4264 => x"8b",
          4265 => x"b0",
          4266 => x"82",
          4267 => x"ff",
          4268 => x"84",
          4269 => x"71",
          4270 => x"04",
          4271 => x"c0",
          4272 => x"04",
          4273 => x"08",
          4274 => x"84",
          4275 => x"3d",
          4276 => x"2b",
          4277 => x"79",
          4278 => x"98",
          4279 => x"13",
          4280 => x"51",
          4281 => x"51",
          4282 => x"82",
          4283 => x"33",
          4284 => x"74",
          4285 => x"82",
          4286 => x"08",
          4287 => x"05",
          4288 => x"71",
          4289 => x"52",
          4290 => x"09",
          4291 => x"38",
          4292 => x"82",
          4293 => x"85",
          4294 => x"fb",
          4295 => x"02",
          4296 => x"05",
          4297 => x"55",
          4298 => x"80",
          4299 => x"82",
          4300 => x"52",
          4301 => x"ac",
          4302 => x"f0",
          4303 => x"a0",
          4304 => x"f1",
          4305 => x"dc",
          4306 => x"51",
          4307 => x"3f",
          4308 => x"05",
          4309 => x"34",
          4310 => x"06",
          4311 => x"77",
          4312 => x"f7",
          4313 => x"34",
          4314 => x"04",
          4315 => x"7c",
          4316 => x"b7",
          4317 => x"88",
          4318 => x"33",
          4319 => x"33",
          4320 => x"82",
          4321 => x"70",
          4322 => x"59",
          4323 => x"74",
          4324 => x"38",
          4325 => x"fb",
          4326 => x"d0",
          4327 => x"29",
          4328 => x"05",
          4329 => x"54",
          4330 => x"9d",
          4331 => x"d4",
          4332 => x"0c",
          4333 => x"33",
          4334 => x"82",
          4335 => x"70",
          4336 => x"5a",
          4337 => x"a7",
          4338 => x"78",
          4339 => x"ff",
          4340 => x"82",
          4341 => x"81",
          4342 => x"82",
          4343 => x"74",
          4344 => x"55",
          4345 => x"87",
          4346 => x"82",
          4347 => x"77",
          4348 => x"38",
          4349 => x"08",
          4350 => x"2e",
          4351 => x"d4",
          4352 => x"74",
          4353 => x"3d",
          4354 => x"76",
          4355 => x"75",
          4356 => x"bf",
          4357 => x"cc",
          4358 => x"51",
          4359 => x"3f",
          4360 => x"08",
          4361 => x"a2",
          4362 => x"0d",
          4363 => x"0d",
          4364 => x"53",
          4365 => x"08",
          4366 => x"2e",
          4367 => x"51",
          4368 => x"80",
          4369 => x"14",
          4370 => x"54",
          4371 => x"e6",
          4372 => x"82",
          4373 => x"82",
          4374 => x"52",
          4375 => x"95",
          4376 => x"80",
          4377 => x"82",
          4378 => x"51",
          4379 => x"80",
          4380 => x"cc",
          4381 => x"0d",
          4382 => x"0d",
          4383 => x"52",
          4384 => x"08",
          4385 => x"a3",
          4386 => x"f8",
          4387 => x"38",
          4388 => x"08",
          4389 => x"52",
          4390 => x"52",
          4391 => x"d3",
          4392 => x"f8",
          4393 => x"ba",
          4394 => x"ff",
          4395 => x"82",
          4396 => x"55",
          4397 => x"d4",
          4398 => x"9d",
          4399 => x"f8",
          4400 => x"70",
          4401 => x"80",
          4402 => x"53",
          4403 => x"17",
          4404 => x"52",
          4405 => x"83",
          4406 => x"2e",
          4407 => x"ff",
          4408 => x"3d",
          4409 => x"3d",
          4410 => x"08",
          4411 => x"5a",
          4412 => x"58",
          4413 => x"82",
          4414 => x"51",
          4415 => x"3f",
          4416 => x"08",
          4417 => x"ff",
          4418 => x"cc",
          4419 => x"80",
          4420 => x"3d",
          4421 => x"81",
          4422 => x"82",
          4423 => x"80",
          4424 => x"75",
          4425 => x"e0",
          4426 => x"f8",
          4427 => x"58",
          4428 => x"82",
          4429 => x"25",
          4430 => x"d4",
          4431 => x"05",
          4432 => x"55",
          4433 => x"74",
          4434 => x"70",
          4435 => x"2a",
          4436 => x"78",
          4437 => x"38",
          4438 => x"38",
          4439 => x"08",
          4440 => x"53",
          4441 => x"c3",
          4442 => x"f8",
          4443 => x"89",
          4444 => x"c0",
          4445 => x"e3",
          4446 => x"2e",
          4447 => x"9b",
          4448 => x"79",
          4449 => x"ee",
          4450 => x"ff",
          4451 => x"ab",
          4452 => x"82",
          4453 => x"74",
          4454 => x"77",
          4455 => x"0c",
          4456 => x"04",
          4457 => x"7c",
          4458 => x"71",
          4459 => x"59",
          4460 => x"a0",
          4461 => x"06",
          4462 => x"33",
          4463 => x"77",
          4464 => x"38",
          4465 => x"5b",
          4466 => x"56",
          4467 => x"a0",
          4468 => x"06",
          4469 => x"75",
          4470 => x"80",
          4471 => x"29",
          4472 => x"05",
          4473 => x"55",
          4474 => x"3f",
          4475 => x"08",
          4476 => x"74",
          4477 => x"b3",
          4478 => x"d4",
          4479 => x"c5",
          4480 => x"33",
          4481 => x"2e",
          4482 => x"82",
          4483 => x"b5",
          4484 => x"3f",
          4485 => x"1a",
          4486 => x"fc",
          4487 => x"05",
          4488 => x"3f",
          4489 => x"08",
          4490 => x"38",
          4491 => x"78",
          4492 => x"fd",
          4493 => x"d4",
          4494 => x"ff",
          4495 => x"85",
          4496 => x"91",
          4497 => x"70",
          4498 => x"51",
          4499 => x"27",
          4500 => x"80",
          4501 => x"d4",
          4502 => x"3d",
          4503 => x"3d",
          4504 => x"08",
          4505 => x"b4",
          4506 => x"5f",
          4507 => x"af",
          4508 => x"d4",
          4509 => x"d4",
          4510 => x"5b",
          4511 => x"38",
          4512 => x"c8",
          4513 => x"73",
          4514 => x"55",
          4515 => x"81",
          4516 => x"70",
          4517 => x"56",
          4518 => x"81",
          4519 => x"51",
          4520 => x"82",
          4521 => x"82",
          4522 => x"82",
          4523 => x"80",
          4524 => x"38",
          4525 => x"52",
          4526 => x"08",
          4527 => x"ae",
          4528 => x"f8",
          4529 => x"8c",
          4530 => x"ec",
          4531 => x"96",
          4532 => x"39",
          4533 => x"08",
          4534 => x"cc",
          4535 => x"f8",
          4536 => x"70",
          4537 => x"99",
          4538 => x"d4",
          4539 => x"82",
          4540 => x"74",
          4541 => x"06",
          4542 => x"82",
          4543 => x"51",
          4544 => x"3f",
          4545 => x"08",
          4546 => x"82",
          4547 => x"25",
          4548 => x"d4",
          4549 => x"05",
          4550 => x"55",
          4551 => x"80",
          4552 => x"ff",
          4553 => x"51",
          4554 => x"81",
          4555 => x"ff",
          4556 => x"93",
          4557 => x"38",
          4558 => x"ff",
          4559 => x"06",
          4560 => x"86",
          4561 => x"d4",
          4562 => x"8c",
          4563 => x"cc",
          4564 => x"84",
          4565 => x"3f",
          4566 => x"ec",
          4567 => x"d4",
          4568 => x"2b",
          4569 => x"51",
          4570 => x"2e",
          4571 => x"81",
          4572 => x"ec",
          4573 => x"98",
          4574 => x"2c",
          4575 => x"33",
          4576 => x"70",
          4577 => x"98",
          4578 => x"84",
          4579 => x"c0",
          4580 => x"15",
          4581 => x"51",
          4582 => x"59",
          4583 => x"58",
          4584 => x"78",
          4585 => x"38",
          4586 => x"b4",
          4587 => x"80",
          4588 => x"ff",
          4589 => x"98",
          4590 => x"80",
          4591 => x"ce",
          4592 => x"74",
          4593 => x"f6",
          4594 => x"d4",
          4595 => x"ff",
          4596 => x"80",
          4597 => x"74",
          4598 => x"34",
          4599 => x"39",
          4600 => x"0a",
          4601 => x"0a",
          4602 => x"2c",
          4603 => x"06",
          4604 => x"73",
          4605 => x"38",
          4606 => x"52",
          4607 => x"ce",
          4608 => x"f8",
          4609 => x"06",
          4610 => x"38",
          4611 => x"56",
          4612 => x"80",
          4613 => x"1c",
          4614 => x"ec",
          4615 => x"98",
          4616 => x"2c",
          4617 => x"33",
          4618 => x"70",
          4619 => x"10",
          4620 => x"2b",
          4621 => x"11",
          4622 => x"51",
          4623 => x"51",
          4624 => x"2e",
          4625 => x"fe",
          4626 => x"c2",
          4627 => x"7d",
          4628 => x"82",
          4629 => x"80",
          4630 => x"b0",
          4631 => x"75",
          4632 => x"34",
          4633 => x"b0",
          4634 => x"3d",
          4635 => x"0c",
          4636 => x"95",
          4637 => x"38",
          4638 => x"82",
          4639 => x"54",
          4640 => x"82",
          4641 => x"54",
          4642 => x"fd",
          4643 => x"ec",
          4644 => x"73",
          4645 => x"38",
          4646 => x"70",
          4647 => x"55",
          4648 => x"9e",
          4649 => x"54",
          4650 => x"15",
          4651 => x"80",
          4652 => x"ff",
          4653 => x"98",
          4654 => x"bc",
          4655 => x"55",
          4656 => x"ec",
          4657 => x"11",
          4658 => x"82",
          4659 => x"73",
          4660 => x"3d",
          4661 => x"82",
          4662 => x"54",
          4663 => x"89",
          4664 => x"54",
          4665 => x"b8",
          4666 => x"bc",
          4667 => x"80",
          4668 => x"ff",
          4669 => x"98",
          4670 => x"b8",
          4671 => x"56",
          4672 => x"25",
          4673 => x"f0",
          4674 => x"74",
          4675 => x"52",
          4676 => x"a1",
          4677 => x"80",
          4678 => x"80",
          4679 => x"98",
          4680 => x"b8",
          4681 => x"55",
          4682 => x"da",
          4683 => x"bc",
          4684 => x"2b",
          4685 => x"82",
          4686 => x"5a",
          4687 => x"74",
          4688 => x"94",
          4689 => x"dc",
          4690 => x"51",
          4691 => x"3f",
          4692 => x"0a",
          4693 => x"0a",
          4694 => x"2c",
          4695 => x"33",
          4696 => x"73",
          4697 => x"38",
          4698 => x"83",
          4699 => x"0b",
          4700 => x"82",
          4701 => x"80",
          4702 => x"dc",
          4703 => x"3f",
          4704 => x"82",
          4705 => x"70",
          4706 => x"55",
          4707 => x"2e",
          4708 => x"82",
          4709 => x"ff",
          4710 => x"82",
          4711 => x"ff",
          4712 => x"82",
          4713 => x"82",
          4714 => x"52",
          4715 => x"a0",
          4716 => x"ec",
          4717 => x"98",
          4718 => x"2c",
          4719 => x"33",
          4720 => x"57",
          4721 => x"ad",
          4722 => x"54",
          4723 => x"74",
          4724 => x"dc",
          4725 => x"33",
          4726 => x"d9",
          4727 => x"80",
          4728 => x"80",
          4729 => x"98",
          4730 => x"b8",
          4731 => x"55",
          4732 => x"d5",
          4733 => x"dc",
          4734 => x"51",
          4735 => x"3f",
          4736 => x"33",
          4737 => x"70",
          4738 => x"ec",
          4739 => x"51",
          4740 => x"74",
          4741 => x"38",
          4742 => x"08",
          4743 => x"ff",
          4744 => x"74",
          4745 => x"29",
          4746 => x"05",
          4747 => x"82",
          4748 => x"58",
          4749 => x"75",
          4750 => x"fa",
          4751 => x"ec",
          4752 => x"05",
          4753 => x"34",
          4754 => x"08",
          4755 => x"ff",
          4756 => x"82",
          4757 => x"79",
          4758 => x"3f",
          4759 => x"08",
          4760 => x"54",
          4761 => x"82",
          4762 => x"54",
          4763 => x"8f",
          4764 => x"73",
          4765 => x"f1",
          4766 => x"39",
          4767 => x"80",
          4768 => x"bc",
          4769 => x"82",
          4770 => x"79",
          4771 => x"0c",
          4772 => x"04",
          4773 => x"33",
          4774 => x"2e",
          4775 => x"82",
          4776 => x"52",
          4777 => x"9e",
          4778 => x"ec",
          4779 => x"05",
          4780 => x"ec",
          4781 => x"81",
          4782 => x"dd",
          4783 => x"bc",
          4784 => x"b8",
          4785 => x"73",
          4786 => x"8c",
          4787 => x"54",
          4788 => x"b8",
          4789 => x"2b",
          4790 => x"75",
          4791 => x"56",
          4792 => x"74",
          4793 => x"74",
          4794 => x"14",
          4795 => x"82",
          4796 => x"52",
          4797 => x"ff",
          4798 => x"74",
          4799 => x"29",
          4800 => x"05",
          4801 => x"82",
          4802 => x"58",
          4803 => x"75",
          4804 => x"82",
          4805 => x"52",
          4806 => x"9d",
          4807 => x"ec",
          4808 => x"98",
          4809 => x"2c",
          4810 => x"33",
          4811 => x"57",
          4812 => x"f8",
          4813 => x"f0",
          4814 => x"88",
          4815 => x"f5",
          4816 => x"80",
          4817 => x"80",
          4818 => x"98",
          4819 => x"b8",
          4820 => x"55",
          4821 => x"de",
          4822 => x"39",
          4823 => x"33",
          4824 => x"06",
          4825 => x"33",
          4826 => x"74",
          4827 => x"e8",
          4828 => x"dc",
          4829 => x"14",
          4830 => x"ec",
          4831 => x"1a",
          4832 => x"54",
          4833 => x"3f",
          4834 => x"33",
          4835 => x"06",
          4836 => x"33",
          4837 => x"75",
          4838 => x"38",
          4839 => x"82",
          4840 => x"80",
          4841 => x"dc",
          4842 => x"3f",
          4843 => x"ec",
          4844 => x"0b",
          4845 => x"34",
          4846 => x"7a",
          4847 => x"d4",
          4848 => x"74",
          4849 => x"38",
          4850 => x"a4",
          4851 => x"d4",
          4852 => x"ec",
          4853 => x"d4",
          4854 => x"ff",
          4855 => x"53",
          4856 => x"51",
          4857 => x"3f",
          4858 => x"c0",
          4859 => x"29",
          4860 => x"05",
          4861 => x"56",
          4862 => x"2e",
          4863 => x"51",
          4864 => x"3f",
          4865 => x"08",
          4866 => x"34",
          4867 => x"08",
          4868 => x"81",
          4869 => x"52",
          4870 => x"a5",
          4871 => x"1b",
          4872 => x"39",
          4873 => x"74",
          4874 => x"ac",
          4875 => x"ff",
          4876 => x"99",
          4877 => x"2e",
          4878 => x"ae",
          4879 => x"f8",
          4880 => x"80",
          4881 => x"74",
          4882 => x"bc",
          4883 => x"f8",
          4884 => x"b8",
          4885 => x"f8",
          4886 => x"06",
          4887 => x"74",
          4888 => x"ff",
          4889 => x"80",
          4890 => x"84",
          4891 => x"fc",
          4892 => x"56",
          4893 => x"2e",
          4894 => x"51",
          4895 => x"3f",
          4896 => x"08",
          4897 => x"34",
          4898 => x"08",
          4899 => x"81",
          4900 => x"52",
          4901 => x"a4",
          4902 => x"1b",
          4903 => x"ff",
          4904 => x"39",
          4905 => x"b8",
          4906 => x"34",
          4907 => x"53",
          4908 => x"33",
          4909 => x"ec",
          4910 => x"9c",
          4911 => x"bc",
          4912 => x"ff",
          4913 => x"b8",
          4914 => x"54",
          4915 => x"f5",
          4916 => x"f0",
          4917 => x"81",
          4918 => x"82",
          4919 => x"74",
          4920 => x"52",
          4921 => x"cd",
          4922 => x"39",
          4923 => x"33",
          4924 => x"2e",
          4925 => x"82",
          4926 => x"52",
          4927 => x"99",
          4928 => x"ec",
          4929 => x"05",
          4930 => x"ec",
          4931 => x"c8",
          4932 => x"0d",
          4933 => x"0b",
          4934 => x"0c",
          4935 => x"82",
          4936 => x"80",
          4937 => x"80",
          4938 => x"f4",
          4939 => x"e4",
          4940 => x"f0",
          4941 => x"58",
          4942 => x"81",
          4943 => x"15",
          4944 => x"f0",
          4945 => x"84",
          4946 => x"85",
          4947 => x"d4",
          4948 => x"77",
          4949 => x"76",
          4950 => x"82",
          4951 => x"82",
          4952 => x"ff",
          4953 => x"80",
          4954 => x"ff",
          4955 => x"88",
          4956 => x"55",
          4957 => x"17",
          4958 => x"17",
          4959 => x"ec",
          4960 => x"29",
          4961 => x"08",
          4962 => x"51",
          4963 => x"82",
          4964 => x"83",
          4965 => x"3d",
          4966 => x"3d",
          4967 => x"81",
          4968 => x"27",
          4969 => x"12",
          4970 => x"11",
          4971 => x"ff",
          4972 => x"51",
          4973 => x"f8",
          4974 => x"0d",
          4975 => x"0d",
          4976 => x"22",
          4977 => x"aa",
          4978 => x"05",
          4979 => x"08",
          4980 => x"71",
          4981 => x"2b",
          4982 => x"33",
          4983 => x"71",
          4984 => x"02",
          4985 => x"05",
          4986 => x"ff",
          4987 => x"70",
          4988 => x"51",
          4989 => x"5b",
          4990 => x"54",
          4991 => x"34",
          4992 => x"34",
          4993 => x"08",
          4994 => x"2a",
          4995 => x"82",
          4996 => x"83",
          4997 => x"d4",
          4998 => x"17",
          4999 => x"12",
          5000 => x"2b",
          5001 => x"2b",
          5002 => x"06",
          5003 => x"52",
          5004 => x"83",
          5005 => x"70",
          5006 => x"54",
          5007 => x"12",
          5008 => x"ff",
          5009 => x"83",
          5010 => x"d4",
          5011 => x"56",
          5012 => x"72",
          5013 => x"89",
          5014 => x"fb",
          5015 => x"d4",
          5016 => x"84",
          5017 => x"22",
          5018 => x"72",
          5019 => x"33",
          5020 => x"71",
          5021 => x"83",
          5022 => x"5b",
          5023 => x"52",
          5024 => x"12",
          5025 => x"33",
          5026 => x"07",
          5027 => x"54",
          5028 => x"70",
          5029 => x"73",
          5030 => x"82",
          5031 => x"70",
          5032 => x"33",
          5033 => x"71",
          5034 => x"83",
          5035 => x"59",
          5036 => x"05",
          5037 => x"87",
          5038 => x"88",
          5039 => x"88",
          5040 => x"56",
          5041 => x"13",
          5042 => x"13",
          5043 => x"f0",
          5044 => x"33",
          5045 => x"71",
          5046 => x"70",
          5047 => x"06",
          5048 => x"53",
          5049 => x"53",
          5050 => x"70",
          5051 => x"87",
          5052 => x"fa",
          5053 => x"a2",
          5054 => x"d4",
          5055 => x"83",
          5056 => x"70",
          5057 => x"33",
          5058 => x"07",
          5059 => x"15",
          5060 => x"12",
          5061 => x"2b",
          5062 => x"07",
          5063 => x"55",
          5064 => x"57",
          5065 => x"80",
          5066 => x"38",
          5067 => x"ab",
          5068 => x"f0",
          5069 => x"70",
          5070 => x"33",
          5071 => x"71",
          5072 => x"74",
          5073 => x"81",
          5074 => x"88",
          5075 => x"83",
          5076 => x"f8",
          5077 => x"54",
          5078 => x"58",
          5079 => x"74",
          5080 => x"52",
          5081 => x"34",
          5082 => x"34",
          5083 => x"08",
          5084 => x"33",
          5085 => x"71",
          5086 => x"83",
          5087 => x"59",
          5088 => x"05",
          5089 => x"12",
          5090 => x"2b",
          5091 => x"ff",
          5092 => x"88",
          5093 => x"52",
          5094 => x"74",
          5095 => x"15",
          5096 => x"0d",
          5097 => x"0d",
          5098 => x"08",
          5099 => x"9e",
          5100 => x"83",
          5101 => x"82",
          5102 => x"12",
          5103 => x"2b",
          5104 => x"07",
          5105 => x"52",
          5106 => x"05",
          5107 => x"13",
          5108 => x"2b",
          5109 => x"05",
          5110 => x"71",
          5111 => x"2a",
          5112 => x"53",
          5113 => x"34",
          5114 => x"34",
          5115 => x"08",
          5116 => x"33",
          5117 => x"71",
          5118 => x"83",
          5119 => x"59",
          5120 => x"05",
          5121 => x"83",
          5122 => x"88",
          5123 => x"88",
          5124 => x"56",
          5125 => x"13",
          5126 => x"13",
          5127 => x"f0",
          5128 => x"11",
          5129 => x"33",
          5130 => x"07",
          5131 => x"0c",
          5132 => x"3d",
          5133 => x"3d",
          5134 => x"d4",
          5135 => x"83",
          5136 => x"ff",
          5137 => x"53",
          5138 => x"a7",
          5139 => x"f0",
          5140 => x"2b",
          5141 => x"11",
          5142 => x"33",
          5143 => x"71",
          5144 => x"75",
          5145 => x"81",
          5146 => x"98",
          5147 => x"2b",
          5148 => x"40",
          5149 => x"58",
          5150 => x"72",
          5151 => x"38",
          5152 => x"52",
          5153 => x"9d",
          5154 => x"39",
          5155 => x"85",
          5156 => x"8b",
          5157 => x"2b",
          5158 => x"79",
          5159 => x"51",
          5160 => x"76",
          5161 => x"75",
          5162 => x"56",
          5163 => x"34",
          5164 => x"08",
          5165 => x"12",
          5166 => x"33",
          5167 => x"07",
          5168 => x"54",
          5169 => x"53",
          5170 => x"34",
          5171 => x"34",
          5172 => x"08",
          5173 => x"0b",
          5174 => x"80",
          5175 => x"34",
          5176 => x"08",
          5177 => x"14",
          5178 => x"14",
          5179 => x"f0",
          5180 => x"33",
          5181 => x"71",
          5182 => x"70",
          5183 => x"07",
          5184 => x"53",
          5185 => x"54",
          5186 => x"72",
          5187 => x"8b",
          5188 => x"ff",
          5189 => x"52",
          5190 => x"08",
          5191 => x"f1",
          5192 => x"2e",
          5193 => x"51",
          5194 => x"83",
          5195 => x"f5",
          5196 => x"7e",
          5197 => x"e2",
          5198 => x"f8",
          5199 => x"ff",
          5200 => x"f0",
          5201 => x"33",
          5202 => x"71",
          5203 => x"70",
          5204 => x"58",
          5205 => x"ff",
          5206 => x"2e",
          5207 => x"75",
          5208 => x"70",
          5209 => x"33",
          5210 => x"07",
          5211 => x"ff",
          5212 => x"70",
          5213 => x"06",
          5214 => x"52",
          5215 => x"59",
          5216 => x"27",
          5217 => x"80",
          5218 => x"75",
          5219 => x"84",
          5220 => x"16",
          5221 => x"2b",
          5222 => x"75",
          5223 => x"81",
          5224 => x"85",
          5225 => x"59",
          5226 => x"83",
          5227 => x"f0",
          5228 => x"33",
          5229 => x"71",
          5230 => x"70",
          5231 => x"06",
          5232 => x"56",
          5233 => x"75",
          5234 => x"81",
          5235 => x"79",
          5236 => x"cc",
          5237 => x"74",
          5238 => x"c4",
          5239 => x"2e",
          5240 => x"89",
          5241 => x"f8",
          5242 => x"ac",
          5243 => x"80",
          5244 => x"75",
          5245 => x"3f",
          5246 => x"08",
          5247 => x"11",
          5248 => x"33",
          5249 => x"71",
          5250 => x"53",
          5251 => x"74",
          5252 => x"70",
          5253 => x"06",
          5254 => x"5c",
          5255 => x"78",
          5256 => x"76",
          5257 => x"57",
          5258 => x"34",
          5259 => x"08",
          5260 => x"71",
          5261 => x"86",
          5262 => x"12",
          5263 => x"2b",
          5264 => x"2a",
          5265 => x"53",
          5266 => x"73",
          5267 => x"75",
          5268 => x"82",
          5269 => x"70",
          5270 => x"33",
          5271 => x"71",
          5272 => x"83",
          5273 => x"5d",
          5274 => x"05",
          5275 => x"15",
          5276 => x"15",
          5277 => x"f0",
          5278 => x"71",
          5279 => x"33",
          5280 => x"71",
          5281 => x"70",
          5282 => x"5a",
          5283 => x"54",
          5284 => x"34",
          5285 => x"34",
          5286 => x"08",
          5287 => x"54",
          5288 => x"f8",
          5289 => x"0d",
          5290 => x"0d",
          5291 => x"d4",
          5292 => x"38",
          5293 => x"71",
          5294 => x"2e",
          5295 => x"51",
          5296 => x"82",
          5297 => x"53",
          5298 => x"f8",
          5299 => x"0d",
          5300 => x"0d",
          5301 => x"5c",
          5302 => x"40",
          5303 => x"08",
          5304 => x"81",
          5305 => x"f4",
          5306 => x"8e",
          5307 => x"ff",
          5308 => x"d4",
          5309 => x"83",
          5310 => x"8b",
          5311 => x"fc",
          5312 => x"54",
          5313 => x"7e",
          5314 => x"3f",
          5315 => x"08",
          5316 => x"06",
          5317 => x"08",
          5318 => x"83",
          5319 => x"ff",
          5320 => x"83",
          5321 => x"70",
          5322 => x"33",
          5323 => x"07",
          5324 => x"70",
          5325 => x"06",
          5326 => x"fc",
          5327 => x"29",
          5328 => x"81",
          5329 => x"88",
          5330 => x"90",
          5331 => x"4e",
          5332 => x"52",
          5333 => x"41",
          5334 => x"5b",
          5335 => x"8f",
          5336 => x"ff",
          5337 => x"31",
          5338 => x"ff",
          5339 => x"82",
          5340 => x"17",
          5341 => x"2b",
          5342 => x"29",
          5343 => x"81",
          5344 => x"98",
          5345 => x"2b",
          5346 => x"45",
          5347 => x"73",
          5348 => x"38",
          5349 => x"70",
          5350 => x"06",
          5351 => x"7b",
          5352 => x"38",
          5353 => x"73",
          5354 => x"81",
          5355 => x"78",
          5356 => x"3f",
          5357 => x"ff",
          5358 => x"e5",
          5359 => x"38",
          5360 => x"89",
          5361 => x"f6",
          5362 => x"a5",
          5363 => x"55",
          5364 => x"80",
          5365 => x"1d",
          5366 => x"83",
          5367 => x"88",
          5368 => x"57",
          5369 => x"3f",
          5370 => x"51",
          5371 => x"82",
          5372 => x"83",
          5373 => x"7e",
          5374 => x"70",
          5375 => x"d4",
          5376 => x"84",
          5377 => x"59",
          5378 => x"3f",
          5379 => x"08",
          5380 => x"75",
          5381 => x"06",
          5382 => x"85",
          5383 => x"54",
          5384 => x"80",
          5385 => x"51",
          5386 => x"82",
          5387 => x"1d",
          5388 => x"83",
          5389 => x"88",
          5390 => x"43",
          5391 => x"3f",
          5392 => x"51",
          5393 => x"82",
          5394 => x"83",
          5395 => x"7e",
          5396 => x"70",
          5397 => x"d4",
          5398 => x"84",
          5399 => x"59",
          5400 => x"3f",
          5401 => x"08",
          5402 => x"60",
          5403 => x"55",
          5404 => x"ff",
          5405 => x"a9",
          5406 => x"52",
          5407 => x"3f",
          5408 => x"08",
          5409 => x"f8",
          5410 => x"93",
          5411 => x"73",
          5412 => x"f8",
          5413 => x"94",
          5414 => x"51",
          5415 => x"7a",
          5416 => x"27",
          5417 => x"53",
          5418 => x"51",
          5419 => x"7a",
          5420 => x"82",
          5421 => x"05",
          5422 => x"f6",
          5423 => x"54",
          5424 => x"f8",
          5425 => x"0d",
          5426 => x"0d",
          5427 => x"70",
          5428 => x"d5",
          5429 => x"f8",
          5430 => x"d4",
          5431 => x"2e",
          5432 => x"53",
          5433 => x"d4",
          5434 => x"ff",
          5435 => x"74",
          5436 => x"0c",
          5437 => x"04",
          5438 => x"02",
          5439 => x"51",
          5440 => x"72",
          5441 => x"82",
          5442 => x"33",
          5443 => x"d4",
          5444 => x"3d",
          5445 => x"3d",
          5446 => x"05",
          5447 => x"05",
          5448 => x"56",
          5449 => x"72",
          5450 => x"e0",
          5451 => x"2b",
          5452 => x"8c",
          5453 => x"88",
          5454 => x"2e",
          5455 => x"88",
          5456 => x"0c",
          5457 => x"8c",
          5458 => x"71",
          5459 => x"87",
          5460 => x"0c",
          5461 => x"08",
          5462 => x"51",
          5463 => x"2e",
          5464 => x"c0",
          5465 => x"51",
          5466 => x"71",
          5467 => x"80",
          5468 => x"92",
          5469 => x"98",
          5470 => x"70",
          5471 => x"38",
          5472 => x"f4",
          5473 => x"d4",
          5474 => x"51",
          5475 => x"f8",
          5476 => x"0d",
          5477 => x"0d",
          5478 => x"02",
          5479 => x"05",
          5480 => x"58",
          5481 => x"52",
          5482 => x"3f",
          5483 => x"08",
          5484 => x"54",
          5485 => x"be",
          5486 => x"75",
          5487 => x"c0",
          5488 => x"87",
          5489 => x"12",
          5490 => x"84",
          5491 => x"40",
          5492 => x"85",
          5493 => x"98",
          5494 => x"7d",
          5495 => x"0c",
          5496 => x"85",
          5497 => x"06",
          5498 => x"71",
          5499 => x"38",
          5500 => x"71",
          5501 => x"05",
          5502 => x"19",
          5503 => x"a2",
          5504 => x"71",
          5505 => x"38",
          5506 => x"83",
          5507 => x"38",
          5508 => x"8a",
          5509 => x"98",
          5510 => x"71",
          5511 => x"c0",
          5512 => x"52",
          5513 => x"87",
          5514 => x"80",
          5515 => x"81",
          5516 => x"c0",
          5517 => x"53",
          5518 => x"82",
          5519 => x"71",
          5520 => x"1a",
          5521 => x"84",
          5522 => x"19",
          5523 => x"06",
          5524 => x"79",
          5525 => x"38",
          5526 => x"80",
          5527 => x"87",
          5528 => x"26",
          5529 => x"73",
          5530 => x"06",
          5531 => x"2e",
          5532 => x"52",
          5533 => x"82",
          5534 => x"8f",
          5535 => x"f3",
          5536 => x"62",
          5537 => x"05",
          5538 => x"57",
          5539 => x"83",
          5540 => x"52",
          5541 => x"3f",
          5542 => x"08",
          5543 => x"54",
          5544 => x"2e",
          5545 => x"81",
          5546 => x"74",
          5547 => x"c0",
          5548 => x"87",
          5549 => x"12",
          5550 => x"84",
          5551 => x"5f",
          5552 => x"0b",
          5553 => x"8c",
          5554 => x"0c",
          5555 => x"80",
          5556 => x"70",
          5557 => x"81",
          5558 => x"54",
          5559 => x"8c",
          5560 => x"81",
          5561 => x"7c",
          5562 => x"58",
          5563 => x"70",
          5564 => x"52",
          5565 => x"8a",
          5566 => x"98",
          5567 => x"71",
          5568 => x"c0",
          5569 => x"52",
          5570 => x"87",
          5571 => x"80",
          5572 => x"81",
          5573 => x"c0",
          5574 => x"53",
          5575 => x"82",
          5576 => x"71",
          5577 => x"19",
          5578 => x"81",
          5579 => x"ff",
          5580 => x"19",
          5581 => x"78",
          5582 => x"38",
          5583 => x"80",
          5584 => x"87",
          5585 => x"26",
          5586 => x"73",
          5587 => x"06",
          5588 => x"2e",
          5589 => x"52",
          5590 => x"82",
          5591 => x"8f",
          5592 => x"fa",
          5593 => x"02",
          5594 => x"05",
          5595 => x"05",
          5596 => x"71",
          5597 => x"57",
          5598 => x"82",
          5599 => x"81",
          5600 => x"54",
          5601 => x"38",
          5602 => x"c0",
          5603 => x"81",
          5604 => x"2e",
          5605 => x"71",
          5606 => x"38",
          5607 => x"87",
          5608 => x"11",
          5609 => x"80",
          5610 => x"80",
          5611 => x"83",
          5612 => x"38",
          5613 => x"72",
          5614 => x"2a",
          5615 => x"51",
          5616 => x"80",
          5617 => x"87",
          5618 => x"08",
          5619 => x"38",
          5620 => x"8c",
          5621 => x"96",
          5622 => x"0c",
          5623 => x"8c",
          5624 => x"08",
          5625 => x"51",
          5626 => x"38",
          5627 => x"56",
          5628 => x"80",
          5629 => x"85",
          5630 => x"77",
          5631 => x"83",
          5632 => x"75",
          5633 => x"d4",
          5634 => x"3d",
          5635 => x"3d",
          5636 => x"11",
          5637 => x"71",
          5638 => x"82",
          5639 => x"53",
          5640 => x"0d",
          5641 => x"0d",
          5642 => x"33",
          5643 => x"71",
          5644 => x"88",
          5645 => x"14",
          5646 => x"07",
          5647 => x"33",
          5648 => x"d4",
          5649 => x"53",
          5650 => x"52",
          5651 => x"04",
          5652 => x"73",
          5653 => x"92",
          5654 => x"52",
          5655 => x"81",
          5656 => x"70",
          5657 => x"70",
          5658 => x"3d",
          5659 => x"3d",
          5660 => x"52",
          5661 => x"70",
          5662 => x"34",
          5663 => x"51",
          5664 => x"81",
          5665 => x"70",
          5666 => x"70",
          5667 => x"05",
          5668 => x"88",
          5669 => x"72",
          5670 => x"0d",
          5671 => x"0d",
          5672 => x"54",
          5673 => x"80",
          5674 => x"71",
          5675 => x"53",
          5676 => x"81",
          5677 => x"ff",
          5678 => x"39",
          5679 => x"04",
          5680 => x"75",
          5681 => x"52",
          5682 => x"70",
          5683 => x"34",
          5684 => x"70",
          5685 => x"3d",
          5686 => x"3d",
          5687 => x"79",
          5688 => x"74",
          5689 => x"56",
          5690 => x"81",
          5691 => x"71",
          5692 => x"16",
          5693 => x"52",
          5694 => x"86",
          5695 => x"2e",
          5696 => x"82",
          5697 => x"86",
          5698 => x"fe",
          5699 => x"76",
          5700 => x"39",
          5701 => x"8a",
          5702 => x"51",
          5703 => x"71",
          5704 => x"33",
          5705 => x"0c",
          5706 => x"04",
          5707 => x"d4",
          5708 => x"fb",
          5709 => x"70",
          5710 => x"81",
          5711 => x"70",
          5712 => x"56",
          5713 => x"55",
          5714 => x"08",
          5715 => x"80",
          5716 => x"83",
          5717 => x"51",
          5718 => x"3f",
          5719 => x"08",
          5720 => x"06",
          5721 => x"2e",
          5722 => x"76",
          5723 => x"74",
          5724 => x"0c",
          5725 => x"04",
          5726 => x"7b",
          5727 => x"83",
          5728 => x"5a",
          5729 => x"80",
          5730 => x"54",
          5731 => x"53",
          5732 => x"53",
          5733 => x"52",
          5734 => x"3f",
          5735 => x"08",
          5736 => x"81",
          5737 => x"82",
          5738 => x"83",
          5739 => x"16",
          5740 => x"18",
          5741 => x"18",
          5742 => x"58",
          5743 => x"9f",
          5744 => x"33",
          5745 => x"2e",
          5746 => x"93",
          5747 => x"76",
          5748 => x"52",
          5749 => x"51",
          5750 => x"83",
          5751 => x"79",
          5752 => x"0c",
          5753 => x"04",
          5754 => x"78",
          5755 => x"80",
          5756 => x"17",
          5757 => x"38",
          5758 => x"fc",
          5759 => x"f8",
          5760 => x"d4",
          5761 => x"38",
          5762 => x"53",
          5763 => x"81",
          5764 => x"f7",
          5765 => x"d4",
          5766 => x"2e",
          5767 => x"55",
          5768 => x"b4",
          5769 => x"82",
          5770 => x"88",
          5771 => x"f8",
          5772 => x"70",
          5773 => x"c0",
          5774 => x"f8",
          5775 => x"d4",
          5776 => x"91",
          5777 => x"55",
          5778 => x"09",
          5779 => x"f0",
          5780 => x"33",
          5781 => x"2e",
          5782 => x"80",
          5783 => x"80",
          5784 => x"f8",
          5785 => x"17",
          5786 => x"fc",
          5787 => x"d4",
          5788 => x"b6",
          5789 => x"d8",
          5790 => x"85",
          5791 => x"75",
          5792 => x"3f",
          5793 => x"e4",
          5794 => x"9c",
          5795 => x"de",
          5796 => x"08",
          5797 => x"17",
          5798 => x"3f",
          5799 => x"52",
          5800 => x"51",
          5801 => x"a4",
          5802 => x"05",
          5803 => x"0c",
          5804 => x"75",
          5805 => x"33",
          5806 => x"3f",
          5807 => x"34",
          5808 => x"52",
          5809 => x"51",
          5810 => x"82",
          5811 => x"80",
          5812 => x"81",
          5813 => x"d4",
          5814 => x"3d",
          5815 => x"3d",
          5816 => x"1a",
          5817 => x"fe",
          5818 => x"54",
          5819 => x"73",
          5820 => x"8a",
          5821 => x"71",
          5822 => x"08",
          5823 => x"75",
          5824 => x"0c",
          5825 => x"04",
          5826 => x"7a",
          5827 => x"56",
          5828 => x"77",
          5829 => x"38",
          5830 => x"08",
          5831 => x"38",
          5832 => x"54",
          5833 => x"2e",
          5834 => x"72",
          5835 => x"38",
          5836 => x"8d",
          5837 => x"39",
          5838 => x"81",
          5839 => x"b6",
          5840 => x"2a",
          5841 => x"2a",
          5842 => x"05",
          5843 => x"55",
          5844 => x"82",
          5845 => x"81",
          5846 => x"83",
          5847 => x"b8",
          5848 => x"17",
          5849 => x"a8",
          5850 => x"55",
          5851 => x"57",
          5852 => x"3f",
          5853 => x"08",
          5854 => x"74",
          5855 => x"14",
          5856 => x"70",
          5857 => x"07",
          5858 => x"71",
          5859 => x"52",
          5860 => x"72",
          5861 => x"75",
          5862 => x"58",
          5863 => x"76",
          5864 => x"15",
          5865 => x"73",
          5866 => x"3f",
          5867 => x"08",
          5868 => x"76",
          5869 => x"06",
          5870 => x"05",
          5871 => x"3f",
          5872 => x"08",
          5873 => x"06",
          5874 => x"76",
          5875 => x"15",
          5876 => x"73",
          5877 => x"3f",
          5878 => x"08",
          5879 => x"82",
          5880 => x"06",
          5881 => x"05",
          5882 => x"3f",
          5883 => x"08",
          5884 => x"58",
          5885 => x"58",
          5886 => x"f8",
          5887 => x"0d",
          5888 => x"0d",
          5889 => x"5a",
          5890 => x"59",
          5891 => x"82",
          5892 => x"9c",
          5893 => x"82",
          5894 => x"33",
          5895 => x"2e",
          5896 => x"72",
          5897 => x"38",
          5898 => x"8d",
          5899 => x"39",
          5900 => x"81",
          5901 => x"f7",
          5902 => x"2a",
          5903 => x"2a",
          5904 => x"05",
          5905 => x"55",
          5906 => x"82",
          5907 => x"59",
          5908 => x"08",
          5909 => x"74",
          5910 => x"16",
          5911 => x"16",
          5912 => x"59",
          5913 => x"53",
          5914 => x"8f",
          5915 => x"2b",
          5916 => x"74",
          5917 => x"71",
          5918 => x"72",
          5919 => x"0b",
          5920 => x"74",
          5921 => x"17",
          5922 => x"75",
          5923 => x"3f",
          5924 => x"08",
          5925 => x"f8",
          5926 => x"38",
          5927 => x"06",
          5928 => x"78",
          5929 => x"54",
          5930 => x"77",
          5931 => x"33",
          5932 => x"71",
          5933 => x"51",
          5934 => x"34",
          5935 => x"76",
          5936 => x"17",
          5937 => x"75",
          5938 => x"3f",
          5939 => x"08",
          5940 => x"f8",
          5941 => x"38",
          5942 => x"ff",
          5943 => x"10",
          5944 => x"76",
          5945 => x"51",
          5946 => x"be",
          5947 => x"2a",
          5948 => x"05",
          5949 => x"f9",
          5950 => x"d4",
          5951 => x"82",
          5952 => x"ab",
          5953 => x"0a",
          5954 => x"2b",
          5955 => x"70",
          5956 => x"70",
          5957 => x"54",
          5958 => x"82",
          5959 => x"8f",
          5960 => x"07",
          5961 => x"f6",
          5962 => x"0b",
          5963 => x"78",
          5964 => x"0c",
          5965 => x"04",
          5966 => x"7a",
          5967 => x"08",
          5968 => x"59",
          5969 => x"a4",
          5970 => x"17",
          5971 => x"38",
          5972 => x"aa",
          5973 => x"73",
          5974 => x"fd",
          5975 => x"d4",
          5976 => x"82",
          5977 => x"80",
          5978 => x"39",
          5979 => x"eb",
          5980 => x"80",
          5981 => x"d4",
          5982 => x"80",
          5983 => x"52",
          5984 => x"84",
          5985 => x"f8",
          5986 => x"d4",
          5987 => x"2e",
          5988 => x"82",
          5989 => x"81",
          5990 => x"82",
          5991 => x"ff",
          5992 => x"80",
          5993 => x"75",
          5994 => x"3f",
          5995 => x"08",
          5996 => x"16",
          5997 => x"94",
          5998 => x"55",
          5999 => x"27",
          6000 => x"15",
          6001 => x"84",
          6002 => x"07",
          6003 => x"17",
          6004 => x"76",
          6005 => x"a6",
          6006 => x"73",
          6007 => x"0c",
          6008 => x"04",
          6009 => x"7c",
          6010 => x"59",
          6011 => x"95",
          6012 => x"08",
          6013 => x"2e",
          6014 => x"17",
          6015 => x"b2",
          6016 => x"ae",
          6017 => x"7a",
          6018 => x"3f",
          6019 => x"82",
          6020 => x"27",
          6021 => x"82",
          6022 => x"55",
          6023 => x"08",
          6024 => x"d2",
          6025 => x"08",
          6026 => x"08",
          6027 => x"38",
          6028 => x"17",
          6029 => x"54",
          6030 => x"82",
          6031 => x"7a",
          6032 => x"06",
          6033 => x"81",
          6034 => x"17",
          6035 => x"83",
          6036 => x"75",
          6037 => x"f9",
          6038 => x"59",
          6039 => x"08",
          6040 => x"81",
          6041 => x"82",
          6042 => x"59",
          6043 => x"08",
          6044 => x"70",
          6045 => x"25",
          6046 => x"82",
          6047 => x"54",
          6048 => x"55",
          6049 => x"38",
          6050 => x"08",
          6051 => x"38",
          6052 => x"54",
          6053 => x"90",
          6054 => x"18",
          6055 => x"38",
          6056 => x"39",
          6057 => x"38",
          6058 => x"16",
          6059 => x"08",
          6060 => x"38",
          6061 => x"78",
          6062 => x"38",
          6063 => x"51",
          6064 => x"82",
          6065 => x"80",
          6066 => x"80",
          6067 => x"f8",
          6068 => x"09",
          6069 => x"38",
          6070 => x"08",
          6071 => x"f8",
          6072 => x"30",
          6073 => x"80",
          6074 => x"07",
          6075 => x"55",
          6076 => x"38",
          6077 => x"09",
          6078 => x"ae",
          6079 => x"80",
          6080 => x"53",
          6081 => x"51",
          6082 => x"82",
          6083 => x"82",
          6084 => x"30",
          6085 => x"f8",
          6086 => x"25",
          6087 => x"79",
          6088 => x"38",
          6089 => x"8f",
          6090 => x"79",
          6091 => x"f9",
          6092 => x"d4",
          6093 => x"74",
          6094 => x"90",
          6095 => x"17",
          6096 => x"94",
          6097 => x"54",
          6098 => x"86",
          6099 => x"94",
          6100 => x"17",
          6101 => x"54",
          6102 => x"34",
          6103 => x"56",
          6104 => x"90",
          6105 => x"80",
          6106 => x"82",
          6107 => x"55",
          6108 => x"56",
          6109 => x"82",
          6110 => x"8c",
          6111 => x"f8",
          6112 => x"70",
          6113 => x"f0",
          6114 => x"f8",
          6115 => x"56",
          6116 => x"08",
          6117 => x"7b",
          6118 => x"f6",
          6119 => x"d4",
          6120 => x"d4",
          6121 => x"17",
          6122 => x"80",
          6123 => x"b8",
          6124 => x"57",
          6125 => x"77",
          6126 => x"81",
          6127 => x"15",
          6128 => x"78",
          6129 => x"81",
          6130 => x"53",
          6131 => x"15",
          6132 => x"ab",
          6133 => x"f8",
          6134 => x"df",
          6135 => x"22",
          6136 => x"30",
          6137 => x"70",
          6138 => x"51",
          6139 => x"82",
          6140 => x"8a",
          6141 => x"f8",
          6142 => x"7c",
          6143 => x"56",
          6144 => x"80",
          6145 => x"f1",
          6146 => x"06",
          6147 => x"e9",
          6148 => x"18",
          6149 => x"08",
          6150 => x"38",
          6151 => x"82",
          6152 => x"38",
          6153 => x"54",
          6154 => x"74",
          6155 => x"82",
          6156 => x"22",
          6157 => x"79",
          6158 => x"38",
          6159 => x"98",
          6160 => x"cd",
          6161 => x"22",
          6162 => x"54",
          6163 => x"26",
          6164 => x"52",
          6165 => x"b0",
          6166 => x"f8",
          6167 => x"d4",
          6168 => x"2e",
          6169 => x"0b",
          6170 => x"08",
          6171 => x"9c",
          6172 => x"d4",
          6173 => x"85",
          6174 => x"bd",
          6175 => x"31",
          6176 => x"73",
          6177 => x"f4",
          6178 => x"d4",
          6179 => x"18",
          6180 => x"18",
          6181 => x"08",
          6182 => x"72",
          6183 => x"38",
          6184 => x"58",
          6185 => x"89",
          6186 => x"18",
          6187 => x"ff",
          6188 => x"05",
          6189 => x"80",
          6190 => x"d4",
          6191 => x"3d",
          6192 => x"3d",
          6193 => x"08",
          6194 => x"a0",
          6195 => x"54",
          6196 => x"77",
          6197 => x"80",
          6198 => x"0c",
          6199 => x"53",
          6200 => x"80",
          6201 => x"38",
          6202 => x"06",
          6203 => x"b5",
          6204 => x"98",
          6205 => x"14",
          6206 => x"92",
          6207 => x"2a",
          6208 => x"56",
          6209 => x"26",
          6210 => x"80",
          6211 => x"16",
          6212 => x"77",
          6213 => x"53",
          6214 => x"38",
          6215 => x"51",
          6216 => x"82",
          6217 => x"53",
          6218 => x"0b",
          6219 => x"08",
          6220 => x"38",
          6221 => x"d4",
          6222 => x"2e",
          6223 => x"9c",
          6224 => x"d4",
          6225 => x"80",
          6226 => x"8a",
          6227 => x"15",
          6228 => x"80",
          6229 => x"14",
          6230 => x"51",
          6231 => x"82",
          6232 => x"53",
          6233 => x"d4",
          6234 => x"2e",
          6235 => x"82",
          6236 => x"f8",
          6237 => x"ba",
          6238 => x"82",
          6239 => x"ff",
          6240 => x"82",
          6241 => x"52",
          6242 => x"f3",
          6243 => x"f8",
          6244 => x"72",
          6245 => x"72",
          6246 => x"f2",
          6247 => x"d4",
          6248 => x"15",
          6249 => x"15",
          6250 => x"b8",
          6251 => x"0c",
          6252 => x"82",
          6253 => x"8a",
          6254 => x"f7",
          6255 => x"7d",
          6256 => x"5b",
          6257 => x"76",
          6258 => x"3f",
          6259 => x"08",
          6260 => x"f8",
          6261 => x"38",
          6262 => x"08",
          6263 => x"08",
          6264 => x"f0",
          6265 => x"d4",
          6266 => x"82",
          6267 => x"80",
          6268 => x"d4",
          6269 => x"18",
          6270 => x"51",
          6271 => x"81",
          6272 => x"81",
          6273 => x"81",
          6274 => x"f8",
          6275 => x"83",
          6276 => x"77",
          6277 => x"72",
          6278 => x"38",
          6279 => x"75",
          6280 => x"81",
          6281 => x"a5",
          6282 => x"f8",
          6283 => x"52",
          6284 => x"8e",
          6285 => x"f8",
          6286 => x"d4",
          6287 => x"2e",
          6288 => x"73",
          6289 => x"81",
          6290 => x"87",
          6291 => x"d4",
          6292 => x"3d",
          6293 => x"3d",
          6294 => x"11",
          6295 => x"ae",
          6296 => x"f8",
          6297 => x"ff",
          6298 => x"33",
          6299 => x"71",
          6300 => x"81",
          6301 => x"94",
          6302 => x"92",
          6303 => x"f8",
          6304 => x"73",
          6305 => x"82",
          6306 => x"85",
          6307 => x"fc",
          6308 => x"79",
          6309 => x"ff",
          6310 => x"12",
          6311 => x"eb",
          6312 => x"70",
          6313 => x"72",
          6314 => x"81",
          6315 => x"73",
          6316 => x"94",
          6317 => x"98",
          6318 => x"0d",
          6319 => x"0d",
          6320 => x"51",
          6321 => x"81",
          6322 => x"80",
          6323 => x"70",
          6324 => x"33",
          6325 => x"81",
          6326 => x"16",
          6327 => x"51",
          6328 => x"70",
          6329 => x"0c",
          6330 => x"04",
          6331 => x"60",
          6332 => x"84",
          6333 => x"5b",
          6334 => x"5d",
          6335 => x"08",
          6336 => x"80",
          6337 => x"08",
          6338 => x"ed",
          6339 => x"d4",
          6340 => x"82",
          6341 => x"82",
          6342 => x"19",
          6343 => x"55",
          6344 => x"38",
          6345 => x"dc",
          6346 => x"33",
          6347 => x"81",
          6348 => x"53",
          6349 => x"34",
          6350 => x"08",
          6351 => x"e5",
          6352 => x"06",
          6353 => x"56",
          6354 => x"08",
          6355 => x"2e",
          6356 => x"83",
          6357 => x"75",
          6358 => x"72",
          6359 => x"d4",
          6360 => x"df",
          6361 => x"72",
          6362 => x"81",
          6363 => x"81",
          6364 => x"2e",
          6365 => x"ff",
          6366 => x"39",
          6367 => x"09",
          6368 => x"ca",
          6369 => x"2a",
          6370 => x"51",
          6371 => x"2e",
          6372 => x"15",
          6373 => x"bf",
          6374 => x"1c",
          6375 => x"0c",
          6376 => x"73",
          6377 => x"81",
          6378 => x"38",
          6379 => x"53",
          6380 => x"09",
          6381 => x"8f",
          6382 => x"08",
          6383 => x"5a",
          6384 => x"82",
          6385 => x"83",
          6386 => x"53",
          6387 => x"38",
          6388 => x"81",
          6389 => x"29",
          6390 => x"54",
          6391 => x"58",
          6392 => x"17",
          6393 => x"51",
          6394 => x"82",
          6395 => x"83",
          6396 => x"56",
          6397 => x"96",
          6398 => x"fe",
          6399 => x"38",
          6400 => x"76",
          6401 => x"73",
          6402 => x"54",
          6403 => x"83",
          6404 => x"09",
          6405 => x"38",
          6406 => x"8c",
          6407 => x"38",
          6408 => x"86",
          6409 => x"06",
          6410 => x"72",
          6411 => x"38",
          6412 => x"26",
          6413 => x"10",
          6414 => x"73",
          6415 => x"70",
          6416 => x"51",
          6417 => x"81",
          6418 => x"5c",
          6419 => x"93",
          6420 => x"fc",
          6421 => x"d4",
          6422 => x"ff",
          6423 => x"7d",
          6424 => x"ff",
          6425 => x"0c",
          6426 => x"52",
          6427 => x"d2",
          6428 => x"f8",
          6429 => x"d4",
          6430 => x"38",
          6431 => x"fd",
          6432 => x"39",
          6433 => x"1a",
          6434 => x"d4",
          6435 => x"3d",
          6436 => x"3d",
          6437 => x"08",
          6438 => x"52",
          6439 => x"d7",
          6440 => x"f8",
          6441 => x"d4",
          6442 => x"a4",
          6443 => x"70",
          6444 => x"0b",
          6445 => x"98",
          6446 => x"7e",
          6447 => x"3f",
          6448 => x"08",
          6449 => x"f8",
          6450 => x"38",
          6451 => x"70",
          6452 => x"75",
          6453 => x"58",
          6454 => x"8b",
          6455 => x"06",
          6456 => x"06",
          6457 => x"86",
          6458 => x"81",
          6459 => x"c3",
          6460 => x"2a",
          6461 => x"51",
          6462 => x"2e",
          6463 => x"82",
          6464 => x"8f",
          6465 => x"06",
          6466 => x"ab",
          6467 => x"86",
          6468 => x"06",
          6469 => x"73",
          6470 => x"75",
          6471 => x"81",
          6472 => x"73",
          6473 => x"38",
          6474 => x"76",
          6475 => x"70",
          6476 => x"ac",
          6477 => x"5d",
          6478 => x"2e",
          6479 => x"81",
          6480 => x"17",
          6481 => x"76",
          6482 => x"06",
          6483 => x"8c",
          6484 => x"18",
          6485 => x"b6",
          6486 => x"f8",
          6487 => x"ff",
          6488 => x"81",
          6489 => x"33",
          6490 => x"8d",
          6491 => x"59",
          6492 => x"5c",
          6493 => x"80",
          6494 => x"05",
          6495 => x"3f",
          6496 => x"08",
          6497 => x"06",
          6498 => x"2e",
          6499 => x"81",
          6500 => x"e6",
          6501 => x"80",
          6502 => x"82",
          6503 => x"78",
          6504 => x"22",
          6505 => x"19",
          6506 => x"df",
          6507 => x"82",
          6508 => x"2e",
          6509 => x"80",
          6510 => x"5a",
          6511 => x"83",
          6512 => x"09",
          6513 => x"38",
          6514 => x"8c",
          6515 => x"a5",
          6516 => x"70",
          6517 => x"81",
          6518 => x"57",
          6519 => x"90",
          6520 => x"2e",
          6521 => x"10",
          6522 => x"51",
          6523 => x"38",
          6524 => x"81",
          6525 => x"54",
          6526 => x"ff",
          6527 => x"bb",
          6528 => x"38",
          6529 => x"b5",
          6530 => x"f8",
          6531 => x"06",
          6532 => x"2e",
          6533 => x"19",
          6534 => x"54",
          6535 => x"8b",
          6536 => x"52",
          6537 => x"51",
          6538 => x"82",
          6539 => x"80",
          6540 => x"81",
          6541 => x"0b",
          6542 => x"80",
          6543 => x"f5",
          6544 => x"d4",
          6545 => x"82",
          6546 => x"80",
          6547 => x"38",
          6548 => x"f8",
          6549 => x"0d",
          6550 => x"0d",
          6551 => x"ab",
          6552 => x"a0",
          6553 => x"5a",
          6554 => x"85",
          6555 => x"8c",
          6556 => x"22",
          6557 => x"73",
          6558 => x"38",
          6559 => x"10",
          6560 => x"51",
          6561 => x"39",
          6562 => x"1a",
          6563 => x"3d",
          6564 => x"59",
          6565 => x"02",
          6566 => x"33",
          6567 => x"73",
          6568 => x"a8",
          6569 => x"0b",
          6570 => x"81",
          6571 => x"08",
          6572 => x"8b",
          6573 => x"78",
          6574 => x"3f",
          6575 => x"80",
          6576 => x"56",
          6577 => x"83",
          6578 => x"55",
          6579 => x"2e",
          6580 => x"83",
          6581 => x"82",
          6582 => x"8f",
          6583 => x"06",
          6584 => x"75",
          6585 => x"90",
          6586 => x"06",
          6587 => x"56",
          6588 => x"87",
          6589 => x"a0",
          6590 => x"ff",
          6591 => x"80",
          6592 => x"c0",
          6593 => x"87",
          6594 => x"bf",
          6595 => x"74",
          6596 => x"06",
          6597 => x"27",
          6598 => x"14",
          6599 => x"34",
          6600 => x"18",
          6601 => x"57",
          6602 => x"e3",
          6603 => x"ec",
          6604 => x"80",
          6605 => x"80",
          6606 => x"38",
          6607 => x"73",
          6608 => x"38",
          6609 => x"33",
          6610 => x"e0",
          6611 => x"f8",
          6612 => x"8c",
          6613 => x"54",
          6614 => x"94",
          6615 => x"55",
          6616 => x"74",
          6617 => x"38",
          6618 => x"33",
          6619 => x"39",
          6620 => x"05",
          6621 => x"78",
          6622 => x"56",
          6623 => x"76",
          6624 => x"38",
          6625 => x"15",
          6626 => x"55",
          6627 => x"34",
          6628 => x"e3",
          6629 => x"f9",
          6630 => x"d4",
          6631 => x"38",
          6632 => x"80",
          6633 => x"fe",
          6634 => x"55",
          6635 => x"2e",
          6636 => x"82",
          6637 => x"55",
          6638 => x"08",
          6639 => x"81",
          6640 => x"38",
          6641 => x"05",
          6642 => x"34",
          6643 => x"05",
          6644 => x"2a",
          6645 => x"51",
          6646 => x"59",
          6647 => x"90",
          6648 => x"8c",
          6649 => x"f8",
          6650 => x"d4",
          6651 => x"59",
          6652 => x"51",
          6653 => x"82",
          6654 => x"57",
          6655 => x"08",
          6656 => x"ff",
          6657 => x"80",
          6658 => x"38",
          6659 => x"90",
          6660 => x"31",
          6661 => x"51",
          6662 => x"82",
          6663 => x"57",
          6664 => x"08",
          6665 => x"a0",
          6666 => x"91",
          6667 => x"f8",
          6668 => x"06",
          6669 => x"08",
          6670 => x"e3",
          6671 => x"d4",
          6672 => x"82",
          6673 => x"81",
          6674 => x"1c",
          6675 => x"08",
          6676 => x"06",
          6677 => x"7c",
          6678 => x"8f",
          6679 => x"34",
          6680 => x"08",
          6681 => x"82",
          6682 => x"52",
          6683 => x"df",
          6684 => x"8d",
          6685 => x"77",
          6686 => x"83",
          6687 => x"8b",
          6688 => x"1b",
          6689 => x"17",
          6690 => x"73",
          6691 => x"80",
          6692 => x"05",
          6693 => x"3f",
          6694 => x"83",
          6695 => x"81",
          6696 => x"77",
          6697 => x"73",
          6698 => x"2e",
          6699 => x"10",
          6700 => x"51",
          6701 => x"38",
          6702 => x"07",
          6703 => x"34",
          6704 => x"1d",
          6705 => x"79",
          6706 => x"3f",
          6707 => x"08",
          6708 => x"f8",
          6709 => x"38",
          6710 => x"78",
          6711 => x"98",
          6712 => x"7b",
          6713 => x"3f",
          6714 => x"08",
          6715 => x"f8",
          6716 => x"a0",
          6717 => x"f8",
          6718 => x"1a",
          6719 => x"c0",
          6720 => x"a0",
          6721 => x"1a",
          6722 => x"91",
          6723 => x"08",
          6724 => x"98",
          6725 => x"73",
          6726 => x"81",
          6727 => x"34",
          6728 => x"82",
          6729 => x"94",
          6730 => x"fa",
          6731 => x"70",
          6732 => x"08",
          6733 => x"56",
          6734 => x"72",
          6735 => x"38",
          6736 => x"51",
          6737 => x"82",
          6738 => x"54",
          6739 => x"08",
          6740 => x"98",
          6741 => x"75",
          6742 => x"3f",
          6743 => x"08",
          6744 => x"f8",
          6745 => x"9c",
          6746 => x"e5",
          6747 => x"0b",
          6748 => x"90",
          6749 => x"27",
          6750 => x"d4",
          6751 => x"74",
          6752 => x"3f",
          6753 => x"08",
          6754 => x"f8",
          6755 => x"c3",
          6756 => x"2e",
          6757 => x"83",
          6758 => x"73",
          6759 => x"0c",
          6760 => x"04",
          6761 => x"7e",
          6762 => x"5f",
          6763 => x"0b",
          6764 => x"98",
          6765 => x"2e",
          6766 => x"ac",
          6767 => x"2e",
          6768 => x"80",
          6769 => x"8c",
          6770 => x"22",
          6771 => x"5c",
          6772 => x"2e",
          6773 => x"78",
          6774 => x"22",
          6775 => x"56",
          6776 => x"38",
          6777 => x"15",
          6778 => x"ff",
          6779 => x"72",
          6780 => x"86",
          6781 => x"80",
          6782 => x"18",
          6783 => x"ff",
          6784 => x"5b",
          6785 => x"52",
          6786 => x"75",
          6787 => x"d5",
          6788 => x"d4",
          6789 => x"ff",
          6790 => x"81",
          6791 => x"95",
          6792 => x"27",
          6793 => x"88",
          6794 => x"7a",
          6795 => x"15",
          6796 => x"9f",
          6797 => x"76",
          6798 => x"07",
          6799 => x"80",
          6800 => x"54",
          6801 => x"2e",
          6802 => x"57",
          6803 => x"7a",
          6804 => x"74",
          6805 => x"5b",
          6806 => x"79",
          6807 => x"22",
          6808 => x"72",
          6809 => x"7a",
          6810 => x"25",
          6811 => x"06",
          6812 => x"77",
          6813 => x"53",
          6814 => x"14",
          6815 => x"89",
          6816 => x"57",
          6817 => x"19",
          6818 => x"1b",
          6819 => x"74",
          6820 => x"38",
          6821 => x"09",
          6822 => x"38",
          6823 => x"78",
          6824 => x"30",
          6825 => x"80",
          6826 => x"54",
          6827 => x"90",
          6828 => x"2e",
          6829 => x"76",
          6830 => x"58",
          6831 => x"57",
          6832 => x"81",
          6833 => x"81",
          6834 => x"79",
          6835 => x"38",
          6836 => x"05",
          6837 => x"81",
          6838 => x"18",
          6839 => x"81",
          6840 => x"8b",
          6841 => x"96",
          6842 => x"57",
          6843 => x"72",
          6844 => x"33",
          6845 => x"72",
          6846 => x"d3",
          6847 => x"89",
          6848 => x"73",
          6849 => x"11",
          6850 => x"99",
          6851 => x"9c",
          6852 => x"11",
          6853 => x"88",
          6854 => x"38",
          6855 => x"53",
          6856 => x"83",
          6857 => x"81",
          6858 => x"80",
          6859 => x"a0",
          6860 => x"ff",
          6861 => x"53",
          6862 => x"81",
          6863 => x"81",
          6864 => x"81",
          6865 => x"56",
          6866 => x"72",
          6867 => x"77",
          6868 => x"53",
          6869 => x"14",
          6870 => x"08",
          6871 => x"51",
          6872 => x"38",
          6873 => x"34",
          6874 => x"53",
          6875 => x"88",
          6876 => x"1c",
          6877 => x"52",
          6878 => x"3f",
          6879 => x"08",
          6880 => x"13",
          6881 => x"3f",
          6882 => x"08",
          6883 => x"98",
          6884 => x"fa",
          6885 => x"f8",
          6886 => x"23",
          6887 => x"04",
          6888 => x"62",
          6889 => x"5e",
          6890 => x"33",
          6891 => x"73",
          6892 => x"38",
          6893 => x"80",
          6894 => x"38",
          6895 => x"8d",
          6896 => x"05",
          6897 => x"0c",
          6898 => x"15",
          6899 => x"70",
          6900 => x"56",
          6901 => x"09",
          6902 => x"38",
          6903 => x"80",
          6904 => x"30",
          6905 => x"78",
          6906 => x"54",
          6907 => x"73",
          6908 => x"63",
          6909 => x"54",
          6910 => x"96",
          6911 => x"0b",
          6912 => x"80",
          6913 => x"e7",
          6914 => x"d4",
          6915 => x"87",
          6916 => x"41",
          6917 => x"11",
          6918 => x"80",
          6919 => x"fc",
          6920 => x"8f",
          6921 => x"f8",
          6922 => x"82",
          6923 => x"ff",
          6924 => x"d4",
          6925 => x"92",
          6926 => x"1a",
          6927 => x"08",
          6928 => x"55",
          6929 => x"81",
          6930 => x"d4",
          6931 => x"ff",
          6932 => x"af",
          6933 => x"9f",
          6934 => x"80",
          6935 => x"51",
          6936 => x"b4",
          6937 => x"dc",
          6938 => x"75",
          6939 => x"91",
          6940 => x"82",
          6941 => x"d9",
          6942 => x"d4",
          6943 => x"de",
          6944 => x"fe",
          6945 => x"38",
          6946 => x"54",
          6947 => x"81",
          6948 => x"89",
          6949 => x"41",
          6950 => x"33",
          6951 => x"73",
          6952 => x"81",
          6953 => x"81",
          6954 => x"dc",
          6955 => x"70",
          6956 => x"07",
          6957 => x"73",
          6958 => x"44",
          6959 => x"82",
          6960 => x"81",
          6961 => x"06",
          6962 => x"22",
          6963 => x"2e",
          6964 => x"d2",
          6965 => x"2e",
          6966 => x"80",
          6967 => x"1a",
          6968 => x"ae",
          6969 => x"06",
          6970 => x"79",
          6971 => x"ae",
          6972 => x"06",
          6973 => x"10",
          6974 => x"74",
          6975 => x"a0",
          6976 => x"ae",
          6977 => x"26",
          6978 => x"54",
          6979 => x"81",
          6980 => x"81",
          6981 => x"78",
          6982 => x"76",
          6983 => x"73",
          6984 => x"84",
          6985 => x"80",
          6986 => x"78",
          6987 => x"05",
          6988 => x"fe",
          6989 => x"a0",
          6990 => x"70",
          6991 => x"51",
          6992 => x"54",
          6993 => x"84",
          6994 => x"38",
          6995 => x"78",
          6996 => x"19",
          6997 => x"56",
          6998 => x"78",
          6999 => x"56",
          7000 => x"76",
          7001 => x"83",
          7002 => x"7a",
          7003 => x"ff",
          7004 => x"56",
          7005 => x"2e",
          7006 => x"93",
          7007 => x"70",
          7008 => x"22",
          7009 => x"73",
          7010 => x"38",
          7011 => x"74",
          7012 => x"06",
          7013 => x"2e",
          7014 => x"85",
          7015 => x"07",
          7016 => x"2e",
          7017 => x"16",
          7018 => x"22",
          7019 => x"ae",
          7020 => x"78",
          7021 => x"05",
          7022 => x"59",
          7023 => x"8f",
          7024 => x"70",
          7025 => x"73",
          7026 => x"81",
          7027 => x"8b",
          7028 => x"a0",
          7029 => x"e8",
          7030 => x"59",
          7031 => x"7c",
          7032 => x"22",
          7033 => x"57",
          7034 => x"2e",
          7035 => x"75",
          7036 => x"38",
          7037 => x"70",
          7038 => x"25",
          7039 => x"7c",
          7040 => x"38",
          7041 => x"89",
          7042 => x"07",
          7043 => x"80",
          7044 => x"7e",
          7045 => x"38",
          7046 => x"79",
          7047 => x"70",
          7048 => x"25",
          7049 => x"51",
          7050 => x"73",
          7051 => x"38",
          7052 => x"fe",
          7053 => x"79",
          7054 => x"76",
          7055 => x"7c",
          7056 => x"be",
          7057 => x"88",
          7058 => x"82",
          7059 => x"06",
          7060 => x"8b",
          7061 => x"76",
          7062 => x"76",
          7063 => x"83",
          7064 => x"51",
          7065 => x"3f",
          7066 => x"08",
          7067 => x"06",
          7068 => x"70",
          7069 => x"55",
          7070 => x"2e",
          7071 => x"80",
          7072 => x"c7",
          7073 => x"57",
          7074 => x"76",
          7075 => x"ff",
          7076 => x"78",
          7077 => x"76",
          7078 => x"59",
          7079 => x"39",
          7080 => x"05",
          7081 => x"55",
          7082 => x"34",
          7083 => x"80",
          7084 => x"80",
          7085 => x"75",
          7086 => x"a8",
          7087 => x"3f",
          7088 => x"08",
          7089 => x"38",
          7090 => x"83",
          7091 => x"a4",
          7092 => x"16",
          7093 => x"26",
          7094 => x"82",
          7095 => x"9f",
          7096 => x"99",
          7097 => x"7b",
          7098 => x"17",
          7099 => x"ff",
          7100 => x"5c",
          7101 => x"05",
          7102 => x"34",
          7103 => x"fd",
          7104 => x"1e",
          7105 => x"81",
          7106 => x"81",
          7107 => x"85",
          7108 => x"34",
          7109 => x"09",
          7110 => x"38",
          7111 => x"81",
          7112 => x"7b",
          7113 => x"73",
          7114 => x"38",
          7115 => x"54",
          7116 => x"09",
          7117 => x"38",
          7118 => x"57",
          7119 => x"70",
          7120 => x"54",
          7121 => x"7b",
          7122 => x"73",
          7123 => x"38",
          7124 => x"57",
          7125 => x"70",
          7126 => x"54",
          7127 => x"85",
          7128 => x"07",
          7129 => x"1f",
          7130 => x"ea",
          7131 => x"d4",
          7132 => x"1f",
          7133 => x"82",
          7134 => x"80",
          7135 => x"82",
          7136 => x"84",
          7137 => x"06",
          7138 => x"74",
          7139 => x"81",
          7140 => x"2a",
          7141 => x"73",
          7142 => x"38",
          7143 => x"54",
          7144 => x"f8",
          7145 => x"80",
          7146 => x"34",
          7147 => x"c2",
          7148 => x"06",
          7149 => x"38",
          7150 => x"39",
          7151 => x"70",
          7152 => x"54",
          7153 => x"86",
          7154 => x"84",
          7155 => x"06",
          7156 => x"73",
          7157 => x"38",
          7158 => x"83",
          7159 => x"05",
          7160 => x"7f",
          7161 => x"3f",
          7162 => x"08",
          7163 => x"f8",
          7164 => x"82",
          7165 => x"92",
          7166 => x"f6",
          7167 => x"5b",
          7168 => x"70",
          7169 => x"59",
          7170 => x"73",
          7171 => x"c6",
          7172 => x"81",
          7173 => x"70",
          7174 => x"52",
          7175 => x"8d",
          7176 => x"38",
          7177 => x"09",
          7178 => x"a5",
          7179 => x"d0",
          7180 => x"ff",
          7181 => x"53",
          7182 => x"91",
          7183 => x"73",
          7184 => x"d0",
          7185 => x"71",
          7186 => x"f7",
          7187 => x"82",
          7188 => x"55",
          7189 => x"55",
          7190 => x"81",
          7191 => x"74",
          7192 => x"56",
          7193 => x"12",
          7194 => x"70",
          7195 => x"38",
          7196 => x"81",
          7197 => x"51",
          7198 => x"51",
          7199 => x"89",
          7200 => x"70",
          7201 => x"53",
          7202 => x"70",
          7203 => x"51",
          7204 => x"09",
          7205 => x"38",
          7206 => x"38",
          7207 => x"77",
          7208 => x"70",
          7209 => x"2a",
          7210 => x"07",
          7211 => x"51",
          7212 => x"8f",
          7213 => x"84",
          7214 => x"83",
          7215 => x"94",
          7216 => x"74",
          7217 => x"38",
          7218 => x"0c",
          7219 => x"86",
          7220 => x"d4",
          7221 => x"82",
          7222 => x"8c",
          7223 => x"fa",
          7224 => x"56",
          7225 => x"17",
          7226 => x"b4",
          7227 => x"52",
          7228 => x"f4",
          7229 => x"82",
          7230 => x"81",
          7231 => x"b6",
          7232 => x"8a",
          7233 => x"f8",
          7234 => x"ff",
          7235 => x"55",
          7236 => x"d5",
          7237 => x"06",
          7238 => x"80",
          7239 => x"33",
          7240 => x"81",
          7241 => x"81",
          7242 => x"81",
          7243 => x"eb",
          7244 => x"70",
          7245 => x"07",
          7246 => x"73",
          7247 => x"81",
          7248 => x"81",
          7249 => x"83",
          7250 => x"b0",
          7251 => x"16",
          7252 => x"3f",
          7253 => x"08",
          7254 => x"f8",
          7255 => x"9d",
          7256 => x"82",
          7257 => x"81",
          7258 => x"ce",
          7259 => x"d4",
          7260 => x"82",
          7261 => x"80",
          7262 => x"82",
          7263 => x"d4",
          7264 => x"3d",
          7265 => x"3d",
          7266 => x"84",
          7267 => x"05",
          7268 => x"80",
          7269 => x"51",
          7270 => x"82",
          7271 => x"58",
          7272 => x"0b",
          7273 => x"08",
          7274 => x"38",
          7275 => x"08",
          7276 => x"ec",
          7277 => x"08",
          7278 => x"56",
          7279 => x"86",
          7280 => x"75",
          7281 => x"fe",
          7282 => x"54",
          7283 => x"2e",
          7284 => x"14",
          7285 => x"a0",
          7286 => x"f8",
          7287 => x"06",
          7288 => x"54",
          7289 => x"38",
          7290 => x"86",
          7291 => x"82",
          7292 => x"06",
          7293 => x"56",
          7294 => x"38",
          7295 => x"80",
          7296 => x"81",
          7297 => x"52",
          7298 => x"51",
          7299 => x"82",
          7300 => x"81",
          7301 => x"81",
          7302 => x"83",
          7303 => x"8f",
          7304 => x"2e",
          7305 => x"82",
          7306 => x"06",
          7307 => x"56",
          7308 => x"38",
          7309 => x"74",
          7310 => x"a3",
          7311 => x"f8",
          7312 => x"06",
          7313 => x"2e",
          7314 => x"80",
          7315 => x"3d",
          7316 => x"83",
          7317 => x"15",
          7318 => x"53",
          7319 => x"8d",
          7320 => x"15",
          7321 => x"3f",
          7322 => x"08",
          7323 => x"70",
          7324 => x"0c",
          7325 => x"16",
          7326 => x"80",
          7327 => x"80",
          7328 => x"54",
          7329 => x"84",
          7330 => x"5b",
          7331 => x"80",
          7332 => x"7a",
          7333 => x"fc",
          7334 => x"d4",
          7335 => x"ff",
          7336 => x"77",
          7337 => x"81",
          7338 => x"76",
          7339 => x"81",
          7340 => x"2e",
          7341 => x"8d",
          7342 => x"26",
          7343 => x"80",
          7344 => x"ca",
          7345 => x"d4",
          7346 => x"ff",
          7347 => x"72",
          7348 => x"09",
          7349 => x"d7",
          7350 => x"14",
          7351 => x"3f",
          7352 => x"08",
          7353 => x"06",
          7354 => x"38",
          7355 => x"51",
          7356 => x"82",
          7357 => x"58",
          7358 => x"0c",
          7359 => x"33",
          7360 => x"80",
          7361 => x"ff",
          7362 => x"ff",
          7363 => x"55",
          7364 => x"81",
          7365 => x"38",
          7366 => x"06",
          7367 => x"80",
          7368 => x"52",
          7369 => x"8a",
          7370 => x"80",
          7371 => x"ff",
          7372 => x"53",
          7373 => x"86",
          7374 => x"83",
          7375 => x"c9",
          7376 => x"ca",
          7377 => x"f8",
          7378 => x"d4",
          7379 => x"15",
          7380 => x"06",
          7381 => x"76",
          7382 => x"80",
          7383 => x"c9",
          7384 => x"d4",
          7385 => x"ff",
          7386 => x"74",
          7387 => x"d8",
          7388 => x"b1",
          7389 => x"f8",
          7390 => x"c6",
          7391 => x"8e",
          7392 => x"f8",
          7393 => x"ff",
          7394 => x"56",
          7395 => x"83",
          7396 => x"14",
          7397 => x"71",
          7398 => x"5a",
          7399 => x"26",
          7400 => x"8a",
          7401 => x"74",
          7402 => x"fe",
          7403 => x"82",
          7404 => x"55",
          7405 => x"08",
          7406 => x"f3",
          7407 => x"f8",
          7408 => x"ff",
          7409 => x"83",
          7410 => x"74",
          7411 => x"26",
          7412 => x"57",
          7413 => x"26",
          7414 => x"57",
          7415 => x"56",
          7416 => x"82",
          7417 => x"15",
          7418 => x"0c",
          7419 => x"0c",
          7420 => x"a8",
          7421 => x"1d",
          7422 => x"54",
          7423 => x"2e",
          7424 => x"af",
          7425 => x"14",
          7426 => x"3f",
          7427 => x"08",
          7428 => x"06",
          7429 => x"72",
          7430 => x"79",
          7431 => x"80",
          7432 => x"c8",
          7433 => x"d4",
          7434 => x"15",
          7435 => x"2b",
          7436 => x"8d",
          7437 => x"2e",
          7438 => x"77",
          7439 => x"0c",
          7440 => x"76",
          7441 => x"38",
          7442 => x"70",
          7443 => x"81",
          7444 => x"53",
          7445 => x"89",
          7446 => x"56",
          7447 => x"08",
          7448 => x"38",
          7449 => x"15",
          7450 => x"90",
          7451 => x"80",
          7452 => x"34",
          7453 => x"09",
          7454 => x"92",
          7455 => x"14",
          7456 => x"3f",
          7457 => x"08",
          7458 => x"06",
          7459 => x"2e",
          7460 => x"80",
          7461 => x"1b",
          7462 => x"ca",
          7463 => x"d4",
          7464 => x"ea",
          7465 => x"f8",
          7466 => x"34",
          7467 => x"51",
          7468 => x"82",
          7469 => x"83",
          7470 => x"53",
          7471 => x"d5",
          7472 => x"06",
          7473 => x"b8",
          7474 => x"d9",
          7475 => x"f8",
          7476 => x"85",
          7477 => x"09",
          7478 => x"38",
          7479 => x"51",
          7480 => x"82",
          7481 => x"86",
          7482 => x"f2",
          7483 => x"06",
          7484 => x"a0",
          7485 => x"ad",
          7486 => x"f8",
          7487 => x"0c",
          7488 => x"51",
          7489 => x"82",
          7490 => x"90",
          7491 => x"74",
          7492 => x"d0",
          7493 => x"53",
          7494 => x"d0",
          7495 => x"15",
          7496 => x"d8",
          7497 => x"0c",
          7498 => x"15",
          7499 => x"75",
          7500 => x"0c",
          7501 => x"04",
          7502 => x"77",
          7503 => x"73",
          7504 => x"38",
          7505 => x"72",
          7506 => x"38",
          7507 => x"71",
          7508 => x"38",
          7509 => x"84",
          7510 => x"52",
          7511 => x"09",
          7512 => x"38",
          7513 => x"51",
          7514 => x"3f",
          7515 => x"08",
          7516 => x"71",
          7517 => x"74",
          7518 => x"83",
          7519 => x"78",
          7520 => x"52",
          7521 => x"f8",
          7522 => x"0d",
          7523 => x"0d",
          7524 => x"33",
          7525 => x"3d",
          7526 => x"56",
          7527 => x"8b",
          7528 => x"82",
          7529 => x"24",
          7530 => x"d4",
          7531 => x"29",
          7532 => x"05",
          7533 => x"55",
          7534 => x"84",
          7535 => x"34",
          7536 => x"80",
          7537 => x"80",
          7538 => x"75",
          7539 => x"75",
          7540 => x"38",
          7541 => x"3d",
          7542 => x"05",
          7543 => x"3f",
          7544 => x"08",
          7545 => x"d4",
          7546 => x"3d",
          7547 => x"3d",
          7548 => x"84",
          7549 => x"05",
          7550 => x"89",
          7551 => x"2e",
          7552 => x"77",
          7553 => x"54",
          7554 => x"05",
          7555 => x"84",
          7556 => x"f6",
          7557 => x"d4",
          7558 => x"82",
          7559 => x"84",
          7560 => x"5c",
          7561 => x"3d",
          7562 => x"ea",
          7563 => x"d4",
          7564 => x"82",
          7565 => x"92",
          7566 => x"d7",
          7567 => x"98",
          7568 => x"73",
          7569 => x"38",
          7570 => x"9c",
          7571 => x"80",
          7572 => x"38",
          7573 => x"95",
          7574 => x"2e",
          7575 => x"aa",
          7576 => x"df",
          7577 => x"d4",
          7578 => x"9e",
          7579 => x"05",
          7580 => x"54",
          7581 => x"38",
          7582 => x"70",
          7583 => x"54",
          7584 => x"8e",
          7585 => x"83",
          7586 => x"88",
          7587 => x"83",
          7588 => x"83",
          7589 => x"06",
          7590 => x"80",
          7591 => x"38",
          7592 => x"51",
          7593 => x"82",
          7594 => x"56",
          7595 => x"0a",
          7596 => x"05",
          7597 => x"3f",
          7598 => x"0b",
          7599 => x"80",
          7600 => x"7a",
          7601 => x"3f",
          7602 => x"9c",
          7603 => x"9e",
          7604 => x"81",
          7605 => x"34",
          7606 => x"80",
          7607 => x"b4",
          7608 => x"54",
          7609 => x"52",
          7610 => x"05",
          7611 => x"3f",
          7612 => x"08",
          7613 => x"f8",
          7614 => x"38",
          7615 => x"82",
          7616 => x"b2",
          7617 => x"84",
          7618 => x"06",
          7619 => x"73",
          7620 => x"38",
          7621 => x"ad",
          7622 => x"2a",
          7623 => x"51",
          7624 => x"2e",
          7625 => x"81",
          7626 => x"80",
          7627 => x"87",
          7628 => x"39",
          7629 => x"51",
          7630 => x"82",
          7631 => x"7b",
          7632 => x"12",
          7633 => x"82",
          7634 => x"81",
          7635 => x"83",
          7636 => x"06",
          7637 => x"80",
          7638 => x"77",
          7639 => x"58",
          7640 => x"08",
          7641 => x"63",
          7642 => x"63",
          7643 => x"57",
          7644 => x"82",
          7645 => x"82",
          7646 => x"88",
          7647 => x"9c",
          7648 => x"c1",
          7649 => x"d4",
          7650 => x"d4",
          7651 => x"1b",
          7652 => x"0c",
          7653 => x"22",
          7654 => x"77",
          7655 => x"80",
          7656 => x"34",
          7657 => x"1a",
          7658 => x"94",
          7659 => x"85",
          7660 => x"06",
          7661 => x"80",
          7662 => x"38",
          7663 => x"08",
          7664 => x"84",
          7665 => x"f8",
          7666 => x"0c",
          7667 => x"70",
          7668 => x"52",
          7669 => x"39",
          7670 => x"51",
          7671 => x"82",
          7672 => x"57",
          7673 => x"08",
          7674 => x"38",
          7675 => x"d4",
          7676 => x"2e",
          7677 => x"83",
          7678 => x"75",
          7679 => x"74",
          7680 => x"07",
          7681 => x"54",
          7682 => x"8a",
          7683 => x"75",
          7684 => x"73",
          7685 => x"98",
          7686 => x"a9",
          7687 => x"ff",
          7688 => x"80",
          7689 => x"76",
          7690 => x"c5",
          7691 => x"d4",
          7692 => x"38",
          7693 => x"39",
          7694 => x"82",
          7695 => x"05",
          7696 => x"84",
          7697 => x"0c",
          7698 => x"82",
          7699 => x"98",
          7700 => x"f2",
          7701 => x"63",
          7702 => x"40",
          7703 => x"7e",
          7704 => x"fc",
          7705 => x"51",
          7706 => x"82",
          7707 => x"55",
          7708 => x"08",
          7709 => x"19",
          7710 => x"80",
          7711 => x"74",
          7712 => x"39",
          7713 => x"81",
          7714 => x"56",
          7715 => x"82",
          7716 => x"39",
          7717 => x"1a",
          7718 => x"82",
          7719 => x"0b",
          7720 => x"81",
          7721 => x"39",
          7722 => x"94",
          7723 => x"55",
          7724 => x"83",
          7725 => x"7b",
          7726 => x"8c",
          7727 => x"08",
          7728 => x"06",
          7729 => x"81",
          7730 => x"8a",
          7731 => x"05",
          7732 => x"06",
          7733 => x"a8",
          7734 => x"38",
          7735 => x"55",
          7736 => x"19",
          7737 => x"51",
          7738 => x"82",
          7739 => x"55",
          7740 => x"ff",
          7741 => x"ff",
          7742 => x"38",
          7743 => x"0c",
          7744 => x"52",
          7745 => x"d6",
          7746 => x"f8",
          7747 => x"ff",
          7748 => x"d4",
          7749 => x"7c",
          7750 => x"57",
          7751 => x"80",
          7752 => x"1a",
          7753 => x"22",
          7754 => x"75",
          7755 => x"38",
          7756 => x"58",
          7757 => x"53",
          7758 => x"1b",
          7759 => x"b8",
          7760 => x"d4",
          7761 => x"d6",
          7762 => x"11",
          7763 => x"74",
          7764 => x"38",
          7765 => x"77",
          7766 => x"78",
          7767 => x"84",
          7768 => x"16",
          7769 => x"08",
          7770 => x"2b",
          7771 => x"ff",
          7772 => x"77",
          7773 => x"ba",
          7774 => x"1a",
          7775 => x"08",
          7776 => x"84",
          7777 => x"57",
          7778 => x"27",
          7779 => x"56",
          7780 => x"52",
          7781 => x"d0",
          7782 => x"f8",
          7783 => x"38",
          7784 => x"19",
          7785 => x"06",
          7786 => x"52",
          7787 => x"bd",
          7788 => x"76",
          7789 => x"17",
          7790 => x"1e",
          7791 => x"18",
          7792 => x"5e",
          7793 => x"39",
          7794 => x"82",
          7795 => x"90",
          7796 => x"f2",
          7797 => x"63",
          7798 => x"40",
          7799 => x"7e",
          7800 => x"fc",
          7801 => x"51",
          7802 => x"82",
          7803 => x"55",
          7804 => x"08",
          7805 => x"18",
          7806 => x"80",
          7807 => x"74",
          7808 => x"39",
          7809 => x"70",
          7810 => x"81",
          7811 => x"56",
          7812 => x"80",
          7813 => x"38",
          7814 => x"0b",
          7815 => x"82",
          7816 => x"39",
          7817 => x"19",
          7818 => x"83",
          7819 => x"18",
          7820 => x"56",
          7821 => x"27",
          7822 => x"09",
          7823 => x"2e",
          7824 => x"94",
          7825 => x"83",
          7826 => x"56",
          7827 => x"38",
          7828 => x"22",
          7829 => x"89",
          7830 => x"55",
          7831 => x"75",
          7832 => x"18",
          7833 => x"9c",
          7834 => x"85",
          7835 => x"08",
          7836 => x"c6",
          7837 => x"d4",
          7838 => x"82",
          7839 => x"80",
          7840 => x"38",
          7841 => x"ff",
          7842 => x"ff",
          7843 => x"38",
          7844 => x"0c",
          7845 => x"85",
          7846 => x"19",
          7847 => x"b4",
          7848 => x"19",
          7849 => x"81",
          7850 => x"74",
          7851 => x"c8",
          7852 => x"f8",
          7853 => x"38",
          7854 => x"52",
          7855 => x"9e",
          7856 => x"f8",
          7857 => x"fe",
          7858 => x"d4",
          7859 => x"7c",
          7860 => x"57",
          7861 => x"80",
          7862 => x"1b",
          7863 => x"22",
          7864 => x"75",
          7865 => x"38",
          7866 => x"59",
          7867 => x"53",
          7868 => x"1a",
          7869 => x"b7",
          7870 => x"d4",
          7871 => x"a4",
          7872 => x"11",
          7873 => x"56",
          7874 => x"27",
          7875 => x"80",
          7876 => x"08",
          7877 => x"2b",
          7878 => x"b8",
          7879 => x"ba",
          7880 => x"55",
          7881 => x"16",
          7882 => x"2b",
          7883 => x"39",
          7884 => x"94",
          7885 => x"94",
          7886 => x"ff",
          7887 => x"82",
          7888 => x"fd",
          7889 => x"77",
          7890 => x"55",
          7891 => x"0c",
          7892 => x"83",
          7893 => x"80",
          7894 => x"55",
          7895 => x"83",
          7896 => x"9c",
          7897 => x"7e",
          7898 => x"fc",
          7899 => x"f8",
          7900 => x"38",
          7901 => x"52",
          7902 => x"83",
          7903 => x"b8",
          7904 => x"ba",
          7905 => x"55",
          7906 => x"16",
          7907 => x"31",
          7908 => x"7f",
          7909 => x"94",
          7910 => x"70",
          7911 => x"8c",
          7912 => x"58",
          7913 => x"76",
          7914 => x"75",
          7915 => x"19",
          7916 => x"39",
          7917 => x"80",
          7918 => x"74",
          7919 => x"80",
          7920 => x"d4",
          7921 => x"3d",
          7922 => x"3d",
          7923 => x"3d",
          7924 => x"70",
          7925 => x"e0",
          7926 => x"f8",
          7927 => x"d4",
          7928 => x"80",
          7929 => x"33",
          7930 => x"70",
          7931 => x"55",
          7932 => x"2e",
          7933 => x"a0",
          7934 => x"78",
          7935 => x"e8",
          7936 => x"f8",
          7937 => x"d4",
          7938 => x"d8",
          7939 => x"08",
          7940 => x"a0",
          7941 => x"73",
          7942 => x"88",
          7943 => x"74",
          7944 => x"51",
          7945 => x"8c",
          7946 => x"9c",
          7947 => x"b8",
          7948 => x"88",
          7949 => x"96",
          7950 => x"b8",
          7951 => x"52",
          7952 => x"ff",
          7953 => x"78",
          7954 => x"83",
          7955 => x"51",
          7956 => x"3f",
          7957 => x"08",
          7958 => x"81",
          7959 => x"57",
          7960 => x"34",
          7961 => x"f8",
          7962 => x"0d",
          7963 => x"0d",
          7964 => x"54",
          7965 => x"82",
          7966 => x"53",
          7967 => x"08",
          7968 => x"3d",
          7969 => x"73",
          7970 => x"3f",
          7971 => x"08",
          7972 => x"f8",
          7973 => x"82",
          7974 => x"74",
          7975 => x"d4",
          7976 => x"3d",
          7977 => x"3d",
          7978 => x"51",
          7979 => x"8b",
          7980 => x"82",
          7981 => x"24",
          7982 => x"d4",
          7983 => x"ec",
          7984 => x"52",
          7985 => x"f8",
          7986 => x"0d",
          7987 => x"0d",
          7988 => x"3d",
          7989 => x"95",
          7990 => x"aa",
          7991 => x"f8",
          7992 => x"d4",
          7993 => x"e0",
          7994 => x"64",
          7995 => x"d0",
          7996 => x"ac",
          7997 => x"f8",
          7998 => x"d4",
          7999 => x"38",
          8000 => x"05",
          8001 => x"2b",
          8002 => x"80",
          8003 => x"76",
          8004 => x"0c",
          8005 => x"02",
          8006 => x"70",
          8007 => x"81",
          8008 => x"56",
          8009 => x"9e",
          8010 => x"53",
          8011 => x"ca",
          8012 => x"d4",
          8013 => x"15",
          8014 => x"82",
          8015 => x"84",
          8016 => x"06",
          8017 => x"55",
          8018 => x"f8",
          8019 => x"0d",
          8020 => x"3d",
          8021 => x"3d",
          8022 => x"3d",
          8023 => x"80",
          8024 => x"53",
          8025 => x"fd",
          8026 => x"80",
          8027 => x"e8",
          8028 => x"d4",
          8029 => x"82",
          8030 => x"83",
          8031 => x"80",
          8032 => x"7a",
          8033 => x"08",
          8034 => x"0c",
          8035 => x"d5",
          8036 => x"73",
          8037 => x"83",
          8038 => x"80",
          8039 => x"52",
          8040 => x"3f",
          8041 => x"08",
          8042 => x"f8",
          8043 => x"38",
          8044 => x"08",
          8045 => x"ff",
          8046 => x"82",
          8047 => x"57",
          8048 => x"08",
          8049 => x"80",
          8050 => x"52",
          8051 => x"86",
          8052 => x"f8",
          8053 => x"3d",
          8054 => x"74",
          8055 => x"3f",
          8056 => x"08",
          8057 => x"f8",
          8058 => x"38",
          8059 => x"51",
          8060 => x"82",
          8061 => x"57",
          8062 => x"08",
          8063 => x"da",
          8064 => x"7b",
          8065 => x"3f",
          8066 => x"f8",
          8067 => x"38",
          8068 => x"51",
          8069 => x"82",
          8070 => x"57",
          8071 => x"08",
          8072 => x"38",
          8073 => x"09",
          8074 => x"38",
          8075 => x"ee",
          8076 => x"ea",
          8077 => x"3d",
          8078 => x"52",
          8079 => x"e4",
          8080 => x"3d",
          8081 => x"11",
          8082 => x"5a",
          8083 => x"2e",
          8084 => x"80",
          8085 => x"81",
          8086 => x"70",
          8087 => x"56",
          8088 => x"81",
          8089 => x"78",
          8090 => x"38",
          8091 => x"9c",
          8092 => x"82",
          8093 => x"18",
          8094 => x"08",
          8095 => x"ff",
          8096 => x"55",
          8097 => x"74",
          8098 => x"38",
          8099 => x"e1",
          8100 => x"55",
          8101 => x"34",
          8102 => x"77",
          8103 => x"81",
          8104 => x"ff",
          8105 => x"3d",
          8106 => x"58",
          8107 => x"80",
          8108 => x"d4",
          8109 => x"29",
          8110 => x"05",
          8111 => x"33",
          8112 => x"56",
          8113 => x"2e",
          8114 => x"16",
          8115 => x"33",
          8116 => x"73",
          8117 => x"16",
          8118 => x"26",
          8119 => x"55",
          8120 => x"91",
          8121 => x"54",
          8122 => x"70",
          8123 => x"34",
          8124 => x"ec",
          8125 => x"70",
          8126 => x"34",
          8127 => x"09",
          8128 => x"38",
          8129 => x"39",
          8130 => x"08",
          8131 => x"59",
          8132 => x"7a",
          8133 => x"5c",
          8134 => x"26",
          8135 => x"7a",
          8136 => x"d4",
          8137 => x"df",
          8138 => x"f7",
          8139 => x"7d",
          8140 => x"05",
          8141 => x"57",
          8142 => x"3f",
          8143 => x"08",
          8144 => x"f8",
          8145 => x"38",
          8146 => x"53",
          8147 => x"38",
          8148 => x"54",
          8149 => x"92",
          8150 => x"33",
          8151 => x"70",
          8152 => x"54",
          8153 => x"38",
          8154 => x"15",
          8155 => x"70",
          8156 => x"58",
          8157 => x"82",
          8158 => x"8a",
          8159 => x"89",
          8160 => x"53",
          8161 => x"b7",
          8162 => x"ff",
          8163 => x"c9",
          8164 => x"d4",
          8165 => x"15",
          8166 => x"53",
          8167 => x"c9",
          8168 => x"d4",
          8169 => x"26",
          8170 => x"30",
          8171 => x"70",
          8172 => x"77",
          8173 => x"18",
          8174 => x"51",
          8175 => x"88",
          8176 => x"73",
          8177 => x"52",
          8178 => x"bc",
          8179 => x"d4",
          8180 => x"82",
          8181 => x"81",
          8182 => x"38",
          8183 => x"08",
          8184 => x"9e",
          8185 => x"f8",
          8186 => x"0c",
          8187 => x"0c",
          8188 => x"81",
          8189 => x"76",
          8190 => x"38",
          8191 => x"94",
          8192 => x"94",
          8193 => x"16",
          8194 => x"2a",
          8195 => x"51",
          8196 => x"72",
          8197 => x"38",
          8198 => x"51",
          8199 => x"3f",
          8200 => x"08",
          8201 => x"f8",
          8202 => x"82",
          8203 => x"56",
          8204 => x"52",
          8205 => x"b5",
          8206 => x"d4",
          8207 => x"73",
          8208 => x"38",
          8209 => x"b0",
          8210 => x"73",
          8211 => x"27",
          8212 => x"98",
          8213 => x"9e",
          8214 => x"08",
          8215 => x"0c",
          8216 => x"06",
          8217 => x"2e",
          8218 => x"52",
          8219 => x"b4",
          8220 => x"d4",
          8221 => x"38",
          8222 => x"16",
          8223 => x"80",
          8224 => x"0b",
          8225 => x"81",
          8226 => x"75",
          8227 => x"d4",
          8228 => x"58",
          8229 => x"54",
          8230 => x"74",
          8231 => x"73",
          8232 => x"90",
          8233 => x"c0",
          8234 => x"90",
          8235 => x"83",
          8236 => x"72",
          8237 => x"38",
          8238 => x"08",
          8239 => x"77",
          8240 => x"80",
          8241 => x"d4",
          8242 => x"3d",
          8243 => x"3d",
          8244 => x"89",
          8245 => x"2e",
          8246 => x"80",
          8247 => x"fc",
          8248 => x"3d",
          8249 => x"e1",
          8250 => x"d4",
          8251 => x"82",
          8252 => x"80",
          8253 => x"76",
          8254 => x"75",
          8255 => x"3f",
          8256 => x"08",
          8257 => x"f8",
          8258 => x"38",
          8259 => x"70",
          8260 => x"57",
          8261 => x"a2",
          8262 => x"33",
          8263 => x"70",
          8264 => x"55",
          8265 => x"2e",
          8266 => x"16",
          8267 => x"51",
          8268 => x"82",
          8269 => x"88",
          8270 => x"54",
          8271 => x"84",
          8272 => x"52",
          8273 => x"bd",
          8274 => x"d4",
          8275 => x"74",
          8276 => x"81",
          8277 => x"85",
          8278 => x"74",
          8279 => x"38",
          8280 => x"74",
          8281 => x"d4",
          8282 => x"3d",
          8283 => x"3d",
          8284 => x"3d",
          8285 => x"70",
          8286 => x"bc",
          8287 => x"f8",
          8288 => x"82",
          8289 => x"73",
          8290 => x"0d",
          8291 => x"0d",
          8292 => x"3d",
          8293 => x"71",
          8294 => x"e7",
          8295 => x"d4",
          8296 => x"82",
          8297 => x"80",
          8298 => x"94",
          8299 => x"f8",
          8300 => x"51",
          8301 => x"3f",
          8302 => x"08",
          8303 => x"39",
          8304 => x"08",
          8305 => x"c2",
          8306 => x"d4",
          8307 => x"82",
          8308 => x"84",
          8309 => x"06",
          8310 => x"53",
          8311 => x"d4",
          8312 => x"38",
          8313 => x"51",
          8314 => x"72",
          8315 => x"ff",
          8316 => x"82",
          8317 => x"84",
          8318 => x"70",
          8319 => x"2c",
          8320 => x"f8",
          8321 => x"51",
          8322 => x"82",
          8323 => x"87",
          8324 => x"ed",
          8325 => x"57",
          8326 => x"3d",
          8327 => x"3d",
          8328 => x"e2",
          8329 => x"f8",
          8330 => x"d4",
          8331 => x"38",
          8332 => x"51",
          8333 => x"82",
          8334 => x"55",
          8335 => x"08",
          8336 => x"80",
          8337 => x"70",
          8338 => x"58",
          8339 => x"85",
          8340 => x"8d",
          8341 => x"2e",
          8342 => x"52",
          8343 => x"c4",
          8344 => x"d4",
          8345 => x"3d",
          8346 => x"3d",
          8347 => x"55",
          8348 => x"92",
          8349 => x"52",
          8350 => x"de",
          8351 => x"d4",
          8352 => x"82",
          8353 => x"82",
          8354 => x"74",
          8355 => x"9c",
          8356 => x"11",
          8357 => x"59",
          8358 => x"75",
          8359 => x"38",
          8360 => x"81",
          8361 => x"5b",
          8362 => x"82",
          8363 => x"39",
          8364 => x"08",
          8365 => x"59",
          8366 => x"09",
          8367 => x"c0",
          8368 => x"5f",
          8369 => x"92",
          8370 => x"51",
          8371 => x"3f",
          8372 => x"08",
          8373 => x"38",
          8374 => x"08",
          8375 => x"38",
          8376 => x"08",
          8377 => x"d4",
          8378 => x"80",
          8379 => x"81",
          8380 => x"59",
          8381 => x"14",
          8382 => x"c9",
          8383 => x"39",
          8384 => x"82",
          8385 => x"57",
          8386 => x"38",
          8387 => x"18",
          8388 => x"ff",
          8389 => x"82",
          8390 => x"5b",
          8391 => x"08",
          8392 => x"7c",
          8393 => x"12",
          8394 => x"52",
          8395 => x"82",
          8396 => x"06",
          8397 => x"14",
          8398 => x"d2",
          8399 => x"f8",
          8400 => x"ff",
          8401 => x"70",
          8402 => x"82",
          8403 => x"51",
          8404 => x"b8",
          8405 => x"a9",
          8406 => x"d4",
          8407 => x"0a",
          8408 => x"70",
          8409 => x"84",
          8410 => x"51",
          8411 => x"ff",
          8412 => x"56",
          8413 => x"38",
          8414 => x"7c",
          8415 => x"0c",
          8416 => x"81",
          8417 => x"74",
          8418 => x"7a",
          8419 => x"0c",
          8420 => x"04",
          8421 => x"79",
          8422 => x"05",
          8423 => x"57",
          8424 => x"82",
          8425 => x"56",
          8426 => x"08",
          8427 => x"91",
          8428 => x"75",
          8429 => x"90",
          8430 => x"81",
          8431 => x"06",
          8432 => x"87",
          8433 => x"2e",
          8434 => x"94",
          8435 => x"73",
          8436 => x"27",
          8437 => x"73",
          8438 => x"d4",
          8439 => x"88",
          8440 => x"76",
          8441 => x"d0",
          8442 => x"f8",
          8443 => x"19",
          8444 => x"ca",
          8445 => x"08",
          8446 => x"ff",
          8447 => x"82",
          8448 => x"ff",
          8449 => x"06",
          8450 => x"56",
          8451 => x"08",
          8452 => x"81",
          8453 => x"82",
          8454 => x"75",
          8455 => x"54",
          8456 => x"08",
          8457 => x"27",
          8458 => x"17",
          8459 => x"d4",
          8460 => x"76",
          8461 => x"80",
          8462 => x"f8",
          8463 => x"17",
          8464 => x"0c",
          8465 => x"80",
          8466 => x"73",
          8467 => x"75",
          8468 => x"38",
          8469 => x"34",
          8470 => x"82",
          8471 => x"89",
          8472 => x"e0",
          8473 => x"53",
          8474 => x"9c",
          8475 => x"3d",
          8476 => x"3f",
          8477 => x"08",
          8478 => x"f8",
          8479 => x"38",
          8480 => x"3d",
          8481 => x"3d",
          8482 => x"ce",
          8483 => x"d4",
          8484 => x"82",
          8485 => x"81",
          8486 => x"80",
          8487 => x"70",
          8488 => x"81",
          8489 => x"56",
          8490 => x"81",
          8491 => x"98",
          8492 => x"74",
          8493 => x"38",
          8494 => x"05",
          8495 => x"06",
          8496 => x"55",
          8497 => x"38",
          8498 => x"51",
          8499 => x"3f",
          8500 => x"08",
          8501 => x"70",
          8502 => x"55",
          8503 => x"2e",
          8504 => x"78",
          8505 => x"f8",
          8506 => x"08",
          8507 => x"38",
          8508 => x"d4",
          8509 => x"76",
          8510 => x"70",
          8511 => x"b5",
          8512 => x"d4",
          8513 => x"82",
          8514 => x"80",
          8515 => x"d4",
          8516 => x"73",
          8517 => x"d4",
          8518 => x"f8",
          8519 => x"d4",
          8520 => x"38",
          8521 => x"d0",
          8522 => x"f8",
          8523 => x"88",
          8524 => x"f8",
          8525 => x"38",
          8526 => x"ef",
          8527 => x"f8",
          8528 => x"f8",
          8529 => x"82",
          8530 => x"07",
          8531 => x"55",
          8532 => x"2e",
          8533 => x"80",
          8534 => x"80",
          8535 => x"77",
          8536 => x"d4",
          8537 => x"f8",
          8538 => x"8c",
          8539 => x"ff",
          8540 => x"82",
          8541 => x"55",
          8542 => x"f8",
          8543 => x"0d",
          8544 => x"0d",
          8545 => x"3d",
          8546 => x"52",
          8547 => x"d7",
          8548 => x"d4",
          8549 => x"82",
          8550 => x"82",
          8551 => x"5e",
          8552 => x"3d",
          8553 => x"cb",
          8554 => x"d4",
          8555 => x"82",
          8556 => x"86",
          8557 => x"82",
          8558 => x"d4",
          8559 => x"2e",
          8560 => x"82",
          8561 => x"80",
          8562 => x"70",
          8563 => x"06",
          8564 => x"54",
          8565 => x"38",
          8566 => x"52",
          8567 => x"52",
          8568 => x"80",
          8569 => x"f8",
          8570 => x"56",
          8571 => x"08",
          8572 => x"54",
          8573 => x"08",
          8574 => x"81",
          8575 => x"82",
          8576 => x"f8",
          8577 => x"09",
          8578 => x"38",
          8579 => x"ba",
          8580 => x"b6",
          8581 => x"f8",
          8582 => x"51",
          8583 => x"3f",
          8584 => x"08",
          8585 => x"f8",
          8586 => x"38",
          8587 => x"52",
          8588 => x"ff",
          8589 => x"78",
          8590 => x"b8",
          8591 => x"54",
          8592 => x"c3",
          8593 => x"88",
          8594 => x"80",
          8595 => x"ff",
          8596 => x"75",
          8597 => x"11",
          8598 => x"b8",
          8599 => x"53",
          8600 => x"53",
          8601 => x"51",
          8602 => x"3f",
          8603 => x"0b",
          8604 => x"34",
          8605 => x"80",
          8606 => x"51",
          8607 => x"3f",
          8608 => x"0b",
          8609 => x"77",
          8610 => x"cd",
          8611 => x"f8",
          8612 => x"d4",
          8613 => x"38",
          8614 => x"0a",
          8615 => x"05",
          8616 => x"ca",
          8617 => x"64",
          8618 => x"ff",
          8619 => x"64",
          8620 => x"8b",
          8621 => x"54",
          8622 => x"15",
          8623 => x"ff",
          8624 => x"82",
          8625 => x"54",
          8626 => x"53",
          8627 => x"51",
          8628 => x"3f",
          8629 => x"f8",
          8630 => x"0d",
          8631 => x"0d",
          8632 => x"05",
          8633 => x"3f",
          8634 => x"3d",
          8635 => x"52",
          8636 => x"d5",
          8637 => x"d4",
          8638 => x"82",
          8639 => x"82",
          8640 => x"4e",
          8641 => x"52",
          8642 => x"52",
          8643 => x"3f",
          8644 => x"08",
          8645 => x"f8",
          8646 => x"38",
          8647 => x"05",
          8648 => x"06",
          8649 => x"73",
          8650 => x"a0",
          8651 => x"08",
          8652 => x"ff",
          8653 => x"ff",
          8654 => x"b0",
          8655 => x"92",
          8656 => x"54",
          8657 => x"3f",
          8658 => x"52",
          8659 => x"d0",
          8660 => x"f8",
          8661 => x"d4",
          8662 => x"38",
          8663 => x"08",
          8664 => x"06",
          8665 => x"a3",
          8666 => x"92",
          8667 => x"81",
          8668 => x"d4",
          8669 => x"2e",
          8670 => x"81",
          8671 => x"51",
          8672 => x"3f",
          8673 => x"08",
          8674 => x"f8",
          8675 => x"38",
          8676 => x"53",
          8677 => x"8d",
          8678 => x"16",
          8679 => x"fd",
          8680 => x"05",
          8681 => x"34",
          8682 => x"70",
          8683 => x"81",
          8684 => x"55",
          8685 => x"74",
          8686 => x"73",
          8687 => x"78",
          8688 => x"83",
          8689 => x"16",
          8690 => x"2a",
          8691 => x"51",
          8692 => x"80",
          8693 => x"38",
          8694 => x"80",
          8695 => x"52",
          8696 => x"b4",
          8697 => x"d4",
          8698 => x"78",
          8699 => x"ee",
          8700 => x"82",
          8701 => x"80",
          8702 => x"38",
          8703 => x"08",
          8704 => x"ff",
          8705 => x"82",
          8706 => x"79",
          8707 => x"58",
          8708 => x"d4",
          8709 => x"c1",
          8710 => x"33",
          8711 => x"2e",
          8712 => x"9a",
          8713 => x"75",
          8714 => x"ff",
          8715 => x"78",
          8716 => x"83",
          8717 => x"39",
          8718 => x"08",
          8719 => x"51",
          8720 => x"82",
          8721 => x"55",
          8722 => x"08",
          8723 => x"51",
          8724 => x"3f",
          8725 => x"08",
          8726 => x"d4",
          8727 => x"3d",
          8728 => x"3d",
          8729 => x"df",
          8730 => x"84",
          8731 => x"05",
          8732 => x"82",
          8733 => x"cc",
          8734 => x"3d",
          8735 => x"3f",
          8736 => x"08",
          8737 => x"f8",
          8738 => x"38",
          8739 => x"52",
          8740 => x"05",
          8741 => x"3f",
          8742 => x"08",
          8743 => x"f8",
          8744 => x"02",
          8745 => x"33",
          8746 => x"54",
          8747 => x"aa",
          8748 => x"06",
          8749 => x"8b",
          8750 => x"06",
          8751 => x"07",
          8752 => x"56",
          8753 => x"34",
          8754 => x"0b",
          8755 => x"78",
          8756 => x"db",
          8757 => x"f8",
          8758 => x"82",
          8759 => x"96",
          8760 => x"ee",
          8761 => x"56",
          8762 => x"3d",
          8763 => x"95",
          8764 => x"92",
          8765 => x"f8",
          8766 => x"d4",
          8767 => x"cb",
          8768 => x"64",
          8769 => x"d0",
          8770 => x"94",
          8771 => x"f8",
          8772 => x"d4",
          8773 => x"38",
          8774 => x"05",
          8775 => x"06",
          8776 => x"73",
          8777 => x"16",
          8778 => x"22",
          8779 => x"07",
          8780 => x"1f",
          8781 => x"b6",
          8782 => x"81",
          8783 => x"34",
          8784 => x"a1",
          8785 => x"d4",
          8786 => x"74",
          8787 => x"0c",
          8788 => x"04",
          8789 => x"6a",
          8790 => x"80",
          8791 => x"cc",
          8792 => x"3d",
          8793 => x"3f",
          8794 => x"08",
          8795 => x"08",
          8796 => x"d4",
          8797 => x"80",
          8798 => x"57",
          8799 => x"81",
          8800 => x"70",
          8801 => x"55",
          8802 => x"80",
          8803 => x"5d",
          8804 => x"52",
          8805 => x"52",
          8806 => x"db",
          8807 => x"f8",
          8808 => x"d4",
          8809 => x"d2",
          8810 => x"73",
          8811 => x"bc",
          8812 => x"f8",
          8813 => x"d4",
          8814 => x"38",
          8815 => x"08",
          8816 => x"08",
          8817 => x"56",
          8818 => x"19",
          8819 => x"59",
          8820 => x"74",
          8821 => x"56",
          8822 => x"ec",
          8823 => x"75",
          8824 => x"74",
          8825 => x"2e",
          8826 => x"16",
          8827 => x"33",
          8828 => x"73",
          8829 => x"38",
          8830 => x"84",
          8831 => x"06",
          8832 => x"7a",
          8833 => x"76",
          8834 => x"07",
          8835 => x"54",
          8836 => x"80",
          8837 => x"80",
          8838 => x"7b",
          8839 => x"53",
          8840 => x"c4",
          8841 => x"f8",
          8842 => x"d4",
          8843 => x"38",
          8844 => x"55",
          8845 => x"56",
          8846 => x"8b",
          8847 => x"56",
          8848 => x"83",
          8849 => x"75",
          8850 => x"51",
          8851 => x"3f",
          8852 => x"08",
          8853 => x"82",
          8854 => x"99",
          8855 => x"e6",
          8856 => x"53",
          8857 => x"b4",
          8858 => x"3d",
          8859 => x"3f",
          8860 => x"08",
          8861 => x"08",
          8862 => x"d4",
          8863 => x"dd",
          8864 => x"a0",
          8865 => x"70",
          8866 => x"9c",
          8867 => x"6d",
          8868 => x"55",
          8869 => x"27",
          8870 => x"77",
          8871 => x"51",
          8872 => x"3f",
          8873 => x"08",
          8874 => x"26",
          8875 => x"82",
          8876 => x"51",
          8877 => x"83",
          8878 => x"d4",
          8879 => x"93",
          8880 => x"d4",
          8881 => x"ff",
          8882 => x"74",
          8883 => x"38",
          8884 => x"c8",
          8885 => x"9c",
          8886 => x"d4",
          8887 => x"38",
          8888 => x"27",
          8889 => x"89",
          8890 => x"8b",
          8891 => x"27",
          8892 => x"55",
          8893 => x"81",
          8894 => x"8f",
          8895 => x"2a",
          8896 => x"70",
          8897 => x"34",
          8898 => x"74",
          8899 => x"05",
          8900 => x"16",
          8901 => x"51",
          8902 => x"9f",
          8903 => x"38",
          8904 => x"54",
          8905 => x"81",
          8906 => x"b1",
          8907 => x"2e",
          8908 => x"a3",
          8909 => x"15",
          8910 => x"54",
          8911 => x"09",
          8912 => x"38",
          8913 => x"75",
          8914 => x"40",
          8915 => x"52",
          8916 => x"52",
          8917 => x"9f",
          8918 => x"f8",
          8919 => x"d4",
          8920 => x"f7",
          8921 => x"74",
          8922 => x"80",
          8923 => x"f8",
          8924 => x"d4",
          8925 => x"38",
          8926 => x"38",
          8927 => x"74",
          8928 => x"39",
          8929 => x"08",
          8930 => x"81",
          8931 => x"38",
          8932 => x"74",
          8933 => x"38",
          8934 => x"51",
          8935 => x"3f",
          8936 => x"08",
          8937 => x"f8",
          8938 => x"a0",
          8939 => x"f8",
          8940 => x"51",
          8941 => x"3f",
          8942 => x"0b",
          8943 => x"8b",
          8944 => x"66",
          8945 => x"d5",
          8946 => x"81",
          8947 => x"34",
          8948 => x"9c",
          8949 => x"d4",
          8950 => x"73",
          8951 => x"d4",
          8952 => x"3d",
          8953 => x"3d",
          8954 => x"02",
          8955 => x"cb",
          8956 => x"3d",
          8957 => x"72",
          8958 => x"5a",
          8959 => x"82",
          8960 => x"58",
          8961 => x"08",
          8962 => x"91",
          8963 => x"77",
          8964 => x"7c",
          8965 => x"38",
          8966 => x"59",
          8967 => x"90",
          8968 => x"81",
          8969 => x"06",
          8970 => x"73",
          8971 => x"54",
          8972 => x"82",
          8973 => x"39",
          8974 => x"8b",
          8975 => x"11",
          8976 => x"2b",
          8977 => x"54",
          8978 => x"fe",
          8979 => x"ff",
          8980 => x"70",
          8981 => x"07",
          8982 => x"d4",
          8983 => x"90",
          8984 => x"40",
          8985 => x"55",
          8986 => x"88",
          8987 => x"08",
          8988 => x"38",
          8989 => x"77",
          8990 => x"56",
          8991 => x"51",
          8992 => x"3f",
          8993 => x"55",
          8994 => x"08",
          8995 => x"38",
          8996 => x"d4",
          8997 => x"2e",
          8998 => x"82",
          8999 => x"ff",
          9000 => x"38",
          9001 => x"08",
          9002 => x"16",
          9003 => x"2e",
          9004 => x"87",
          9005 => x"74",
          9006 => x"74",
          9007 => x"81",
          9008 => x"38",
          9009 => x"ff",
          9010 => x"2e",
          9011 => x"7b",
          9012 => x"80",
          9013 => x"81",
          9014 => x"81",
          9015 => x"06",
          9016 => x"56",
          9017 => x"52",
          9018 => x"9e",
          9019 => x"d4",
          9020 => x"82",
          9021 => x"80",
          9022 => x"81",
          9023 => x"56",
          9024 => x"d3",
          9025 => x"ff",
          9026 => x"7c",
          9027 => x"55",
          9028 => x"b3",
          9029 => x"1b",
          9030 => x"1b",
          9031 => x"33",
          9032 => x"54",
          9033 => x"34",
          9034 => x"fe",
          9035 => x"08",
          9036 => x"74",
          9037 => x"75",
          9038 => x"16",
          9039 => x"33",
          9040 => x"73",
          9041 => x"77",
          9042 => x"d4",
          9043 => x"3d",
          9044 => x"3d",
          9045 => x"02",
          9046 => x"eb",
          9047 => x"3d",
          9048 => x"59",
          9049 => x"8b",
          9050 => x"82",
          9051 => x"24",
          9052 => x"82",
          9053 => x"84",
          9054 => x"c0",
          9055 => x"51",
          9056 => x"2e",
          9057 => x"75",
          9058 => x"f8",
          9059 => x"06",
          9060 => x"7e",
          9061 => x"fe",
          9062 => x"f8",
          9063 => x"06",
          9064 => x"56",
          9065 => x"74",
          9066 => x"76",
          9067 => x"81",
          9068 => x"8a",
          9069 => x"b2",
          9070 => x"fc",
          9071 => x"52",
          9072 => x"93",
          9073 => x"d4",
          9074 => x"38",
          9075 => x"80",
          9076 => x"74",
          9077 => x"26",
          9078 => x"15",
          9079 => x"74",
          9080 => x"38",
          9081 => x"80",
          9082 => x"84",
          9083 => x"92",
          9084 => x"80",
          9085 => x"38",
          9086 => x"06",
          9087 => x"2e",
          9088 => x"56",
          9089 => x"78",
          9090 => x"89",
          9091 => x"2b",
          9092 => x"43",
          9093 => x"38",
          9094 => x"30",
          9095 => x"77",
          9096 => x"91",
          9097 => x"c2",
          9098 => x"f8",
          9099 => x"52",
          9100 => x"92",
          9101 => x"56",
          9102 => x"08",
          9103 => x"77",
          9104 => x"77",
          9105 => x"f8",
          9106 => x"45",
          9107 => x"bf",
          9108 => x"8e",
          9109 => x"26",
          9110 => x"74",
          9111 => x"48",
          9112 => x"75",
          9113 => x"38",
          9114 => x"81",
          9115 => x"fa",
          9116 => x"2a",
          9117 => x"56",
          9118 => x"2e",
          9119 => x"87",
          9120 => x"82",
          9121 => x"38",
          9122 => x"55",
          9123 => x"83",
          9124 => x"81",
          9125 => x"56",
          9126 => x"80",
          9127 => x"38",
          9128 => x"83",
          9129 => x"06",
          9130 => x"78",
          9131 => x"91",
          9132 => x"0b",
          9133 => x"22",
          9134 => x"80",
          9135 => x"74",
          9136 => x"38",
          9137 => x"56",
          9138 => x"17",
          9139 => x"57",
          9140 => x"2e",
          9141 => x"75",
          9142 => x"79",
          9143 => x"fe",
          9144 => x"82",
          9145 => x"84",
          9146 => x"05",
          9147 => x"5e",
          9148 => x"80",
          9149 => x"f8",
          9150 => x"8a",
          9151 => x"fd",
          9152 => x"75",
          9153 => x"38",
          9154 => x"78",
          9155 => x"8c",
          9156 => x"0b",
          9157 => x"22",
          9158 => x"80",
          9159 => x"74",
          9160 => x"38",
          9161 => x"56",
          9162 => x"17",
          9163 => x"57",
          9164 => x"2e",
          9165 => x"75",
          9166 => x"79",
          9167 => x"fe",
          9168 => x"82",
          9169 => x"10",
          9170 => x"82",
          9171 => x"9f",
          9172 => x"38",
          9173 => x"d4",
          9174 => x"82",
          9175 => x"05",
          9176 => x"2a",
          9177 => x"56",
          9178 => x"17",
          9179 => x"81",
          9180 => x"60",
          9181 => x"65",
          9182 => x"12",
          9183 => x"30",
          9184 => x"74",
          9185 => x"59",
          9186 => x"7d",
          9187 => x"81",
          9188 => x"76",
          9189 => x"41",
          9190 => x"76",
          9191 => x"90",
          9192 => x"62",
          9193 => x"51",
          9194 => x"26",
          9195 => x"75",
          9196 => x"31",
          9197 => x"65",
          9198 => x"fe",
          9199 => x"82",
          9200 => x"58",
          9201 => x"09",
          9202 => x"38",
          9203 => x"08",
          9204 => x"26",
          9205 => x"78",
          9206 => x"79",
          9207 => x"78",
          9208 => x"86",
          9209 => x"82",
          9210 => x"06",
          9211 => x"83",
          9212 => x"82",
          9213 => x"27",
          9214 => x"8f",
          9215 => x"55",
          9216 => x"26",
          9217 => x"59",
          9218 => x"62",
          9219 => x"74",
          9220 => x"38",
          9221 => x"88",
          9222 => x"f8",
          9223 => x"26",
          9224 => x"86",
          9225 => x"1a",
          9226 => x"79",
          9227 => x"38",
          9228 => x"80",
          9229 => x"2e",
          9230 => x"83",
          9231 => x"9f",
          9232 => x"8b",
          9233 => x"06",
          9234 => x"74",
          9235 => x"84",
          9236 => x"52",
          9237 => x"90",
          9238 => x"53",
          9239 => x"52",
          9240 => x"90",
          9241 => x"80",
          9242 => x"51",
          9243 => x"3f",
          9244 => x"34",
          9245 => x"ff",
          9246 => x"1b",
          9247 => x"d0",
          9248 => x"90",
          9249 => x"83",
          9250 => x"70",
          9251 => x"80",
          9252 => x"55",
          9253 => x"ff",
          9254 => x"66",
          9255 => x"ff",
          9256 => x"38",
          9257 => x"ff",
          9258 => x"1b",
          9259 => x"a0",
          9260 => x"74",
          9261 => x"51",
          9262 => x"3f",
          9263 => x"1c",
          9264 => x"98",
          9265 => x"8f",
          9266 => x"ff",
          9267 => x"51",
          9268 => x"3f",
          9269 => x"1b",
          9270 => x"92",
          9271 => x"2e",
          9272 => x"80",
          9273 => x"88",
          9274 => x"80",
          9275 => x"ff",
          9276 => x"7c",
          9277 => x"51",
          9278 => x"3f",
          9279 => x"1b",
          9280 => x"ea",
          9281 => x"b0",
          9282 => x"8e",
          9283 => x"52",
          9284 => x"ff",
          9285 => x"ff",
          9286 => x"c0",
          9287 => x"0b",
          9288 => x"34",
          9289 => x"c6",
          9290 => x"c7",
          9291 => x"39",
          9292 => x"0a",
          9293 => x"51",
          9294 => x"3f",
          9295 => x"ff",
          9296 => x"1b",
          9297 => x"88",
          9298 => x"0b",
          9299 => x"a9",
          9300 => x"34",
          9301 => x"c6",
          9302 => x"1b",
          9303 => x"bd",
          9304 => x"d5",
          9305 => x"1b",
          9306 => x"ff",
          9307 => x"81",
          9308 => x"7a",
          9309 => x"ff",
          9310 => x"81",
          9311 => x"f8",
          9312 => x"38",
          9313 => x"09",
          9314 => x"ee",
          9315 => x"60",
          9316 => x"7a",
          9317 => x"ff",
          9318 => x"84",
          9319 => x"52",
          9320 => x"8e",
          9321 => x"8b",
          9322 => x"52",
          9323 => x"8d",
          9324 => x"8a",
          9325 => x"52",
          9326 => x"51",
          9327 => x"3f",
          9328 => x"83",
          9329 => x"ff",
          9330 => x"82",
          9331 => x"1b",
          9332 => x"9a",
          9333 => x"d5",
          9334 => x"ff",
          9335 => x"75",
          9336 => x"05",
          9337 => x"7e",
          9338 => x"93",
          9339 => x"60",
          9340 => x"52",
          9341 => x"89",
          9342 => x"53",
          9343 => x"51",
          9344 => x"3f",
          9345 => x"58",
          9346 => x"09",
          9347 => x"38",
          9348 => x"51",
          9349 => x"3f",
          9350 => x"1b",
          9351 => x"ce",
          9352 => x"52",
          9353 => x"91",
          9354 => x"ff",
          9355 => x"81",
          9356 => x"f8",
          9357 => x"7a",
          9358 => x"b2",
          9359 => x"61",
          9360 => x"26",
          9361 => x"57",
          9362 => x"53",
          9363 => x"51",
          9364 => x"3f",
          9365 => x"08",
          9366 => x"84",
          9367 => x"d4",
          9368 => x"7a",
          9369 => x"d8",
          9370 => x"75",
          9371 => x"56",
          9372 => x"81",
          9373 => x"80",
          9374 => x"38",
          9375 => x"83",
          9376 => x"63",
          9377 => x"74",
          9378 => x"38",
          9379 => x"54",
          9380 => x"52",
          9381 => x"87",
          9382 => x"d4",
          9383 => x"c1",
          9384 => x"75",
          9385 => x"56",
          9386 => x"8c",
          9387 => x"2e",
          9388 => x"56",
          9389 => x"ff",
          9390 => x"84",
          9391 => x"2e",
          9392 => x"56",
          9393 => x"58",
          9394 => x"38",
          9395 => x"77",
          9396 => x"ff",
          9397 => x"82",
          9398 => x"78",
          9399 => x"f0",
          9400 => x"1b",
          9401 => x"34",
          9402 => x"16",
          9403 => x"82",
          9404 => x"83",
          9405 => x"84",
          9406 => x"67",
          9407 => x"fd",
          9408 => x"51",
          9409 => x"3f",
          9410 => x"16",
          9411 => x"f8",
          9412 => x"bf",
          9413 => x"86",
          9414 => x"d4",
          9415 => x"16",
          9416 => x"83",
          9417 => x"ff",
          9418 => x"66",
          9419 => x"1b",
          9420 => x"ba",
          9421 => x"77",
          9422 => x"7e",
          9423 => x"bf",
          9424 => x"82",
          9425 => x"a2",
          9426 => x"80",
          9427 => x"ff",
          9428 => x"81",
          9429 => x"f8",
          9430 => x"89",
          9431 => x"8a",
          9432 => x"86",
          9433 => x"f8",
          9434 => x"82",
          9435 => x"99",
          9436 => x"f5",
          9437 => x"60",
          9438 => x"79",
          9439 => x"5a",
          9440 => x"78",
          9441 => x"8d",
          9442 => x"55",
          9443 => x"fc",
          9444 => x"51",
          9445 => x"7a",
          9446 => x"81",
          9447 => x"8c",
          9448 => x"74",
          9449 => x"38",
          9450 => x"81",
          9451 => x"81",
          9452 => x"8a",
          9453 => x"06",
          9454 => x"76",
          9455 => x"76",
          9456 => x"55",
          9457 => x"f8",
          9458 => x"0d",
          9459 => x"0d",
          9460 => x"05",
          9461 => x"59",
          9462 => x"2e",
          9463 => x"87",
          9464 => x"76",
          9465 => x"84",
          9466 => x"80",
          9467 => x"38",
          9468 => x"77",
          9469 => x"56",
          9470 => x"34",
          9471 => x"bb",
          9472 => x"38",
          9473 => x"05",
          9474 => x"8c",
          9475 => x"08",
          9476 => x"3f",
          9477 => x"70",
          9478 => x"07",
          9479 => x"30",
          9480 => x"56",
          9481 => x"0c",
          9482 => x"18",
          9483 => x"0d",
          9484 => x"0d",
          9485 => x"08",
          9486 => x"75",
          9487 => x"89",
          9488 => x"54",
          9489 => x"16",
          9490 => x"51",
          9491 => x"82",
          9492 => x"91",
          9493 => x"08",
          9494 => x"81",
          9495 => x"88",
          9496 => x"83",
          9497 => x"74",
          9498 => x"0c",
          9499 => x"04",
          9500 => x"75",
          9501 => x"53",
          9502 => x"51",
          9503 => x"3f",
          9504 => x"85",
          9505 => x"ea",
          9506 => x"80",
          9507 => x"6a",
          9508 => x"70",
          9509 => x"d8",
          9510 => x"72",
          9511 => x"3f",
          9512 => x"8d",
          9513 => x"0d",
          9514 => x"0d",
          9515 => x"05",
          9516 => x"55",
          9517 => x"72",
          9518 => x"8a",
          9519 => x"ff",
          9520 => x"80",
          9521 => x"ff",
          9522 => x"51",
          9523 => x"2e",
          9524 => x"b4",
          9525 => x"2e",
          9526 => x"c8",
          9527 => x"72",
          9528 => x"38",
          9529 => x"83",
          9530 => x"53",
          9531 => x"ff",
          9532 => x"71",
          9533 => x"c4",
          9534 => x"51",
          9535 => x"81",
          9536 => x"81",
          9537 => x"51",
          9538 => x"f8",
          9539 => x"0d",
          9540 => x"0d",
          9541 => x"22",
          9542 => x"96",
          9543 => x"51",
          9544 => x"80",
          9545 => x"38",
          9546 => x"39",
          9547 => x"2e",
          9548 => x"91",
          9549 => x"ff",
          9550 => x"70",
          9551 => x"c4",
          9552 => x"54",
          9553 => x"d4",
          9554 => x"3d",
          9555 => x"3d",
          9556 => x"70",
          9557 => x"26",
          9558 => x"70",
          9559 => x"06",
          9560 => x"57",
          9561 => x"72",
          9562 => x"82",
          9563 => x"75",
          9564 => x"57",
          9565 => x"70",
          9566 => x"75",
          9567 => x"52",
          9568 => x"fb",
          9569 => x"82",
          9570 => x"70",
          9571 => x"81",
          9572 => x"18",
          9573 => x"53",
          9574 => x"80",
          9575 => x"88",
          9576 => x"38",
          9577 => x"82",
          9578 => x"51",
          9579 => x"71",
          9580 => x"76",
          9581 => x"54",
          9582 => x"c3",
          9583 => x"31",
          9584 => x"71",
          9585 => x"a4",
          9586 => x"51",
          9587 => x"12",
          9588 => x"d0",
          9589 => x"39",
          9590 => x"90",
          9591 => x"51",
          9592 => x"b0",
          9593 => x"39",
          9594 => x"51",
          9595 => x"ff",
          9596 => x"39",
          9597 => x"38",
          9598 => x"56",
          9599 => x"71",
          9600 => x"d4",
          9601 => x"3d",
          9602 => x"00",
          9603 => x"ff",
          9604 => x"ff",
          9605 => x"ff",
          9606 => x"00",
          9607 => x"00",
          9608 => x"00",
          9609 => x"00",
          9610 => x"00",
          9611 => x"00",
          9612 => x"00",
          9613 => x"00",
          9614 => x"00",
          9615 => x"00",
          9616 => x"00",
          9617 => x"00",
          9618 => x"00",
          9619 => x"00",
          9620 => x"00",
          9621 => x"00",
          9622 => x"00",
          9623 => x"00",
          9624 => x"00",
          9625 => x"00",
          9626 => x"00",
          9627 => x"00",
          9628 => x"00",
          9629 => x"00",
          9630 => x"00",
          9631 => x"00",
          9632 => x"00",
          9633 => x"00",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"00",
          9638 => x"00",
          9639 => x"00",
          9640 => x"00",
          9641 => x"00",
          9642 => x"00",
          9643 => x"00",
          9644 => x"00",
          9645 => x"00",
          9646 => x"00",
          9647 => x"00",
          9648 => x"00",
          9649 => x"00",
          9650 => x"00",
          9651 => x"00",
          9652 => x"00",
          9653 => x"00",
          9654 => x"00",
          9655 => x"00",
          9656 => x"00",
          9657 => x"00",
          9658 => x"00",
          9659 => x"00",
          9660 => x"00",
          9661 => x"00",
          9662 => x"00",
          9663 => x"00",
          9664 => x"00",
          9665 => x"00",
          9666 => x"00",
          9667 => x"00",
          9668 => x"00",
          9669 => x"00",
          9670 => x"00",
          9671 => x"00",
          9672 => x"00",
          9673 => x"00",
          9674 => x"00",
          9675 => x"00",
          9676 => x"00",
          9677 => x"00",
          9678 => x"00",
          9679 => x"00",
          9680 => x"00",
          9681 => x"00",
          9682 => x"00",
          9683 => x"00",
          9684 => x"00",
          9685 => x"00",
          9686 => x"00",
          9687 => x"00",
          9688 => x"00",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"00",
          9693 => x"00",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"00",
          9721 => x"00",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"00",
          9726 => x"00",
          9727 => x"00",
          9728 => x"00",
          9729 => x"00",
          9730 => x"00",
          9731 => x"00",
          9732 => x"00",
          9733 => x"00",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"64",
          9752 => x"74",
          9753 => x"64",
          9754 => x"74",
          9755 => x"66",
          9756 => x"74",
          9757 => x"66",
          9758 => x"64",
          9759 => x"66",
          9760 => x"63",
          9761 => x"6d",
          9762 => x"61",
          9763 => x"6d",
          9764 => x"79",
          9765 => x"6d",
          9766 => x"66",
          9767 => x"6d",
          9768 => x"70",
          9769 => x"6d",
          9770 => x"6d",
          9771 => x"6d",
          9772 => x"68",
          9773 => x"68",
          9774 => x"68",
          9775 => x"68",
          9776 => x"63",
          9777 => x"00",
          9778 => x"6a",
          9779 => x"72",
          9780 => x"61",
          9781 => x"72",
          9782 => x"74",
          9783 => x"69",
          9784 => x"00",
          9785 => x"74",
          9786 => x"00",
          9787 => x"74",
          9788 => x"69",
          9789 => x"6d",
          9790 => x"69",
          9791 => x"6b",
          9792 => x"00",
          9793 => x"65",
          9794 => x"44",
          9795 => x"20",
          9796 => x"6f",
          9797 => x"49",
          9798 => x"72",
          9799 => x"20",
          9800 => x"6f",
          9801 => x"44",
          9802 => x"20",
          9803 => x"20",
          9804 => x"64",
          9805 => x"4e",
          9806 => x"69",
          9807 => x"66",
          9808 => x"64",
          9809 => x"4e",
          9810 => x"61",
          9811 => x"66",
          9812 => x"64",
          9813 => x"49",
          9814 => x"6c",
          9815 => x"66",
          9816 => x"6e",
          9817 => x"2e",
          9818 => x"41",
          9819 => x"73",
          9820 => x"65",
          9821 => x"64",
          9822 => x"46",
          9823 => x"20",
          9824 => x"65",
          9825 => x"20",
          9826 => x"73",
          9827 => x"00",
          9828 => x"46",
          9829 => x"20",
          9830 => x"64",
          9831 => x"69",
          9832 => x"6c",
          9833 => x"00",
          9834 => x"53",
          9835 => x"73",
          9836 => x"69",
          9837 => x"70",
          9838 => x"65",
          9839 => x"64",
          9840 => x"44",
          9841 => x"65",
          9842 => x"6d",
          9843 => x"20",
          9844 => x"69",
          9845 => x"6c",
          9846 => x"00",
          9847 => x"44",
          9848 => x"20",
          9849 => x"20",
          9850 => x"62",
          9851 => x"2e",
          9852 => x"4e",
          9853 => x"6f",
          9854 => x"74",
          9855 => x"65",
          9856 => x"6c",
          9857 => x"73",
          9858 => x"20",
          9859 => x"6e",
          9860 => x"6e",
          9861 => x"73",
          9862 => x"46",
          9863 => x"61",
          9864 => x"62",
          9865 => x"65",
          9866 => x"54",
          9867 => x"6f",
          9868 => x"20",
          9869 => x"72",
          9870 => x"6f",
          9871 => x"61",
          9872 => x"6c",
          9873 => x"2e",
          9874 => x"46",
          9875 => x"20",
          9876 => x"6c",
          9877 => x"65",
          9878 => x"49",
          9879 => x"66",
          9880 => x"69",
          9881 => x"20",
          9882 => x"6f",
          9883 => x"00",
          9884 => x"54",
          9885 => x"6d",
          9886 => x"20",
          9887 => x"6e",
          9888 => x"6c",
          9889 => x"00",
          9890 => x"50",
          9891 => x"6d",
          9892 => x"72",
          9893 => x"6e",
          9894 => x"72",
          9895 => x"2e",
          9896 => x"53",
          9897 => x"65",
          9898 => x"00",
          9899 => x"55",
          9900 => x"6f",
          9901 => x"65",
          9902 => x"72",
          9903 => x"0a",
          9904 => x"20",
          9905 => x"65",
          9906 => x"73",
          9907 => x"20",
          9908 => x"20",
          9909 => x"65",
          9910 => x"65",
          9911 => x"00",
          9912 => x"72",
          9913 => x"00",
          9914 => x"30",
          9915 => x"38",
          9916 => x"20",
          9917 => x"30",
          9918 => x"2c",
          9919 => x"25",
          9920 => x"78",
          9921 => x"49",
          9922 => x"25",
          9923 => x"78",
          9924 => x"38",
          9925 => x"25",
          9926 => x"78",
          9927 => x"25",
          9928 => x"58",
          9929 => x"3a",
          9930 => x"25",
          9931 => x"00",
          9932 => x"20",
          9933 => x"20",
          9934 => x"00",
          9935 => x"25",
          9936 => x"00",
          9937 => x"20",
          9938 => x"20",
          9939 => x"7c",
          9940 => x"7a",
          9941 => x"0a",
          9942 => x"25",
          9943 => x"00",
          9944 => x"30",
          9945 => x"32",
          9946 => x"32",
          9947 => x"76",
          9948 => x"34",
          9949 => x"20",
          9950 => x"2c",
          9951 => x"76",
          9952 => x"32",
          9953 => x"25",
          9954 => x"73",
          9955 => x"0a",
          9956 => x"5a",
          9957 => x"49",
          9958 => x"72",
          9959 => x"74",
          9960 => x"6e",
          9961 => x"72",
          9962 => x"54",
          9963 => x"72",
          9964 => x"74",
          9965 => x"75",
          9966 => x"50",
          9967 => x"69",
          9968 => x"72",
          9969 => x"74",
          9970 => x"49",
          9971 => x"4c",
          9972 => x"20",
          9973 => x"65",
          9974 => x"70",
          9975 => x"49",
          9976 => x"4c",
          9977 => x"20",
          9978 => x"65",
          9979 => x"70",
          9980 => x"55",
          9981 => x"30",
          9982 => x"20",
          9983 => x"65",
          9984 => x"70",
          9985 => x"55",
          9986 => x"30",
          9987 => x"20",
          9988 => x"65",
          9989 => x"70",
          9990 => x"55",
          9991 => x"31",
          9992 => x"20",
          9993 => x"65",
          9994 => x"70",
          9995 => x"55",
          9996 => x"31",
          9997 => x"20",
          9998 => x"65",
          9999 => x"70",
         10000 => x"53",
         10001 => x"69",
         10002 => x"75",
         10003 => x"69",
         10004 => x"2e",
         10005 => x"45",
         10006 => x"6c",
         10007 => x"20",
         10008 => x"65",
         10009 => x"2e",
         10010 => x"61",
         10011 => x"65",
         10012 => x"2e",
         10013 => x"00",
         10014 => x"7a",
         10015 => x"68",
         10016 => x"30",
         10017 => x"46",
         10018 => x"65",
         10019 => x"6f",
         10020 => x"69",
         10021 => x"6c",
         10022 => x"20",
         10023 => x"63",
         10024 => x"20",
         10025 => x"70",
         10026 => x"73",
         10027 => x"6e",
         10028 => x"6d",
         10029 => x"61",
         10030 => x"2e",
         10031 => x"2a",
         10032 => x"43",
         10033 => x"72",
         10034 => x"2e",
         10035 => x"00",
         10036 => x"43",
         10037 => x"69",
         10038 => x"2e",
         10039 => x"43",
         10040 => x"61",
         10041 => x"67",
         10042 => x"00",
         10043 => x"25",
         10044 => x"78",
         10045 => x"38",
         10046 => x"3e",
         10047 => x"6c",
         10048 => x"30",
         10049 => x"0a",
         10050 => x"44",
         10051 => x"20",
         10052 => x"6f",
         10053 => x"0a",
         10054 => x"70",
         10055 => x"65",
         10056 => x"25",
         10057 => x"58",
         10058 => x"32",
         10059 => x"3f",
         10060 => x"25",
         10061 => x"58",
         10062 => x"34",
         10063 => x"25",
         10064 => x"58",
         10065 => x"38",
         10066 => x"00",
         10067 => x"45",
         10068 => x"75",
         10069 => x"67",
         10070 => x"64",
         10071 => x"20",
         10072 => x"6c",
         10073 => x"2e",
         10074 => x"43",
         10075 => x"69",
         10076 => x"63",
         10077 => x"20",
         10078 => x"30",
         10079 => x"20",
         10080 => x"0a",
         10081 => x"43",
         10082 => x"20",
         10083 => x"75",
         10084 => x"64",
         10085 => x"64",
         10086 => x"25",
         10087 => x"0a",
         10088 => x"52",
         10089 => x"61",
         10090 => x"6e",
         10091 => x"70",
         10092 => x"63",
         10093 => x"6f",
         10094 => x"2e",
         10095 => x"43",
         10096 => x"20",
         10097 => x"6f",
         10098 => x"6e",
         10099 => x"2e",
         10100 => x"5a",
         10101 => x"62",
         10102 => x"25",
         10103 => x"25",
         10104 => x"73",
         10105 => x"00",
         10106 => x"25",
         10107 => x"25",
         10108 => x"73",
         10109 => x"25",
         10110 => x"25",
         10111 => x"42",
         10112 => x"63",
         10113 => x"61",
         10114 => x"00",
         10115 => x"4d",
         10116 => x"72",
         10117 => x"78",
         10118 => x"73",
         10119 => x"2c",
         10120 => x"6e",
         10121 => x"20",
         10122 => x"63",
         10123 => x"20",
         10124 => x"6d",
         10125 => x"2e",
         10126 => x"52",
         10127 => x"69",
         10128 => x"2e",
         10129 => x"45",
         10130 => x"6c",
         10131 => x"20",
         10132 => x"65",
         10133 => x"70",
         10134 => x"2e",
         10135 => x"25",
         10136 => x"64",
         10137 => x"20",
         10138 => x"25",
         10139 => x"64",
         10140 => x"25",
         10141 => x"53",
         10142 => x"43",
         10143 => x"69",
         10144 => x"61",
         10145 => x"6e",
         10146 => x"20",
         10147 => x"6f",
         10148 => x"6f",
         10149 => x"6f",
         10150 => x"67",
         10151 => x"3a",
         10152 => x"76",
         10153 => x"73",
         10154 => x"70",
         10155 => x"65",
         10156 => x"64",
         10157 => x"20",
         10158 => x"57",
         10159 => x"44",
         10160 => x"20",
         10161 => x"30",
         10162 => x"25",
         10163 => x"29",
         10164 => x"20",
         10165 => x"53",
         10166 => x"4d",
         10167 => x"20",
         10168 => x"30",
         10169 => x"25",
         10170 => x"29",
         10171 => x"20",
         10172 => x"49",
         10173 => x"20",
         10174 => x"4d",
         10175 => x"30",
         10176 => x"25",
         10177 => x"29",
         10178 => x"20",
         10179 => x"42",
         10180 => x"20",
         10181 => x"20",
         10182 => x"30",
         10183 => x"25",
         10184 => x"29",
         10185 => x"20",
         10186 => x"52",
         10187 => x"20",
         10188 => x"20",
         10189 => x"30",
         10190 => x"25",
         10191 => x"29",
         10192 => x"20",
         10193 => x"53",
         10194 => x"41",
         10195 => x"20",
         10196 => x"65",
         10197 => x"65",
         10198 => x"25",
         10199 => x"29",
         10200 => x"20",
         10201 => x"54",
         10202 => x"52",
         10203 => x"20",
         10204 => x"69",
         10205 => x"73",
         10206 => x"25",
         10207 => x"29",
         10208 => x"20",
         10209 => x"49",
         10210 => x"20",
         10211 => x"4c",
         10212 => x"68",
         10213 => x"65",
         10214 => x"25",
         10215 => x"29",
         10216 => x"20",
         10217 => x"57",
         10218 => x"42",
         10219 => x"20",
         10220 => x"00",
         10221 => x"20",
         10222 => x"57",
         10223 => x"32",
         10224 => x"20",
         10225 => x"49",
         10226 => x"4c",
         10227 => x"20",
         10228 => x"50",
         10229 => x"20",
         10230 => x"53",
         10231 => x"41",
         10232 => x"65",
         10233 => x"73",
         10234 => x"20",
         10235 => x"43",
         10236 => x"52",
         10237 => x"74",
         10238 => x"63",
         10239 => x"20",
         10240 => x"72",
         10241 => x"20",
         10242 => x"30",
         10243 => x"00",
         10244 => x"20",
         10245 => x"43",
         10246 => x"4d",
         10247 => x"72",
         10248 => x"74",
         10249 => x"20",
         10250 => x"72",
         10251 => x"20",
         10252 => x"30",
         10253 => x"00",
         10254 => x"20",
         10255 => x"53",
         10256 => x"6b",
         10257 => x"61",
         10258 => x"41",
         10259 => x"65",
         10260 => x"20",
         10261 => x"20",
         10262 => x"30",
         10263 => x"00",
         10264 => x"4d",
         10265 => x"3a",
         10266 => x"20",
         10267 => x"5a",
         10268 => x"49",
         10269 => x"20",
         10270 => x"20",
         10271 => x"20",
         10272 => x"20",
         10273 => x"20",
         10274 => x"30",
         10275 => x"00",
         10276 => x"20",
         10277 => x"53",
         10278 => x"65",
         10279 => x"6c",
         10280 => x"20",
         10281 => x"71",
         10282 => x"20",
         10283 => x"20",
         10284 => x"64",
         10285 => x"34",
         10286 => x"7a",
         10287 => x"20",
         10288 => x"53",
         10289 => x"4d",
         10290 => x"6f",
         10291 => x"46",
         10292 => x"20",
         10293 => x"20",
         10294 => x"20",
         10295 => x"64",
         10296 => x"34",
         10297 => x"7a",
         10298 => x"20",
         10299 => x"57",
         10300 => x"62",
         10301 => x"20",
         10302 => x"41",
         10303 => x"6c",
         10304 => x"20",
         10305 => x"71",
         10306 => x"64",
         10307 => x"34",
         10308 => x"7a",
         10309 => x"53",
         10310 => x"6c",
         10311 => x"4d",
         10312 => x"75",
         10313 => x"46",
         10314 => x"00",
         10315 => x"45",
         10316 => x"45",
         10317 => x"00",
         10318 => x"55",
         10319 => x"6f",
         10320 => x"00",
         10321 => x"01",
         10322 => x"00",
         10323 => x"00",
         10324 => x"01",
         10325 => x"00",
         10326 => x"00",
         10327 => x"01",
         10328 => x"00",
         10329 => x"00",
         10330 => x"01",
         10331 => x"00",
         10332 => x"00",
         10333 => x"01",
         10334 => x"00",
         10335 => x"00",
         10336 => x"01",
         10337 => x"00",
         10338 => x"00",
         10339 => x"01",
         10340 => x"00",
         10341 => x"00",
         10342 => x"01",
         10343 => x"00",
         10344 => x"00",
         10345 => x"01",
         10346 => x"00",
         10347 => x"00",
         10348 => x"01",
         10349 => x"00",
         10350 => x"00",
         10351 => x"01",
         10352 => x"00",
         10353 => x"00",
         10354 => x"04",
         10355 => x"00",
         10356 => x"00",
         10357 => x"04",
         10358 => x"00",
         10359 => x"00",
         10360 => x"04",
         10361 => x"00",
         10362 => x"00",
         10363 => x"03",
         10364 => x"00",
         10365 => x"00",
         10366 => x"04",
         10367 => x"00",
         10368 => x"00",
         10369 => x"04",
         10370 => x"00",
         10371 => x"00",
         10372 => x"04",
         10373 => x"00",
         10374 => x"00",
         10375 => x"03",
         10376 => x"00",
         10377 => x"00",
         10378 => x"03",
         10379 => x"00",
         10380 => x"00",
         10381 => x"03",
         10382 => x"00",
         10383 => x"00",
         10384 => x"03",
         10385 => x"00",
         10386 => x"1b",
         10387 => x"1b",
         10388 => x"1b",
         10389 => x"1b",
         10390 => x"1b",
         10391 => x"1b",
         10392 => x"1b",
         10393 => x"1b",
         10394 => x"1b",
         10395 => x"1b",
         10396 => x"1b",
         10397 => x"10",
         10398 => x"0e",
         10399 => x"0d",
         10400 => x"0b",
         10401 => x"08",
         10402 => x"06",
         10403 => x"05",
         10404 => x"04",
         10405 => x"03",
         10406 => x"02",
         10407 => x"01",
         10408 => x"68",
         10409 => x"6f",
         10410 => x"68",
         10411 => x"00",
         10412 => x"21",
         10413 => x"25",
         10414 => x"75",
         10415 => x"73",
         10416 => x"46",
         10417 => x"65",
         10418 => x"6f",
         10419 => x"73",
         10420 => x"74",
         10421 => x"68",
         10422 => x"6f",
         10423 => x"66",
         10424 => x"20",
         10425 => x"45",
         10426 => x"00",
         10427 => x"43",
         10428 => x"6f",
         10429 => x"70",
         10430 => x"63",
         10431 => x"74",
         10432 => x"69",
         10433 => x"72",
         10434 => x"69",
         10435 => x"20",
         10436 => x"61",
         10437 => x"6e",
         10438 => x"53",
         10439 => x"22",
         10440 => x"3e",
         10441 => x"00",
         10442 => x"2b",
         10443 => x"5b",
         10444 => x"46",
         10445 => x"46",
         10446 => x"32",
         10447 => x"eb",
         10448 => x"53",
         10449 => x"35",
         10450 => x"4e",
         10451 => x"41",
         10452 => x"20",
         10453 => x"41",
         10454 => x"20",
         10455 => x"4e",
         10456 => x"41",
         10457 => x"20",
         10458 => x"41",
         10459 => x"20",
         10460 => x"00",
         10461 => x"00",
         10462 => x"00",
         10463 => x"00",
         10464 => x"01",
         10465 => x"09",
         10466 => x"14",
         10467 => x"1e",
         10468 => x"80",
         10469 => x"8e",
         10470 => x"45",
         10471 => x"49",
         10472 => x"90",
         10473 => x"99",
         10474 => x"59",
         10475 => x"9c",
         10476 => x"41",
         10477 => x"a5",
         10478 => x"a8",
         10479 => x"ac",
         10480 => x"b0",
         10481 => x"b4",
         10482 => x"b8",
         10483 => x"bc",
         10484 => x"c0",
         10485 => x"c4",
         10486 => x"c8",
         10487 => x"cc",
         10488 => x"d0",
         10489 => x"d4",
         10490 => x"d8",
         10491 => x"dc",
         10492 => x"e0",
         10493 => x"e4",
         10494 => x"e8",
         10495 => x"ec",
         10496 => x"f0",
         10497 => x"f4",
         10498 => x"f8",
         10499 => x"fc",
         10500 => x"2b",
         10501 => x"3d",
         10502 => x"5c",
         10503 => x"3c",
         10504 => x"7f",
         10505 => x"00",
         10506 => x"00",
         10507 => x"01",
         10508 => x"00",
         10509 => x"00",
         10510 => x"00",
         10511 => x"00",
         10512 => x"00",
         10513 => x"00",
         10514 => x"00",
         10515 => x"00",
         10516 => x"00",
         10517 => x"00",
         10518 => x"00",
         10519 => x"00",
         10520 => x"00",
         10521 => x"00",
         10522 => x"00",
         10523 => x"00",
         10524 => x"00",
         10525 => x"00",
         10526 => x"00",
         10527 => x"00",
         10528 => x"20",
         10529 => x"00",
         10530 => x"00",
         10531 => x"00",
         10532 => x"00",
         10533 => x"00",
         10534 => x"00",
         10535 => x"00",
         10536 => x"00",
         10537 => x"25",
         10538 => x"25",
         10539 => x"25",
         10540 => x"25",
         10541 => x"25",
         10542 => x"25",
         10543 => x"25",
         10544 => x"25",
         10545 => x"25",
         10546 => x"25",
         10547 => x"25",
         10548 => x"25",
         10549 => x"25",
         10550 => x"25",
         10551 => x"25",
         10552 => x"25",
         10553 => x"25",
         10554 => x"25",
         10555 => x"25",
         10556 => x"25",
         10557 => x"25",
         10558 => x"25",
         10559 => x"25",
         10560 => x"25",
         10561 => x"03",
         10562 => x"03",
         10563 => x"03",
         10564 => x"00",
         10565 => x"03",
         10566 => x"03",
         10567 => x"22",
         10568 => x"03",
         10569 => x"22",
         10570 => x"22",
         10571 => x"23",
         10572 => x"00",
         10573 => x"00",
         10574 => x"00",
         10575 => x"20",
         10576 => x"25",
         10577 => x"00",
         10578 => x"00",
         10579 => x"00",
         10580 => x"00",
         10581 => x"01",
         10582 => x"01",
         10583 => x"01",
         10584 => x"01",
         10585 => x"01",
         10586 => x"01",
         10587 => x"00",
         10588 => x"01",
         10589 => x"01",
         10590 => x"01",
         10591 => x"01",
         10592 => x"01",
         10593 => x"01",
         10594 => x"01",
         10595 => x"01",
         10596 => x"01",
         10597 => x"01",
         10598 => x"01",
         10599 => x"01",
         10600 => x"01",
         10601 => x"01",
         10602 => x"01",
         10603 => x"01",
         10604 => x"01",
         10605 => x"01",
         10606 => x"01",
         10607 => x"01",
         10608 => x"01",
         10609 => x"01",
         10610 => x"01",
         10611 => x"01",
         10612 => x"01",
         10613 => x"01",
         10614 => x"01",
         10615 => x"01",
         10616 => x"01",
         10617 => x"01",
         10618 => x"01",
         10619 => x"01",
         10620 => x"01",
         10621 => x"01",
         10622 => x"01",
         10623 => x"01",
         10624 => x"01",
         10625 => x"01",
         10626 => x"01",
         10627 => x"01",
         10628 => x"01",
         10629 => x"01",
         10630 => x"00",
         10631 => x"01",
         10632 => x"01",
         10633 => x"02",
         10634 => x"02",
         10635 => x"2c",
         10636 => x"02",
         10637 => x"2c",
         10638 => x"02",
         10639 => x"02",
         10640 => x"01",
         10641 => x"00",
         10642 => x"01",
         10643 => x"01",
         10644 => x"02",
         10645 => x"02",
         10646 => x"02",
         10647 => x"02",
         10648 => x"01",
         10649 => x"02",
         10650 => x"02",
         10651 => x"02",
         10652 => x"01",
         10653 => x"02",
         10654 => x"02",
         10655 => x"02",
         10656 => x"02",
         10657 => x"01",
         10658 => x"02",
         10659 => x"02",
         10660 => x"02",
         10661 => x"02",
         10662 => x"02",
         10663 => x"02",
         10664 => x"01",
         10665 => x"02",
         10666 => x"02",
         10667 => x"02",
         10668 => x"01",
         10669 => x"01",
         10670 => x"02",
         10671 => x"02",
         10672 => x"02",
         10673 => x"01",
         10674 => x"00",
         10675 => x"03",
         10676 => x"03",
         10677 => x"03",
         10678 => x"03",
         10679 => x"03",
         10680 => x"03",
         10681 => x"03",
         10682 => x"03",
         10683 => x"03",
         10684 => x"03",
         10685 => x"03",
         10686 => x"01",
         10687 => x"00",
         10688 => x"03",
         10689 => x"03",
         10690 => x"03",
         10691 => x"03",
         10692 => x"03",
         10693 => x"03",
         10694 => x"07",
         10695 => x"01",
         10696 => x"01",
         10697 => x"01",
         10698 => x"00",
         10699 => x"04",
         10700 => x"05",
         10701 => x"00",
         10702 => x"1d",
         10703 => x"2c",
         10704 => x"01",
         10705 => x"01",
         10706 => x"06",
         10707 => x"06",
         10708 => x"06",
         10709 => x"06",
         10710 => x"06",
         10711 => x"00",
         10712 => x"1f",
         10713 => x"1f",
         10714 => x"1f",
         10715 => x"1f",
         10716 => x"1f",
         10717 => x"1f",
         10718 => x"1f",
         10719 => x"1f",
         10720 => x"1f",
         10721 => x"1f",
         10722 => x"1f",
         10723 => x"1f",
         10724 => x"1f",
         10725 => x"1f",
         10726 => x"1f",
         10727 => x"1f",
         10728 => x"1f",
         10729 => x"1f",
         10730 => x"1f",
         10731 => x"1f",
         10732 => x"06",
         10733 => x"06",
         10734 => x"00",
         10735 => x"1f",
         10736 => x"1f",
         10737 => x"00",
         10738 => x"21",
         10739 => x"21",
         10740 => x"21",
         10741 => x"05",
         10742 => x"04",
         10743 => x"01",
         10744 => x"01",
         10745 => x"01",
         10746 => x"01",
         10747 => x"08",
         10748 => x"03",
         10749 => x"00",
         10750 => x"00",
         10751 => x"01",
         10752 => x"00",
         10753 => x"00",
         10754 => x"00",
         10755 => x"01",
         10756 => x"00",
         10757 => x"00",
         10758 => x"00",
         10759 => x"01",
         10760 => x"00",
         10761 => x"00",
         10762 => x"00",
         10763 => x"01",
         10764 => x"00",
         10765 => x"00",
         10766 => x"00",
         10767 => x"01",
         10768 => x"00",
         10769 => x"00",
         10770 => x"00",
         10771 => x"01",
         10772 => x"00",
         10773 => x"00",
         10774 => x"00",
         10775 => x"01",
         10776 => x"00",
         10777 => x"00",
         10778 => x"00",
         10779 => x"01",
         10780 => x"00",
         10781 => x"00",
         10782 => x"00",
         10783 => x"01",
         10784 => x"00",
         10785 => x"00",
         10786 => x"00",
         10787 => x"01",
         10788 => x"00",
         10789 => x"00",
         10790 => x"00",
         10791 => x"01",
         10792 => x"00",
         10793 => x"00",
         10794 => x"00",
         10795 => x"01",
         10796 => x"00",
         10797 => x"00",
         10798 => x"00",
         10799 => x"01",
         10800 => x"00",
         10801 => x"00",
         10802 => x"00",
         10803 => x"01",
         10804 => x"00",
         10805 => x"00",
         10806 => x"00",
         10807 => x"01",
         10808 => x"00",
         10809 => x"00",
         10810 => x"00",
         10811 => x"01",
         10812 => x"00",
         10813 => x"00",
         10814 => x"00",
         10815 => x"01",
         10816 => x"00",
         10817 => x"00",
         10818 => x"00",
         10819 => x"01",
         10820 => x"00",
         10821 => x"00",
         10822 => x"00",
         10823 => x"01",
         10824 => x"00",
         10825 => x"00",
         10826 => x"00",
         10827 => x"01",
         10828 => x"00",
         10829 => x"00",
         10830 => x"00",
         10831 => x"01",
         10832 => x"00",
         10833 => x"00",
         10834 => x"00",
         10835 => x"01",
         10836 => x"00",
         10837 => x"00",
         10838 => x"00",
         10839 => x"01",
         10840 => x"00",
         10841 => x"00",
         10842 => x"00",
         10843 => x"01",
         10844 => x"00",
         10845 => x"00",
         10846 => x"00",
         10847 => x"01",
         10848 => x"00",
         10849 => x"00",
         10850 => x"00",
         10851 => x"01",
         10852 => x"00",
         10853 => x"00",
         10854 => x"00",
         10855 => x"00",
         10856 => x"00",
         10857 => x"00",
         10858 => x"00",
         10859 => x"00",
         10860 => x"00",
         10861 => x"00",
         10862 => x"00",
         10863 => x"01",
         10864 => x"01",
         10865 => x"00",
         10866 => x"00",
         10867 => x"00",
         10868 => x"00",
         10869 => x"05",
         10870 => x"05",
         10871 => x"05",
         10872 => x"00",
         10873 => x"01",
         10874 => x"01",
         10875 => x"01",
         10876 => x"01",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"00",
         10884 => x"00",
         10885 => x"00",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"00",
         10890 => x"00",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"00",
         10895 => x"00",
         10896 => x"00",
         10897 => x"00",
         10898 => x"00",
         10899 => x"00",
         10900 => x"00",
         10901 => x"00",
         10902 => x"01",
         10903 => x"00",
         10904 => x"01",
         10905 => x"00",
         10906 => x"02",
         10907 => x"00",
         10908 => x"00",
         10909 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
