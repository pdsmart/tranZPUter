-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.softZPU_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"b0",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"be",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"ac",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"ab",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8f",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"90",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"91",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"92",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"98",
           386 => x"f6",
           387 => x"98",
           388 => x"80",
           389 => x"ba",
           390 => x"ee",
           391 => x"98",
           392 => x"80",
           393 => x"ba",
           394 => x"f3",
           395 => x"98",
           396 => x"80",
           397 => x"ba",
           398 => x"e0",
           399 => x"98",
           400 => x"80",
           401 => x"ba",
           402 => x"a3",
           403 => x"98",
           404 => x"80",
           405 => x"ba",
           406 => x"f6",
           407 => x"98",
           408 => x"80",
           409 => x"ba",
           410 => x"86",
           411 => x"98",
           412 => x"80",
           413 => x"ba",
           414 => x"82",
           415 => x"98",
           416 => x"80",
           417 => x"ba",
           418 => x"88",
           419 => x"98",
           420 => x"80",
           421 => x"ba",
           422 => x"a8",
           423 => x"98",
           424 => x"80",
           425 => x"ba",
           426 => x"d1",
           427 => x"98",
           428 => x"80",
           429 => x"ba",
           430 => x"8a",
           431 => x"98",
           432 => x"80",
           433 => x"ba",
           434 => x"d4",
           435 => x"ba",
           436 => x"c0",
           437 => x"84",
           438 => x"80",
           439 => x"84",
           440 => x"80",
           441 => x"04",
           442 => x"0c",
           443 => x"2d",
           444 => x"08",
           445 => x"90",
           446 => x"98",
           447 => x"ca",
           448 => x"98",
           449 => x"80",
           450 => x"ba",
           451 => x"c9",
           452 => x"ba",
           453 => x"c0",
           454 => x"84",
           455 => x"82",
           456 => x"84",
           457 => x"80",
           458 => x"04",
           459 => x"0c",
           460 => x"2d",
           461 => x"08",
           462 => x"90",
           463 => x"98",
           464 => x"89",
           465 => x"98",
           466 => x"80",
           467 => x"ba",
           468 => x"ed",
           469 => x"ba",
           470 => x"c0",
           471 => x"84",
           472 => x"82",
           473 => x"84",
           474 => x"80",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"90",
           480 => x"98",
           481 => x"87",
           482 => x"98",
           483 => x"80",
           484 => x"ba",
           485 => x"f3",
           486 => x"ba",
           487 => x"c0",
           488 => x"84",
           489 => x"82",
           490 => x"84",
           491 => x"80",
           492 => x"04",
           493 => x"0c",
           494 => x"2d",
           495 => x"08",
           496 => x"90",
           497 => x"98",
           498 => x"b0",
           499 => x"98",
           500 => x"80",
           501 => x"ba",
           502 => x"8b",
           503 => x"ba",
           504 => x"c0",
           505 => x"84",
           506 => x"82",
           507 => x"84",
           508 => x"80",
           509 => x"04",
           510 => x"0c",
           511 => x"2d",
           512 => x"08",
           513 => x"90",
           514 => x"98",
           515 => x"d1",
           516 => x"98",
           517 => x"80",
           518 => x"ba",
           519 => x"e6",
           520 => x"ba",
           521 => x"c0",
           522 => x"84",
           523 => x"82",
           524 => x"84",
           525 => x"80",
           526 => x"04",
           527 => x"0c",
           528 => x"2d",
           529 => x"08",
           530 => x"90",
           531 => x"98",
           532 => x"f0",
           533 => x"98",
           534 => x"80",
           535 => x"ba",
           536 => x"96",
           537 => x"ba",
           538 => x"c0",
           539 => x"84",
           540 => x"83",
           541 => x"84",
           542 => x"80",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"90",
           548 => x"98",
           549 => x"c8",
           550 => x"98",
           551 => x"80",
           552 => x"ba",
           553 => x"a4",
           554 => x"ba",
           555 => x"c0",
           556 => x"84",
           557 => x"83",
           558 => x"84",
           559 => x"80",
           560 => x"04",
           561 => x"0c",
           562 => x"2d",
           563 => x"08",
           564 => x"90",
           565 => x"98",
           566 => x"ac",
           567 => x"98",
           568 => x"80",
           569 => x"ba",
           570 => x"f5",
           571 => x"ba",
           572 => x"c0",
           573 => x"84",
           574 => x"81",
           575 => x"84",
           576 => x"80",
           577 => x"04",
           578 => x"0c",
           579 => x"2d",
           580 => x"08",
           581 => x"90",
           582 => x"98",
           583 => x"e9",
           584 => x"98",
           585 => x"80",
           586 => x"ba",
           587 => x"d7",
           588 => x"ba",
           589 => x"c0",
           590 => x"84",
           591 => x"b1",
           592 => x"ba",
           593 => x"c0",
           594 => x"84",
           595 => x"81",
           596 => x"84",
           597 => x"80",
           598 => x"04",
           599 => x"0c",
           600 => x"2d",
           601 => x"08",
           602 => x"90",
           603 => x"98",
           604 => x"86",
           605 => x"98",
           606 => x"80",
           607 => x"ba",
           608 => x"d5",
           609 => x"ba",
           610 => x"c0",
           611 => x"3c",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"00",
           621 => x"ff",
           622 => x"06",
           623 => x"83",
           624 => x"10",
           625 => x"fc",
           626 => x"51",
           627 => x"80",
           628 => x"ff",
           629 => x"06",
           630 => x"52",
           631 => x"0a",
           632 => x"38",
           633 => x"51",
           634 => x"8c",
           635 => x"f8",
           636 => x"80",
           637 => x"05",
           638 => x"0b",
           639 => x"04",
           640 => x"80",
           641 => x"00",
           642 => x"87",
           643 => x"84",
           644 => x"56",
           645 => x"84",
           646 => x"51",
           647 => x"86",
           648 => x"fa",
           649 => x"7a",
           650 => x"33",
           651 => x"06",
           652 => x"07",
           653 => x"57",
           654 => x"72",
           655 => x"06",
           656 => x"ff",
           657 => x"8a",
           658 => x"70",
           659 => x"2a",
           660 => x"56",
           661 => x"25",
           662 => x"80",
           663 => x"75",
           664 => x"3f",
           665 => x"08",
           666 => x"8c",
           667 => x"ae",
           668 => x"8c",
           669 => x"81",
           670 => x"ff",
           671 => x"32",
           672 => x"72",
           673 => x"51",
           674 => x"73",
           675 => x"38",
           676 => x"76",
           677 => x"ba",
           678 => x"3d",
           679 => x"0b",
           680 => x"0c",
           681 => x"04",
           682 => x"7d",
           683 => x"84",
           684 => x"34",
           685 => x"0a",
           686 => x"88",
           687 => x"52",
           688 => x"05",
           689 => x"73",
           690 => x"74",
           691 => x"0d",
           692 => x"0d",
           693 => x"05",
           694 => x"75",
           695 => x"85",
           696 => x"f1",
           697 => x"63",
           698 => x"5d",
           699 => x"1f",
           700 => x"33",
           701 => x"81",
           702 => x"55",
           703 => x"54",
           704 => x"09",
           705 => x"d2",
           706 => x"57",
           707 => x"80",
           708 => x"1c",
           709 => x"54",
           710 => x"2e",
           711 => x"d0",
           712 => x"89",
           713 => x"38",
           714 => x"70",
           715 => x"25",
           716 => x"78",
           717 => x"80",
           718 => x"7a",
           719 => x"81",
           720 => x"40",
           721 => x"2e",
           722 => x"82",
           723 => x"7b",
           724 => x"ff",
           725 => x"1d",
           726 => x"84",
           727 => x"91",
           728 => x"7a",
           729 => x"78",
           730 => x"79",
           731 => x"98",
           732 => x"2c",
           733 => x"80",
           734 => x"0a",
           735 => x"2c",
           736 => x"56",
           737 => x"24",
           738 => x"73",
           739 => x"72",
           740 => x"78",
           741 => x"58",
           742 => x"38",
           743 => x"76",
           744 => x"81",
           745 => x"81",
           746 => x"5a",
           747 => x"33",
           748 => x"fe",
           749 => x"9e",
           750 => x"76",
           751 => x"3f",
           752 => x"76",
           753 => x"ff",
           754 => x"83",
           755 => x"06",
           756 => x"8a",
           757 => x"74",
           758 => x"7e",
           759 => x"17",
           760 => x"d8",
           761 => x"72",
           762 => x"ca",
           763 => x"73",
           764 => x"e0",
           765 => x"80",
           766 => x"eb",
           767 => x"76",
           768 => x"3f",
           769 => x"58",
           770 => x"86",
           771 => x"39",
           772 => x"fe",
           773 => x"5a",
           774 => x"05",
           775 => x"83",
           776 => x"5e",
           777 => x"84",
           778 => x"79",
           779 => x"93",
           780 => x"ba",
           781 => x"ff",
           782 => x"8c",
           783 => x"05",
           784 => x"89",
           785 => x"84",
           786 => x"b0",
           787 => x"7e",
           788 => x"40",
           789 => x"75",
           790 => x"3f",
           791 => x"08",
           792 => x"8c",
           793 => x"7d",
           794 => x"31",
           795 => x"b2",
           796 => x"7e",
           797 => x"38",
           798 => x"80",
           799 => x"80",
           800 => x"2c",
           801 => x"86",
           802 => x"06",
           803 => x"80",
           804 => x"77",
           805 => x"29",
           806 => x"05",
           807 => x"2e",
           808 => x"84",
           809 => x"fc",
           810 => x"53",
           811 => x"58",
           812 => x"70",
           813 => x"55",
           814 => x"9e",
           815 => x"2c",
           816 => x"06",
           817 => x"73",
           818 => x"38",
           819 => x"f7",
           820 => x"2a",
           821 => x"41",
           822 => x"81",
           823 => x"80",
           824 => x"38",
           825 => x"90",
           826 => x"2c",
           827 => x"06",
           828 => x"73",
           829 => x"96",
           830 => x"2a",
           831 => x"73",
           832 => x"7a",
           833 => x"06",
           834 => x"98",
           835 => x"2a",
           836 => x"73",
           837 => x"7e",
           838 => x"73",
           839 => x"7a",
           840 => x"06",
           841 => x"2e",
           842 => x"78",
           843 => x"29",
           844 => x"05",
           845 => x"5a",
           846 => x"74",
           847 => x"7c",
           848 => x"88",
           849 => x"78",
           850 => x"29",
           851 => x"05",
           852 => x"5a",
           853 => x"80",
           854 => x"74",
           855 => x"72",
           856 => x"38",
           857 => x"80",
           858 => x"ff",
           859 => x"98",
           860 => x"55",
           861 => x"9d",
           862 => x"b0",
           863 => x"3f",
           864 => x"80",
           865 => x"ff",
           866 => x"98",
           867 => x"55",
           868 => x"e5",
           869 => x"2a",
           870 => x"5c",
           871 => x"2e",
           872 => x"76",
           873 => x"84",
           874 => x"80",
           875 => x"ca",
           876 => x"d3",
           877 => x"38",
           878 => x"9c",
           879 => x"7c",
           880 => x"70",
           881 => x"87",
           882 => x"84",
           883 => x"09",
           884 => x"38",
           885 => x"5b",
           886 => x"fc",
           887 => x"78",
           888 => x"29",
           889 => x"05",
           890 => x"5a",
           891 => x"75",
           892 => x"38",
           893 => x"51",
           894 => x"e2",
           895 => x"07",
           896 => x"07",
           897 => x"5b",
           898 => x"38",
           899 => x"7a",
           900 => x"5b",
           901 => x"90",
           902 => x"05",
           903 => x"83",
           904 => x"5f",
           905 => x"5a",
           906 => x"7f",
           907 => x"77",
           908 => x"06",
           909 => x"70",
           910 => x"07",
           911 => x"80",
           912 => x"80",
           913 => x"2c",
           914 => x"56",
           915 => x"7a",
           916 => x"81",
           917 => x"7a",
           918 => x"77",
           919 => x"80",
           920 => x"80",
           921 => x"2c",
           922 => x"80",
           923 => x"b3",
           924 => x"a0",
           925 => x"3f",
           926 => x"1a",
           927 => x"ff",
           928 => x"79",
           929 => x"2e",
           930 => x"7c",
           931 => x"81",
           932 => x"51",
           933 => x"e2",
           934 => x"70",
           935 => x"06",
           936 => x"83",
           937 => x"fe",
           938 => x"52",
           939 => x"05",
           940 => x"85",
           941 => x"39",
           942 => x"06",
           943 => x"07",
           944 => x"80",
           945 => x"80",
           946 => x"2c",
           947 => x"80",
           948 => x"2a",
           949 => x"5d",
           950 => x"fd",
           951 => x"fb",
           952 => x"84",
           953 => x"70",
           954 => x"56",
           955 => x"82",
           956 => x"83",
           957 => x"5b",
           958 => x"5e",
           959 => x"7a",
           960 => x"33",
           961 => x"f8",
           962 => x"ca",
           963 => x"07",
           964 => x"33",
           965 => x"f7",
           966 => x"ba",
           967 => x"84",
           968 => x"77",
           969 => x"58",
           970 => x"82",
           971 => x"51",
           972 => x"84",
           973 => x"83",
           974 => x"78",
           975 => x"2b",
           976 => x"90",
           977 => x"87",
           978 => x"c0",
           979 => x"58",
           980 => x"be",
           981 => x"39",
           982 => x"05",
           983 => x"81",
           984 => x"41",
           985 => x"cf",
           986 => x"87",
           987 => x"ba",
           988 => x"ff",
           989 => x"71",
           990 => x"54",
           991 => x"7a",
           992 => x"7c",
           993 => x"76",
           994 => x"f7",
           995 => x"78",
           996 => x"29",
           997 => x"05",
           998 => x"5a",
           999 => x"74",
          1000 => x"38",
          1001 => x"51",
          1002 => x"e2",
          1003 => x"b0",
          1004 => x"3f",
          1005 => x"09",
          1006 => x"e3",
          1007 => x"76",
          1008 => x"3f",
          1009 => x"81",
          1010 => x"80",
          1011 => x"38",
          1012 => x"75",
          1013 => x"71",
          1014 => x"70",
          1015 => x"83",
          1016 => x"5a",
          1017 => x"fa",
          1018 => x"a2",
          1019 => x"ad",
          1020 => x"3f",
          1021 => x"54",
          1022 => x"fa",
          1023 => x"ad",
          1024 => x"75",
          1025 => x"82",
          1026 => x"81",
          1027 => x"80",
          1028 => x"38",
          1029 => x"78",
          1030 => x"2b",
          1031 => x"5a",
          1032 => x"39",
          1033 => x"51",
          1034 => x"c8",
          1035 => x"a0",
          1036 => x"3f",
          1037 => x"78",
          1038 => x"88",
          1039 => x"ba",
          1040 => x"ff",
          1041 => x"71",
          1042 => x"54",
          1043 => x"39",
          1044 => x"7e",
          1045 => x"ff",
          1046 => x"57",
          1047 => x"39",
          1048 => x"84",
          1049 => x"53",
          1050 => x"51",
          1051 => x"84",
          1052 => x"fa",
          1053 => x"55",
          1054 => x"d5",
          1055 => x"11",
          1056 => x"2a",
          1057 => x"81",
          1058 => x"58",
          1059 => x"56",
          1060 => x"09",
          1061 => x"d5",
          1062 => x"81",
          1063 => x"53",
          1064 => x"b0",
          1065 => x"f0",
          1066 => x"51",
          1067 => x"53",
          1068 => x"ba",
          1069 => x"2e",
          1070 => x"57",
          1071 => x"05",
          1072 => x"72",
          1073 => x"38",
          1074 => x"08",
          1075 => x"84",
          1076 => x"54",
          1077 => x"08",
          1078 => x"90",
          1079 => x"74",
          1080 => x"8c",
          1081 => x"83",
          1082 => x"76",
          1083 => x"ba",
          1084 => x"3d",
          1085 => x"3d",
          1086 => x"56",
          1087 => x"85",
          1088 => x"81",
          1089 => x"70",
          1090 => x"55",
          1091 => x"56",
          1092 => x"09",
          1093 => x"38",
          1094 => x"05",
          1095 => x"72",
          1096 => x"81",
          1097 => x"76",
          1098 => x"ba",
          1099 => x"3d",
          1100 => x"70",
          1101 => x"33",
          1102 => x"2e",
          1103 => x"52",
          1104 => x"15",
          1105 => x"2d",
          1106 => x"08",
          1107 => x"38",
          1108 => x"81",
          1109 => x"54",
          1110 => x"38",
          1111 => x"3d",
          1112 => x"f0",
          1113 => x"51",
          1114 => x"3d",
          1115 => x"3d",
          1116 => x"85",
          1117 => x"81",
          1118 => x"81",
          1119 => x"56",
          1120 => x"72",
          1121 => x"82",
          1122 => x"54",
          1123 => x"ac",
          1124 => x"08",
          1125 => x"16",
          1126 => x"38",
          1127 => x"76",
          1128 => x"08",
          1129 => x"0c",
          1130 => x"53",
          1131 => x"16",
          1132 => x"75",
          1133 => x"0c",
          1134 => x"04",
          1135 => x"81",
          1136 => x"90",
          1137 => x"73",
          1138 => x"84",
          1139 => x"e3",
          1140 => x"08",
          1141 => x"16",
          1142 => x"d7",
          1143 => x"0d",
          1144 => x"33",
          1145 => x"06",
          1146 => x"81",
          1147 => x"56",
          1148 => x"71",
          1149 => x"86",
          1150 => x"52",
          1151 => x"72",
          1152 => x"06",
          1153 => x"2e",
          1154 => x"75",
          1155 => x"53",
          1156 => x"2e",
          1157 => x"81",
          1158 => x"8c",
          1159 => x"05",
          1160 => x"71",
          1161 => x"54",
          1162 => x"8c",
          1163 => x"0d",
          1164 => x"bf",
          1165 => x"85",
          1166 => x"16",
          1167 => x"8c",
          1168 => x"16",
          1169 => x"8c",
          1170 => x"0d",
          1171 => x"94",
          1172 => x"74",
          1173 => x"8c",
          1174 => x"ba",
          1175 => x"25",
          1176 => x"85",
          1177 => x"90",
          1178 => x"84",
          1179 => x"ff",
          1180 => x"71",
          1181 => x"72",
          1182 => x"ff",
          1183 => x"ba",
          1184 => x"3d",
          1185 => x"a0",
          1186 => x"85",
          1187 => x"54",
          1188 => x"3d",
          1189 => x"71",
          1190 => x"71",
          1191 => x"53",
          1192 => x"f7",
          1193 => x"52",
          1194 => x"05",
          1195 => x"70",
          1196 => x"05",
          1197 => x"f0",
          1198 => x"ba",
          1199 => x"3d",
          1200 => x"3d",
          1201 => x"71",
          1202 => x"52",
          1203 => x"2e",
          1204 => x"72",
          1205 => x"70",
          1206 => x"38",
          1207 => x"05",
          1208 => x"70",
          1209 => x"34",
          1210 => x"70",
          1211 => x"84",
          1212 => x"86",
          1213 => x"70",
          1214 => x"75",
          1215 => x"70",
          1216 => x"53",
          1217 => x"13",
          1218 => x"33",
          1219 => x"11",
          1220 => x"2e",
          1221 => x"13",
          1222 => x"53",
          1223 => x"34",
          1224 => x"70",
          1225 => x"39",
          1226 => x"74",
          1227 => x"71",
          1228 => x"53",
          1229 => x"f7",
          1230 => x"70",
          1231 => x"ba",
          1232 => x"84",
          1233 => x"fd",
          1234 => x"77",
          1235 => x"54",
          1236 => x"05",
          1237 => x"70",
          1238 => x"05",
          1239 => x"f0",
          1240 => x"ba",
          1241 => x"3d",
          1242 => x"3d",
          1243 => x"71",
          1244 => x"52",
          1245 => x"2e",
          1246 => x"70",
          1247 => x"33",
          1248 => x"05",
          1249 => x"11",
          1250 => x"38",
          1251 => x"8c",
          1252 => x"0d",
          1253 => x"0d",
          1254 => x"55",
          1255 => x"80",
          1256 => x"73",
          1257 => x"81",
          1258 => x"52",
          1259 => x"2e",
          1260 => x"9a",
          1261 => x"54",
          1262 => x"b7",
          1263 => x"53",
          1264 => x"80",
          1265 => x"ba",
          1266 => x"3d",
          1267 => x"80",
          1268 => x"73",
          1269 => x"51",
          1270 => x"e9",
          1271 => x"33",
          1272 => x"71",
          1273 => x"38",
          1274 => x"84",
          1275 => x"86",
          1276 => x"71",
          1277 => x"0c",
          1278 => x"04",
          1279 => x"77",
          1280 => x"52",
          1281 => x"3f",
          1282 => x"08",
          1283 => x"08",
          1284 => x"55",
          1285 => x"3f",
          1286 => x"08",
          1287 => x"8c",
          1288 => x"9b",
          1289 => x"8c",
          1290 => x"80",
          1291 => x"53",
          1292 => x"ba",
          1293 => x"fe",
          1294 => x"ba",
          1295 => x"73",
          1296 => x"0c",
          1297 => x"04",
          1298 => x"75",
          1299 => x"54",
          1300 => x"71",
          1301 => x"38",
          1302 => x"05",
          1303 => x"70",
          1304 => x"38",
          1305 => x"71",
          1306 => x"81",
          1307 => x"ff",
          1308 => x"31",
          1309 => x"84",
          1310 => x"85",
          1311 => x"fd",
          1312 => x"77",
          1313 => x"53",
          1314 => x"80",
          1315 => x"72",
          1316 => x"05",
          1317 => x"11",
          1318 => x"38",
          1319 => x"8c",
          1320 => x"0d",
          1321 => x"0d",
          1322 => x"54",
          1323 => x"80",
          1324 => x"76",
          1325 => x"3f",
          1326 => x"08",
          1327 => x"53",
          1328 => x"8d",
          1329 => x"80",
          1330 => x"84",
          1331 => x"31",
          1332 => x"72",
          1333 => x"cb",
          1334 => x"72",
          1335 => x"c3",
          1336 => x"74",
          1337 => x"72",
          1338 => x"2b",
          1339 => x"55",
          1340 => x"76",
          1341 => x"72",
          1342 => x"2a",
          1343 => x"77",
          1344 => x"31",
          1345 => x"2c",
          1346 => x"7b",
          1347 => x"71",
          1348 => x"5c",
          1349 => x"55",
          1350 => x"74",
          1351 => x"10",
          1352 => x"71",
          1353 => x"0c",
          1354 => x"04",
          1355 => x"76",
          1356 => x"80",
          1357 => x"70",
          1358 => x"25",
          1359 => x"90",
          1360 => x"71",
          1361 => x"fe",
          1362 => x"30",
          1363 => x"83",
          1364 => x"31",
          1365 => x"70",
          1366 => x"70",
          1367 => x"25",
          1368 => x"71",
          1369 => x"2a",
          1370 => x"1b",
          1371 => x"06",
          1372 => x"80",
          1373 => x"71",
          1374 => x"2a",
          1375 => x"81",
          1376 => x"06",
          1377 => x"74",
          1378 => x"19",
          1379 => x"8c",
          1380 => x"54",
          1381 => x"56",
          1382 => x"55",
          1383 => x"56",
          1384 => x"58",
          1385 => x"86",
          1386 => x"fd",
          1387 => x"77",
          1388 => x"53",
          1389 => x"94",
          1390 => x"8c",
          1391 => x"74",
          1392 => x"ba",
          1393 => x"85",
          1394 => x"fa",
          1395 => x"7a",
          1396 => x"53",
          1397 => x"8b",
          1398 => x"fe",
          1399 => x"ba",
          1400 => x"e0",
          1401 => x"80",
          1402 => x"73",
          1403 => x"3f",
          1404 => x"8c",
          1405 => x"73",
          1406 => x"26",
          1407 => x"80",
          1408 => x"2e",
          1409 => x"12",
          1410 => x"a0",
          1411 => x"71",
          1412 => x"54",
          1413 => x"74",
          1414 => x"38",
          1415 => x"9f",
          1416 => x"10",
          1417 => x"72",
          1418 => x"9f",
          1419 => x"06",
          1420 => x"75",
          1421 => x"1c",
          1422 => x"52",
          1423 => x"53",
          1424 => x"72",
          1425 => x"0c",
          1426 => x"04",
          1427 => x"78",
          1428 => x"9f",
          1429 => x"2c",
          1430 => x"9f",
          1431 => x"73",
          1432 => x"74",
          1433 => x"75",
          1434 => x"56",
          1435 => x"fc",
          1436 => x"ba",
          1437 => x"32",
          1438 => x"ba",
          1439 => x"3d",
          1440 => x"3d",
          1441 => x"5b",
          1442 => x"7b",
          1443 => x"70",
          1444 => x"59",
          1445 => x"09",
          1446 => x"38",
          1447 => x"78",
          1448 => x"55",
          1449 => x"2e",
          1450 => x"ad",
          1451 => x"38",
          1452 => x"81",
          1453 => x"14",
          1454 => x"77",
          1455 => x"db",
          1456 => x"80",
          1457 => x"27",
          1458 => x"80",
          1459 => x"89",
          1460 => x"70",
          1461 => x"55",
          1462 => x"70",
          1463 => x"51",
          1464 => x"27",
          1465 => x"13",
          1466 => x"06",
          1467 => x"73",
          1468 => x"38",
          1469 => x"81",
          1470 => x"76",
          1471 => x"16",
          1472 => x"70",
          1473 => x"56",
          1474 => x"ff",
          1475 => x"80",
          1476 => x"75",
          1477 => x"7a",
          1478 => x"75",
          1479 => x"0c",
          1480 => x"04",
          1481 => x"70",
          1482 => x"33",
          1483 => x"73",
          1484 => x"81",
          1485 => x"38",
          1486 => x"78",
          1487 => x"55",
          1488 => x"e2",
          1489 => x"90",
          1490 => x"f8",
          1491 => x"81",
          1492 => x"27",
          1493 => x"14",
          1494 => x"88",
          1495 => x"27",
          1496 => x"75",
          1497 => x"0c",
          1498 => x"04",
          1499 => x"15",
          1500 => x"70",
          1501 => x"80",
          1502 => x"39",
          1503 => x"ba",
          1504 => x"3d",
          1505 => x"3d",
          1506 => x"5b",
          1507 => x"7b",
          1508 => x"70",
          1509 => x"59",
          1510 => x"09",
          1511 => x"38",
          1512 => x"78",
          1513 => x"55",
          1514 => x"2e",
          1515 => x"ad",
          1516 => x"38",
          1517 => x"81",
          1518 => x"14",
          1519 => x"77",
          1520 => x"db",
          1521 => x"80",
          1522 => x"27",
          1523 => x"80",
          1524 => x"89",
          1525 => x"70",
          1526 => x"55",
          1527 => x"70",
          1528 => x"51",
          1529 => x"27",
          1530 => x"13",
          1531 => x"06",
          1532 => x"73",
          1533 => x"38",
          1534 => x"81",
          1535 => x"76",
          1536 => x"16",
          1537 => x"70",
          1538 => x"56",
          1539 => x"ff",
          1540 => x"80",
          1541 => x"75",
          1542 => x"7a",
          1543 => x"75",
          1544 => x"0c",
          1545 => x"04",
          1546 => x"70",
          1547 => x"33",
          1548 => x"73",
          1549 => x"81",
          1550 => x"38",
          1551 => x"78",
          1552 => x"55",
          1553 => x"e2",
          1554 => x"90",
          1555 => x"f8",
          1556 => x"81",
          1557 => x"27",
          1558 => x"14",
          1559 => x"88",
          1560 => x"27",
          1561 => x"75",
          1562 => x"0c",
          1563 => x"04",
          1564 => x"15",
          1565 => x"70",
          1566 => x"80",
          1567 => x"39",
          1568 => x"ba",
          1569 => x"3d",
          1570 => x"d6",
          1571 => x"ba",
          1572 => x"ff",
          1573 => x"8c",
          1574 => x"3d",
          1575 => x"71",
          1576 => x"38",
          1577 => x"83",
          1578 => x"52",
          1579 => x"83",
          1580 => x"ef",
          1581 => x"3d",
          1582 => x"ce",
          1583 => x"b3",
          1584 => x"0d",
          1585 => x"8c",
          1586 => x"3f",
          1587 => x"04",
          1588 => x"51",
          1589 => x"83",
          1590 => x"83",
          1591 => x"ef",
          1592 => x"3d",
          1593 => x"cf",
          1594 => x"87",
          1595 => x"0d",
          1596 => x"ec",
          1597 => x"3f",
          1598 => x"04",
          1599 => x"51",
          1600 => x"83",
          1601 => x"83",
          1602 => x"ee",
          1603 => x"3d",
          1604 => x"d0",
          1605 => x"db",
          1606 => x"0d",
          1607 => x"d4",
          1608 => x"3f",
          1609 => x"04",
          1610 => x"51",
          1611 => x"83",
          1612 => x"83",
          1613 => x"ee",
          1614 => x"3d",
          1615 => x"d1",
          1616 => x"af",
          1617 => x"0d",
          1618 => x"ac",
          1619 => x"3f",
          1620 => x"04",
          1621 => x"51",
          1622 => x"83",
          1623 => x"83",
          1624 => x"ee",
          1625 => x"3d",
          1626 => x"d1",
          1627 => x"83",
          1628 => x"0d",
          1629 => x"f0",
          1630 => x"3f",
          1631 => x"04",
          1632 => x"51",
          1633 => x"83",
          1634 => x"83",
          1635 => x"ed",
          1636 => x"3d",
          1637 => x"3d",
          1638 => x"84",
          1639 => x"05",
          1640 => x"80",
          1641 => x"70",
          1642 => x"25",
          1643 => x"59",
          1644 => x"87",
          1645 => x"38",
          1646 => x"77",
          1647 => x"ff",
          1648 => x"93",
          1649 => x"e2",
          1650 => x"77",
          1651 => x"70",
          1652 => x"96",
          1653 => x"ba",
          1654 => x"84",
          1655 => x"80",
          1656 => x"38",
          1657 => x"af",
          1658 => x"30",
          1659 => x"80",
          1660 => x"70",
          1661 => x"06",
          1662 => x"58",
          1663 => x"aa",
          1664 => x"98",
          1665 => x"74",
          1666 => x"80",
          1667 => x"52",
          1668 => x"29",
          1669 => x"3f",
          1670 => x"08",
          1671 => x"bc",
          1672 => x"83",
          1673 => x"df",
          1674 => x"84",
          1675 => x"96",
          1676 => x"84",
          1677 => x"87",
          1678 => x"0c",
          1679 => x"08",
          1680 => x"d4",
          1681 => x"80",
          1682 => x"77",
          1683 => x"97",
          1684 => x"8c",
          1685 => x"ba",
          1686 => x"88",
          1687 => x"74",
          1688 => x"80",
          1689 => x"75",
          1690 => x"d5",
          1691 => x"52",
          1692 => x"b1",
          1693 => x"8c",
          1694 => x"51",
          1695 => x"84",
          1696 => x"54",
          1697 => x"53",
          1698 => x"d2",
          1699 => x"f8",
          1700 => x"39",
          1701 => x"7c",
          1702 => x"b7",
          1703 => x"59",
          1704 => x"53",
          1705 => x"51",
          1706 => x"84",
          1707 => x"8b",
          1708 => x"2e",
          1709 => x"81",
          1710 => x"77",
          1711 => x"0c",
          1712 => x"04",
          1713 => x"d5",
          1714 => x"55",
          1715 => x"ba",
          1716 => x"52",
          1717 => x"2d",
          1718 => x"08",
          1719 => x"0c",
          1720 => x"04",
          1721 => x"7f",
          1722 => x"8c",
          1723 => x"05",
          1724 => x"15",
          1725 => x"5c",
          1726 => x"5e",
          1727 => x"83",
          1728 => x"52",
          1729 => x"51",
          1730 => x"83",
          1731 => x"dd",
          1732 => x"54",
          1733 => x"b2",
          1734 => x"2e",
          1735 => x"7c",
          1736 => x"a8",
          1737 => x"53",
          1738 => x"81",
          1739 => x"33",
          1740 => x"d0",
          1741 => x"3f",
          1742 => x"d5",
          1743 => x"54",
          1744 => x"aa",
          1745 => x"26",
          1746 => x"d2",
          1747 => x"b8",
          1748 => x"75",
          1749 => x"c0",
          1750 => x"70",
          1751 => x"80",
          1752 => x"27",
          1753 => x"55",
          1754 => x"74",
          1755 => x"81",
          1756 => x"06",
          1757 => x"06",
          1758 => x"80",
          1759 => x"80",
          1760 => x"81",
          1761 => x"d5",
          1762 => x"a0",
          1763 => x"3f",
          1764 => x"78",
          1765 => x"38",
          1766 => x"51",
          1767 => x"78",
          1768 => x"5c",
          1769 => x"9d",
          1770 => x"ba",
          1771 => x"2b",
          1772 => x"58",
          1773 => x"2e",
          1774 => x"76",
          1775 => x"c3",
          1776 => x"57",
          1777 => x"fe",
          1778 => x"0b",
          1779 => x"0c",
          1780 => x"04",
          1781 => x"51",
          1782 => x"81",
          1783 => x"f0",
          1784 => x"a0",
          1785 => x"3f",
          1786 => x"fe",
          1787 => x"da",
          1788 => x"f0",
          1789 => x"3f",
          1790 => x"d5",
          1791 => x"54",
          1792 => x"ea",
          1793 => x"27",
          1794 => x"73",
          1795 => x"7a",
          1796 => x"72",
          1797 => x"d2",
          1798 => x"ec",
          1799 => x"84",
          1800 => x"53",
          1801 => x"ea",
          1802 => x"74",
          1803 => x"fe",
          1804 => x"d2",
          1805 => x"d0",
          1806 => x"84",
          1807 => x"53",
          1808 => x"ea",
          1809 => x"79",
          1810 => x"38",
          1811 => x"72",
          1812 => x"38",
          1813 => x"83",
          1814 => x"db",
          1815 => x"14",
          1816 => x"08",
          1817 => x"51",
          1818 => x"78",
          1819 => x"38",
          1820 => x"84",
          1821 => x"52",
          1822 => x"f2",
          1823 => x"56",
          1824 => x"80",
          1825 => x"84",
          1826 => x"81",
          1827 => x"88",
          1828 => x"2e",
          1829 => x"a0",
          1830 => x"d0",
          1831 => x"06",
          1832 => x"90",
          1833 => x"39",
          1834 => x"af",
          1835 => x"8c",
          1836 => x"70",
          1837 => x"a0",
          1838 => x"72",
          1839 => x"30",
          1840 => x"73",
          1841 => x"51",
          1842 => x"57",
          1843 => x"80",
          1844 => x"38",
          1845 => x"83",
          1846 => x"8c",
          1847 => x"70",
          1848 => x"a0",
          1849 => x"72",
          1850 => x"30",
          1851 => x"73",
          1852 => x"51",
          1853 => x"57",
          1854 => x"73",
          1855 => x"38",
          1856 => x"80",
          1857 => x"8c",
          1858 => x"0d",
          1859 => x"0d",
          1860 => x"80",
          1861 => x"d1",
          1862 => x"9c",
          1863 => x"d3",
          1864 => x"88",
          1865 => x"9c",
          1866 => x"81",
          1867 => x"06",
          1868 => x"82",
          1869 => x"82",
          1870 => x"06",
          1871 => x"82",
          1872 => x"83",
          1873 => x"06",
          1874 => x"81",
          1875 => x"84",
          1876 => x"06",
          1877 => x"81",
          1878 => x"85",
          1879 => x"06",
          1880 => x"80",
          1881 => x"86",
          1882 => x"06",
          1883 => x"80",
          1884 => x"87",
          1885 => x"06",
          1886 => x"a9",
          1887 => x"2a",
          1888 => x"72",
          1889 => x"e9",
          1890 => x"0d",
          1891 => x"9c",
          1892 => x"d3",
          1893 => x"94",
          1894 => x"9b",
          1895 => x"d1",
          1896 => x"0d",
          1897 => x"9b",
          1898 => x"d3",
          1899 => x"fc",
          1900 => x"9b",
          1901 => x"88",
          1902 => x"53",
          1903 => x"c6",
          1904 => x"81",
          1905 => x"3f",
          1906 => x"51",
          1907 => x"80",
          1908 => x"3f",
          1909 => x"70",
          1910 => x"52",
          1911 => x"ff",
          1912 => x"39",
          1913 => x"ac",
          1914 => x"88",
          1915 => x"3f",
          1916 => x"a0",
          1917 => x"2a",
          1918 => x"51",
          1919 => x"2e",
          1920 => x"ff",
          1921 => x"51",
          1922 => x"83",
          1923 => x"9b",
          1924 => x"51",
          1925 => x"72",
          1926 => x"81",
          1927 => x"71",
          1928 => x"c2",
          1929 => x"39",
          1930 => x"e8",
          1931 => x"b0",
          1932 => x"3f",
          1933 => x"dc",
          1934 => x"2a",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"ff",
          1938 => x"51",
          1939 => x"83",
          1940 => x"9a",
          1941 => x"51",
          1942 => x"72",
          1943 => x"81",
          1944 => x"71",
          1945 => x"e6",
          1946 => x"39",
          1947 => x"a4",
          1948 => x"d4",
          1949 => x"3f",
          1950 => x"98",
          1951 => x"2a",
          1952 => x"51",
          1953 => x"2e",
          1954 => x"ff",
          1955 => x"3d",
          1956 => x"41",
          1957 => x"84",
          1958 => x"42",
          1959 => x"51",
          1960 => x"3f",
          1961 => x"08",
          1962 => x"9b",
          1963 => x"78",
          1964 => x"b1",
          1965 => x"a8",
          1966 => x"3f",
          1967 => x"83",
          1968 => x"d6",
          1969 => x"48",
          1970 => x"80",
          1971 => x"eb",
          1972 => x"0b",
          1973 => x"33",
          1974 => x"06",
          1975 => x"80",
          1976 => x"38",
          1977 => x"83",
          1978 => x"81",
          1979 => x"7d",
          1980 => x"c1",
          1981 => x"5a",
          1982 => x"2e",
          1983 => x"79",
          1984 => x"a0",
          1985 => x"06",
          1986 => x"1a",
          1987 => x"5a",
          1988 => x"f6",
          1989 => x"7b",
          1990 => x"38",
          1991 => x"83",
          1992 => x"70",
          1993 => x"e7",
          1994 => x"ba",
          1995 => x"ba",
          1996 => x"7a",
          1997 => x"52",
          1998 => x"3f",
          1999 => x"08",
          2000 => x"1b",
          2001 => x"81",
          2002 => x"38",
          2003 => x"81",
          2004 => x"5b",
          2005 => x"c4",
          2006 => x"33",
          2007 => x"2e",
          2008 => x"80",
          2009 => x"51",
          2010 => x"84",
          2011 => x"5e",
          2012 => x"08",
          2013 => x"d3",
          2014 => x"8c",
          2015 => x"3d",
          2016 => x"51",
          2017 => x"84",
          2018 => x"60",
          2019 => x"5c",
          2020 => x"81",
          2021 => x"ba",
          2022 => x"e7",
          2023 => x"ba",
          2024 => x"26",
          2025 => x"81",
          2026 => x"5e",
          2027 => x"2e",
          2028 => x"7a",
          2029 => x"ec",
          2030 => x"2e",
          2031 => x"7b",
          2032 => x"83",
          2033 => x"7c",
          2034 => x"3f",
          2035 => x"58",
          2036 => x"57",
          2037 => x"55",
          2038 => x"80",
          2039 => x"80",
          2040 => x"51",
          2041 => x"84",
          2042 => x"84",
          2043 => x"09",
          2044 => x"72",
          2045 => x"51",
          2046 => x"80",
          2047 => x"26",
          2048 => x"5a",
          2049 => x"59",
          2050 => x"8d",
          2051 => x"70",
          2052 => x"5c",
          2053 => x"95",
          2054 => x"32",
          2055 => x"07",
          2056 => x"f8",
          2057 => x"2e",
          2058 => x"7d",
          2059 => x"aa",
          2060 => x"e0",
          2061 => x"3f",
          2062 => x"f8",
          2063 => x"7e",
          2064 => x"3f",
          2065 => x"ef",
          2066 => x"81",
          2067 => x"59",
          2068 => x"38",
          2069 => x"d5",
          2070 => x"d1",
          2071 => x"89",
          2072 => x"ba",
          2073 => x"c5",
          2074 => x"0b",
          2075 => x"80",
          2076 => x"9c",
          2077 => x"52",
          2078 => x"f7",
          2079 => x"ba",
          2080 => x"2e",
          2081 => x"ba",
          2082 => x"df",
          2083 => x"0b",
          2084 => x"33",
          2085 => x"06",
          2086 => x"82",
          2087 => x"06",
          2088 => x"91",
          2089 => x"9c",
          2090 => x"9d",
          2091 => x"0b",
          2092 => x"80",
          2093 => x"9c",
          2094 => x"52",
          2095 => x"ce",
          2096 => x"5a",
          2097 => x"b7",
          2098 => x"7c",
          2099 => x"85",
          2100 => x"78",
          2101 => x"fd",
          2102 => x"10",
          2103 => x"9c",
          2104 => x"08",
          2105 => x"ec",
          2106 => x"3f",
          2107 => x"83",
          2108 => x"80",
          2109 => x"e4",
          2110 => x"53",
          2111 => x"bb",
          2112 => x"85",
          2113 => x"ba",
          2114 => x"2e",
          2115 => x"fb",
          2116 => x"70",
          2117 => x"41",
          2118 => x"39",
          2119 => x"51",
          2120 => x"7d",
          2121 => x"b2",
          2122 => x"39",
          2123 => x"56",
          2124 => x"d6",
          2125 => x"53",
          2126 => x"52",
          2127 => x"e8",
          2128 => x"39",
          2129 => x"3f",
          2130 => x"9a",
          2131 => x"ef",
          2132 => x"83",
          2133 => x"3f",
          2134 => x"81",
          2135 => x"fa",
          2136 => x"d6",
          2137 => x"8b",
          2138 => x"78",
          2139 => x"c0",
          2140 => x"3f",
          2141 => x"fa",
          2142 => x"3d",
          2143 => x"53",
          2144 => x"51",
          2145 => x"84",
          2146 => x"80",
          2147 => x"38",
          2148 => x"d6",
          2149 => x"f0",
          2150 => x"79",
          2151 => x"8c",
          2152 => x"fa",
          2153 => x"ba",
          2154 => x"83",
          2155 => x"d0",
          2156 => x"8b",
          2157 => x"ff",
          2158 => x"ff",
          2159 => x"eb",
          2160 => x"ba",
          2161 => x"2e",
          2162 => x"68",
          2163 => x"94",
          2164 => x"3f",
          2165 => x"04",
          2166 => x"f4",
          2167 => x"80",
          2168 => x"9e",
          2169 => x"8c",
          2170 => x"f9",
          2171 => x"3d",
          2172 => x"53",
          2173 => x"51",
          2174 => x"84",
          2175 => x"86",
          2176 => x"59",
          2177 => x"78",
          2178 => x"b0",
          2179 => x"3f",
          2180 => x"08",
          2181 => x"52",
          2182 => x"87",
          2183 => x"7e",
          2184 => x"ae",
          2185 => x"38",
          2186 => x"87",
          2187 => x"84",
          2188 => x"59",
          2189 => x"3d",
          2190 => x"53",
          2191 => x"51",
          2192 => x"84",
          2193 => x"80",
          2194 => x"38",
          2195 => x"f0",
          2196 => x"80",
          2197 => x"aa",
          2198 => x"8c",
          2199 => x"38",
          2200 => x"22",
          2201 => x"83",
          2202 => x"cf",
          2203 => x"d5",
          2204 => x"80",
          2205 => x"51",
          2206 => x"7e",
          2207 => x"59",
          2208 => x"f8",
          2209 => x"9f",
          2210 => x"38",
          2211 => x"70",
          2212 => x"39",
          2213 => x"84",
          2214 => x"80",
          2215 => x"e6",
          2216 => x"8c",
          2217 => x"f8",
          2218 => x"3d",
          2219 => x"53",
          2220 => x"51",
          2221 => x"84",
          2222 => x"80",
          2223 => x"38",
          2224 => x"f8",
          2225 => x"80",
          2226 => x"ba",
          2227 => x"8c",
          2228 => x"f7",
          2229 => x"d7",
          2230 => x"ac",
          2231 => x"5d",
          2232 => x"27",
          2233 => x"65",
          2234 => x"33",
          2235 => x"7a",
          2236 => x"38",
          2237 => x"54",
          2238 => x"78",
          2239 => x"dc",
          2240 => x"3f",
          2241 => x"5c",
          2242 => x"1b",
          2243 => x"39",
          2244 => x"84",
          2245 => x"80",
          2246 => x"ea",
          2247 => x"8c",
          2248 => x"f7",
          2249 => x"3d",
          2250 => x"53",
          2251 => x"51",
          2252 => x"84",
          2253 => x"80",
          2254 => x"38",
          2255 => x"f8",
          2256 => x"80",
          2257 => x"be",
          2258 => x"8c",
          2259 => x"f6",
          2260 => x"d7",
          2261 => x"b0",
          2262 => x"79",
          2263 => x"93",
          2264 => x"79",
          2265 => x"5b",
          2266 => x"65",
          2267 => x"eb",
          2268 => x"ff",
          2269 => x"ff",
          2270 => x"e8",
          2271 => x"ba",
          2272 => x"2e",
          2273 => x"b8",
          2274 => x"11",
          2275 => x"05",
          2276 => x"3f",
          2277 => x"08",
          2278 => x"70",
          2279 => x"83",
          2280 => x"cc",
          2281 => x"d5",
          2282 => x"80",
          2283 => x"51",
          2284 => x"7e",
          2285 => x"59",
          2286 => x"f6",
          2287 => x"9f",
          2288 => x"38",
          2289 => x"49",
          2290 => x"59",
          2291 => x"05",
          2292 => x"68",
          2293 => x"b8",
          2294 => x"11",
          2295 => x"05",
          2296 => x"3f",
          2297 => x"08",
          2298 => x"d3",
          2299 => x"02",
          2300 => x"33",
          2301 => x"81",
          2302 => x"3d",
          2303 => x"53",
          2304 => x"51",
          2305 => x"84",
          2306 => x"ff",
          2307 => x"af",
          2308 => x"ff",
          2309 => x"ff",
          2310 => x"e6",
          2311 => x"ba",
          2312 => x"2e",
          2313 => x"b8",
          2314 => x"11",
          2315 => x"05",
          2316 => x"3f",
          2317 => x"08",
          2318 => x"83",
          2319 => x"fe",
          2320 => x"ff",
          2321 => x"e6",
          2322 => x"ba",
          2323 => x"38",
          2324 => x"08",
          2325 => x"90",
          2326 => x"3f",
          2327 => x"59",
          2328 => x"8f",
          2329 => x"7a",
          2330 => x"05",
          2331 => x"79",
          2332 => x"8a",
          2333 => x"3f",
          2334 => x"b8",
          2335 => x"05",
          2336 => x"3f",
          2337 => x"08",
          2338 => x"80",
          2339 => x"88",
          2340 => x"53",
          2341 => x"08",
          2342 => x"e9",
          2343 => x"ba",
          2344 => x"2e",
          2345 => x"84",
          2346 => x"51",
          2347 => x"f4",
          2348 => x"3d",
          2349 => x"53",
          2350 => x"51",
          2351 => x"84",
          2352 => x"91",
          2353 => x"90",
          2354 => x"80",
          2355 => x"38",
          2356 => x"08",
          2357 => x"fe",
          2358 => x"ff",
          2359 => x"e5",
          2360 => x"ba",
          2361 => x"38",
          2362 => x"33",
          2363 => x"2e",
          2364 => x"83",
          2365 => x"47",
          2366 => x"f8",
          2367 => x"80",
          2368 => x"82",
          2369 => x"8c",
          2370 => x"a5",
          2371 => x"5c",
          2372 => x"2e",
          2373 => x"5c",
          2374 => x"70",
          2375 => x"07",
          2376 => x"06",
          2377 => x"79",
          2378 => x"38",
          2379 => x"83",
          2380 => x"83",
          2381 => x"d6",
          2382 => x"55",
          2383 => x"53",
          2384 => x"51",
          2385 => x"83",
          2386 => x"d6",
          2387 => x"ef",
          2388 => x"71",
          2389 => x"84",
          2390 => x"3d",
          2391 => x"53",
          2392 => x"51",
          2393 => x"84",
          2394 => x"80",
          2395 => x"38",
          2396 => x"0c",
          2397 => x"05",
          2398 => x"fe",
          2399 => x"ff",
          2400 => x"e1",
          2401 => x"ba",
          2402 => x"38",
          2403 => x"64",
          2404 => x"ce",
          2405 => x"70",
          2406 => x"23",
          2407 => x"3d",
          2408 => x"53",
          2409 => x"51",
          2410 => x"84",
          2411 => x"80",
          2412 => x"38",
          2413 => x"80",
          2414 => x"7e",
          2415 => x"40",
          2416 => x"b8",
          2417 => x"11",
          2418 => x"05",
          2419 => x"3f",
          2420 => x"08",
          2421 => x"f1",
          2422 => x"3d",
          2423 => x"53",
          2424 => x"51",
          2425 => x"84",
          2426 => x"80",
          2427 => x"38",
          2428 => x"80",
          2429 => x"7c",
          2430 => x"05",
          2431 => x"39",
          2432 => x"f0",
          2433 => x"80",
          2434 => x"f6",
          2435 => x"8c",
          2436 => x"81",
          2437 => x"64",
          2438 => x"64",
          2439 => x"46",
          2440 => x"39",
          2441 => x"09",
          2442 => x"93",
          2443 => x"83",
          2444 => x"80",
          2445 => x"b8",
          2446 => x"c8",
          2447 => x"8c",
          2448 => x"7c",
          2449 => x"3f",
          2450 => x"83",
          2451 => x"d4",
          2452 => x"eb",
          2453 => x"fe",
          2454 => x"ff",
          2455 => x"e0",
          2456 => x"ba",
          2457 => x"2e",
          2458 => x"59",
          2459 => x"05",
          2460 => x"82",
          2461 => x"78",
          2462 => x"39",
          2463 => x"33",
          2464 => x"2e",
          2465 => x"83",
          2466 => x"47",
          2467 => x"83",
          2468 => x"5c",
          2469 => x"a1",
          2470 => x"d0",
          2471 => x"b5",
          2472 => x"f0",
          2473 => x"3f",
          2474 => x"b6",
          2475 => x"f0",
          2476 => x"3f",
          2477 => x"cc",
          2478 => x"92",
          2479 => x"80",
          2480 => x"83",
          2481 => x"49",
          2482 => x"83",
          2483 => x"d3",
          2484 => x"c6",
          2485 => x"92",
          2486 => x"80",
          2487 => x"83",
          2488 => x"47",
          2489 => x"83",
          2490 => x"5e",
          2491 => x"9b",
          2492 => x"e0",
          2493 => x"dd",
          2494 => x"93",
          2495 => x"80",
          2496 => x"83",
          2497 => x"47",
          2498 => x"83",
          2499 => x"5d",
          2500 => x"9b",
          2501 => x"e8",
          2502 => x"b9",
          2503 => x"8e",
          2504 => x"80",
          2505 => x"83",
          2506 => x"47",
          2507 => x"83",
          2508 => x"fc",
          2509 => x"fb",
          2510 => x"f2",
          2511 => x"05",
          2512 => x"39",
          2513 => x"80",
          2514 => x"bc",
          2515 => x"94",
          2516 => x"56",
          2517 => x"80",
          2518 => x"da",
          2519 => x"ba",
          2520 => x"2b",
          2521 => x"55",
          2522 => x"52",
          2523 => x"b5",
          2524 => x"ba",
          2525 => x"77",
          2526 => x"94",
          2527 => x"56",
          2528 => x"80",
          2529 => x"da",
          2530 => x"ba",
          2531 => x"2b",
          2532 => x"55",
          2533 => x"52",
          2534 => x"89",
          2535 => x"ba",
          2536 => x"77",
          2537 => x"83",
          2538 => x"94",
          2539 => x"80",
          2540 => x"c0",
          2541 => x"81",
          2542 => x"81",
          2543 => x"83",
          2544 => x"a1",
          2545 => x"5e",
          2546 => x"0b",
          2547 => x"88",
          2548 => x"72",
          2549 => x"f0",
          2550 => x"f5",
          2551 => x"3f",
          2552 => x"ba",
          2553 => x"fc",
          2554 => x"f8",
          2555 => x"fc",
          2556 => x"3f",
          2557 => x"70",
          2558 => x"94",
          2559 => x"d3",
          2560 => x"d3",
          2561 => x"15",
          2562 => x"d3",
          2563 => x"f8",
          2564 => x"3f",
          2565 => x"80",
          2566 => x"0d",
          2567 => x"56",
          2568 => x"52",
          2569 => x"2e",
          2570 => x"74",
          2571 => x"ff",
          2572 => x"70",
          2573 => x"81",
          2574 => x"81",
          2575 => x"70",
          2576 => x"53",
          2577 => x"a0",
          2578 => x"71",
          2579 => x"54",
          2580 => x"81",
          2581 => x"52",
          2582 => x"80",
          2583 => x"72",
          2584 => x"ff",
          2585 => x"54",
          2586 => x"83",
          2587 => x"70",
          2588 => x"38",
          2589 => x"86",
          2590 => x"52",
          2591 => x"73",
          2592 => x"52",
          2593 => x"2e",
          2594 => x"83",
          2595 => x"70",
          2596 => x"30",
          2597 => x"76",
          2598 => x"53",
          2599 => x"88",
          2600 => x"70",
          2601 => x"34",
          2602 => x"74",
          2603 => x"ba",
          2604 => x"3d",
          2605 => x"80",
          2606 => x"73",
          2607 => x"be",
          2608 => x"52",
          2609 => x"70",
          2610 => x"53",
          2611 => x"a2",
          2612 => x"81",
          2613 => x"81",
          2614 => x"75",
          2615 => x"81",
          2616 => x"06",
          2617 => x"dc",
          2618 => x"0d",
          2619 => x"08",
          2620 => x"0b",
          2621 => x"0c",
          2622 => x"04",
          2623 => x"05",
          2624 => x"da",
          2625 => x"ba",
          2626 => x"2e",
          2627 => x"84",
          2628 => x"86",
          2629 => x"fc",
          2630 => x"82",
          2631 => x"05",
          2632 => x"52",
          2633 => x"81",
          2634 => x"13",
          2635 => x"54",
          2636 => x"9e",
          2637 => x"38",
          2638 => x"51",
          2639 => x"97",
          2640 => x"38",
          2641 => x"54",
          2642 => x"bb",
          2643 => x"38",
          2644 => x"55",
          2645 => x"bb",
          2646 => x"38",
          2647 => x"55",
          2648 => x"87",
          2649 => x"d9",
          2650 => x"22",
          2651 => x"73",
          2652 => x"80",
          2653 => x"0b",
          2654 => x"9c",
          2655 => x"87",
          2656 => x"0c",
          2657 => x"87",
          2658 => x"0c",
          2659 => x"87",
          2660 => x"0c",
          2661 => x"87",
          2662 => x"0c",
          2663 => x"87",
          2664 => x"0c",
          2665 => x"87",
          2666 => x"0c",
          2667 => x"98",
          2668 => x"87",
          2669 => x"0c",
          2670 => x"c0",
          2671 => x"80",
          2672 => x"ba",
          2673 => x"3d",
          2674 => x"3d",
          2675 => x"87",
          2676 => x"5d",
          2677 => x"87",
          2678 => x"08",
          2679 => x"23",
          2680 => x"b8",
          2681 => x"82",
          2682 => x"c0",
          2683 => x"5a",
          2684 => x"34",
          2685 => x"b0",
          2686 => x"84",
          2687 => x"c0",
          2688 => x"5a",
          2689 => x"34",
          2690 => x"a8",
          2691 => x"86",
          2692 => x"c0",
          2693 => x"5c",
          2694 => x"23",
          2695 => x"a0",
          2696 => x"8a",
          2697 => x"7d",
          2698 => x"ff",
          2699 => x"7b",
          2700 => x"06",
          2701 => x"33",
          2702 => x"33",
          2703 => x"33",
          2704 => x"33",
          2705 => x"33",
          2706 => x"ff",
          2707 => x"83",
          2708 => x"ff",
          2709 => x"8f",
          2710 => x"fe",
          2711 => x"93",
          2712 => x"72",
          2713 => x"38",
          2714 => x"e8",
          2715 => x"ba",
          2716 => x"2b",
          2717 => x"51",
          2718 => x"2e",
          2719 => x"86",
          2720 => x"2e",
          2721 => x"84",
          2722 => x"84",
          2723 => x"72",
          2724 => x"8a",
          2725 => x"8c",
          2726 => x"70",
          2727 => x"52",
          2728 => x"09",
          2729 => x"38",
          2730 => x"e7",
          2731 => x"ba",
          2732 => x"2b",
          2733 => x"51",
          2734 => x"2e",
          2735 => x"39",
          2736 => x"80",
          2737 => x"71",
          2738 => x"81",
          2739 => x"ce",
          2740 => x"8c",
          2741 => x"70",
          2742 => x"52",
          2743 => x"eb",
          2744 => x"07",
          2745 => x"52",
          2746 => x"db",
          2747 => x"ba",
          2748 => x"3d",
          2749 => x"3d",
          2750 => x"05",
          2751 => x"c4",
          2752 => x"ff",
          2753 => x"55",
          2754 => x"80",
          2755 => x"c0",
          2756 => x"70",
          2757 => x"81",
          2758 => x"52",
          2759 => x"8c",
          2760 => x"2a",
          2761 => x"51",
          2762 => x"38",
          2763 => x"81",
          2764 => x"80",
          2765 => x"71",
          2766 => x"06",
          2767 => x"38",
          2768 => x"06",
          2769 => x"94",
          2770 => x"80",
          2771 => x"87",
          2772 => x"52",
          2773 => x"74",
          2774 => x"0c",
          2775 => x"04",
          2776 => x"70",
          2777 => x"51",
          2778 => x"72",
          2779 => x"06",
          2780 => x"2e",
          2781 => x"93",
          2782 => x"52",
          2783 => x"c0",
          2784 => x"94",
          2785 => x"96",
          2786 => x"06",
          2787 => x"70",
          2788 => x"39",
          2789 => x"02",
          2790 => x"70",
          2791 => x"2a",
          2792 => x"70",
          2793 => x"34",
          2794 => x"04",
          2795 => x"78",
          2796 => x"33",
          2797 => x"57",
          2798 => x"80",
          2799 => x"15",
          2800 => x"33",
          2801 => x"06",
          2802 => x"71",
          2803 => x"ff",
          2804 => x"94",
          2805 => x"96",
          2806 => x"06",
          2807 => x"70",
          2808 => x"38",
          2809 => x"70",
          2810 => x"51",
          2811 => x"72",
          2812 => x"06",
          2813 => x"2e",
          2814 => x"93",
          2815 => x"52",
          2816 => x"75",
          2817 => x"51",
          2818 => x"80",
          2819 => x"2e",
          2820 => x"c0",
          2821 => x"73",
          2822 => x"17",
          2823 => x"57",
          2824 => x"38",
          2825 => x"8c",
          2826 => x"0d",
          2827 => x"2a",
          2828 => x"51",
          2829 => x"38",
          2830 => x"81",
          2831 => x"80",
          2832 => x"71",
          2833 => x"06",
          2834 => x"2e",
          2835 => x"87",
          2836 => x"08",
          2837 => x"70",
          2838 => x"54",
          2839 => x"38",
          2840 => x"3d",
          2841 => x"9e",
          2842 => x"9c",
          2843 => x"52",
          2844 => x"2e",
          2845 => x"87",
          2846 => x"08",
          2847 => x"0c",
          2848 => x"a8",
          2849 => x"cc",
          2850 => x"9e",
          2851 => x"f2",
          2852 => x"c0",
          2853 => x"83",
          2854 => x"87",
          2855 => x"08",
          2856 => x"0c",
          2857 => x"a0",
          2858 => x"dc",
          2859 => x"9e",
          2860 => x"f2",
          2861 => x"c0",
          2862 => x"83",
          2863 => x"87",
          2864 => x"08",
          2865 => x"0c",
          2866 => x"b8",
          2867 => x"ec",
          2868 => x"9e",
          2869 => x"f2",
          2870 => x"c0",
          2871 => x"83",
          2872 => x"87",
          2873 => x"08",
          2874 => x"0c",
          2875 => x"80",
          2876 => x"83",
          2877 => x"87",
          2878 => x"08",
          2879 => x"0c",
          2880 => x"88",
          2881 => x"84",
          2882 => x"9e",
          2883 => x"f3",
          2884 => x"0b",
          2885 => x"34",
          2886 => x"c0",
          2887 => x"70",
          2888 => x"06",
          2889 => x"70",
          2890 => x"71",
          2891 => x"34",
          2892 => x"c0",
          2893 => x"70",
          2894 => x"06",
          2895 => x"70",
          2896 => x"38",
          2897 => x"83",
          2898 => x"80",
          2899 => x"9e",
          2900 => x"90",
          2901 => x"51",
          2902 => x"80",
          2903 => x"81",
          2904 => x"f3",
          2905 => x"0b",
          2906 => x"90",
          2907 => x"80",
          2908 => x"52",
          2909 => x"2e",
          2910 => x"52",
          2911 => x"90",
          2912 => x"87",
          2913 => x"08",
          2914 => x"80",
          2915 => x"52",
          2916 => x"83",
          2917 => x"71",
          2918 => x"34",
          2919 => x"c0",
          2920 => x"70",
          2921 => x"06",
          2922 => x"70",
          2923 => x"38",
          2924 => x"83",
          2925 => x"80",
          2926 => x"9e",
          2927 => x"84",
          2928 => x"51",
          2929 => x"80",
          2930 => x"81",
          2931 => x"f3",
          2932 => x"0b",
          2933 => x"90",
          2934 => x"80",
          2935 => x"52",
          2936 => x"2e",
          2937 => x"52",
          2938 => x"94",
          2939 => x"87",
          2940 => x"08",
          2941 => x"80",
          2942 => x"52",
          2943 => x"83",
          2944 => x"71",
          2945 => x"34",
          2946 => x"c0",
          2947 => x"70",
          2948 => x"06",
          2949 => x"70",
          2950 => x"38",
          2951 => x"83",
          2952 => x"80",
          2953 => x"9e",
          2954 => x"a0",
          2955 => x"52",
          2956 => x"2e",
          2957 => x"52",
          2958 => x"97",
          2959 => x"9e",
          2960 => x"80",
          2961 => x"2a",
          2962 => x"83",
          2963 => x"80",
          2964 => x"9e",
          2965 => x"84",
          2966 => x"52",
          2967 => x"2e",
          2968 => x"52",
          2969 => x"99",
          2970 => x"9e",
          2971 => x"f0",
          2972 => x"2a",
          2973 => x"83",
          2974 => x"80",
          2975 => x"9e",
          2976 => x"88",
          2977 => x"52",
          2978 => x"83",
          2979 => x"71",
          2980 => x"34",
          2981 => x"90",
          2982 => x"51",
          2983 => x"9c",
          2984 => x"0d",
          2985 => x"fd",
          2986 => x"3d",
          2987 => x"8c",
          2988 => x"d4",
          2989 => x"8c",
          2990 => x"86",
          2991 => x"d9",
          2992 => x"af",
          2993 => x"8e",
          2994 => x"85",
          2995 => x"f3",
          2996 => x"73",
          2997 => x"83",
          2998 => x"56",
          2999 => x"38",
          3000 => x"33",
          3001 => x"ff",
          3002 => x"92",
          3003 => x"84",
          3004 => x"f3",
          3005 => x"75",
          3006 => x"83",
          3007 => x"54",
          3008 => x"38",
          3009 => x"33",
          3010 => x"ed",
          3011 => x"8d",
          3012 => x"83",
          3013 => x"f3",
          3014 => x"73",
          3015 => x"83",
          3016 => x"55",
          3017 => x"38",
          3018 => x"33",
          3019 => x"f4",
          3020 => x"96",
          3021 => x"81",
          3022 => x"d9",
          3023 => x"b3",
          3024 => x"f0",
          3025 => x"d9",
          3026 => x"b5",
          3027 => x"f2",
          3028 => x"83",
          3029 => x"ff",
          3030 => x"83",
          3031 => x"52",
          3032 => x"51",
          3033 => x"3f",
          3034 => x"51",
          3035 => x"83",
          3036 => x"52",
          3037 => x"51",
          3038 => x"3f",
          3039 => x"08",
          3040 => x"c0",
          3041 => x"ca",
          3042 => x"ba",
          3043 => x"84",
          3044 => x"71",
          3045 => x"84",
          3046 => x"52",
          3047 => x"51",
          3048 => x"3f",
          3049 => x"33",
          3050 => x"c3",
          3051 => x"8e",
          3052 => x"8a",
          3053 => x"c3",
          3054 => x"3d",
          3055 => x"f3",
          3056 => x"bd",
          3057 => x"75",
          3058 => x"3f",
          3059 => x"08",
          3060 => x"29",
          3061 => x"54",
          3062 => x"8c",
          3063 => x"db",
          3064 => x"b4",
          3065 => x"51",
          3066 => x"87",
          3067 => x"83",
          3068 => x"56",
          3069 => x"52",
          3070 => x"a9",
          3071 => x"8c",
          3072 => x"c0",
          3073 => x"31",
          3074 => x"ba",
          3075 => x"83",
          3076 => x"ff",
          3077 => x"83",
          3078 => x"55",
          3079 => x"ff",
          3080 => x"9a",
          3081 => x"f0",
          3082 => x"3f",
          3083 => x"51",
          3084 => x"83",
          3085 => x"52",
          3086 => x"51",
          3087 => x"3f",
          3088 => x"08",
          3089 => x"ec",
          3090 => x"bc",
          3091 => x"f8",
          3092 => x"da",
          3093 => x"b3",
          3094 => x"da",
          3095 => x"93",
          3096 => x"fc",
          3097 => x"da",
          3098 => x"b3",
          3099 => x"f3",
          3100 => x"bd",
          3101 => x"75",
          3102 => x"3f",
          3103 => x"08",
          3104 => x"29",
          3105 => x"54",
          3106 => x"8c",
          3107 => x"da",
          3108 => x"b2",
          3109 => x"f3",
          3110 => x"74",
          3111 => x"8d",
          3112 => x"39",
          3113 => x"51",
          3114 => x"3f",
          3115 => x"33",
          3116 => x"2e",
          3117 => x"fe",
          3118 => x"dc",
          3119 => x"bf",
          3120 => x"f3",
          3121 => x"75",
          3122 => x"e5",
          3123 => x"83",
          3124 => x"ff",
          3125 => x"83",
          3126 => x"55",
          3127 => x"fc",
          3128 => x"39",
          3129 => x"51",
          3130 => x"3f",
          3131 => x"33",
          3132 => x"2e",
          3133 => x"d7",
          3134 => x"9a",
          3135 => x"dc",
          3136 => x"b2",
          3137 => x"f3",
          3138 => x"75",
          3139 => x"86",
          3140 => x"83",
          3141 => x"52",
          3142 => x"51",
          3143 => x"3f",
          3144 => x"33",
          3145 => x"2e",
          3146 => x"cd",
          3147 => x"98",
          3148 => x"dc",
          3149 => x"b1",
          3150 => x"f3",
          3151 => x"73",
          3152 => x"c0",
          3153 => x"83",
          3154 => x"83",
          3155 => x"11",
          3156 => x"dd",
          3157 => x"b1",
          3158 => x"f3",
          3159 => x"75",
          3160 => x"97",
          3161 => x"83",
          3162 => x"83",
          3163 => x"11",
          3164 => x"dd",
          3165 => x"b1",
          3166 => x"f3",
          3167 => x"73",
          3168 => x"ee",
          3169 => x"83",
          3170 => x"83",
          3171 => x"11",
          3172 => x"dd",
          3173 => x"b0",
          3174 => x"f3",
          3175 => x"74",
          3176 => x"c5",
          3177 => x"83",
          3178 => x"83",
          3179 => x"11",
          3180 => x"dd",
          3181 => x"b0",
          3182 => x"f3",
          3183 => x"75",
          3184 => x"9c",
          3185 => x"83",
          3186 => x"83",
          3187 => x"11",
          3188 => x"dd",
          3189 => x"b0",
          3190 => x"f3",
          3191 => x"73",
          3192 => x"f3",
          3193 => x"83",
          3194 => x"ff",
          3195 => x"83",
          3196 => x"ff",
          3197 => x"83",
          3198 => x"55",
          3199 => x"f9",
          3200 => x"39",
          3201 => x"02",
          3202 => x"52",
          3203 => x"8c",
          3204 => x"10",
          3205 => x"05",
          3206 => x"04",
          3207 => x"51",
          3208 => x"3f",
          3209 => x"04",
          3210 => x"51",
          3211 => x"3f",
          3212 => x"04",
          3213 => x"51",
          3214 => x"3f",
          3215 => x"04",
          3216 => x"51",
          3217 => x"3f",
          3218 => x"04",
          3219 => x"51",
          3220 => x"3f",
          3221 => x"04",
          3222 => x"51",
          3223 => x"3f",
          3224 => x"04",
          3225 => x"0c",
          3226 => x"87",
          3227 => x"0c",
          3228 => x"a0",
          3229 => x"96",
          3230 => x"d9",
          3231 => x"3d",
          3232 => x"08",
          3233 => x"70",
          3234 => x"52",
          3235 => x"08",
          3236 => x"d2",
          3237 => x"8c",
          3238 => x"38",
          3239 => x"ff",
          3240 => x"f8",
          3241 => x"80",
          3242 => x"51",
          3243 => x"3f",
          3244 => x"08",
          3245 => x"38",
          3246 => x"ec",
          3247 => x"8c",
          3248 => x"57",
          3249 => x"84",
          3250 => x"25",
          3251 => x"ba",
          3252 => x"05",
          3253 => x"55",
          3254 => x"74",
          3255 => x"70",
          3256 => x"2a",
          3257 => x"78",
          3258 => x"38",
          3259 => x"38",
          3260 => x"08",
          3261 => x"53",
          3262 => x"ea",
          3263 => x"8c",
          3264 => x"78",
          3265 => x"38",
          3266 => x"8c",
          3267 => x"0d",
          3268 => x"84",
          3269 => x"f0",
          3270 => x"2e",
          3271 => x"e8",
          3272 => x"79",
          3273 => x"3f",
          3274 => x"bf",
          3275 => x"3d",
          3276 => x"ba",
          3277 => x"34",
          3278 => x"e2",
          3279 => x"ad",
          3280 => x"0b",
          3281 => x"0c",
          3282 => x"04",
          3283 => x"ab",
          3284 => x"3d",
          3285 => x"5d",
          3286 => x"57",
          3287 => x"a0",
          3288 => x"38",
          3289 => x"3d",
          3290 => x"10",
          3291 => x"f4",
          3292 => x"08",
          3293 => x"bf",
          3294 => x"ba",
          3295 => x"79",
          3296 => x"51",
          3297 => x"84",
          3298 => x"90",
          3299 => x"33",
          3300 => x"2e",
          3301 => x"73",
          3302 => x"38",
          3303 => x"81",
          3304 => x"54",
          3305 => x"c2",
          3306 => x"73",
          3307 => x"0c",
          3308 => x"04",
          3309 => x"aa",
          3310 => x"11",
          3311 => x"05",
          3312 => x"3f",
          3313 => x"08",
          3314 => x"38",
          3315 => x"78",
          3316 => x"fd",
          3317 => x"ba",
          3318 => x"ff",
          3319 => x"80",
          3320 => x"81",
          3321 => x"ff",
          3322 => x"82",
          3323 => x"fa",
          3324 => x"39",
          3325 => x"05",
          3326 => x"27",
          3327 => x"81",
          3328 => x"70",
          3329 => x"73",
          3330 => x"81",
          3331 => x"38",
          3332 => x"eb",
          3333 => x"8d",
          3334 => x"fe",
          3335 => x"84",
          3336 => x"53",
          3337 => x"08",
          3338 => x"85",
          3339 => x"ba",
          3340 => x"d0",
          3341 => x"f8",
          3342 => x"f8",
          3343 => x"82",
          3344 => x"84",
          3345 => x"80",
          3346 => x"77",
          3347 => x"d8",
          3348 => x"8c",
          3349 => x"0b",
          3350 => x"08",
          3351 => x"84",
          3352 => x"ff",
          3353 => x"58",
          3354 => x"34",
          3355 => x"52",
          3356 => x"e1",
          3357 => x"ff",
          3358 => x"74",
          3359 => x"81",
          3360 => x"38",
          3361 => x"ba",
          3362 => x"3d",
          3363 => x"3d",
          3364 => x"08",
          3365 => x"b9",
          3366 => x"41",
          3367 => x"b4",
          3368 => x"f3",
          3369 => x"f3",
          3370 => x"5d",
          3371 => x"74",
          3372 => x"33",
          3373 => x"80",
          3374 => x"38",
          3375 => x"91",
          3376 => x"70",
          3377 => x"57",
          3378 => x"38",
          3379 => x"90",
          3380 => x"3d",
          3381 => x"5f",
          3382 => x"ff",
          3383 => x"8c",
          3384 => x"70",
          3385 => x"56",
          3386 => x"ec",
          3387 => x"ff",
          3388 => x"c8",
          3389 => x"2b",
          3390 => x"84",
          3391 => x"70",
          3392 => x"97",
          3393 => x"2c",
          3394 => x"10",
          3395 => x"05",
          3396 => x"70",
          3397 => x"5c",
          3398 => x"5b",
          3399 => x"81",
          3400 => x"2e",
          3401 => x"78",
          3402 => x"87",
          3403 => x"80",
          3404 => x"ff",
          3405 => x"98",
          3406 => x"80",
          3407 => x"cb",
          3408 => x"16",
          3409 => x"56",
          3410 => x"83",
          3411 => x"33",
          3412 => x"61",
          3413 => x"83",
          3414 => x"08",
          3415 => x"56",
          3416 => x"2e",
          3417 => x"76",
          3418 => x"38",
          3419 => x"c4",
          3420 => x"76",
          3421 => x"99",
          3422 => x"70",
          3423 => x"98",
          3424 => x"c4",
          3425 => x"2b",
          3426 => x"71",
          3427 => x"70",
          3428 => x"de",
          3429 => x"5f",
          3430 => x"58",
          3431 => x"7a",
          3432 => x"90",
          3433 => x"d1",
          3434 => x"ac",
          3435 => x"76",
          3436 => x"75",
          3437 => x"29",
          3438 => x"05",
          3439 => x"70",
          3440 => x"59",
          3441 => x"95",
          3442 => x"38",
          3443 => x"70",
          3444 => x"55",
          3445 => x"de",
          3446 => x"42",
          3447 => x"25",
          3448 => x"de",
          3449 => x"18",
          3450 => x"55",
          3451 => x"ff",
          3452 => x"80",
          3453 => x"38",
          3454 => x"81",
          3455 => x"2e",
          3456 => x"fe",
          3457 => x"56",
          3458 => x"80",
          3459 => x"e9",
          3460 => x"d1",
          3461 => x"84",
          3462 => x"79",
          3463 => x"7f",
          3464 => x"74",
          3465 => x"b0",
          3466 => x"10",
          3467 => x"05",
          3468 => x"04",
          3469 => x"15",
          3470 => x"80",
          3471 => x"c8",
          3472 => x"84",
          3473 => x"d9",
          3474 => x"d0",
          3475 => x"80",
          3476 => x"38",
          3477 => x"08",
          3478 => x"ff",
          3479 => x"84",
          3480 => x"ff",
          3481 => x"84",
          3482 => x"fc",
          3483 => x"d1",
          3484 => x"81",
          3485 => x"d1",
          3486 => x"57",
          3487 => x"27",
          3488 => x"84",
          3489 => x"52",
          3490 => x"77",
          3491 => x"34",
          3492 => x"33",
          3493 => x"b5",
          3494 => x"bc",
          3495 => x"2e",
          3496 => x"7c",
          3497 => x"f3",
          3498 => x"08",
          3499 => x"8f",
          3500 => x"84",
          3501 => x"75",
          3502 => x"d1",
          3503 => x"d1",
          3504 => x"56",
          3505 => x"b6",
          3506 => x"f0",
          3507 => x"51",
          3508 => x"3f",
          3509 => x"08",
          3510 => x"ff",
          3511 => x"84",
          3512 => x"52",
          3513 => x"b5",
          3514 => x"d1",
          3515 => x"05",
          3516 => x"d1",
          3517 => x"81",
          3518 => x"74",
          3519 => x"51",
          3520 => x"3f",
          3521 => x"d0",
          3522 => x"39",
          3523 => x"83",
          3524 => x"56",
          3525 => x"38",
          3526 => x"83",
          3527 => x"fc",
          3528 => x"55",
          3529 => x"38",
          3530 => x"75",
          3531 => x"a8",
          3532 => x"ff",
          3533 => x"84",
          3534 => x"84",
          3535 => x"84",
          3536 => x"81",
          3537 => x"05",
          3538 => x"7b",
          3539 => x"9a",
          3540 => x"cc",
          3541 => x"d0",
          3542 => x"74",
          3543 => x"9e",
          3544 => x"f0",
          3545 => x"51",
          3546 => x"3f",
          3547 => x"08",
          3548 => x"ff",
          3549 => x"84",
          3550 => x"52",
          3551 => x"b3",
          3552 => x"d1",
          3553 => x"05",
          3554 => x"d1",
          3555 => x"81",
          3556 => x"c7",
          3557 => x"d0",
          3558 => x"ff",
          3559 => x"cc",
          3560 => x"55",
          3561 => x"fa",
          3562 => x"d5",
          3563 => x"81",
          3564 => x"84",
          3565 => x"7b",
          3566 => x"52",
          3567 => x"ae",
          3568 => x"d0",
          3569 => x"ff",
          3570 => x"cc",
          3571 => x"55",
          3572 => x"fa",
          3573 => x"d5",
          3574 => x"81",
          3575 => x"84",
          3576 => x"7b",
          3577 => x"52",
          3578 => x"82",
          3579 => x"d0",
          3580 => x"ff",
          3581 => x"cc",
          3582 => x"55",
          3583 => x"ff",
          3584 => x"d4",
          3585 => x"d0",
          3586 => x"cc",
          3587 => x"74",
          3588 => x"c4",
          3589 => x"5b",
          3590 => x"cc",
          3591 => x"2b",
          3592 => x"7c",
          3593 => x"43",
          3594 => x"76",
          3595 => x"38",
          3596 => x"08",
          3597 => x"ff",
          3598 => x"84",
          3599 => x"70",
          3600 => x"98",
          3601 => x"cc",
          3602 => x"57",
          3603 => x"24",
          3604 => x"84",
          3605 => x"52",
          3606 => x"b2",
          3607 => x"81",
          3608 => x"81",
          3609 => x"70",
          3610 => x"d1",
          3611 => x"56",
          3612 => x"24",
          3613 => x"84",
          3614 => x"52",
          3615 => x"b1",
          3616 => x"81",
          3617 => x"81",
          3618 => x"70",
          3619 => x"d1",
          3620 => x"56",
          3621 => x"25",
          3622 => x"f8",
          3623 => x"16",
          3624 => x"33",
          3625 => x"d5",
          3626 => x"77",
          3627 => x"b1",
          3628 => x"81",
          3629 => x"81",
          3630 => x"70",
          3631 => x"d1",
          3632 => x"57",
          3633 => x"25",
          3634 => x"7b",
          3635 => x"18",
          3636 => x"84",
          3637 => x"52",
          3638 => x"ff",
          3639 => x"75",
          3640 => x"29",
          3641 => x"05",
          3642 => x"84",
          3643 => x"5b",
          3644 => x"76",
          3645 => x"38",
          3646 => x"84",
          3647 => x"55",
          3648 => x"f7",
          3649 => x"d5",
          3650 => x"88",
          3651 => x"de",
          3652 => x"d0",
          3653 => x"57",
          3654 => x"d0",
          3655 => x"ff",
          3656 => x"39",
          3657 => x"33",
          3658 => x"80",
          3659 => x"d5",
          3660 => x"8a",
          3661 => x"b6",
          3662 => x"cc",
          3663 => x"f4",
          3664 => x"ba",
          3665 => x"ff",
          3666 => x"89",
          3667 => x"d1",
          3668 => x"76",
          3669 => x"d8",
          3670 => x"fc",
          3671 => x"10",
          3672 => x"05",
          3673 => x"5e",
          3674 => x"a0",
          3675 => x"2b",
          3676 => x"83",
          3677 => x"81",
          3678 => x"57",
          3679 => x"ca",
          3680 => x"8c",
          3681 => x"83",
          3682 => x"70",
          3683 => x"f3",
          3684 => x"08",
          3685 => x"74",
          3686 => x"83",
          3687 => x"56",
          3688 => x"8c",
          3689 => x"f4",
          3690 => x"80",
          3691 => x"38",
          3692 => x"d1",
          3693 => x"0b",
          3694 => x"34",
          3695 => x"8c",
          3696 => x"0d",
          3697 => x"d0",
          3698 => x"80",
          3699 => x"84",
          3700 => x"52",
          3701 => x"af",
          3702 => x"d5",
          3703 => x"a0",
          3704 => x"8a",
          3705 => x"f0",
          3706 => x"51",
          3707 => x"3f",
          3708 => x"33",
          3709 => x"75",
          3710 => x"34",
          3711 => x"06",
          3712 => x"38",
          3713 => x"51",
          3714 => x"3f",
          3715 => x"d1",
          3716 => x"0b",
          3717 => x"34",
          3718 => x"83",
          3719 => x"0b",
          3720 => x"84",
          3721 => x"55",
          3722 => x"b6",
          3723 => x"f0",
          3724 => x"51",
          3725 => x"3f",
          3726 => x"08",
          3727 => x"ff",
          3728 => x"84",
          3729 => x"52",
          3730 => x"ae",
          3731 => x"d1",
          3732 => x"05",
          3733 => x"d1",
          3734 => x"81",
          3735 => x"74",
          3736 => x"d2",
          3737 => x"9f",
          3738 => x"0b",
          3739 => x"34",
          3740 => x"d1",
          3741 => x"84",
          3742 => x"b4",
          3743 => x"84",
          3744 => x"70",
          3745 => x"5c",
          3746 => x"2e",
          3747 => x"84",
          3748 => x"ff",
          3749 => x"84",
          3750 => x"ff",
          3751 => x"84",
          3752 => x"84",
          3753 => x"52",
          3754 => x"ad",
          3755 => x"d1",
          3756 => x"98",
          3757 => x"2c",
          3758 => x"33",
          3759 => x"56",
          3760 => x"80",
          3761 => x"d5",
          3762 => x"a0",
          3763 => x"9e",
          3764 => x"d0",
          3765 => x"2b",
          3766 => x"84",
          3767 => x"5d",
          3768 => x"74",
          3769 => x"f0",
          3770 => x"f0",
          3771 => x"51",
          3772 => x"3f",
          3773 => x"0a",
          3774 => x"0a",
          3775 => x"2c",
          3776 => x"33",
          3777 => x"74",
          3778 => x"cc",
          3779 => x"f0",
          3780 => x"51",
          3781 => x"3f",
          3782 => x"0a",
          3783 => x"0a",
          3784 => x"2c",
          3785 => x"33",
          3786 => x"78",
          3787 => x"b9",
          3788 => x"39",
          3789 => x"81",
          3790 => x"34",
          3791 => x"08",
          3792 => x"51",
          3793 => x"3f",
          3794 => x"0a",
          3795 => x"0a",
          3796 => x"2c",
          3797 => x"33",
          3798 => x"75",
          3799 => x"e6",
          3800 => x"57",
          3801 => x"77",
          3802 => x"f0",
          3803 => x"33",
          3804 => x"fa",
          3805 => x"80",
          3806 => x"80",
          3807 => x"98",
          3808 => x"cc",
          3809 => x"5b",
          3810 => x"ff",
          3811 => x"b6",
          3812 => x"d0",
          3813 => x"ff",
          3814 => x"76",
          3815 => x"b8",
          3816 => x"cc",
          3817 => x"75",
          3818 => x"74",
          3819 => x"98",
          3820 => x"76",
          3821 => x"38",
          3822 => x"7a",
          3823 => x"34",
          3824 => x"0a",
          3825 => x"0a",
          3826 => x"2c",
          3827 => x"33",
          3828 => x"75",
          3829 => x"38",
          3830 => x"74",
          3831 => x"34",
          3832 => x"06",
          3833 => x"b3",
          3834 => x"34",
          3835 => x"33",
          3836 => x"25",
          3837 => x"17",
          3838 => x"d1",
          3839 => x"57",
          3840 => x"33",
          3841 => x"0a",
          3842 => x"0a",
          3843 => x"2c",
          3844 => x"06",
          3845 => x"58",
          3846 => x"81",
          3847 => x"98",
          3848 => x"2c",
          3849 => x"06",
          3850 => x"75",
          3851 => x"a8",
          3852 => x"f0",
          3853 => x"51",
          3854 => x"3f",
          3855 => x"0a",
          3856 => x"0a",
          3857 => x"2c",
          3858 => x"33",
          3859 => x"75",
          3860 => x"84",
          3861 => x"f0",
          3862 => x"51",
          3863 => x"3f",
          3864 => x"0a",
          3865 => x"0a",
          3866 => x"2c",
          3867 => x"33",
          3868 => x"74",
          3869 => x"b9",
          3870 => x"39",
          3871 => x"08",
          3872 => x"2e",
          3873 => x"75",
          3874 => x"9c",
          3875 => x"8c",
          3876 => x"cc",
          3877 => x"8c",
          3878 => x"06",
          3879 => x"75",
          3880 => x"ff",
          3881 => x"84",
          3882 => x"84",
          3883 => x"56",
          3884 => x"2e",
          3885 => x"84",
          3886 => x"52",
          3887 => x"a9",
          3888 => x"d5",
          3889 => x"a0",
          3890 => x"a2",
          3891 => x"f0",
          3892 => x"51",
          3893 => x"3f",
          3894 => x"33",
          3895 => x"7a",
          3896 => x"34",
          3897 => x"06",
          3898 => x"a8",
          3899 => x"da",
          3900 => x"8c",
          3901 => x"f8",
          3902 => x"8c",
          3903 => x"38",
          3904 => x"f4",
          3905 => x"ca",
          3906 => x"39",
          3907 => x"08",
          3908 => x"70",
          3909 => x"ff",
          3910 => x"75",
          3911 => x"29",
          3912 => x"05",
          3913 => x"84",
          3914 => x"52",
          3915 => x"76",
          3916 => x"84",
          3917 => x"70",
          3918 => x"98",
          3919 => x"ff",
          3920 => x"5a",
          3921 => x"25",
          3922 => x"fd",
          3923 => x"f3",
          3924 => x"2e",
          3925 => x"83",
          3926 => x"93",
          3927 => x"55",
          3928 => x"ff",
          3929 => x"58",
          3930 => x"25",
          3931 => x"0b",
          3932 => x"34",
          3933 => x"08",
          3934 => x"2e",
          3935 => x"74",
          3936 => x"c5",
          3937 => x"f8",
          3938 => x"da",
          3939 => x"0b",
          3940 => x"0c",
          3941 => x"3d",
          3942 => x"bc",
          3943 => x"80",
          3944 => x"80",
          3945 => x"16",
          3946 => x"56",
          3947 => x"ff",
          3948 => x"ba",
          3949 => x"ff",
          3950 => x"84",
          3951 => x"84",
          3952 => x"84",
          3953 => x"81",
          3954 => x"05",
          3955 => x"7b",
          3956 => x"96",
          3957 => x"84",
          3958 => x"84",
          3959 => x"57",
          3960 => x"80",
          3961 => x"38",
          3962 => x"08",
          3963 => x"ff",
          3964 => x"84",
          3965 => x"52",
          3966 => x"a6",
          3967 => x"d5",
          3968 => x"88",
          3969 => x"e6",
          3970 => x"d0",
          3971 => x"5a",
          3972 => x"d0",
          3973 => x"ff",
          3974 => x"39",
          3975 => x"80",
          3976 => x"d0",
          3977 => x"84",
          3978 => x"7b",
          3979 => x"0c",
          3980 => x"04",
          3981 => x"a9",
          3982 => x"ba",
          3983 => x"d1",
          3984 => x"ba",
          3985 => x"ff",
          3986 => x"53",
          3987 => x"51",
          3988 => x"3f",
          3989 => x"81",
          3990 => x"d1",
          3991 => x"d1",
          3992 => x"52",
          3993 => x"80",
          3994 => x"38",
          3995 => x"08",
          3996 => x"ff",
          3997 => x"84",
          3998 => x"52",
          3999 => x"a5",
          4000 => x"d5",
          4001 => x"88",
          4002 => x"e2",
          4003 => x"d0",
          4004 => x"57",
          4005 => x"d0",
          4006 => x"ff",
          4007 => x"39",
          4008 => x"a9",
          4009 => x"ba",
          4010 => x"d1",
          4011 => x"ba",
          4012 => x"ff",
          4013 => x"53",
          4014 => x"51",
          4015 => x"3f",
          4016 => x"81",
          4017 => x"d1",
          4018 => x"d1",
          4019 => x"58",
          4020 => x"80",
          4021 => x"38",
          4022 => x"08",
          4023 => x"ff",
          4024 => x"84",
          4025 => x"52",
          4026 => x"a5",
          4027 => x"d5",
          4028 => x"88",
          4029 => x"f6",
          4030 => x"d0",
          4031 => x"41",
          4032 => x"d0",
          4033 => x"ff",
          4034 => x"39",
          4035 => x"d7",
          4036 => x"f3",
          4037 => x"82",
          4038 => x"06",
          4039 => x"05",
          4040 => x"54",
          4041 => x"80",
          4042 => x"84",
          4043 => x"7b",
          4044 => x"fc",
          4045 => x"10",
          4046 => x"05",
          4047 => x"41",
          4048 => x"2e",
          4049 => x"75",
          4050 => x"74",
          4051 => x"9a",
          4052 => x"fc",
          4053 => x"70",
          4054 => x"5a",
          4055 => x"27",
          4056 => x"77",
          4057 => x"34",
          4058 => x"b4",
          4059 => x"05",
          4060 => x"7b",
          4061 => x"81",
          4062 => x"83",
          4063 => x"52",
          4064 => x"ba",
          4065 => x"f3",
          4066 => x"81",
          4067 => x"80",
          4068 => x"d0",
          4069 => x"84",
          4070 => x"7b",
          4071 => x"0c",
          4072 => x"04",
          4073 => x"52",
          4074 => x"08",
          4075 => x"c7",
          4076 => x"8c",
          4077 => x"38",
          4078 => x"08",
          4079 => x"5d",
          4080 => x"08",
          4081 => x"52",
          4082 => x"b8",
          4083 => x"ba",
          4084 => x"84",
          4085 => x"7b",
          4086 => x"06",
          4087 => x"84",
          4088 => x"51",
          4089 => x"3f",
          4090 => x"08",
          4091 => x"84",
          4092 => x"25",
          4093 => x"84",
          4094 => x"ff",
          4095 => x"58",
          4096 => x"34",
          4097 => x"06",
          4098 => x"33",
          4099 => x"83",
          4100 => x"70",
          4101 => x"58",
          4102 => x"f2",
          4103 => x"2b",
          4104 => x"83",
          4105 => x"81",
          4106 => x"58",
          4107 => x"9a",
          4108 => x"8c",
          4109 => x"83",
          4110 => x"70",
          4111 => x"f3",
          4112 => x"08",
          4113 => x"74",
          4114 => x"1d",
          4115 => x"06",
          4116 => x"7d",
          4117 => x"80",
          4118 => x"2e",
          4119 => x"fe",
          4120 => x"e8",
          4121 => x"e6",
          4122 => x"79",
          4123 => x"ff",
          4124 => x"83",
          4125 => x"81",
          4126 => x"ff",
          4127 => x"93",
          4128 => x"c8",
          4129 => x"83",
          4130 => x"ff",
          4131 => x"51",
          4132 => x"3f",
          4133 => x"33",
          4134 => x"87",
          4135 => x"f3",
          4136 => x"1b",
          4137 => x"56",
          4138 => x"9e",
          4139 => x"8c",
          4140 => x"83",
          4141 => x"70",
          4142 => x"f3",
          4143 => x"08",
          4144 => x"74",
          4145 => x"82",
          4146 => x"39",
          4147 => x"fc",
          4148 => x"39",
          4149 => x"fc",
          4150 => x"39",
          4151 => x"51",
          4152 => x"3f",
          4153 => x"38",
          4154 => x"f2",
          4155 => x"80",
          4156 => x"02",
          4157 => x"c7",
          4158 => x"53",
          4159 => x"81",
          4160 => x"81",
          4161 => x"38",
          4162 => x"83",
          4163 => x"82",
          4164 => x"38",
          4165 => x"80",
          4166 => x"b0",
          4167 => x"57",
          4168 => x"a0",
          4169 => x"2e",
          4170 => x"83",
          4171 => x"75",
          4172 => x"34",
          4173 => x"ba",
          4174 => x"b8",
          4175 => x"2b",
          4176 => x"07",
          4177 => x"07",
          4178 => x"7f",
          4179 => x"5b",
          4180 => x"94",
          4181 => x"70",
          4182 => x"0c",
          4183 => x"84",
          4184 => x"76",
          4185 => x"38",
          4186 => x"a2",
          4187 => x"b8",
          4188 => x"de",
          4189 => x"31",
          4190 => x"a0",
          4191 => x"15",
          4192 => x"70",
          4193 => x"34",
          4194 => x"72",
          4195 => x"3d",
          4196 => x"a3",
          4197 => x"83",
          4198 => x"70",
          4199 => x"83",
          4200 => x"71",
          4201 => x"74",
          4202 => x"58",
          4203 => x"a3",
          4204 => x"84",
          4205 => x"70",
          4206 => x"84",
          4207 => x"70",
          4208 => x"83",
          4209 => x"70",
          4210 => x"06",
          4211 => x"5d",
          4212 => x"5e",
          4213 => x"73",
          4214 => x"38",
          4215 => x"75",
          4216 => x"81",
          4217 => x"81",
          4218 => x"81",
          4219 => x"83",
          4220 => x"62",
          4221 => x"70",
          4222 => x"5d",
          4223 => x"5b",
          4224 => x"26",
          4225 => x"f9",
          4226 => x"76",
          4227 => x"7d",
          4228 => x"5f",
          4229 => x"5c",
          4230 => x"fe",
          4231 => x"7d",
          4232 => x"77",
          4233 => x"38",
          4234 => x"81",
          4235 => x"83",
          4236 => x"74",
          4237 => x"56",
          4238 => x"87",
          4239 => x"59",
          4240 => x"80",
          4241 => x"80",
          4242 => x"ff",
          4243 => x"ff",
          4244 => x"ff",
          4245 => x"ba",
          4246 => x"29",
          4247 => x"57",
          4248 => x"57",
          4249 => x"81",
          4250 => x"81",
          4251 => x"81",
          4252 => x"71",
          4253 => x"54",
          4254 => x"2e",
          4255 => x"80",
          4256 => x"bc",
          4257 => x"83",
          4258 => x"83",
          4259 => x"70",
          4260 => x"90",
          4261 => x"88",
          4262 => x"07",
          4263 => x"56",
          4264 => x"79",
          4265 => x"38",
          4266 => x"72",
          4267 => x"83",
          4268 => x"70",
          4269 => x"70",
          4270 => x"83",
          4271 => x"71",
          4272 => x"87",
          4273 => x"11",
          4274 => x"56",
          4275 => x"a3",
          4276 => x"14",
          4277 => x"33",
          4278 => x"06",
          4279 => x"33",
          4280 => x"06",
          4281 => x"22",
          4282 => x"ff",
          4283 => x"29",
          4284 => x"5a",
          4285 => x"5f",
          4286 => x"79",
          4287 => x"38",
          4288 => x"15",
          4289 => x"19",
          4290 => x"81",
          4291 => x"81",
          4292 => x"71",
          4293 => x"ff",
          4294 => x"81",
          4295 => x"75",
          4296 => x"5b",
          4297 => x"7b",
          4298 => x"38",
          4299 => x"53",
          4300 => x"16",
          4301 => x"5b",
          4302 => x"e2",
          4303 => x"06",
          4304 => x"da",
          4305 => x"39",
          4306 => x"7b",
          4307 => x"9a",
          4308 => x"0d",
          4309 => x"9c",
          4310 => x"74",
          4311 => x"74",
          4312 => x"80",
          4313 => x"73",
          4314 => x"34",
          4315 => x"94",
          4316 => x"34",
          4317 => x"ff",
          4318 => x"86",
          4319 => x"55",
          4320 => x"34",
          4321 => x"85",
          4322 => x"75",
          4323 => x"83",
          4324 => x"3f",
          4325 => x"e0",
          4326 => x"54",
          4327 => x"87",
          4328 => x"73",
          4329 => x"07",
          4330 => x"75",
          4331 => x"70",
          4332 => x"80",
          4333 => x"53",
          4334 => x"87",
          4335 => x"08",
          4336 => x"81",
          4337 => x"72",
          4338 => x"f3",
          4339 => x"81",
          4340 => x"07",
          4341 => x"34",
          4342 => x"84",
          4343 => x"80",
          4344 => x"8c",
          4345 => x"0d",
          4346 => x"80",
          4347 => x"8c",
          4348 => x"3d",
          4349 => x"05",
          4350 => x"05",
          4351 => x"84",
          4352 => x"5b",
          4353 => x"53",
          4354 => x"82",
          4355 => x"b8",
          4356 => x"f9",
          4357 => x"f9",
          4358 => x"71",
          4359 => x"a3",
          4360 => x"83",
          4361 => x"5f",
          4362 => x"71",
          4363 => x"70",
          4364 => x"06",
          4365 => x"33",
          4366 => x"53",
          4367 => x"83",
          4368 => x"f9",
          4369 => x"05",
          4370 => x"f9",
          4371 => x"f9",
          4372 => x"05",
          4373 => x"06",
          4374 => x"06",
          4375 => x"72",
          4376 => x"8c",
          4377 => x"53",
          4378 => x"bc",
          4379 => x"ba",
          4380 => x"ff",
          4381 => x"b7",
          4382 => x"55",
          4383 => x"26",
          4384 => x"84",
          4385 => x"76",
          4386 => x"58",
          4387 => x"9f",
          4388 => x"38",
          4389 => x"70",
          4390 => x"e0",
          4391 => x"e0",
          4392 => x"72",
          4393 => x"54",
          4394 => x"81",
          4395 => x"81",
          4396 => x"b7",
          4397 => x"e3",
          4398 => x"9f",
          4399 => x"83",
          4400 => x"84",
          4401 => x"54",
          4402 => x"e0",
          4403 => x"74",
          4404 => x"05",
          4405 => x"14",
          4406 => x"74",
          4407 => x"84",
          4408 => x"ff",
          4409 => x"83",
          4410 => x"75",
          4411 => x"ff",
          4412 => x"ff",
          4413 => x"54",
          4414 => x"81",
          4415 => x"74",
          4416 => x"84",
          4417 => x"71",
          4418 => x"55",
          4419 => x"87",
          4420 => x"58",
          4421 => x"80",
          4422 => x"06",
          4423 => x"06",
          4424 => x"19",
          4425 => x"57",
          4426 => x"b9",
          4427 => x"de",
          4428 => x"e0",
          4429 => x"84",
          4430 => x"33",
          4431 => x"05",
          4432 => x"70",
          4433 => x"33",
          4434 => x"05",
          4435 => x"15",
          4436 => x"33",
          4437 => x"33",
          4438 => x"19",
          4439 => x"55",
          4440 => x"ce",
          4441 => x"72",
          4442 => x"0c",
          4443 => x"04",
          4444 => x"bc",
          4445 => x"ba",
          4446 => x"ff",
          4447 => x"b7",
          4448 => x"55",
          4449 => x"27",
          4450 => x"77",
          4451 => x"dd",
          4452 => x"ff",
          4453 => x"83",
          4454 => x"56",
          4455 => x"2e",
          4456 => x"fe",
          4457 => x"76",
          4458 => x"84",
          4459 => x"71",
          4460 => x"72",
          4461 => x"52",
          4462 => x"73",
          4463 => x"38",
          4464 => x"33",
          4465 => x"15",
          4466 => x"55",
          4467 => x"0b",
          4468 => x"34",
          4469 => x"81",
          4470 => x"ff",
          4471 => x"80",
          4472 => x"38",
          4473 => x"e0",
          4474 => x"75",
          4475 => x"57",
          4476 => x"53",
          4477 => x"fd",
          4478 => x"0b",
          4479 => x"33",
          4480 => x"89",
          4481 => x"be",
          4482 => x"84",
          4483 => x"33",
          4484 => x"b7",
          4485 => x"fc",
          4486 => x"3d",
          4487 => x"84",
          4488 => x"33",
          4489 => x"86",
          4490 => x"70",
          4491 => x"c4",
          4492 => x"70",
          4493 => x"b8",
          4494 => x"71",
          4495 => x"38",
          4496 => x"bd",
          4497 => x"84",
          4498 => x"86",
          4499 => x"80",
          4500 => x"bd",
          4501 => x"bc",
          4502 => x"ff",
          4503 => x"72",
          4504 => x"38",
          4505 => x"70",
          4506 => x"34",
          4507 => x"ba",
          4508 => x"3d",
          4509 => x"f9",
          4510 => x"73",
          4511 => x"70",
          4512 => x"06",
          4513 => x"54",
          4514 => x"bc",
          4515 => x"83",
          4516 => x"72",
          4517 => x"ff",
          4518 => x"55",
          4519 => x"75",
          4520 => x"70",
          4521 => x"f9",
          4522 => x"0b",
          4523 => x"0c",
          4524 => x"04",
          4525 => x"33",
          4526 => x"70",
          4527 => x"2c",
          4528 => x"56",
          4529 => x"83",
          4530 => x"80",
          4531 => x"8c",
          4532 => x"0d",
          4533 => x"bd",
          4534 => x"84",
          4535 => x"ff",
          4536 => x"51",
          4537 => x"83",
          4538 => x"72",
          4539 => x"34",
          4540 => x"ba",
          4541 => x"3d",
          4542 => x"0b",
          4543 => x"34",
          4544 => x"33",
          4545 => x"33",
          4546 => x"52",
          4547 => x"fe",
          4548 => x"12",
          4549 => x"f9",
          4550 => x"d0",
          4551 => x"0d",
          4552 => x"33",
          4553 => x"26",
          4554 => x"10",
          4555 => x"d0",
          4556 => x"08",
          4557 => x"b8",
          4558 => x"f0",
          4559 => x"2b",
          4560 => x"70",
          4561 => x"07",
          4562 => x"51",
          4563 => x"2e",
          4564 => x"9c",
          4565 => x"0b",
          4566 => x"34",
          4567 => x"ba",
          4568 => x"3d",
          4569 => x"f9",
          4570 => x"9f",
          4571 => x"51",
          4572 => x"b8",
          4573 => x"84",
          4574 => x"83",
          4575 => x"83",
          4576 => x"80",
          4577 => x"70",
          4578 => x"34",
          4579 => x"f9",
          4580 => x"fe",
          4581 => x"51",
          4582 => x"b8",
          4583 => x"80",
          4584 => x"f9",
          4585 => x"0b",
          4586 => x"0c",
          4587 => x"04",
          4588 => x"33",
          4589 => x"84",
          4590 => x"83",
          4591 => x"ff",
          4592 => x"f9",
          4593 => x"07",
          4594 => x"f9",
          4595 => x"a5",
          4596 => x"b8",
          4597 => x"06",
          4598 => x"70",
          4599 => x"34",
          4600 => x"83",
          4601 => x"81",
          4602 => x"07",
          4603 => x"f9",
          4604 => x"81",
          4605 => x"b8",
          4606 => x"06",
          4607 => x"70",
          4608 => x"34",
          4609 => x"83",
          4610 => x"81",
          4611 => x"70",
          4612 => x"34",
          4613 => x"83",
          4614 => x"81",
          4615 => x"d0",
          4616 => x"83",
          4617 => x"fe",
          4618 => x"f9",
          4619 => x"bf",
          4620 => x"51",
          4621 => x"b8",
          4622 => x"39",
          4623 => x"33",
          4624 => x"80",
          4625 => x"70",
          4626 => x"34",
          4627 => x"83",
          4628 => x"81",
          4629 => x"c0",
          4630 => x"83",
          4631 => x"fe",
          4632 => x"f9",
          4633 => x"af",
          4634 => x"51",
          4635 => x"b8",
          4636 => x"39",
          4637 => x"33",
          4638 => x"51",
          4639 => x"b8",
          4640 => x"39",
          4641 => x"33",
          4642 => x"82",
          4643 => x"83",
          4644 => x"fd",
          4645 => x"3d",
          4646 => x"05",
          4647 => x"05",
          4648 => x"33",
          4649 => x"33",
          4650 => x"33",
          4651 => x"33",
          4652 => x"33",
          4653 => x"5d",
          4654 => x"82",
          4655 => x"38",
          4656 => x"a5",
          4657 => x"2e",
          4658 => x"7d",
          4659 => x"34",
          4660 => x"b8",
          4661 => x"83",
          4662 => x"7b",
          4663 => x"23",
          4664 => x"bd",
          4665 => x"0d",
          4666 => x"2e",
          4667 => x"db",
          4668 => x"84",
          4669 => x"81",
          4670 => x"84",
          4671 => x"83",
          4672 => x"a8",
          4673 => x"bd",
          4674 => x"83",
          4675 => x"79",
          4676 => x"80",
          4677 => x"b7",
          4678 => x"84",
          4679 => x"55",
          4680 => x"53",
          4681 => x"e3",
          4682 => x"81",
          4683 => x"84",
          4684 => x"80",
          4685 => x"84",
          4686 => x"f9",
          4687 => x"83",
          4688 => x"7c",
          4689 => x"34",
          4690 => x"04",
          4691 => x"b8",
          4692 => x"0b",
          4693 => x"34",
          4694 => x"f9",
          4695 => x"0b",
          4696 => x"34",
          4697 => x"f9",
          4698 => x"b9",
          4699 => x"84",
          4700 => x"57",
          4701 => x"33",
          4702 => x"7b",
          4703 => x"7a",
          4704 => x"e0",
          4705 => x"80",
          4706 => x"84",
          4707 => x"5a",
          4708 => x"27",
          4709 => x"10",
          4710 => x"05",
          4711 => x"59",
          4712 => x"51",
          4713 => x"3f",
          4714 => x"81",
          4715 => x"b9",
          4716 => x"5b",
          4717 => x"26",
          4718 => x"d2",
          4719 => x"80",
          4720 => x"84",
          4721 => x"80",
          4722 => x"84",
          4723 => x"f9",
          4724 => x"83",
          4725 => x"7c",
          4726 => x"34",
          4727 => x"04",
          4728 => x"b8",
          4729 => x"0b",
          4730 => x"34",
          4731 => x"f9",
          4732 => x"0b",
          4733 => x"34",
          4734 => x"f9",
          4735 => x"f7",
          4736 => x"92",
          4737 => x"ba",
          4738 => x"83",
          4739 => x"fe",
          4740 => x"80",
          4741 => x"f0",
          4742 => x"8c",
          4743 => x"ba",
          4744 => x"fd",
          4745 => x"f7",
          4746 => x"52",
          4747 => x"51",
          4748 => x"3f",
          4749 => x"81",
          4750 => x"5a",
          4751 => x"3d",
          4752 => x"84",
          4753 => x"33",
          4754 => x"33",
          4755 => x"33",
          4756 => x"33",
          4757 => x"12",
          4758 => x"80",
          4759 => x"ba",
          4760 => x"59",
          4761 => x"29",
          4762 => x"ff",
          4763 => x"f8",
          4764 => x"59",
          4765 => x"57",
          4766 => x"81",
          4767 => x"89",
          4768 => x"38",
          4769 => x"81",
          4770 => x"81",
          4771 => x"38",
          4772 => x"82",
          4773 => x"b8",
          4774 => x"f9",
          4775 => x"f9",
          4776 => x"72",
          4777 => x"56",
          4778 => x"88",
          4779 => x"a3",
          4780 => x"34",
          4781 => x"33",
          4782 => x"33",
          4783 => x"22",
          4784 => x"12",
          4785 => x"53",
          4786 => x"be",
          4787 => x"f9",
          4788 => x"71",
          4789 => x"54",
          4790 => x"33",
          4791 => x"80",
          4792 => x"b8",
          4793 => x"81",
          4794 => x"f9",
          4795 => x"f9",
          4796 => x"72",
          4797 => x"5b",
          4798 => x"83",
          4799 => x"84",
          4800 => x"34",
          4801 => x"81",
          4802 => x"55",
          4803 => x"81",
          4804 => x"b8",
          4805 => x"77",
          4806 => x"ff",
          4807 => x"83",
          4808 => x"84",
          4809 => x"53",
          4810 => x"8c",
          4811 => x"84",
          4812 => x"80",
          4813 => x"38",
          4814 => x"ba",
          4815 => x"3d",
          4816 => x"8d",
          4817 => x"75",
          4818 => x"f7",
          4819 => x"2e",
          4820 => x"fe",
          4821 => x"52",
          4822 => x"96",
          4823 => x"83",
          4824 => x"ff",
          4825 => x"f9",
          4826 => x"53",
          4827 => x"13",
          4828 => x"75",
          4829 => x"81",
          4830 => x"38",
          4831 => x"52",
          4832 => x"ba",
          4833 => x"70",
          4834 => x"54",
          4835 => x"26",
          4836 => x"76",
          4837 => x"fd",
          4838 => x"13",
          4839 => x"06",
          4840 => x"73",
          4841 => x"fe",
          4842 => x"83",
          4843 => x"fe",
          4844 => x"52",
          4845 => x"de",
          4846 => x"84",
          4847 => x"89",
          4848 => x"75",
          4849 => x"09",
          4850 => x"ca",
          4851 => x"bd",
          4852 => x"ff",
          4853 => x"05",
          4854 => x"38",
          4855 => x"83",
          4856 => x"76",
          4857 => x"fc",
          4858 => x"f9",
          4859 => x"81",
          4860 => x"ff",
          4861 => x"fe",
          4862 => x"53",
          4863 => x"bd",
          4864 => x"39",
          4865 => x"f9",
          4866 => x"52",
          4867 => x"e2",
          4868 => x"39",
          4869 => x"51",
          4870 => x"fe",
          4871 => x"3d",
          4872 => x"f3",
          4873 => x"b9",
          4874 => x"59",
          4875 => x"81",
          4876 => x"82",
          4877 => x"38",
          4878 => x"84",
          4879 => x"8a",
          4880 => x"38",
          4881 => x"84",
          4882 => x"89",
          4883 => x"38",
          4884 => x"33",
          4885 => x"33",
          4886 => x"33",
          4887 => x"05",
          4888 => x"84",
          4889 => x"33",
          4890 => x"80",
          4891 => x"b8",
          4892 => x"f9",
          4893 => x"f9",
          4894 => x"71",
          4895 => x"5a",
          4896 => x"83",
          4897 => x"34",
          4898 => x"33",
          4899 => x"62",
          4900 => x"83",
          4901 => x"7f",
          4902 => x"80",
          4903 => x"b8",
          4904 => x"81",
          4905 => x"f9",
          4906 => x"f9",
          4907 => x"72",
          4908 => x"40",
          4909 => x"83",
          4910 => x"84",
          4911 => x"34",
          4912 => x"81",
          4913 => x"58",
          4914 => x"81",
          4915 => x"b8",
          4916 => x"79",
          4917 => x"ff",
          4918 => x"83",
          4919 => x"80",
          4920 => x"8c",
          4921 => x"0d",
          4922 => x"2e",
          4923 => x"b7",
          4924 => x"fd",
          4925 => x"2e",
          4926 => x"78",
          4927 => x"89",
          4928 => x"0b",
          4929 => x"0c",
          4930 => x"33",
          4931 => x"33",
          4932 => x"33",
          4933 => x"05",
          4934 => x"84",
          4935 => x"33",
          4936 => x"80",
          4937 => x"b8",
          4938 => x"f9",
          4939 => x"f9",
          4940 => x"71",
          4941 => x"5f",
          4942 => x"83",
          4943 => x"34",
          4944 => x"33",
          4945 => x"19",
          4946 => x"f9",
          4947 => x"a3",
          4948 => x"34",
          4949 => x"33",
          4950 => x"06",
          4951 => x"22",
          4952 => x"33",
          4953 => x"11",
          4954 => x"58",
          4955 => x"b8",
          4956 => x"98",
          4957 => x"81",
          4958 => x"81",
          4959 => x"60",
          4960 => x"ca",
          4961 => x"f9",
          4962 => x"0b",
          4963 => x"0c",
          4964 => x"04",
          4965 => x"82",
          4966 => x"9b",
          4967 => x"38",
          4968 => x"09",
          4969 => x"a8",
          4970 => x"83",
          4971 => x"80",
          4972 => x"8c",
          4973 => x"0d",
          4974 => x"2e",
          4975 => x"d0",
          4976 => x"89",
          4977 => x"38",
          4978 => x"33",
          4979 => x"57",
          4980 => x"8c",
          4981 => x"b9",
          4982 => x"77",
          4983 => x"59",
          4984 => x"b9",
          4985 => x"80",
          4986 => x"8c",
          4987 => x"0d",
          4988 => x"2e",
          4989 => x"80",
          4990 => x"88",
          4991 => x"80",
          4992 => x"bc",
          4993 => x"bd",
          4994 => x"29",
          4995 => x"40",
          4996 => x"19",
          4997 => x"a0",
          4998 => x"84",
          4999 => x"83",
          5000 => x"83",
          5001 => x"72",
          5002 => x"41",
          5003 => x"78",
          5004 => x"1f",
          5005 => x"bc",
          5006 => x"29",
          5007 => x"83",
          5008 => x"87",
          5009 => x"1b",
          5010 => x"80",
          5011 => x"ff",
          5012 => x"ba",
          5013 => x"bd",
          5014 => x"29",
          5015 => x"43",
          5016 => x"f9",
          5017 => x"84",
          5018 => x"34",
          5019 => x"fe",
          5020 => x"52",
          5021 => x"fa",
          5022 => x"83",
          5023 => x"fe",
          5024 => x"b8",
          5025 => x"f9",
          5026 => x"81",
          5027 => x"f9",
          5028 => x"71",
          5029 => x"a3",
          5030 => x"83",
          5031 => x"40",
          5032 => x"7e",
          5033 => x"83",
          5034 => x"83",
          5035 => x"5a",
          5036 => x"5c",
          5037 => x"86",
          5038 => x"81",
          5039 => x"1a",
          5040 => x"fc",
          5041 => x"56",
          5042 => x"bd",
          5043 => x"39",
          5044 => x"b9",
          5045 => x"0b",
          5046 => x"34",
          5047 => x"b9",
          5048 => x"0b",
          5049 => x"34",
          5050 => x"b9",
          5051 => x"0b",
          5052 => x"0c",
          5053 => x"04",
          5054 => x"33",
          5055 => x"34",
          5056 => x"33",
          5057 => x"34",
          5058 => x"33",
          5059 => x"34",
          5060 => x"b9",
          5061 => x"0b",
          5062 => x"0c",
          5063 => x"04",
          5064 => x"2e",
          5065 => x"fa",
          5066 => x"f9",
          5067 => x"b8",
          5068 => x"81",
          5069 => x"f9",
          5070 => x"81",
          5071 => x"75",
          5072 => x"a3",
          5073 => x"83",
          5074 => x"5c",
          5075 => x"29",
          5076 => x"ff",
          5077 => x"f8",
          5078 => x"5c",
          5079 => x"5b",
          5080 => x"2e",
          5081 => x"78",
          5082 => x"ff",
          5083 => x"75",
          5084 => x"57",
          5085 => x"bd",
          5086 => x"ff",
          5087 => x"ff",
          5088 => x"ff",
          5089 => x"29",
          5090 => x"5b",
          5091 => x"33",
          5092 => x"80",
          5093 => x"b8",
          5094 => x"f9",
          5095 => x"f9",
          5096 => x"71",
          5097 => x"5e",
          5098 => x"0b",
          5099 => x"18",
          5100 => x"bc",
          5101 => x"29",
          5102 => x"56",
          5103 => x"33",
          5104 => x"80",
          5105 => x"b8",
          5106 => x"81",
          5107 => x"f9",
          5108 => x"f9",
          5109 => x"72",
          5110 => x"5d",
          5111 => x"83",
          5112 => x"7f",
          5113 => x"05",
          5114 => x"70",
          5115 => x"5c",
          5116 => x"26",
          5117 => x"84",
          5118 => x"5a",
          5119 => x"38",
          5120 => x"77",
          5121 => x"34",
          5122 => x"33",
          5123 => x"06",
          5124 => x"56",
          5125 => x"78",
          5126 => x"d8",
          5127 => x"2e",
          5128 => x"78",
          5129 => x"a8",
          5130 => x"8c",
          5131 => x"83",
          5132 => x"bf",
          5133 => x"b4",
          5134 => x"38",
          5135 => x"83",
          5136 => x"58",
          5137 => x"80",
          5138 => x"bd",
          5139 => x"81",
          5140 => x"3f",
          5141 => x"ba",
          5142 => x"3d",
          5143 => x"f9",
          5144 => x"b8",
          5145 => x"81",
          5146 => x"f9",
          5147 => x"81",
          5148 => x"75",
          5149 => x"a3",
          5150 => x"83",
          5151 => x"5c",
          5152 => x"29",
          5153 => x"ff",
          5154 => x"f8",
          5155 => x"53",
          5156 => x"5b",
          5157 => x"2e",
          5158 => x"80",
          5159 => x"ff",
          5160 => x"ff",
          5161 => x"ff",
          5162 => x"29",
          5163 => x"40",
          5164 => x"33",
          5165 => x"80",
          5166 => x"b8",
          5167 => x"f9",
          5168 => x"f9",
          5169 => x"71",
          5170 => x"41",
          5171 => x"0b",
          5172 => x"1c",
          5173 => x"bc",
          5174 => x"29",
          5175 => x"83",
          5176 => x"87",
          5177 => x"1a",
          5178 => x"80",
          5179 => x"ff",
          5180 => x"ba",
          5181 => x"bd",
          5182 => x"29",
          5183 => x"5a",
          5184 => x"f9",
          5185 => x"98",
          5186 => x"60",
          5187 => x"81",
          5188 => x"58",
          5189 => x"81",
          5190 => x"b8",
          5191 => x"77",
          5192 => x"ff",
          5193 => x"83",
          5194 => x"81",
          5195 => x"ff",
          5196 => x"7b",
          5197 => x"a7",
          5198 => x"bc",
          5199 => x"80",
          5200 => x"bd",
          5201 => x"ff",
          5202 => x"ff",
          5203 => x"ff",
          5204 => x"29",
          5205 => x"43",
          5206 => x"84",
          5207 => x"87",
          5208 => x"1b",
          5209 => x"80",
          5210 => x"bd",
          5211 => x"ba",
          5212 => x"29",
          5213 => x"5e",
          5214 => x"83",
          5215 => x"34",
          5216 => x"33",
          5217 => x"1e",
          5218 => x"f9",
          5219 => x"a3",
          5220 => x"34",
          5221 => x"33",
          5222 => x"06",
          5223 => x"22",
          5224 => x"33",
          5225 => x"11",
          5226 => x"40",
          5227 => x"b8",
          5228 => x"de",
          5229 => x"81",
          5230 => x"ff",
          5231 => x"79",
          5232 => x"d6",
          5233 => x"f9",
          5234 => x"df",
          5235 => x"84",
          5236 => x"80",
          5237 => x"8c",
          5238 => x"0d",
          5239 => x"be",
          5240 => x"84",
          5241 => x"33",
          5242 => x"f9",
          5243 => x"81",
          5244 => x"ff",
          5245 => x"ca",
          5246 => x"84",
          5247 => x"80",
          5248 => x"8c",
          5249 => x"0d",
          5250 => x"be",
          5251 => x"84",
          5252 => x"33",
          5253 => x"f9",
          5254 => x"b8",
          5255 => x"f9",
          5256 => x"5b",
          5257 => x"fc",
          5258 => x"b9",
          5259 => x"3d",
          5260 => x"d8",
          5261 => x"8a",
          5262 => x"ba",
          5263 => x"2e",
          5264 => x"84",
          5265 => x"81",
          5266 => x"75",
          5267 => x"34",
          5268 => x"fe",
          5269 => x"80",
          5270 => x"61",
          5271 => x"05",
          5272 => x"39",
          5273 => x"17",
          5274 => x"b8",
          5275 => x"7b",
          5276 => x"bc",
          5277 => x"80",
          5278 => x"bd",
          5279 => x"5c",
          5280 => x"84",
          5281 => x"83",
          5282 => x"83",
          5283 => x"72",
          5284 => x"41",
          5285 => x"b8",
          5286 => x"7f",
          5287 => x"80",
          5288 => x"b8",
          5289 => x"f9",
          5290 => x"f9",
          5291 => x"71",
          5292 => x"43",
          5293 => x"83",
          5294 => x"34",
          5295 => x"33",
          5296 => x"1b",
          5297 => x"f9",
          5298 => x"87",
          5299 => x"05",
          5300 => x"80",
          5301 => x"ff",
          5302 => x"ba",
          5303 => x"bd",
          5304 => x"29",
          5305 => x"5a",
          5306 => x"f9",
          5307 => x"98",
          5308 => x"81",
          5309 => x"ff",
          5310 => x"60",
          5311 => x"a2",
          5312 => x"81",
          5313 => x"90",
          5314 => x"1a",
          5315 => x"f9",
          5316 => x"0b",
          5317 => x"0c",
          5318 => x"33",
          5319 => x"2e",
          5320 => x"84",
          5321 => x"56",
          5322 => x"38",
          5323 => x"51",
          5324 => x"80",
          5325 => x"8c",
          5326 => x"0d",
          5327 => x"f4",
          5328 => x"bc",
          5329 => x"f5",
          5330 => x"bd",
          5331 => x"f6",
          5332 => x"83",
          5333 => x"ff",
          5334 => x"f9",
          5335 => x"b9",
          5336 => x"f9",
          5337 => x"b9",
          5338 => x"f9",
          5339 => x"b9",
          5340 => x"9e",
          5341 => x"8d",
          5342 => x"80",
          5343 => x"38",
          5344 => x"22",
          5345 => x"2e",
          5346 => x"ff",
          5347 => x"f9",
          5348 => x"05",
          5349 => x"bc",
          5350 => x"54",
          5351 => x"e4",
          5352 => x"3d",
          5353 => x"fe",
          5354 => x"76",
          5355 => x"f8",
          5356 => x"8c",
          5357 => x"06",
          5358 => x"33",
          5359 => x"41",
          5360 => x"fe",
          5361 => x"52",
          5362 => x"51",
          5363 => x"3f",
          5364 => x"80",
          5365 => x"8d",
          5366 => x"79",
          5367 => x"5b",
          5368 => x"fe",
          5369 => x"10",
          5370 => x"05",
          5371 => x"57",
          5372 => x"26",
          5373 => x"75",
          5374 => x"c7",
          5375 => x"7e",
          5376 => x"b9",
          5377 => x"7d",
          5378 => x"a4",
          5379 => x"bc",
          5380 => x"e1",
          5381 => x"31",
          5382 => x"9f",
          5383 => x"5a",
          5384 => x"5c",
          5385 => x"bc",
          5386 => x"39",
          5387 => x"33",
          5388 => x"2e",
          5389 => x"84",
          5390 => x"ff",
          5391 => x"ff",
          5392 => x"80",
          5393 => x"5f",
          5394 => x"fd",
          5395 => x"83",
          5396 => x"fd",
          5397 => x"0b",
          5398 => x"34",
          5399 => x"33",
          5400 => x"06",
          5401 => x"80",
          5402 => x"38",
          5403 => x"75",
          5404 => x"34",
          5405 => x"80",
          5406 => x"bd",
          5407 => x"bc",
          5408 => x"ff",
          5409 => x"57",
          5410 => x"25",
          5411 => x"81",
          5412 => x"83",
          5413 => x"fc",
          5414 => x"b9",
          5415 => x"7f",
          5416 => x"e0",
          5417 => x"bd",
          5418 => x"e1",
          5419 => x"31",
          5420 => x"9f",
          5421 => x"5a",
          5422 => x"5a",
          5423 => x"bd",
          5424 => x"39",
          5425 => x"33",
          5426 => x"2e",
          5427 => x"84",
          5428 => x"41",
          5429 => x"09",
          5430 => x"b6",
          5431 => x"80",
          5432 => x"bd",
          5433 => x"bc",
          5434 => x"29",
          5435 => x"a0",
          5436 => x"f9",
          5437 => x"51",
          5438 => x"60",
          5439 => x"83",
          5440 => x"83",
          5441 => x"87",
          5442 => x"06",
          5443 => x"5d",
          5444 => x"80",
          5445 => x"38",
          5446 => x"f8",
          5447 => x"f2",
          5448 => x"8d",
          5449 => x"80",
          5450 => x"38",
          5451 => x"22",
          5452 => x"2e",
          5453 => x"fb",
          5454 => x"0b",
          5455 => x"34",
          5456 => x"84",
          5457 => x"56",
          5458 => x"90",
          5459 => x"b9",
          5460 => x"f9",
          5461 => x"7c",
          5462 => x"80",
          5463 => x"59",
          5464 => x"7d",
          5465 => x"75",
          5466 => x"f9",
          5467 => x"a2",
          5468 => x"8d",
          5469 => x"80",
          5470 => x"38",
          5471 => x"33",
          5472 => x"33",
          5473 => x"84",
          5474 => x"ff",
          5475 => x"56",
          5476 => x"83",
          5477 => x"76",
          5478 => x"34",
          5479 => x"83",
          5480 => x"fe",
          5481 => x"80",
          5482 => x"8d",
          5483 => x"76",
          5484 => x"c7",
          5485 => x"84",
          5486 => x"70",
          5487 => x"83",
          5488 => x"fe",
          5489 => x"81",
          5490 => x"ff",
          5491 => x"8d",
          5492 => x"58",
          5493 => x"0b",
          5494 => x"33",
          5495 => x"80",
          5496 => x"84",
          5497 => x"56",
          5498 => x"83",
          5499 => x"81",
          5500 => x"ff",
          5501 => x"f3",
          5502 => x"39",
          5503 => x"33",
          5504 => x"27",
          5505 => x"84",
          5506 => x"ff",
          5507 => x"ff",
          5508 => x"e1",
          5509 => x"70",
          5510 => x"84",
          5511 => x"70",
          5512 => x"ff",
          5513 => x"52",
          5514 => x"5c",
          5515 => x"83",
          5516 => x"79",
          5517 => x"23",
          5518 => x"06",
          5519 => x"5f",
          5520 => x"83",
          5521 => x"76",
          5522 => x"34",
          5523 => x"33",
          5524 => x"40",
          5525 => x"f9",
          5526 => x"56",
          5527 => x"bd",
          5528 => x"39",
          5529 => x"33",
          5530 => x"2e",
          5531 => x"84",
          5532 => x"84",
          5533 => x"40",
          5534 => x"26",
          5535 => x"83",
          5536 => x"84",
          5537 => x"70",
          5538 => x"83",
          5539 => x"71",
          5540 => x"87",
          5541 => x"05",
          5542 => x"22",
          5543 => x"7e",
          5544 => x"83",
          5545 => x"83",
          5546 => x"46",
          5547 => x"5f",
          5548 => x"2e",
          5549 => x"79",
          5550 => x"06",
          5551 => x"5d",
          5552 => x"24",
          5553 => x"84",
          5554 => x"56",
          5555 => x"8e",
          5556 => x"16",
          5557 => x"f9",
          5558 => x"81",
          5559 => x"7c",
          5560 => x"80",
          5561 => x"e5",
          5562 => x"ff",
          5563 => x"76",
          5564 => x"38",
          5565 => x"75",
          5566 => x"34",
          5567 => x"06",
          5568 => x"22",
          5569 => x"5a",
          5570 => x"90",
          5571 => x"31",
          5572 => x"81",
          5573 => x"71",
          5574 => x"5b",
          5575 => x"a3",
          5576 => x"87",
          5577 => x"7f",
          5578 => x"7f",
          5579 => x"71",
          5580 => x"42",
          5581 => x"79",
          5582 => x"d6",
          5583 => x"de",
          5584 => x"e0",
          5585 => x"84",
          5586 => x"33",
          5587 => x"05",
          5588 => x"70",
          5589 => x"33",
          5590 => x"05",
          5591 => x"18",
          5592 => x"33",
          5593 => x"33",
          5594 => x"1d",
          5595 => x"58",
          5596 => x"f7",
          5597 => x"e0",
          5598 => x"84",
          5599 => x"33",
          5600 => x"05",
          5601 => x"70",
          5602 => x"33",
          5603 => x"05",
          5604 => x"18",
          5605 => x"33",
          5606 => x"33",
          5607 => x"1d",
          5608 => x"58",
          5609 => x"ff",
          5610 => x"e6",
          5611 => x"8d",
          5612 => x"80",
          5613 => x"38",
          5614 => x"b9",
          5615 => x"d8",
          5616 => x"ce",
          5617 => x"84",
          5618 => x"ff",
          5619 => x"8d",
          5620 => x"40",
          5621 => x"2e",
          5622 => x"b9",
          5623 => x"75",
          5624 => x"81",
          5625 => x"38",
          5626 => x"33",
          5627 => x"ff",
          5628 => x"bc",
          5629 => x"5c",
          5630 => x"2e",
          5631 => x"84",
          5632 => x"40",
          5633 => x"f6",
          5634 => x"81",
          5635 => x"60",
          5636 => x"fe",
          5637 => x"26",
          5638 => x"07",
          5639 => x"f2",
          5640 => x"10",
          5641 => x"29",
          5642 => x"a3",
          5643 => x"70",
          5644 => x"87",
          5645 => x"05",
          5646 => x"58",
          5647 => x"8b",
          5648 => x"83",
          5649 => x"8b",
          5650 => x"f9",
          5651 => x"98",
          5652 => x"2b",
          5653 => x"2b",
          5654 => x"79",
          5655 => x"5f",
          5656 => x"27",
          5657 => x"77",
          5658 => x"59",
          5659 => x"70",
          5660 => x"0c",
          5661 => x"ee",
          5662 => x"80",
          5663 => x"ff",
          5664 => x"7e",
          5665 => x"60",
          5666 => x"83",
          5667 => x"7d",
          5668 => x"05",
          5669 => x"5a",
          5670 => x"8c",
          5671 => x"31",
          5672 => x"29",
          5673 => x"40",
          5674 => x"57",
          5675 => x"26",
          5676 => x"83",
          5677 => x"84",
          5678 => x"59",
          5679 => x"e0",
          5680 => x"79",
          5681 => x"05",
          5682 => x"17",
          5683 => x"26",
          5684 => x"a0",
          5685 => x"19",
          5686 => x"70",
          5687 => x"34",
          5688 => x"75",
          5689 => x"38",
          5690 => x"ff",
          5691 => x"ff",
          5692 => x"fe",
          5693 => x"f9",
          5694 => x"80",
          5695 => x"84",
          5696 => x"06",
          5697 => x"07",
          5698 => x"7b",
          5699 => x"09",
          5700 => x"38",
          5701 => x"83",
          5702 => x"81",
          5703 => x"ff",
          5704 => x"f5",
          5705 => x"f9",
          5706 => x"5e",
          5707 => x"1e",
          5708 => x"83",
          5709 => x"84",
          5710 => x"83",
          5711 => x"84",
          5712 => x"42",
          5713 => x"fa",
          5714 => x"f9",
          5715 => x"07",
          5716 => x"f9",
          5717 => x"18",
          5718 => x"06",
          5719 => x"fb",
          5720 => x"b8",
          5721 => x"06",
          5722 => x"75",
          5723 => x"34",
          5724 => x"f9",
          5725 => x"fb",
          5726 => x"56",
          5727 => x"b8",
          5728 => x"83",
          5729 => x"81",
          5730 => x"07",
          5731 => x"f9",
          5732 => x"39",
          5733 => x"33",
          5734 => x"90",
          5735 => x"83",
          5736 => x"ff",
          5737 => x"f1",
          5738 => x"b8",
          5739 => x"70",
          5740 => x"59",
          5741 => x"39",
          5742 => x"33",
          5743 => x"56",
          5744 => x"b8",
          5745 => x"39",
          5746 => x"33",
          5747 => x"90",
          5748 => x"83",
          5749 => x"fe",
          5750 => x"f9",
          5751 => x"ef",
          5752 => x"07",
          5753 => x"f9",
          5754 => x"ea",
          5755 => x"b8",
          5756 => x"06",
          5757 => x"56",
          5758 => x"b8",
          5759 => x"39",
          5760 => x"33",
          5761 => x"a0",
          5762 => x"83",
          5763 => x"fe",
          5764 => x"f9",
          5765 => x"fe",
          5766 => x"56",
          5767 => x"b8",
          5768 => x"39",
          5769 => x"33",
          5770 => x"84",
          5771 => x"83",
          5772 => x"fe",
          5773 => x"f9",
          5774 => x"fa",
          5775 => x"56",
          5776 => x"b8",
          5777 => x"39",
          5778 => x"33",
          5779 => x"56",
          5780 => x"b8",
          5781 => x"39",
          5782 => x"33",
          5783 => x"56",
          5784 => x"b8",
          5785 => x"39",
          5786 => x"33",
          5787 => x"56",
          5788 => x"b8",
          5789 => x"39",
          5790 => x"33",
          5791 => x"80",
          5792 => x"75",
          5793 => x"34",
          5794 => x"83",
          5795 => x"81",
          5796 => x"07",
          5797 => x"f9",
          5798 => x"ba",
          5799 => x"83",
          5800 => x"80",
          5801 => x"d2",
          5802 => x"ff",
          5803 => x"f4",
          5804 => x"bc",
          5805 => x"f5",
          5806 => x"bd",
          5807 => x"f6",
          5808 => x"83",
          5809 => x"80",
          5810 => x"88",
          5811 => x"39",
          5812 => x"b9",
          5813 => x"0b",
          5814 => x"0c",
          5815 => x"04",
          5816 => x"bd",
          5817 => x"bd",
          5818 => x"ff",
          5819 => x"05",
          5820 => x"39",
          5821 => x"42",
          5822 => x"11",
          5823 => x"51",
          5824 => x"3f",
          5825 => x"08",
          5826 => x"ba",
          5827 => x"b9",
          5828 => x"0b",
          5829 => x"34",
          5830 => x"ba",
          5831 => x"3d",
          5832 => x"83",
          5833 => x"ef",
          5834 => x"b9",
          5835 => x"11",
          5836 => x"84",
          5837 => x"7b",
          5838 => x"06",
          5839 => x"ca",
          5840 => x"b9",
          5841 => x"80",
          5842 => x"8c",
          5843 => x"80",
          5844 => x"bd",
          5845 => x"81",
          5846 => x"3f",
          5847 => x"33",
          5848 => x"06",
          5849 => x"56",
          5850 => x"80",
          5851 => x"bd",
          5852 => x"81",
          5853 => x"3f",
          5854 => x"8a",
          5855 => x"de",
          5856 => x"39",
          5857 => x"33",
          5858 => x"09",
          5859 => x"72",
          5860 => x"57",
          5861 => x"75",
          5862 => x"d9",
          5863 => x"80",
          5864 => x"60",
          5865 => x"38",
          5866 => x"bd",
          5867 => x"39",
          5868 => x"33",
          5869 => x"09",
          5870 => x"72",
          5871 => x"57",
          5872 => x"83",
          5873 => x"81",
          5874 => x"ff",
          5875 => x"59",
          5876 => x"78",
          5877 => x"38",
          5878 => x"bb",
          5879 => x"ff",
          5880 => x"ff",
          5881 => x"81",
          5882 => x"a6",
          5883 => x"bc",
          5884 => x"80",
          5885 => x"ff",
          5886 => x"bd",
          5887 => x"29",
          5888 => x"a0",
          5889 => x"f9",
          5890 => x"5f",
          5891 => x"05",
          5892 => x"ff",
          5893 => x"92",
          5894 => x"44",
          5895 => x"77",
          5896 => x"f5",
          5897 => x"ff",
          5898 => x"11",
          5899 => x"7b",
          5900 => x"38",
          5901 => x"33",
          5902 => x"27",
          5903 => x"ff",
          5904 => x"83",
          5905 => x"7c",
          5906 => x"ff",
          5907 => x"80",
          5908 => x"df",
          5909 => x"ff",
          5910 => x"76",
          5911 => x"38",
          5912 => x"75",
          5913 => x"34",
          5914 => x"06",
          5915 => x"22",
          5916 => x"5a",
          5917 => x"90",
          5918 => x"31",
          5919 => x"81",
          5920 => x"71",
          5921 => x"5f",
          5922 => x"a3",
          5923 => x"87",
          5924 => x"7c",
          5925 => x"7f",
          5926 => x"71",
          5927 => x"41",
          5928 => x"79",
          5929 => x"ea",
          5930 => x"de",
          5931 => x"e0",
          5932 => x"84",
          5933 => x"33",
          5934 => x"05",
          5935 => x"70",
          5936 => x"33",
          5937 => x"05",
          5938 => x"18",
          5939 => x"33",
          5940 => x"33",
          5941 => x"1d",
          5942 => x"58",
          5943 => x"ec",
          5944 => x"e0",
          5945 => x"84",
          5946 => x"33",
          5947 => x"05",
          5948 => x"70",
          5949 => x"33",
          5950 => x"05",
          5951 => x"18",
          5952 => x"33",
          5953 => x"33",
          5954 => x"1d",
          5955 => x"58",
          5956 => x"ff",
          5957 => x"fa",
          5958 => x"be",
          5959 => x"84",
          5960 => x"33",
          5961 => x"f9",
          5962 => x"b8",
          5963 => x"f9",
          5964 => x"b7",
          5965 => x"5c",
          5966 => x"e9",
          5967 => x"d2",
          5968 => x"ff",
          5969 => x"ff",
          5970 => x"5c",
          5971 => x"61",
          5972 => x"76",
          5973 => x"f9",
          5974 => x"81",
          5975 => x"19",
          5976 => x"7a",
          5977 => x"80",
          5978 => x"f9",
          5979 => x"b8",
          5980 => x"81",
          5981 => x"12",
          5982 => x"80",
          5983 => x"8d",
          5984 => x"75",
          5985 => x"34",
          5986 => x"83",
          5987 => x"81",
          5988 => x"80",
          5989 => x"59",
          5990 => x"7f",
          5991 => x"38",
          5992 => x"c5",
          5993 => x"2e",
          5994 => x"f4",
          5995 => x"f9",
          5996 => x"81",
          5997 => x"f9",
          5998 => x"44",
          5999 => x"76",
          6000 => x"81",
          6001 => x"38",
          6002 => x"ff",
          6003 => x"83",
          6004 => x"fd",
          6005 => x"1a",
          6006 => x"f9",
          6007 => x"e7",
          6008 => x"31",
          6009 => x"f9",
          6010 => x"90",
          6011 => x"58",
          6012 => x"26",
          6013 => x"80",
          6014 => x"05",
          6015 => x"f9",
          6016 => x"70",
          6017 => x"34",
          6018 => x"f4",
          6019 => x"76",
          6020 => x"58",
          6021 => x"b8",
          6022 => x"81",
          6023 => x"79",
          6024 => x"38",
          6025 => x"79",
          6026 => x"75",
          6027 => x"23",
          6028 => x"80",
          6029 => x"bc",
          6030 => x"39",
          6031 => x"ba",
          6032 => x"39",
          6033 => x"f9",
          6034 => x"8e",
          6035 => x"83",
          6036 => x"f1",
          6037 => x"f9",
          6038 => x"5a",
          6039 => x"1a",
          6040 => x"80",
          6041 => x"91",
          6042 => x"39",
          6043 => x"02",
          6044 => x"84",
          6045 => x"54",
          6046 => x"2e",
          6047 => x"51",
          6048 => x"80",
          6049 => x"8c",
          6050 => x"0d",
          6051 => x"73",
          6052 => x"3f",
          6053 => x"ba",
          6054 => x"3d",
          6055 => x"3d",
          6056 => x"05",
          6057 => x"0b",
          6058 => x"33",
          6059 => x"06",
          6060 => x"11",
          6061 => x"55",
          6062 => x"2e",
          6063 => x"81",
          6064 => x"83",
          6065 => x"74",
          6066 => x"ba",
          6067 => x"3d",
          6068 => x"f7",
          6069 => x"82",
          6070 => x"2e",
          6071 => x"73",
          6072 => x"71",
          6073 => x"70",
          6074 => x"5d",
          6075 => x"83",
          6076 => x"ff",
          6077 => x"7b",
          6078 => x"81",
          6079 => x"7b",
          6080 => x"32",
          6081 => x"80",
          6082 => x"5c",
          6083 => x"80",
          6084 => x"38",
          6085 => x"33",
          6086 => x"33",
          6087 => x"33",
          6088 => x"12",
          6089 => x"80",
          6090 => x"ba",
          6091 => x"5d",
          6092 => x"05",
          6093 => x"ff",
          6094 => x"91",
          6095 => x"55",
          6096 => x"2e",
          6097 => x"81",
          6098 => x"86",
          6099 => x"34",
          6100 => x"c0",
          6101 => x"87",
          6102 => x"08",
          6103 => x"2e",
          6104 => x"ee",
          6105 => x"57",
          6106 => x"bc",
          6107 => x"14",
          6108 => x"06",
          6109 => x"f9",
          6110 => x"38",
          6111 => x"f7",
          6112 => x"70",
          6113 => x"83",
          6114 => x"33",
          6115 => x"72",
          6116 => x"c1",
          6117 => x"ff",
          6118 => x"38",
          6119 => x"c0",
          6120 => x"81",
          6121 => x"79",
          6122 => x"85",
          6123 => x"83",
          6124 => x"34",
          6125 => x"14",
          6126 => x"b6",
          6127 => x"14",
          6128 => x"06",
          6129 => x"74",
          6130 => x"38",
          6131 => x"33",
          6132 => x"70",
          6133 => x"56",
          6134 => x"f7",
          6135 => x"81",
          6136 => x"86",
          6137 => x"70",
          6138 => x"54",
          6139 => x"2e",
          6140 => x"81",
          6141 => x"e5",
          6142 => x"81",
          6143 => x"80",
          6144 => x"38",
          6145 => x"f7",
          6146 => x"0b",
          6147 => x"33",
          6148 => x"08",
          6149 => x"33",
          6150 => x"e8",
          6151 => x"e7",
          6152 => x"42",
          6153 => x"56",
          6154 => x"16",
          6155 => x"81",
          6156 => x"38",
          6157 => x"16",
          6158 => x"80",
          6159 => x"38",
          6160 => x"16",
          6161 => x"81",
          6162 => x"38",
          6163 => x"16",
          6164 => x"81",
          6165 => x"81",
          6166 => x"73",
          6167 => x"8d",
          6168 => x"d4",
          6169 => x"72",
          6170 => x"da",
          6171 => x"ff",
          6172 => x"81",
          6173 => x"8c",
          6174 => x"d4",
          6175 => x"81",
          6176 => x"80",
          6177 => x"e0",
          6178 => x"05",
          6179 => x"9c",
          6180 => x"73",
          6181 => x"ec",
          6182 => x"87",
          6183 => x"08",
          6184 => x"0c",
          6185 => x"70",
          6186 => x"57",
          6187 => x"27",
          6188 => x"76",
          6189 => x"34",
          6190 => x"e8",
          6191 => x"19",
          6192 => x"26",
          6193 => x"72",
          6194 => x"c9",
          6195 => x"79",
          6196 => x"f8",
          6197 => x"73",
          6198 => x"38",
          6199 => x"87",
          6200 => x"08",
          6201 => x"7d",
          6202 => x"38",
          6203 => x"f8",
          6204 => x"54",
          6205 => x"83",
          6206 => x"73",
          6207 => x"34",
          6208 => x"9c",
          6209 => x"94",
          6210 => x"ff",
          6211 => x"81",
          6212 => x"83",
          6213 => x"33",
          6214 => x"88",
          6215 => x"34",
          6216 => x"fc",
          6217 => x"f7",
          6218 => x"72",
          6219 => x"9c",
          6220 => x"2e",
          6221 => x"80",
          6222 => x"81",
          6223 => x"8a",
          6224 => x"fe",
          6225 => x"74",
          6226 => x"59",
          6227 => x"9b",
          6228 => x"2e",
          6229 => x"83",
          6230 => x"81",
          6231 => x"38",
          6232 => x"80",
          6233 => x"81",
          6234 => x"87",
          6235 => x"98",
          6236 => x"72",
          6237 => x"38",
          6238 => x"9c",
          6239 => x"70",
          6240 => x"76",
          6241 => x"06",
          6242 => x"71",
          6243 => x"53",
          6244 => x"80",
          6245 => x"38",
          6246 => x"10",
          6247 => x"76",
          6248 => x"78",
          6249 => x"9c",
          6250 => x"5b",
          6251 => x"87",
          6252 => x"08",
          6253 => x"0c",
          6254 => x"39",
          6255 => x"81",
          6256 => x"38",
          6257 => x"06",
          6258 => x"39",
          6259 => x"9b",
          6260 => x"2e",
          6261 => x"80",
          6262 => x"82",
          6263 => x"72",
          6264 => x"e8",
          6265 => x"32",
          6266 => x"80",
          6267 => x"40",
          6268 => x"8a",
          6269 => x"2e",
          6270 => x"f9",
          6271 => x"ff",
          6272 => x"38",
          6273 => x"10",
          6274 => x"f8",
          6275 => x"33",
          6276 => x"7c",
          6277 => x"38",
          6278 => x"81",
          6279 => x"57",
          6280 => x"e2",
          6281 => x"83",
          6282 => x"80",
          6283 => x"38",
          6284 => x"33",
          6285 => x"91",
          6286 => x"ff",
          6287 => x"51",
          6288 => x"78",
          6289 => x"0c",
          6290 => x"04",
          6291 => x"81",
          6292 => x"f6",
          6293 => x"ff",
          6294 => x"83",
          6295 => x"33",
          6296 => x"7a",
          6297 => x"15",
          6298 => x"39",
          6299 => x"f7",
          6300 => x"ff",
          6301 => x"c0",
          6302 => x"0b",
          6303 => x"15",
          6304 => x"39",
          6305 => x"06",
          6306 => x"ff",
          6307 => x"38",
          6308 => x"16",
          6309 => x"75",
          6310 => x"38",
          6311 => x"06",
          6312 => x"2e",
          6313 => x"fb",
          6314 => x"f7",
          6315 => x"fa",
          6316 => x"98",
          6317 => x"55",
          6318 => x"fb",
          6319 => x"c0",
          6320 => x"83",
          6321 => x"76",
          6322 => x"59",
          6323 => x"ff",
          6324 => x"c0",
          6325 => x"ca",
          6326 => x"f7",
          6327 => x"09",
          6328 => x"72",
          6329 => x"72",
          6330 => x"34",
          6331 => x"f7",
          6332 => x"f7",
          6333 => x"f7",
          6334 => x"83",
          6335 => x"83",
          6336 => x"5d",
          6337 => x"5c",
          6338 => x"9c",
          6339 => x"2e",
          6340 => x"fc",
          6341 => x"59",
          6342 => x"fc",
          6343 => x"81",
          6344 => x"06",
          6345 => x"fd",
          6346 => x"76",
          6347 => x"54",
          6348 => x"80",
          6349 => x"83",
          6350 => x"75",
          6351 => x"54",
          6352 => x"83",
          6353 => x"f7",
          6354 => x"0b",
          6355 => x"33",
          6356 => x"83",
          6357 => x"73",
          6358 => x"34",
          6359 => x"95",
          6360 => x"83",
          6361 => x"84",
          6362 => x"38",
          6363 => x"f7",
          6364 => x"ff",
          6365 => x"ff",
          6366 => x"ff",
          6367 => x"57",
          6368 => x"79",
          6369 => x"80",
          6370 => x"f9",
          6371 => x"81",
          6372 => x"15",
          6373 => x"73",
          6374 => x"80",
          6375 => x"f9",
          6376 => x"b8",
          6377 => x"81",
          6378 => x"ff",
          6379 => x"75",
          6380 => x"80",
          6381 => x"f9",
          6382 => x"59",
          6383 => x"81",
          6384 => x"ff",
          6385 => x"ff",
          6386 => x"39",
          6387 => x"95",
          6388 => x"08",
          6389 => x"f0",
          6390 => x"eb",
          6391 => x"83",
          6392 => x"83",
          6393 => x"59",
          6394 => x"80",
          6395 => x"51",
          6396 => x"82",
          6397 => x"f9",
          6398 => x"0b",
          6399 => x"08",
          6400 => x"a7",
          6401 => x"14",
          6402 => x"98",
          6403 => x"e0",
          6404 => x"0b",
          6405 => x"08",
          6406 => x"0b",
          6407 => x"80",
          6408 => x"80",
          6409 => x"c0",
          6410 => x"83",
          6411 => x"56",
          6412 => x"05",
          6413 => x"98",
          6414 => x"87",
          6415 => x"08",
          6416 => x"2e",
          6417 => x"15",
          6418 => x"98",
          6419 => x"53",
          6420 => x"87",
          6421 => x"fe",
          6422 => x"87",
          6423 => x"08",
          6424 => x"71",
          6425 => x"cd",
          6426 => x"72",
          6427 => x"c5",
          6428 => x"98",
          6429 => x"ce",
          6430 => x"87",
          6431 => x"08",
          6432 => x"98",
          6433 => x"75",
          6434 => x"38",
          6435 => x"87",
          6436 => x"08",
          6437 => x"74",
          6438 => x"72",
          6439 => x"db",
          6440 => x"98",
          6441 => x"ff",
          6442 => x"27",
          6443 => x"56",
          6444 => x"9d",
          6445 => x"2e",
          6446 => x"81",
          6447 => x"72",
          6448 => x"75",
          6449 => x"38",
          6450 => x"8c",
          6451 => x"0d",
          6452 => x"70",
          6453 => x"58",
          6454 => x"38",
          6455 => x"e4",
          6456 => x"fe",
          6457 => x"77",
          6458 => x"0c",
          6459 => x"04",
          6460 => x"7a",
          6461 => x"a7",
          6462 => x"53",
          6463 => x"f4",
          6464 => x"88",
          6465 => x"80",
          6466 => x"76",
          6467 => x"51",
          6468 => x"72",
          6469 => x"73",
          6470 => x"71",
          6471 => x"72",
          6472 => x"76",
          6473 => x"73",
          6474 => x"83",
          6475 => x"53",
          6476 => x"34",
          6477 => x"08",
          6478 => x"72",
          6479 => x"83",
          6480 => x"56",
          6481 => x"81",
          6482 => x"0b",
          6483 => x"e8",
          6484 => x"98",
          6485 => x"f4",
          6486 => x"80",
          6487 => x"54",
          6488 => x"9c",
          6489 => x"c0",
          6490 => x"52",
          6491 => x"f6",
          6492 => x"33",
          6493 => x"9c",
          6494 => x"75",
          6495 => x"38",
          6496 => x"2e",
          6497 => x"c0",
          6498 => x"52",
          6499 => x"74",
          6500 => x"38",
          6501 => x"ff",
          6502 => x"38",
          6503 => x"9c",
          6504 => x"90",
          6505 => x"c0",
          6506 => x"53",
          6507 => x"9c",
          6508 => x"73",
          6509 => x"81",
          6510 => x"c0",
          6511 => x"53",
          6512 => x"27",
          6513 => x"81",
          6514 => x"38",
          6515 => x"a4",
          6516 => x"56",
          6517 => x"80",
          6518 => x"56",
          6519 => x"80",
          6520 => x"80",
          6521 => x"38",
          6522 => x"06",
          6523 => x"d5",
          6524 => x"71",
          6525 => x"57",
          6526 => x"80",
          6527 => x"84",
          6528 => x"53",
          6529 => x"27",
          6530 => x"70",
          6531 => x"33",
          6532 => x"05",
          6533 => x"72",
          6534 => x"77",
          6535 => x"0c",
          6536 => x"04",
          6537 => x"e4",
          6538 => x"fe",
          6539 => x"77",
          6540 => x"0c",
          6541 => x"04",
          6542 => x"81",
          6543 => x"54",
          6544 => x"38",
          6545 => x"ab",
          6546 => x"0d",
          6547 => x"05",
          6548 => x"57",
          6549 => x"83",
          6550 => x"78",
          6551 => x"fc",
          6552 => x"70",
          6553 => x"07",
          6554 => x"58",
          6555 => x"34",
          6556 => x"52",
          6557 => x"34",
          6558 => x"53",
          6559 => x"34",
          6560 => x"34",
          6561 => x"98",
          6562 => x"11",
          6563 => x"57",
          6564 => x"71",
          6565 => x"38",
          6566 => x"05",
          6567 => x"70",
          6568 => x"34",
          6569 => x"f0",
          6570 => x"98",
          6571 => x"82",
          6572 => x"f4",
          6573 => x"80",
          6574 => x"85",
          6575 => x"98",
          6576 => x"fe",
          6577 => x"34",
          6578 => x"f0",
          6579 => x"87",
          6580 => x"08",
          6581 => x"08",
          6582 => x"90",
          6583 => x"c0",
          6584 => x"53",
          6585 => x"9c",
          6586 => x"73",
          6587 => x"81",
          6588 => x"c0",
          6589 => x"57",
          6590 => x"27",
          6591 => x"81",
          6592 => x"38",
          6593 => x"a4",
          6594 => x"56",
          6595 => x"80",
          6596 => x"56",
          6597 => x"80",
          6598 => x"c0",
          6599 => x"80",
          6600 => x"54",
          6601 => x"9c",
          6602 => x"c0",
          6603 => x"56",
          6604 => x"f6",
          6605 => x"33",
          6606 => x"9c",
          6607 => x"71",
          6608 => x"38",
          6609 => x"2e",
          6610 => x"c0",
          6611 => x"52",
          6612 => x"74",
          6613 => x"72",
          6614 => x"2e",
          6615 => x"80",
          6616 => x"75",
          6617 => x"53",
          6618 => x"38",
          6619 => x"ff",
          6620 => x"74",
          6621 => x"84",
          6622 => x"89",
          6623 => x"ff",
          6624 => x"ff",
          6625 => x"76",
          6626 => x"70",
          6627 => x"56",
          6628 => x"2e",
          6629 => x"0b",
          6630 => x"52",
          6631 => x"d3",
          6632 => x"ba",
          6633 => x"3d",
          6634 => x"3d",
          6635 => x"98",
          6636 => x"d0",
          6637 => x"0b",
          6638 => x"08",
          6639 => x"0b",
          6640 => x"80",
          6641 => x"80",
          6642 => x"c0",
          6643 => x"83",
          6644 => x"56",
          6645 => x"05",
          6646 => x"98",
          6647 => x"87",
          6648 => x"08",
          6649 => x"2e",
          6650 => x"15",
          6651 => x"98",
          6652 => x"52",
          6653 => x"87",
          6654 => x"fe",
          6655 => x"87",
          6656 => x"08",
          6657 => x"70",
          6658 => x"cd",
          6659 => x"71",
          6660 => x"c5",
          6661 => x"98",
          6662 => x"ce",
          6663 => x"87",
          6664 => x"08",
          6665 => x"98",
          6666 => x"72",
          6667 => x"38",
          6668 => x"87",
          6669 => x"08",
          6670 => x"74",
          6671 => x"71",
          6672 => x"db",
          6673 => x"98",
          6674 => x"ff",
          6675 => x"27",
          6676 => x"53",
          6677 => x"91",
          6678 => x"2e",
          6679 => x"81",
          6680 => x"71",
          6681 => x"ff",
          6682 => x"70",
          6683 => x"57",
          6684 => x"80",
          6685 => x"e5",
          6686 => x"cf",
          6687 => x"3d",
          6688 => x"3d",
          6689 => x"fc",
          6690 => x"31",
          6691 => x"83",
          6692 => x"70",
          6693 => x"11",
          6694 => x"12",
          6695 => x"2b",
          6696 => x"07",
          6697 => x"33",
          6698 => x"71",
          6699 => x"90",
          6700 => x"54",
          6701 => x"5d",
          6702 => x"56",
          6703 => x"71",
          6704 => x"38",
          6705 => x"11",
          6706 => x"33",
          6707 => x"71",
          6708 => x"76",
          6709 => x"81",
          6710 => x"98",
          6711 => x"2b",
          6712 => x"5c",
          6713 => x"52",
          6714 => x"83",
          6715 => x"13",
          6716 => x"33",
          6717 => x"71",
          6718 => x"75",
          6719 => x"2a",
          6720 => x"57",
          6721 => x"34",
          6722 => x"06",
          6723 => x"13",
          6724 => x"fc",
          6725 => x"84",
          6726 => x"13",
          6727 => x"2b",
          6728 => x"2a",
          6729 => x"54",
          6730 => x"14",
          6731 => x"14",
          6732 => x"fc",
          6733 => x"80",
          6734 => x"34",
          6735 => x"13",
          6736 => x"fc",
          6737 => x"84",
          6738 => x"85",
          6739 => x"b9",
          6740 => x"70",
          6741 => x"33",
          6742 => x"07",
          6743 => x"07",
          6744 => x"58",
          6745 => x"74",
          6746 => x"81",
          6747 => x"3d",
          6748 => x"12",
          6749 => x"33",
          6750 => x"71",
          6751 => x"75",
          6752 => x"33",
          6753 => x"71",
          6754 => x"70",
          6755 => x"58",
          6756 => x"58",
          6757 => x"12",
          6758 => x"12",
          6759 => x"fc",
          6760 => x"84",
          6761 => x"12",
          6762 => x"2b",
          6763 => x"07",
          6764 => x"52",
          6765 => x"12",
          6766 => x"33",
          6767 => x"07",
          6768 => x"52",
          6769 => x"77",
          6770 => x"72",
          6771 => x"84",
          6772 => x"15",
          6773 => x"12",
          6774 => x"2b",
          6775 => x"ff",
          6776 => x"2a",
          6777 => x"52",
          6778 => x"77",
          6779 => x"84",
          6780 => x"70",
          6781 => x"81",
          6782 => x"8b",
          6783 => x"2b",
          6784 => x"70",
          6785 => x"33",
          6786 => x"07",
          6787 => x"8f",
          6788 => x"77",
          6789 => x"2a",
          6790 => x"54",
          6791 => x"54",
          6792 => x"14",
          6793 => x"14",
          6794 => x"fc",
          6795 => x"70",
          6796 => x"33",
          6797 => x"71",
          6798 => x"74",
          6799 => x"81",
          6800 => x"88",
          6801 => x"ff",
          6802 => x"88",
          6803 => x"53",
          6804 => x"54",
          6805 => x"34",
          6806 => x"34",
          6807 => x"08",
          6808 => x"11",
          6809 => x"33",
          6810 => x"71",
          6811 => x"74",
          6812 => x"81",
          6813 => x"98",
          6814 => x"2b",
          6815 => x"5d",
          6816 => x"53",
          6817 => x"25",
          6818 => x"71",
          6819 => x"33",
          6820 => x"07",
          6821 => x"07",
          6822 => x"59",
          6823 => x"75",
          6824 => x"16",
          6825 => x"fc",
          6826 => x"70",
          6827 => x"33",
          6828 => x"71",
          6829 => x"74",
          6830 => x"33",
          6831 => x"71",
          6832 => x"70",
          6833 => x"5c",
          6834 => x"56",
          6835 => x"82",
          6836 => x"83",
          6837 => x"3d",
          6838 => x"3d",
          6839 => x"b9",
          6840 => x"58",
          6841 => x"8f",
          6842 => x"2e",
          6843 => x"51",
          6844 => x"89",
          6845 => x"84",
          6846 => x"84",
          6847 => x"a0",
          6848 => x"b9",
          6849 => x"80",
          6850 => x"52",
          6851 => x"51",
          6852 => x"3f",
          6853 => x"08",
          6854 => x"34",
          6855 => x"16",
          6856 => x"fc",
          6857 => x"84",
          6858 => x"0b",
          6859 => x"84",
          6860 => x"56",
          6861 => x"34",
          6862 => x"17",
          6863 => x"fc",
          6864 => x"f8",
          6865 => x"fe",
          6866 => x"70",
          6867 => x"06",
          6868 => x"58",
          6869 => x"74",
          6870 => x"73",
          6871 => x"84",
          6872 => x"70",
          6873 => x"84",
          6874 => x"05",
          6875 => x"55",
          6876 => x"34",
          6877 => x"15",
          6878 => x"39",
          6879 => x"7b",
          6880 => x"81",
          6881 => x"27",
          6882 => x"12",
          6883 => x"05",
          6884 => x"ff",
          6885 => x"70",
          6886 => x"06",
          6887 => x"08",
          6888 => x"85",
          6889 => x"88",
          6890 => x"52",
          6891 => x"55",
          6892 => x"54",
          6893 => x"80",
          6894 => x"10",
          6895 => x"70",
          6896 => x"33",
          6897 => x"07",
          6898 => x"ff",
          6899 => x"70",
          6900 => x"06",
          6901 => x"56",
          6902 => x"54",
          6903 => x"27",
          6904 => x"80",
          6905 => x"75",
          6906 => x"84",
          6907 => x"13",
          6908 => x"2b",
          6909 => x"75",
          6910 => x"81",
          6911 => x"85",
          6912 => x"54",
          6913 => x"83",
          6914 => x"70",
          6915 => x"33",
          6916 => x"07",
          6917 => x"ff",
          6918 => x"5d",
          6919 => x"70",
          6920 => x"38",
          6921 => x"51",
          6922 => x"82",
          6923 => x"51",
          6924 => x"82",
          6925 => x"75",
          6926 => x"38",
          6927 => x"83",
          6928 => x"74",
          6929 => x"07",
          6930 => x"5b",
          6931 => x"5a",
          6932 => x"78",
          6933 => x"84",
          6934 => x"15",
          6935 => x"53",
          6936 => x"14",
          6937 => x"14",
          6938 => x"fc",
          6939 => x"70",
          6940 => x"33",
          6941 => x"07",
          6942 => x"8f",
          6943 => x"74",
          6944 => x"ff",
          6945 => x"88",
          6946 => x"53",
          6947 => x"52",
          6948 => x"34",
          6949 => x"06",
          6950 => x"12",
          6951 => x"fc",
          6952 => x"75",
          6953 => x"81",
          6954 => x"b9",
          6955 => x"19",
          6956 => x"87",
          6957 => x"8b",
          6958 => x"2b",
          6959 => x"58",
          6960 => x"57",
          6961 => x"34",
          6962 => x"34",
          6963 => x"08",
          6964 => x"78",
          6965 => x"33",
          6966 => x"71",
          6967 => x"70",
          6968 => x"54",
          6969 => x"86",
          6970 => x"87",
          6971 => x"b9",
          6972 => x"19",
          6973 => x"85",
          6974 => x"8b",
          6975 => x"2b",
          6976 => x"58",
          6977 => x"52",
          6978 => x"34",
          6979 => x"34",
          6980 => x"08",
          6981 => x"78",
          6982 => x"33",
          6983 => x"71",
          6984 => x"70",
          6985 => x"5c",
          6986 => x"84",
          6987 => x"85",
          6988 => x"b9",
          6989 => x"84",
          6990 => x"84",
          6991 => x"8b",
          6992 => x"86",
          6993 => x"15",
          6994 => x"2b",
          6995 => x"07",
          6996 => x"17",
          6997 => x"33",
          6998 => x"07",
          6999 => x"5a",
          7000 => x"54",
          7001 => x"12",
          7002 => x"12",
          7003 => x"fc",
          7004 => x"84",
          7005 => x"12",
          7006 => x"2b",
          7007 => x"07",
          7008 => x"14",
          7009 => x"33",
          7010 => x"07",
          7011 => x"58",
          7012 => x"56",
          7013 => x"70",
          7014 => x"76",
          7015 => x"84",
          7016 => x"18",
          7017 => x"12",
          7018 => x"2b",
          7019 => x"ff",
          7020 => x"2a",
          7021 => x"57",
          7022 => x"74",
          7023 => x"84",
          7024 => x"18",
          7025 => x"fe",
          7026 => x"3d",
          7027 => x"b9",
          7028 => x"58",
          7029 => x"a0",
          7030 => x"77",
          7031 => x"84",
          7032 => x"89",
          7033 => x"77",
          7034 => x"3f",
          7035 => x"08",
          7036 => x"0c",
          7037 => x"04",
          7038 => x"0b",
          7039 => x"0c",
          7040 => x"84",
          7041 => x"82",
          7042 => x"76",
          7043 => x"f4",
          7044 => x"eb",
          7045 => x"fc",
          7046 => x"75",
          7047 => x"81",
          7048 => x"b9",
          7049 => x"76",
          7050 => x"81",
          7051 => x"34",
          7052 => x"08",
          7053 => x"17",
          7054 => x"87",
          7055 => x"b9",
          7056 => x"b9",
          7057 => x"05",
          7058 => x"07",
          7059 => x"ff",
          7060 => x"2a",
          7061 => x"56",
          7062 => x"34",
          7063 => x"34",
          7064 => x"22",
          7065 => x"10",
          7066 => x"08",
          7067 => x"55",
          7068 => x"15",
          7069 => x"83",
          7070 => x"54",
          7071 => x"fe",
          7072 => x"e3",
          7073 => x"0d",
          7074 => x"5f",
          7075 => x"b9",
          7076 => x"45",
          7077 => x"2e",
          7078 => x"7e",
          7079 => x"af",
          7080 => x"2e",
          7081 => x"81",
          7082 => x"27",
          7083 => x"fb",
          7084 => x"82",
          7085 => x"ff",
          7086 => x"58",
          7087 => x"ff",
          7088 => x"31",
          7089 => x"83",
          7090 => x"70",
          7091 => x"11",
          7092 => x"12",
          7093 => x"2b",
          7094 => x"31",
          7095 => x"ff",
          7096 => x"10",
          7097 => x"73",
          7098 => x"11",
          7099 => x"12",
          7100 => x"2b",
          7101 => x"2b",
          7102 => x"53",
          7103 => x"44",
          7104 => x"44",
          7105 => x"52",
          7106 => x"80",
          7107 => x"fd",
          7108 => x"33",
          7109 => x"71",
          7110 => x"70",
          7111 => x"19",
          7112 => x"12",
          7113 => x"2b",
          7114 => x"07",
          7115 => x"56",
          7116 => x"74",
          7117 => x"38",
          7118 => x"82",
          7119 => x"1b",
          7120 => x"2e",
          7121 => x"60",
          7122 => x"f9",
          7123 => x"58",
          7124 => x"87",
          7125 => x"18",
          7126 => x"24",
          7127 => x"76",
          7128 => x"81",
          7129 => x"8b",
          7130 => x"2b",
          7131 => x"70",
          7132 => x"33",
          7133 => x"71",
          7134 => x"47",
          7135 => x"53",
          7136 => x"80",
          7137 => x"ba",
          7138 => x"82",
          7139 => x"12",
          7140 => x"2b",
          7141 => x"07",
          7142 => x"11",
          7143 => x"33",
          7144 => x"71",
          7145 => x"7e",
          7146 => x"33",
          7147 => x"71",
          7148 => x"70",
          7149 => x"57",
          7150 => x"41",
          7151 => x"59",
          7152 => x"1d",
          7153 => x"1d",
          7154 => x"fc",
          7155 => x"84",
          7156 => x"12",
          7157 => x"2b",
          7158 => x"07",
          7159 => x"14",
          7160 => x"33",
          7161 => x"07",
          7162 => x"5f",
          7163 => x"40",
          7164 => x"77",
          7165 => x"7b",
          7166 => x"84",
          7167 => x"16",
          7168 => x"12",
          7169 => x"2b",
          7170 => x"ff",
          7171 => x"2a",
          7172 => x"59",
          7173 => x"79",
          7174 => x"84",
          7175 => x"70",
          7176 => x"33",
          7177 => x"71",
          7178 => x"83",
          7179 => x"05",
          7180 => x"15",
          7181 => x"2b",
          7182 => x"2a",
          7183 => x"5d",
          7184 => x"55",
          7185 => x"75",
          7186 => x"84",
          7187 => x"70",
          7188 => x"81",
          7189 => x"8b",
          7190 => x"2b",
          7191 => x"82",
          7192 => x"15",
          7193 => x"2b",
          7194 => x"2a",
          7195 => x"5d",
          7196 => x"55",
          7197 => x"34",
          7198 => x"34",
          7199 => x"08",
          7200 => x"11",
          7201 => x"33",
          7202 => x"07",
          7203 => x"56",
          7204 => x"42",
          7205 => x"7e",
          7206 => x"51",
          7207 => x"3f",
          7208 => x"08",
          7209 => x"61",
          7210 => x"70",
          7211 => x"06",
          7212 => x"7a",
          7213 => x"b6",
          7214 => x"73",
          7215 => x"0c",
          7216 => x"04",
          7217 => x"0b",
          7218 => x"0c",
          7219 => x"84",
          7220 => x"82",
          7221 => x"60",
          7222 => x"f4",
          7223 => x"9f",
          7224 => x"fc",
          7225 => x"7e",
          7226 => x"81",
          7227 => x"b9",
          7228 => x"60",
          7229 => x"81",
          7230 => x"34",
          7231 => x"08",
          7232 => x"1d",
          7233 => x"87",
          7234 => x"b9",
          7235 => x"b9",
          7236 => x"05",
          7237 => x"07",
          7238 => x"ff",
          7239 => x"2a",
          7240 => x"57",
          7241 => x"34",
          7242 => x"34",
          7243 => x"22",
          7244 => x"10",
          7245 => x"08",
          7246 => x"55",
          7247 => x"15",
          7248 => x"83",
          7249 => x"b9",
          7250 => x"7e",
          7251 => x"76",
          7252 => x"8c",
          7253 => x"7f",
          7254 => x"df",
          7255 => x"f4",
          7256 => x"ba",
          7257 => x"ba",
          7258 => x"3d",
          7259 => x"1c",
          7260 => x"08",
          7261 => x"71",
          7262 => x"7f",
          7263 => x"81",
          7264 => x"88",
          7265 => x"ff",
          7266 => x"88",
          7267 => x"5b",
          7268 => x"7b",
          7269 => x"1c",
          7270 => x"b9",
          7271 => x"7c",
          7272 => x"58",
          7273 => x"34",
          7274 => x"34",
          7275 => x"08",
          7276 => x"33",
          7277 => x"71",
          7278 => x"70",
          7279 => x"ff",
          7280 => x"05",
          7281 => x"ff",
          7282 => x"2a",
          7283 => x"57",
          7284 => x"63",
          7285 => x"34",
          7286 => x"06",
          7287 => x"83",
          7288 => x"b9",
          7289 => x"5b",
          7290 => x"60",
          7291 => x"61",
          7292 => x"08",
          7293 => x"51",
          7294 => x"7e",
          7295 => x"39",
          7296 => x"70",
          7297 => x"06",
          7298 => x"ac",
          7299 => x"ff",
          7300 => x"31",
          7301 => x"ff",
          7302 => x"33",
          7303 => x"71",
          7304 => x"70",
          7305 => x"1b",
          7306 => x"12",
          7307 => x"2b",
          7308 => x"07",
          7309 => x"54",
          7310 => x"54",
          7311 => x"f9",
          7312 => x"bc",
          7313 => x"24",
          7314 => x"80",
          7315 => x"8f",
          7316 => x"ff",
          7317 => x"61",
          7318 => x"dd",
          7319 => x"39",
          7320 => x"0b",
          7321 => x"0c",
          7322 => x"84",
          7323 => x"82",
          7324 => x"7e",
          7325 => x"f4",
          7326 => x"83",
          7327 => x"fc",
          7328 => x"7a",
          7329 => x"81",
          7330 => x"b9",
          7331 => x"7e",
          7332 => x"81",
          7333 => x"34",
          7334 => x"08",
          7335 => x"19",
          7336 => x"87",
          7337 => x"b9",
          7338 => x"b9",
          7339 => x"05",
          7340 => x"07",
          7341 => x"ff",
          7342 => x"2a",
          7343 => x"44",
          7344 => x"05",
          7345 => x"89",
          7346 => x"b9",
          7347 => x"10",
          7348 => x"b9",
          7349 => x"f8",
          7350 => x"7e",
          7351 => x"34",
          7352 => x"05",
          7353 => x"39",
          7354 => x"83",
          7355 => x"83",
          7356 => x"5b",
          7357 => x"fb",
          7358 => x"f2",
          7359 => x"2e",
          7360 => x"7e",
          7361 => x"3f",
          7362 => x"84",
          7363 => x"95",
          7364 => x"76",
          7365 => x"33",
          7366 => x"71",
          7367 => x"83",
          7368 => x"11",
          7369 => x"87",
          7370 => x"8b",
          7371 => x"2b",
          7372 => x"84",
          7373 => x"15",
          7374 => x"2b",
          7375 => x"2a",
          7376 => x"56",
          7377 => x"53",
          7378 => x"78",
          7379 => x"34",
          7380 => x"05",
          7381 => x"fc",
          7382 => x"84",
          7383 => x"12",
          7384 => x"2b",
          7385 => x"07",
          7386 => x"14",
          7387 => x"33",
          7388 => x"07",
          7389 => x"5b",
          7390 => x"5d",
          7391 => x"73",
          7392 => x"34",
          7393 => x"05",
          7394 => x"fc",
          7395 => x"33",
          7396 => x"71",
          7397 => x"81",
          7398 => x"70",
          7399 => x"5c",
          7400 => x"7d",
          7401 => x"1e",
          7402 => x"fc",
          7403 => x"82",
          7404 => x"12",
          7405 => x"2b",
          7406 => x"07",
          7407 => x"33",
          7408 => x"71",
          7409 => x"70",
          7410 => x"5c",
          7411 => x"57",
          7412 => x"7c",
          7413 => x"1d",
          7414 => x"fc",
          7415 => x"70",
          7416 => x"33",
          7417 => x"71",
          7418 => x"74",
          7419 => x"33",
          7420 => x"71",
          7421 => x"70",
          7422 => x"47",
          7423 => x"5c",
          7424 => x"82",
          7425 => x"83",
          7426 => x"b9",
          7427 => x"1f",
          7428 => x"83",
          7429 => x"88",
          7430 => x"57",
          7431 => x"83",
          7432 => x"58",
          7433 => x"84",
          7434 => x"bd",
          7435 => x"b9",
          7436 => x"84",
          7437 => x"ff",
          7438 => x"5f",
          7439 => x"84",
          7440 => x"84",
          7441 => x"a0",
          7442 => x"b9",
          7443 => x"80",
          7444 => x"52",
          7445 => x"51",
          7446 => x"3f",
          7447 => x"08",
          7448 => x"34",
          7449 => x"17",
          7450 => x"fc",
          7451 => x"84",
          7452 => x"0b",
          7453 => x"84",
          7454 => x"54",
          7455 => x"34",
          7456 => x"15",
          7457 => x"fc",
          7458 => x"f8",
          7459 => x"fe",
          7460 => x"70",
          7461 => x"06",
          7462 => x"45",
          7463 => x"61",
          7464 => x"60",
          7465 => x"84",
          7466 => x"70",
          7467 => x"84",
          7468 => x"05",
          7469 => x"5d",
          7470 => x"34",
          7471 => x"1c",
          7472 => x"e7",
          7473 => x"54",
          7474 => x"86",
          7475 => x"1a",
          7476 => x"2b",
          7477 => x"07",
          7478 => x"1c",
          7479 => x"33",
          7480 => x"07",
          7481 => x"5c",
          7482 => x"59",
          7483 => x"84",
          7484 => x"61",
          7485 => x"84",
          7486 => x"70",
          7487 => x"33",
          7488 => x"71",
          7489 => x"83",
          7490 => x"05",
          7491 => x"87",
          7492 => x"88",
          7493 => x"88",
          7494 => x"48",
          7495 => x"59",
          7496 => x"86",
          7497 => x"64",
          7498 => x"84",
          7499 => x"1d",
          7500 => x"12",
          7501 => x"2b",
          7502 => x"ff",
          7503 => x"2a",
          7504 => x"58",
          7505 => x"7f",
          7506 => x"84",
          7507 => x"70",
          7508 => x"81",
          7509 => x"8b",
          7510 => x"2b",
          7511 => x"70",
          7512 => x"33",
          7513 => x"07",
          7514 => x"8f",
          7515 => x"77",
          7516 => x"2a",
          7517 => x"5a",
          7518 => x"44",
          7519 => x"17",
          7520 => x"17",
          7521 => x"fc",
          7522 => x"70",
          7523 => x"33",
          7524 => x"71",
          7525 => x"74",
          7526 => x"81",
          7527 => x"88",
          7528 => x"ff",
          7529 => x"88",
          7530 => x"5e",
          7531 => x"41",
          7532 => x"34",
          7533 => x"05",
          7534 => x"ff",
          7535 => x"fa",
          7536 => x"15",
          7537 => x"33",
          7538 => x"71",
          7539 => x"79",
          7540 => x"33",
          7541 => x"71",
          7542 => x"70",
          7543 => x"5e",
          7544 => x"5d",
          7545 => x"34",
          7546 => x"34",
          7547 => x"08",
          7548 => x"11",
          7549 => x"33",
          7550 => x"71",
          7551 => x"74",
          7552 => x"33",
          7553 => x"71",
          7554 => x"70",
          7555 => x"56",
          7556 => x"42",
          7557 => x"60",
          7558 => x"75",
          7559 => x"34",
          7560 => x"08",
          7561 => x"81",
          7562 => x"88",
          7563 => x"ff",
          7564 => x"88",
          7565 => x"58",
          7566 => x"34",
          7567 => x"34",
          7568 => x"08",
          7569 => x"33",
          7570 => x"71",
          7571 => x"83",
          7572 => x"05",
          7573 => x"12",
          7574 => x"2b",
          7575 => x"2b",
          7576 => x"06",
          7577 => x"88",
          7578 => x"5f",
          7579 => x"42",
          7580 => x"82",
          7581 => x"83",
          7582 => x"b9",
          7583 => x"1f",
          7584 => x"12",
          7585 => x"2b",
          7586 => x"07",
          7587 => x"33",
          7588 => x"71",
          7589 => x"81",
          7590 => x"70",
          7591 => x"54",
          7592 => x"59",
          7593 => x"7c",
          7594 => x"1d",
          7595 => x"fc",
          7596 => x"82",
          7597 => x"12",
          7598 => x"2b",
          7599 => x"07",
          7600 => x"11",
          7601 => x"33",
          7602 => x"71",
          7603 => x"78",
          7604 => x"33",
          7605 => x"71",
          7606 => x"70",
          7607 => x"57",
          7608 => x"42",
          7609 => x"5a",
          7610 => x"84",
          7611 => x"85",
          7612 => x"b9",
          7613 => x"17",
          7614 => x"85",
          7615 => x"8b",
          7616 => x"2b",
          7617 => x"86",
          7618 => x"15",
          7619 => x"2b",
          7620 => x"2a",
          7621 => x"52",
          7622 => x"57",
          7623 => x"34",
          7624 => x"34",
          7625 => x"08",
          7626 => x"81",
          7627 => x"88",
          7628 => x"ff",
          7629 => x"88",
          7630 => x"5e",
          7631 => x"34",
          7632 => x"34",
          7633 => x"08",
          7634 => x"11",
          7635 => x"33",
          7636 => x"71",
          7637 => x"74",
          7638 => x"81",
          7639 => x"88",
          7640 => x"88",
          7641 => x"45",
          7642 => x"55",
          7643 => x"34",
          7644 => x"34",
          7645 => x"08",
          7646 => x"33",
          7647 => x"71",
          7648 => x"83",
          7649 => x"05",
          7650 => x"83",
          7651 => x"88",
          7652 => x"88",
          7653 => x"45",
          7654 => x"55",
          7655 => x"1a",
          7656 => x"1a",
          7657 => x"fc",
          7658 => x"82",
          7659 => x"12",
          7660 => x"2b",
          7661 => x"62",
          7662 => x"2b",
          7663 => x"5d",
          7664 => x"05",
          7665 => x"fa",
          7666 => x"fc",
          7667 => x"05",
          7668 => x"1c",
          7669 => x"ff",
          7670 => x"5f",
          7671 => x"86",
          7672 => x"1a",
          7673 => x"2b",
          7674 => x"07",
          7675 => x"1c",
          7676 => x"33",
          7677 => x"07",
          7678 => x"40",
          7679 => x"41",
          7680 => x"84",
          7681 => x"61",
          7682 => x"84",
          7683 => x"70",
          7684 => x"33",
          7685 => x"71",
          7686 => x"83",
          7687 => x"05",
          7688 => x"87",
          7689 => x"88",
          7690 => x"88",
          7691 => x"5f",
          7692 => x"41",
          7693 => x"86",
          7694 => x"64",
          7695 => x"84",
          7696 => x"1d",
          7697 => x"12",
          7698 => x"2b",
          7699 => x"ff",
          7700 => x"2a",
          7701 => x"55",
          7702 => x"7c",
          7703 => x"84",
          7704 => x"70",
          7705 => x"81",
          7706 => x"8b",
          7707 => x"2b",
          7708 => x"70",
          7709 => x"33",
          7710 => x"07",
          7711 => x"8f",
          7712 => x"77",
          7713 => x"2a",
          7714 => x"49",
          7715 => x"58",
          7716 => x"1e",
          7717 => x"1e",
          7718 => x"fc",
          7719 => x"70",
          7720 => x"33",
          7721 => x"71",
          7722 => x"74",
          7723 => x"81",
          7724 => x"88",
          7725 => x"ff",
          7726 => x"88",
          7727 => x"49",
          7728 => x"5e",
          7729 => x"34",
          7730 => x"34",
          7731 => x"ff",
          7732 => x"83",
          7733 => x"52",
          7734 => x"3f",
          7735 => x"08",
          7736 => x"8c",
          7737 => x"93",
          7738 => x"73",
          7739 => x"8c",
          7740 => x"b4",
          7741 => x"51",
          7742 => x"61",
          7743 => x"27",
          7744 => x"f0",
          7745 => x"3d",
          7746 => x"29",
          7747 => x"08",
          7748 => x"80",
          7749 => x"77",
          7750 => x"38",
          7751 => x"8c",
          7752 => x"0d",
          7753 => x"e4",
          7754 => x"ba",
          7755 => x"84",
          7756 => x"80",
          7757 => x"77",
          7758 => x"84",
          7759 => x"51",
          7760 => x"3f",
          7761 => x"8c",
          7762 => x"0d",
          7763 => x"f4",
          7764 => x"fc",
          7765 => x"0b",
          7766 => x"23",
          7767 => x"53",
          7768 => x"ff",
          7769 => x"b6",
          7770 => x"b9",
          7771 => x"76",
          7772 => x"0b",
          7773 => x"84",
          7774 => x"54",
          7775 => x"34",
          7776 => x"15",
          7777 => x"fc",
          7778 => x"86",
          7779 => x"0b",
          7780 => x"84",
          7781 => x"84",
          7782 => x"ff",
          7783 => x"80",
          7784 => x"ff",
          7785 => x"88",
          7786 => x"55",
          7787 => x"17",
          7788 => x"17",
          7789 => x"f8",
          7790 => x"10",
          7791 => x"fc",
          7792 => x"05",
          7793 => x"82",
          7794 => x"0b",
          7795 => x"77",
          7796 => x"2e",
          7797 => x"fe",
          7798 => x"3d",
          7799 => x"05",
          7800 => x"52",
          7801 => x"87",
          7802 => x"88",
          7803 => x"71",
          7804 => x"0c",
          7805 => x"04",
          7806 => x"02",
          7807 => x"52",
          7808 => x"81",
          7809 => x"71",
          7810 => x"3f",
          7811 => x"08",
          7812 => x"53",
          7813 => x"72",
          7814 => x"13",
          7815 => x"88",
          7816 => x"72",
          7817 => x"0c",
          7818 => x"04",
          7819 => x"7c",
          7820 => x"8c",
          7821 => x"33",
          7822 => x"59",
          7823 => x"74",
          7824 => x"84",
          7825 => x"33",
          7826 => x"06",
          7827 => x"73",
          7828 => x"58",
          7829 => x"c0",
          7830 => x"78",
          7831 => x"76",
          7832 => x"3f",
          7833 => x"08",
          7834 => x"55",
          7835 => x"a7",
          7836 => x"98",
          7837 => x"73",
          7838 => x"78",
          7839 => x"74",
          7840 => x"06",
          7841 => x"2e",
          7842 => x"54",
          7843 => x"84",
          7844 => x"8b",
          7845 => x"84",
          7846 => x"19",
          7847 => x"06",
          7848 => x"79",
          7849 => x"ac",
          7850 => x"f7",
          7851 => x"7e",
          7852 => x"05",
          7853 => x"5a",
          7854 => x"81",
          7855 => x"26",
          7856 => x"ba",
          7857 => x"54",
          7858 => x"54",
          7859 => x"bd",
          7860 => x"85",
          7861 => x"98",
          7862 => x"53",
          7863 => x"51",
          7864 => x"84",
          7865 => x"81",
          7866 => x"74",
          7867 => x"38",
          7868 => x"8c",
          7869 => x"e2",
          7870 => x"26",
          7871 => x"fc",
          7872 => x"54",
          7873 => x"83",
          7874 => x"73",
          7875 => x"ba",
          7876 => x"3d",
          7877 => x"80",
          7878 => x"70",
          7879 => x"5a",
          7880 => x"78",
          7881 => x"38",
          7882 => x"3d",
          7883 => x"84",
          7884 => x"33",
          7885 => x"9f",
          7886 => x"53",
          7887 => x"71",
          7888 => x"38",
          7889 => x"12",
          7890 => x"81",
          7891 => x"53",
          7892 => x"85",
          7893 => x"98",
          7894 => x"53",
          7895 => x"96",
          7896 => x"25",
          7897 => x"83",
          7898 => x"84",
          7899 => x"ba",
          7900 => x"3d",
          7901 => x"80",
          7902 => x"73",
          7903 => x"0c",
          7904 => x"04",
          7905 => x"0c",
          7906 => x"ba",
          7907 => x"3d",
          7908 => x"84",
          7909 => x"92",
          7910 => x"54",
          7911 => x"71",
          7912 => x"2a",
          7913 => x"51",
          7914 => x"8a",
          7915 => x"98",
          7916 => x"74",
          7917 => x"c0",
          7918 => x"51",
          7919 => x"81",
          7920 => x"c0",
          7921 => x"52",
          7922 => x"06",
          7923 => x"2e",
          7924 => x"71",
          7925 => x"54",
          7926 => x"ff",
          7927 => x"3d",
          7928 => x"80",
          7929 => x"33",
          7930 => x"57",
          7931 => x"09",
          7932 => x"38",
          7933 => x"75",
          7934 => x"87",
          7935 => x"80",
          7936 => x"33",
          7937 => x"3f",
          7938 => x"08",
          7939 => x"38",
          7940 => x"84",
          7941 => x"8c",
          7942 => x"81",
          7943 => x"08",
          7944 => x"70",
          7945 => x"33",
          7946 => x"ff",
          7947 => x"84",
          7948 => x"77",
          7949 => x"06",
          7950 => x"ba",
          7951 => x"19",
          7952 => x"08",
          7953 => x"08",
          7954 => x"08",
          7955 => x"08",
          7956 => x"5b",
          7957 => x"ff",
          7958 => x"18",
          7959 => x"82",
          7960 => x"06",
          7961 => x"81",
          7962 => x"53",
          7963 => x"18",
          7964 => x"b7",
          7965 => x"33",
          7966 => x"83",
          7967 => x"06",
          7968 => x"84",
          7969 => x"76",
          7970 => x"81",
          7971 => x"38",
          7972 => x"84",
          7973 => x"57",
          7974 => x"81",
          7975 => x"ff",
          7976 => x"f4",
          7977 => x"0b",
          7978 => x"34",
          7979 => x"84",
          7980 => x"80",
          7981 => x"80",
          7982 => x"19",
          7983 => x"0b",
          7984 => x"80",
          7985 => x"19",
          7986 => x"0b",
          7987 => x"34",
          7988 => x"84",
          7989 => x"80",
          7990 => x"9e",
          7991 => x"e1",
          7992 => x"19",
          7993 => x"08",
          7994 => x"a0",
          7995 => x"88",
          7996 => x"84",
          7997 => x"74",
          7998 => x"75",
          7999 => x"34",
          8000 => x"5b",
          8001 => x"19",
          8002 => x"08",
          8003 => x"a4",
          8004 => x"88",
          8005 => x"84",
          8006 => x"7a",
          8007 => x"75",
          8008 => x"34",
          8009 => x"55",
          8010 => x"19",
          8011 => x"08",
          8012 => x"b4",
          8013 => x"81",
          8014 => x"79",
          8015 => x"33",
          8016 => x"3f",
          8017 => x"34",
          8018 => x"52",
          8019 => x"51",
          8020 => x"84",
          8021 => x"80",
          8022 => x"38",
          8023 => x"f3",
          8024 => x"60",
          8025 => x"56",
          8026 => x"27",
          8027 => x"17",
          8028 => x"8c",
          8029 => x"77",
          8030 => x"0c",
          8031 => x"04",
          8032 => x"56",
          8033 => x"2e",
          8034 => x"74",
          8035 => x"a5",
          8036 => x"2e",
          8037 => x"dd",
          8038 => x"2a",
          8039 => x"2a",
          8040 => x"05",
          8041 => x"5b",
          8042 => x"79",
          8043 => x"83",
          8044 => x"7b",
          8045 => x"81",
          8046 => x"38",
          8047 => x"53",
          8048 => x"81",
          8049 => x"f8",
          8050 => x"ba",
          8051 => x"2e",
          8052 => x"59",
          8053 => x"b4",
          8054 => x"ff",
          8055 => x"83",
          8056 => x"b8",
          8057 => x"1c",
          8058 => x"a8",
          8059 => x"53",
          8060 => x"b4",
          8061 => x"2e",
          8062 => x"0b",
          8063 => x"71",
          8064 => x"74",
          8065 => x"81",
          8066 => x"38",
          8067 => x"53",
          8068 => x"81",
          8069 => x"f8",
          8070 => x"ba",
          8071 => x"2e",
          8072 => x"59",
          8073 => x"b4",
          8074 => x"fe",
          8075 => x"83",
          8076 => x"b8",
          8077 => x"88",
          8078 => x"78",
          8079 => x"84",
          8080 => x"59",
          8081 => x"fe",
          8082 => x"9f",
          8083 => x"ba",
          8084 => x"3d",
          8085 => x"88",
          8086 => x"08",
          8087 => x"17",
          8088 => x"b5",
          8089 => x"83",
          8090 => x"5c",
          8091 => x"7b",
          8092 => x"06",
          8093 => x"81",
          8094 => x"b8",
          8095 => x"17",
          8096 => x"a8",
          8097 => x"8c",
          8098 => x"85",
          8099 => x"81",
          8100 => x"18",
          8101 => x"df",
          8102 => x"83",
          8103 => x"05",
          8104 => x"11",
          8105 => x"71",
          8106 => x"84",
          8107 => x"57",
          8108 => x"0d",
          8109 => x"2e",
          8110 => x"fd",
          8111 => x"87",
          8112 => x"08",
          8113 => x"17",
          8114 => x"b5",
          8115 => x"83",
          8116 => x"5c",
          8117 => x"7b",
          8118 => x"06",
          8119 => x"81",
          8120 => x"b8",
          8121 => x"17",
          8122 => x"c0",
          8123 => x"8c",
          8124 => x"85",
          8125 => x"81",
          8126 => x"18",
          8127 => x"f7",
          8128 => x"2b",
          8129 => x"77",
          8130 => x"83",
          8131 => x"12",
          8132 => x"2b",
          8133 => x"07",
          8134 => x"70",
          8135 => x"2b",
          8136 => x"80",
          8137 => x"80",
          8138 => x"ba",
          8139 => x"5c",
          8140 => x"56",
          8141 => x"04",
          8142 => x"17",
          8143 => x"17",
          8144 => x"18",
          8145 => x"f6",
          8146 => x"5a",
          8147 => x"08",
          8148 => x"81",
          8149 => x"38",
          8150 => x"08",
          8151 => x"b4",
          8152 => x"18",
          8153 => x"ba",
          8154 => x"5e",
          8155 => x"08",
          8156 => x"38",
          8157 => x"55",
          8158 => x"09",
          8159 => x"f7",
          8160 => x"b4",
          8161 => x"18",
          8162 => x"7b",
          8163 => x"33",
          8164 => x"3f",
          8165 => x"df",
          8166 => x"b4",
          8167 => x"b8",
          8168 => x"81",
          8169 => x"5c",
          8170 => x"84",
          8171 => x"7b",
          8172 => x"06",
          8173 => x"84",
          8174 => x"83",
          8175 => x"17",
          8176 => x"08",
          8177 => x"a0",
          8178 => x"8b",
          8179 => x"33",
          8180 => x"2e",
          8181 => x"84",
          8182 => x"5b",
          8183 => x"81",
          8184 => x"08",
          8185 => x"70",
          8186 => x"33",
          8187 => x"bb",
          8188 => x"84",
          8189 => x"7b",
          8190 => x"06",
          8191 => x"84",
          8192 => x"83",
          8193 => x"17",
          8194 => x"08",
          8195 => x"8c",
          8196 => x"7d",
          8197 => x"27",
          8198 => x"82",
          8199 => x"74",
          8200 => x"81",
          8201 => x"38",
          8202 => x"17",
          8203 => x"08",
          8204 => x"52",
          8205 => x"51",
          8206 => x"7a",
          8207 => x"39",
          8208 => x"17",
          8209 => x"17",
          8210 => x"18",
          8211 => x"f4",
          8212 => x"5a",
          8213 => x"08",
          8214 => x"81",
          8215 => x"38",
          8216 => x"08",
          8217 => x"b4",
          8218 => x"18",
          8219 => x"ba",
          8220 => x"55",
          8221 => x"08",
          8222 => x"38",
          8223 => x"55",
          8224 => x"09",
          8225 => x"84",
          8226 => x"b4",
          8227 => x"18",
          8228 => x"7d",
          8229 => x"33",
          8230 => x"3f",
          8231 => x"ec",
          8232 => x"b4",
          8233 => x"18",
          8234 => x"7b",
          8235 => x"33",
          8236 => x"3f",
          8237 => x"81",
          8238 => x"bb",
          8239 => x"39",
          8240 => x"60",
          8241 => x"57",
          8242 => x"81",
          8243 => x"38",
          8244 => x"08",
          8245 => x"78",
          8246 => x"78",
          8247 => x"74",
          8248 => x"80",
          8249 => x"2e",
          8250 => x"77",
          8251 => x"0c",
          8252 => x"04",
          8253 => x"a8",
          8254 => x"58",
          8255 => x"1a",
          8256 => x"76",
          8257 => x"b6",
          8258 => x"33",
          8259 => x"7c",
          8260 => x"81",
          8261 => x"38",
          8262 => x"53",
          8263 => x"81",
          8264 => x"f2",
          8265 => x"ba",
          8266 => x"2e",
          8267 => x"58",
          8268 => x"b4",
          8269 => x"58",
          8270 => x"38",
          8271 => x"fe",
          8272 => x"7b",
          8273 => x"06",
          8274 => x"b8",
          8275 => x"88",
          8276 => x"b9",
          8277 => x"0b",
          8278 => x"77",
          8279 => x"0c",
          8280 => x"04",
          8281 => x"09",
          8282 => x"ff",
          8283 => x"2a",
          8284 => x"05",
          8285 => x"b4",
          8286 => x"5c",
          8287 => x"85",
          8288 => x"19",
          8289 => x"5d",
          8290 => x"09",
          8291 => x"bd",
          8292 => x"77",
          8293 => x"52",
          8294 => x"51",
          8295 => x"84",
          8296 => x"80",
          8297 => x"ff",
          8298 => x"77",
          8299 => x"79",
          8300 => x"b7",
          8301 => x"2b",
          8302 => x"79",
          8303 => x"83",
          8304 => x"98",
          8305 => x"06",
          8306 => x"06",
          8307 => x"5e",
          8308 => x"34",
          8309 => x"56",
          8310 => x"34",
          8311 => x"5a",
          8312 => x"34",
          8313 => x"5b",
          8314 => x"34",
          8315 => x"1a",
          8316 => x"39",
          8317 => x"16",
          8318 => x"a8",
          8319 => x"b4",
          8320 => x"59",
          8321 => x"2e",
          8322 => x"0b",
          8323 => x"71",
          8324 => x"74",
          8325 => x"81",
          8326 => x"38",
          8327 => x"53",
          8328 => x"81",
          8329 => x"f0",
          8330 => x"ba",
          8331 => x"2e",
          8332 => x"58",
          8333 => x"b4",
          8334 => x"58",
          8335 => x"38",
          8336 => x"06",
          8337 => x"81",
          8338 => x"06",
          8339 => x"7a",
          8340 => x"2e",
          8341 => x"84",
          8342 => x"06",
          8343 => x"06",
          8344 => x"5a",
          8345 => x"81",
          8346 => x"34",
          8347 => x"a8",
          8348 => x"56",
          8349 => x"1a",
          8350 => x"74",
          8351 => x"dd",
          8352 => x"74",
          8353 => x"70",
          8354 => x"33",
          8355 => x"9b",
          8356 => x"84",
          8357 => x"7f",
          8358 => x"06",
          8359 => x"84",
          8360 => x"83",
          8361 => x"19",
          8362 => x"1b",
          8363 => x"1b",
          8364 => x"8c",
          8365 => x"56",
          8366 => x"27",
          8367 => x"19",
          8368 => x"82",
          8369 => x"38",
          8370 => x"53",
          8371 => x"19",
          8372 => x"d8",
          8373 => x"8c",
          8374 => x"85",
          8375 => x"81",
          8376 => x"1a",
          8377 => x"83",
          8378 => x"ff",
          8379 => x"05",
          8380 => x"56",
          8381 => x"38",
          8382 => x"76",
          8383 => x"06",
          8384 => x"07",
          8385 => x"76",
          8386 => x"83",
          8387 => x"cb",
          8388 => x"76",
          8389 => x"70",
          8390 => x"33",
          8391 => x"8b",
          8392 => x"84",
          8393 => x"7c",
          8394 => x"06",
          8395 => x"84",
          8396 => x"83",
          8397 => x"19",
          8398 => x"1b",
          8399 => x"1b",
          8400 => x"8c",
          8401 => x"40",
          8402 => x"27",
          8403 => x"82",
          8404 => x"74",
          8405 => x"81",
          8406 => x"38",
          8407 => x"1e",
          8408 => x"81",
          8409 => x"ee",
          8410 => x"5a",
          8411 => x"81",
          8412 => x"b8",
          8413 => x"81",
          8414 => x"57",
          8415 => x"81",
          8416 => x"8c",
          8417 => x"09",
          8418 => x"ae",
          8419 => x"8c",
          8420 => x"34",
          8421 => x"70",
          8422 => x"31",
          8423 => x"84",
          8424 => x"5f",
          8425 => x"74",
          8426 => x"f0",
          8427 => x"33",
          8428 => x"2e",
          8429 => x"fc",
          8430 => x"54",
          8431 => x"76",
          8432 => x"33",
          8433 => x"3f",
          8434 => x"d0",
          8435 => x"76",
          8436 => x"70",
          8437 => x"33",
          8438 => x"cf",
          8439 => x"84",
          8440 => x"7c",
          8441 => x"06",
          8442 => x"84",
          8443 => x"83",
          8444 => x"19",
          8445 => x"1b",
          8446 => x"1b",
          8447 => x"8c",
          8448 => x"40",
          8449 => x"27",
          8450 => x"82",
          8451 => x"74",
          8452 => x"81",
          8453 => x"38",
          8454 => x"1e",
          8455 => x"81",
          8456 => x"ed",
          8457 => x"5a",
          8458 => x"81",
          8459 => x"53",
          8460 => x"19",
          8461 => x"f3",
          8462 => x"fd",
          8463 => x"76",
          8464 => x"06",
          8465 => x"83",
          8466 => x"59",
          8467 => x"b8",
          8468 => x"88",
          8469 => x"b9",
          8470 => x"fa",
          8471 => x"fd",
          8472 => x"76",
          8473 => x"fc",
          8474 => x"b8",
          8475 => x"33",
          8476 => x"8f",
          8477 => x"f0",
          8478 => x"42",
          8479 => x"58",
          8480 => x"7d",
          8481 => x"75",
          8482 => x"7d",
          8483 => x"79",
          8484 => x"7d",
          8485 => x"7a",
          8486 => x"fa",
          8487 => x"3d",
          8488 => x"71",
          8489 => x"5a",
          8490 => x"38",
          8491 => x"57",
          8492 => x"80",
          8493 => x"9c",
          8494 => x"80",
          8495 => x"19",
          8496 => x"54",
          8497 => x"80",
          8498 => x"7b",
          8499 => x"38",
          8500 => x"16",
          8501 => x"08",
          8502 => x"38",
          8503 => x"77",
          8504 => x"38",
          8505 => x"51",
          8506 => x"84",
          8507 => x"80",
          8508 => x"38",
          8509 => x"ba",
          8510 => x"2e",
          8511 => x"ba",
          8512 => x"70",
          8513 => x"07",
          8514 => x"7b",
          8515 => x"55",
          8516 => x"aa",
          8517 => x"2e",
          8518 => x"ff",
          8519 => x"55",
          8520 => x"8c",
          8521 => x"0d",
          8522 => x"ff",
          8523 => x"ba",
          8524 => x"ca",
          8525 => x"79",
          8526 => x"3f",
          8527 => x"84",
          8528 => x"27",
          8529 => x"ba",
          8530 => x"84",
          8531 => x"ff",
          8532 => x"9c",
          8533 => x"ba",
          8534 => x"c4",
          8535 => x"fe",
          8536 => x"1b",
          8537 => x"08",
          8538 => x"38",
          8539 => x"52",
          8540 => x"eb",
          8541 => x"84",
          8542 => x"81",
          8543 => x"38",
          8544 => x"08",
          8545 => x"70",
          8546 => x"25",
          8547 => x"84",
          8548 => x"54",
          8549 => x"55",
          8550 => x"38",
          8551 => x"08",
          8552 => x"38",
          8553 => x"54",
          8554 => x"fe",
          8555 => x"9c",
          8556 => x"fe",
          8557 => x"70",
          8558 => x"96",
          8559 => x"2e",
          8560 => x"ff",
          8561 => x"78",
          8562 => x"3f",
          8563 => x"08",
          8564 => x"08",
          8565 => x"ba",
          8566 => x"80",
          8567 => x"55",
          8568 => x"38",
          8569 => x"38",
          8570 => x"0c",
          8571 => x"fe",
          8572 => x"08",
          8573 => x"78",
          8574 => x"ff",
          8575 => x"0c",
          8576 => x"81",
          8577 => x"84",
          8578 => x"55",
          8579 => x"8c",
          8580 => x"0d",
          8581 => x"84",
          8582 => x"8c",
          8583 => x"84",
          8584 => x"58",
          8585 => x"73",
          8586 => x"b8",
          8587 => x"7a",
          8588 => x"f5",
          8589 => x"ba",
          8590 => x"ff",
          8591 => x"ba",
          8592 => x"ba",
          8593 => x"3d",
          8594 => x"56",
          8595 => x"ff",
          8596 => x"55",
          8597 => x"f8",
          8598 => x"7c",
          8599 => x"55",
          8600 => x"80",
          8601 => x"df",
          8602 => x"06",
          8603 => x"d7",
          8604 => x"19",
          8605 => x"08",
          8606 => x"df",
          8607 => x"56",
          8608 => x"80",
          8609 => x"85",
          8610 => x"0b",
          8611 => x"5a",
          8612 => x"27",
          8613 => x"17",
          8614 => x"0c",
          8615 => x"0c",
          8616 => x"53",
          8617 => x"80",
          8618 => x"73",
          8619 => x"98",
          8620 => x"83",
          8621 => x"b8",
          8622 => x"0c",
          8623 => x"84",
          8624 => x"8a",
          8625 => x"82",
          8626 => x"8c",
          8627 => x"0d",
          8628 => x"08",
          8629 => x"2e",
          8630 => x"8a",
          8631 => x"89",
          8632 => x"73",
          8633 => x"38",
          8634 => x"53",
          8635 => x"14",
          8636 => x"59",
          8637 => x"8d",
          8638 => x"22",
          8639 => x"b0",
          8640 => x"5a",
          8641 => x"19",
          8642 => x"39",
          8643 => x"51",
          8644 => x"84",
          8645 => x"55",
          8646 => x"08",
          8647 => x"38",
          8648 => x"ba",
          8649 => x"ff",
          8650 => x"17",
          8651 => x"ba",
          8652 => x"27",
          8653 => x"73",
          8654 => x"73",
          8655 => x"38",
          8656 => x"81",
          8657 => x"8c",
          8658 => x"0d",
          8659 => x"0d",
          8660 => x"90",
          8661 => x"05",
          8662 => x"f0",
          8663 => x"27",
          8664 => x"0b",
          8665 => x"98",
          8666 => x"84",
          8667 => x"2e",
          8668 => x"83",
          8669 => x"7a",
          8670 => x"15",
          8671 => x"57",
          8672 => x"38",
          8673 => x"88",
          8674 => x"55",
          8675 => x"81",
          8676 => x"98",
          8677 => x"90",
          8678 => x"1b",
          8679 => x"18",
          8680 => x"75",
          8681 => x"0c",
          8682 => x"04",
          8683 => x"0c",
          8684 => x"ff",
          8685 => x"2a",
          8686 => x"da",
          8687 => x"76",
          8688 => x"3f",
          8689 => x"08",
          8690 => x"81",
          8691 => x"8c",
          8692 => x"38",
          8693 => x"ba",
          8694 => x"2e",
          8695 => x"19",
          8696 => x"8c",
          8697 => x"91",
          8698 => x"2e",
          8699 => x"94",
          8700 => x"76",
          8701 => x"3f",
          8702 => x"08",
          8703 => x"84",
          8704 => x"80",
          8705 => x"38",
          8706 => x"ba",
          8707 => x"2e",
          8708 => x"81",
          8709 => x"8c",
          8710 => x"ff",
          8711 => x"ba",
          8712 => x"1a",
          8713 => x"7d",
          8714 => x"fe",
          8715 => x"08",
          8716 => x"56",
          8717 => x"78",
          8718 => x"8a",
          8719 => x"71",
          8720 => x"08",
          8721 => x"7b",
          8722 => x"b8",
          8723 => x"80",
          8724 => x"80",
          8725 => x"05",
          8726 => x"15",
          8727 => x"38",
          8728 => x"19",
          8729 => x"75",
          8730 => x"38",
          8731 => x"1c",
          8732 => x"81",
          8733 => x"e4",
          8734 => x"ba",
          8735 => x"e7",
          8736 => x"56",
          8737 => x"98",
          8738 => x"0b",
          8739 => x"0c",
          8740 => x"04",
          8741 => x"19",
          8742 => x"19",
          8743 => x"1a",
          8744 => x"e4",
          8745 => x"ba",
          8746 => x"f3",
          8747 => x"8c",
          8748 => x"34",
          8749 => x"a8",
          8750 => x"55",
          8751 => x"08",
          8752 => x"38",
          8753 => x"5c",
          8754 => x"09",
          8755 => x"db",
          8756 => x"b4",
          8757 => x"1a",
          8758 => x"75",
          8759 => x"33",
          8760 => x"3f",
          8761 => x"8a",
          8762 => x"74",
          8763 => x"06",
          8764 => x"2e",
          8765 => x"a7",
          8766 => x"18",
          8767 => x"9c",
          8768 => x"05",
          8769 => x"58",
          8770 => x"fd",
          8771 => x"19",
          8772 => x"29",
          8773 => x"05",
          8774 => x"5c",
          8775 => x"81",
          8776 => x"8c",
          8777 => x"0d",
          8778 => x"0d",
          8779 => x"5c",
          8780 => x"5a",
          8781 => x"70",
          8782 => x"58",
          8783 => x"80",
          8784 => x"38",
          8785 => x"75",
          8786 => x"b4",
          8787 => x"2e",
          8788 => x"83",
          8789 => x"58",
          8790 => x"2e",
          8791 => x"81",
          8792 => x"54",
          8793 => x"19",
          8794 => x"33",
          8795 => x"3f",
          8796 => x"08",
          8797 => x"38",
          8798 => x"57",
          8799 => x"0c",
          8800 => x"82",
          8801 => x"1c",
          8802 => x"58",
          8803 => x"2e",
          8804 => x"8b",
          8805 => x"06",
          8806 => x"06",
          8807 => x"86",
          8808 => x"81",
          8809 => x"30",
          8810 => x"70",
          8811 => x"25",
          8812 => x"07",
          8813 => x"57",
          8814 => x"38",
          8815 => x"06",
          8816 => x"88",
          8817 => x"38",
          8818 => x"81",
          8819 => x"ff",
          8820 => x"7b",
          8821 => x"3f",
          8822 => x"08",
          8823 => x"8c",
          8824 => x"38",
          8825 => x"56",
          8826 => x"38",
          8827 => x"8c",
          8828 => x"0d",
          8829 => x"b4",
          8830 => x"7e",
          8831 => x"33",
          8832 => x"3f",
          8833 => x"ba",
          8834 => x"2e",
          8835 => x"fe",
          8836 => x"ba",
          8837 => x"1a",
          8838 => x"08",
          8839 => x"31",
          8840 => x"08",
          8841 => x"a0",
          8842 => x"fe",
          8843 => x"19",
          8844 => x"82",
          8845 => x"06",
          8846 => x"81",
          8847 => x"08",
          8848 => x"05",
          8849 => x"81",
          8850 => x"e0",
          8851 => x"57",
          8852 => x"79",
          8853 => x"81",
          8854 => x"38",
          8855 => x"81",
          8856 => x"80",
          8857 => x"8d",
          8858 => x"81",
          8859 => x"90",
          8860 => x"ac",
          8861 => x"5e",
          8862 => x"2e",
          8863 => x"ff",
          8864 => x"fe",
          8865 => x"56",
          8866 => x"09",
          8867 => x"be",
          8868 => x"84",
          8869 => x"98",
          8870 => x"84",
          8871 => x"94",
          8872 => x"77",
          8873 => x"39",
          8874 => x"57",
          8875 => x"09",
          8876 => x"38",
          8877 => x"9b",
          8878 => x"1a",
          8879 => x"2b",
          8880 => x"41",
          8881 => x"38",
          8882 => x"81",
          8883 => x"29",
          8884 => x"5a",
          8885 => x"5b",
          8886 => x"17",
          8887 => x"81",
          8888 => x"33",
          8889 => x"07",
          8890 => x"7a",
          8891 => x"c5",
          8892 => x"fe",
          8893 => x"38",
          8894 => x"05",
          8895 => x"75",
          8896 => x"1a",
          8897 => x"57",
          8898 => x"cc",
          8899 => x"70",
          8900 => x"06",
          8901 => x"80",
          8902 => x"79",
          8903 => x"fe",
          8904 => x"10",
          8905 => x"80",
          8906 => x"1d",
          8907 => x"06",
          8908 => x"9d",
          8909 => x"ff",
          8910 => x"38",
          8911 => x"fe",
          8912 => x"a8",
          8913 => x"8b",
          8914 => x"2a",
          8915 => x"29",
          8916 => x"81",
          8917 => x"40",
          8918 => x"81",
          8919 => x"19",
          8920 => x"76",
          8921 => x"7e",
          8922 => x"38",
          8923 => x"1d",
          8924 => x"ba",
          8925 => x"3d",
          8926 => x"3d",
          8927 => x"08",
          8928 => x"52",
          8929 => x"cf",
          8930 => x"8c",
          8931 => x"ba",
          8932 => x"80",
          8933 => x"70",
          8934 => x"0b",
          8935 => x"b8",
          8936 => x"1c",
          8937 => x"58",
          8938 => x"76",
          8939 => x"38",
          8940 => x"78",
          8941 => x"78",
          8942 => x"06",
          8943 => x"81",
          8944 => x"b8",
          8945 => x"1b",
          8946 => x"e0",
          8947 => x"8c",
          8948 => x"85",
          8949 => x"81",
          8950 => x"1c",
          8951 => x"76",
          8952 => x"9c",
          8953 => x"33",
          8954 => x"80",
          8955 => x"38",
          8956 => x"bf",
          8957 => x"ff",
          8958 => x"77",
          8959 => x"76",
          8960 => x"80",
          8961 => x"83",
          8962 => x"55",
          8963 => x"81",
          8964 => x"80",
          8965 => x"8f",
          8966 => x"38",
          8967 => x"78",
          8968 => x"8b",
          8969 => x"2a",
          8970 => x"29",
          8971 => x"81",
          8972 => x"57",
          8973 => x"81",
          8974 => x"19",
          8975 => x"76",
          8976 => x"7f",
          8977 => x"38",
          8978 => x"81",
          8979 => x"a7",
          8980 => x"a0",
          8981 => x"78",
          8982 => x"5a",
          8983 => x"81",
          8984 => x"71",
          8985 => x"1a",
          8986 => x"40",
          8987 => x"81",
          8988 => x"80",
          8989 => x"81",
          8990 => x"0b",
          8991 => x"80",
          8992 => x"f5",
          8993 => x"ba",
          8994 => x"84",
          8995 => x"80",
          8996 => x"38",
          8997 => x"8c",
          8998 => x"0d",
          8999 => x"b4",
          9000 => x"7d",
          9001 => x"33",
          9002 => x"3f",
          9003 => x"ba",
          9004 => x"2e",
          9005 => x"fe",
          9006 => x"ba",
          9007 => x"1c",
          9008 => x"08",
          9009 => x"31",
          9010 => x"08",
          9011 => x"a0",
          9012 => x"fd",
          9013 => x"1b",
          9014 => x"82",
          9015 => x"06",
          9016 => x"81",
          9017 => x"08",
          9018 => x"05",
          9019 => x"81",
          9020 => x"db",
          9021 => x"57",
          9022 => x"77",
          9023 => x"39",
          9024 => x"70",
          9025 => x"06",
          9026 => x"fe",
          9027 => x"86",
          9028 => x"5a",
          9029 => x"93",
          9030 => x"33",
          9031 => x"06",
          9032 => x"08",
          9033 => x"0c",
          9034 => x"76",
          9035 => x"38",
          9036 => x"74",
          9037 => x"7b",
          9038 => x"3f",
          9039 => x"08",
          9040 => x"8c",
          9041 => x"fc",
          9042 => x"c8",
          9043 => x"2e",
          9044 => x"81",
          9045 => x"0b",
          9046 => x"fe",
          9047 => x"19",
          9048 => x"77",
          9049 => x"06",
          9050 => x"1b",
          9051 => x"33",
          9052 => x"71",
          9053 => x"59",
          9054 => x"ff",
          9055 => x"33",
          9056 => x"8d",
          9057 => x"5b",
          9058 => x"59",
          9059 => x"8c",
          9060 => x"05",
          9061 => x"71",
          9062 => x"2b",
          9063 => x"57",
          9064 => x"80",
          9065 => x"81",
          9066 => x"84",
          9067 => x"81",
          9068 => x"84",
          9069 => x"7a",
          9070 => x"70",
          9071 => x"81",
          9072 => x"81",
          9073 => x"75",
          9074 => x"08",
          9075 => x"06",
          9076 => x"76",
          9077 => x"58",
          9078 => x"ff",
          9079 => x"33",
          9080 => x"81",
          9081 => x"75",
          9082 => x"38",
          9083 => x"8d",
          9084 => x"60",
          9085 => x"41",
          9086 => x"b4",
          9087 => x"70",
          9088 => x"5e",
          9089 => x"39",
          9090 => x"ba",
          9091 => x"3d",
          9092 => x"83",
          9093 => x"ff",
          9094 => x"ff",
          9095 => x"39",
          9096 => x"68",
          9097 => x"ab",
          9098 => x"a0",
          9099 => x"5d",
          9100 => x"74",
          9101 => x"74",
          9102 => x"70",
          9103 => x"5d",
          9104 => x"8e",
          9105 => x"70",
          9106 => x"22",
          9107 => x"74",
          9108 => x"3d",
          9109 => x"40",
          9110 => x"58",
          9111 => x"70",
          9112 => x"33",
          9113 => x"05",
          9114 => x"15",
          9115 => x"38",
          9116 => x"05",
          9117 => x"06",
          9118 => x"80",
          9119 => x"38",
          9120 => x"ab",
          9121 => x"0b",
          9122 => x"5b",
          9123 => x"7b",
          9124 => x"7a",
          9125 => x"55",
          9126 => x"05",
          9127 => x"70",
          9128 => x"34",
          9129 => x"74",
          9130 => x"7b",
          9131 => x"38",
          9132 => x"56",
          9133 => x"2e",
          9134 => x"82",
          9135 => x"8f",
          9136 => x"06",
          9137 => x"76",
          9138 => x"83",
          9139 => x"72",
          9140 => x"06",
          9141 => x"57",
          9142 => x"87",
          9143 => x"a0",
          9144 => x"ff",
          9145 => x"80",
          9146 => x"78",
          9147 => x"ca",
          9148 => x"84",
          9149 => x"05",
          9150 => x"b0",
          9151 => x"55",
          9152 => x"84",
          9153 => x"55",
          9154 => x"ff",
          9155 => x"78",
          9156 => x"59",
          9157 => x"38",
          9158 => x"80",
          9159 => x"76",
          9160 => x"80",
          9161 => x"38",
          9162 => x"74",
          9163 => x"38",
          9164 => x"75",
          9165 => x"a2",
          9166 => x"70",
          9167 => x"74",
          9168 => x"81",
          9169 => x"81",
          9170 => x"55",
          9171 => x"8e",
          9172 => x"78",
          9173 => x"81",
          9174 => x"57",
          9175 => x"77",
          9176 => x"27",
          9177 => x"7d",
          9178 => x"3f",
          9179 => x"08",
          9180 => x"1b",
          9181 => x"7b",
          9182 => x"38",
          9183 => x"80",
          9184 => x"e7",
          9185 => x"8c",
          9186 => x"ba",
          9187 => x"2e",
          9188 => x"82",
          9189 => x"80",
          9190 => x"ab",
          9191 => x"08",
          9192 => x"80",
          9193 => x"57",
          9194 => x"2a",
          9195 => x"81",
          9196 => x"2e",
          9197 => x"52",
          9198 => x"fe",
          9199 => x"84",
          9200 => x"1b",
          9201 => x"7d",
          9202 => x"3f",
          9203 => x"08",
          9204 => x"8c",
          9205 => x"38",
          9206 => x"08",
          9207 => x"59",
          9208 => x"56",
          9209 => x"18",
          9210 => x"85",
          9211 => x"18",
          9212 => x"77",
          9213 => x"06",
          9214 => x"81",
          9215 => x"b8",
          9216 => x"18",
          9217 => x"a4",
          9218 => x"8c",
          9219 => x"85",
          9220 => x"81",
          9221 => x"19",
          9222 => x"76",
          9223 => x"1e",
          9224 => x"56",
          9225 => x"e5",
          9226 => x"38",
          9227 => x"80",
          9228 => x"56",
          9229 => x"2e",
          9230 => x"81",
          9231 => x"7b",
          9232 => x"38",
          9233 => x"51",
          9234 => x"84",
          9235 => x"56",
          9236 => x"08",
          9237 => x"88",
          9238 => x"75",
          9239 => x"89",
          9240 => x"75",
          9241 => x"ff",
          9242 => x"81",
          9243 => x"1e",
          9244 => x"1c",
          9245 => x"af",
          9246 => x"33",
          9247 => x"7f",
          9248 => x"81",
          9249 => x"b8",
          9250 => x"1c",
          9251 => x"9c",
          9252 => x"8c",
          9253 => x"85",
          9254 => x"81",
          9255 => x"1d",
          9256 => x"75",
          9257 => x"a0",
          9258 => x"08",
          9259 => x"76",
          9260 => x"58",
          9261 => x"55",
          9262 => x"8b",
          9263 => x"08",
          9264 => x"55",
          9265 => x"05",
          9266 => x"70",
          9267 => x"34",
          9268 => x"74",
          9269 => x"1e",
          9270 => x"33",
          9271 => x"5a",
          9272 => x"34",
          9273 => x"1d",
          9274 => x"75",
          9275 => x"0c",
          9276 => x"04",
          9277 => x"70",
          9278 => x"07",
          9279 => x"74",
          9280 => x"74",
          9281 => x"7d",
          9282 => x"3f",
          9283 => x"08",
          9284 => x"8c",
          9285 => x"fd",
          9286 => x"bd",
          9287 => x"b4",
          9288 => x"7c",
          9289 => x"33",
          9290 => x"3f",
          9291 => x"08",
          9292 => x"81",
          9293 => x"38",
          9294 => x"08",
          9295 => x"b4",
          9296 => x"19",
          9297 => x"74",
          9298 => x"27",
          9299 => x"18",
          9300 => x"82",
          9301 => x"38",
          9302 => x"08",
          9303 => x"39",
          9304 => x"90",
          9305 => x"31",
          9306 => x"51",
          9307 => x"84",
          9308 => x"58",
          9309 => x"08",
          9310 => x"79",
          9311 => x"08",
          9312 => x"57",
          9313 => x"75",
          9314 => x"05",
          9315 => x"05",
          9316 => x"76",
          9317 => x"ff",
          9318 => x"59",
          9319 => x"e4",
          9320 => x"ff",
          9321 => x"43",
          9322 => x"08",
          9323 => x"b4",
          9324 => x"2e",
          9325 => x"1c",
          9326 => x"76",
          9327 => x"06",
          9328 => x"81",
          9329 => x"b8",
          9330 => x"1c",
          9331 => x"dc",
          9332 => x"8c",
          9333 => x"85",
          9334 => x"81",
          9335 => x"1d",
          9336 => x"75",
          9337 => x"8c",
          9338 => x"1f",
          9339 => x"ff",
          9340 => x"5f",
          9341 => x"34",
          9342 => x"1c",
          9343 => x"1c",
          9344 => x"1c",
          9345 => x"1c",
          9346 => x"29",
          9347 => x"77",
          9348 => x"76",
          9349 => x"2e",
          9350 => x"10",
          9351 => x"81",
          9352 => x"56",
          9353 => x"18",
          9354 => x"55",
          9355 => x"81",
          9356 => x"76",
          9357 => x"75",
          9358 => x"85",
          9359 => x"ff",
          9360 => x"58",
          9361 => x"cb",
          9362 => x"ff",
          9363 => x"b3",
          9364 => x"1f",
          9365 => x"58",
          9366 => x"81",
          9367 => x"7b",
          9368 => x"83",
          9369 => x"52",
          9370 => x"e1",
          9371 => x"8c",
          9372 => x"ba",
          9373 => x"f1",
          9374 => x"05",
          9375 => x"a9",
          9376 => x"39",
          9377 => x"1c",
          9378 => x"1c",
          9379 => x"1d",
          9380 => x"d0",
          9381 => x"56",
          9382 => x"08",
          9383 => x"84",
          9384 => x"83",
          9385 => x"1c",
          9386 => x"08",
          9387 => x"8c",
          9388 => x"60",
          9389 => x"27",
          9390 => x"82",
          9391 => x"61",
          9392 => x"81",
          9393 => x"38",
          9394 => x"1c",
          9395 => x"08",
          9396 => x"52",
          9397 => x"51",
          9398 => x"77",
          9399 => x"39",
          9400 => x"08",
          9401 => x"43",
          9402 => x"e5",
          9403 => x"06",
          9404 => x"fb",
          9405 => x"70",
          9406 => x"80",
          9407 => x"38",
          9408 => x"7c",
          9409 => x"5d",
          9410 => x"81",
          9411 => x"08",
          9412 => x"81",
          9413 => x"cf",
          9414 => x"ba",
          9415 => x"2e",
          9416 => x"bc",
          9417 => x"8c",
          9418 => x"34",
          9419 => x"a8",
          9420 => x"55",
          9421 => x"08",
          9422 => x"82",
          9423 => x"7e",
          9424 => x"38",
          9425 => x"08",
          9426 => x"39",
          9427 => x"41",
          9428 => x"2e",
          9429 => x"fc",
          9430 => x"1a",
          9431 => x"39",
          9432 => x"56",
          9433 => x"fc",
          9434 => x"fd",
          9435 => x"b4",
          9436 => x"1d",
          9437 => x"61",
          9438 => x"33",
          9439 => x"3f",
          9440 => x"81",
          9441 => x"08",
          9442 => x"05",
          9443 => x"81",
          9444 => x"ce",
          9445 => x"e3",
          9446 => x"0d",
          9447 => x"08",
          9448 => x"80",
          9449 => x"34",
          9450 => x"80",
          9451 => x"38",
          9452 => x"ff",
          9453 => x"38",
          9454 => x"60",
          9455 => x"70",
          9456 => x"5b",
          9457 => x"78",
          9458 => x"77",
          9459 => x"70",
          9460 => x"5b",
          9461 => x"82",
          9462 => x"d0",
          9463 => x"83",
          9464 => x"58",
          9465 => x"ff",
          9466 => x"38",
          9467 => x"76",
          9468 => x"5d",
          9469 => x"79",
          9470 => x"30",
          9471 => x"70",
          9472 => x"5a",
          9473 => x"18",
          9474 => x"80",
          9475 => x"34",
          9476 => x"1f",
          9477 => x"9c",
          9478 => x"70",
          9479 => x"58",
          9480 => x"a0",
          9481 => x"74",
          9482 => x"bc",
          9483 => x"32",
          9484 => x"72",
          9485 => x"55",
          9486 => x"8b",
          9487 => x"72",
          9488 => x"38",
          9489 => x"81",
          9490 => x"81",
          9491 => x"77",
          9492 => x"59",
          9493 => x"58",
          9494 => x"ff",
          9495 => x"18",
          9496 => x"80",
          9497 => x"34",
          9498 => x"53",
          9499 => x"77",
          9500 => x"bf",
          9501 => x"34",
          9502 => x"17",
          9503 => x"80",
          9504 => x"34",
          9505 => x"8c",
          9506 => x"53",
          9507 => x"73",
          9508 => x"9c",
          9509 => x"8b",
          9510 => x"1e",
          9511 => x"08",
          9512 => x"11",
          9513 => x"33",
          9514 => x"71",
          9515 => x"81",
          9516 => x"72",
          9517 => x"75",
          9518 => x"64",
          9519 => x"16",
          9520 => x"33",
          9521 => x"07",
          9522 => x"40",
          9523 => x"55",
          9524 => x"23",
          9525 => x"98",
          9526 => x"88",
          9527 => x"54",
          9528 => x"23",
          9529 => x"04",
          9530 => x"fe",
          9531 => x"1d",
          9532 => x"ff",
          9533 => x"5b",
          9534 => x"52",
          9535 => x"74",
          9536 => x"91",
          9537 => x"ba",
          9538 => x"ff",
          9539 => x"81",
          9540 => x"ad",
          9541 => x"27",
          9542 => x"74",
          9543 => x"73",
          9544 => x"97",
          9545 => x"78",
          9546 => x"0b",
          9547 => x"56",
          9548 => x"75",
          9549 => x"5c",
          9550 => x"fd",
          9551 => x"ba",
          9552 => x"76",
          9553 => x"07",
          9554 => x"80",
          9555 => x"55",
          9556 => x"f9",
          9557 => x"34",
          9558 => x"58",
          9559 => x"1f",
          9560 => x"cd",
          9561 => x"89",
          9562 => x"57",
          9563 => x"2e",
          9564 => x"7c",
          9565 => x"57",
          9566 => x"14",
          9567 => x"11",
          9568 => x"99",
          9569 => x"9c",
          9570 => x"11",
          9571 => x"88",
          9572 => x"38",
          9573 => x"53",
          9574 => x"5e",
          9575 => x"8a",
          9576 => x"70",
          9577 => x"06",
          9578 => x"78",
          9579 => x"5a",
          9580 => x"81",
          9581 => x"71",
          9582 => x"5e",
          9583 => x"56",
          9584 => x"38",
          9585 => x"72",
          9586 => x"cc",
          9587 => x"30",
          9588 => x"70",
          9589 => x"53",
          9590 => x"fc",
          9591 => x"3d",
          9592 => x"08",
          9593 => x"5c",
          9594 => x"33",
          9595 => x"74",
          9596 => x"38",
          9597 => x"80",
          9598 => x"df",
          9599 => x"2e",
          9600 => x"98",
          9601 => x"1d",
          9602 => x"96",
          9603 => x"41",
          9604 => x"75",
          9605 => x"38",
          9606 => x"16",
          9607 => x"57",
          9608 => x"81",
          9609 => x"55",
          9610 => x"df",
          9611 => x"0c",
          9612 => x"81",
          9613 => x"ff",
          9614 => x"8b",
          9615 => x"18",
          9616 => x"23",
          9617 => x"73",
          9618 => x"06",
          9619 => x"70",
          9620 => x"27",
          9621 => x"07",
          9622 => x"55",
          9623 => x"38",
          9624 => x"2e",
          9625 => x"74",
          9626 => x"b2",
          9627 => x"a8",
          9628 => x"a8",
          9629 => x"ff",
          9630 => x"56",
          9631 => x"81",
          9632 => x"75",
          9633 => x"81",
          9634 => x"70",
          9635 => x"56",
          9636 => x"ee",
          9637 => x"ff",
          9638 => x"81",
          9639 => x"81",
          9640 => x"fd",
          9641 => x"18",
          9642 => x"23",
          9643 => x"70",
          9644 => x"52",
          9645 => x"57",
          9646 => x"fe",
          9647 => x"cb",
          9648 => x"80",
          9649 => x"30",
          9650 => x"73",
          9651 => x"58",
          9652 => x"2e",
          9653 => x"14",
          9654 => x"80",
          9655 => x"55",
          9656 => x"dd",
          9657 => x"dc",
          9658 => x"70",
          9659 => x"07",
          9660 => x"72",
          9661 => x"88",
          9662 => x"33",
          9663 => x"3d",
          9664 => x"74",
          9665 => x"90",
          9666 => x"83",
          9667 => x"51",
          9668 => x"3f",
          9669 => x"08",
          9670 => x"06",
          9671 => x"8d",
          9672 => x"73",
          9673 => x"0c",
          9674 => x"04",
          9675 => x"33",
          9676 => x"06",
          9677 => x"80",
          9678 => x"38",
          9679 => x"80",
          9680 => x"34",
          9681 => x"51",
          9682 => x"84",
          9683 => x"84",
          9684 => x"93",
          9685 => x"81",
          9686 => x"32",
          9687 => x"80",
          9688 => x"41",
          9689 => x"7d",
          9690 => x"38",
          9691 => x"80",
          9692 => x"55",
          9693 => x"af",
          9694 => x"72",
          9695 => x"70",
          9696 => x"25",
          9697 => x"54",
          9698 => x"38",
          9699 => x"9f",
          9700 => x"2b",
          9701 => x"2e",
          9702 => x"76",
          9703 => x"d1",
          9704 => x"59",
          9705 => x"a7",
          9706 => x"78",
          9707 => x"70",
          9708 => x"32",
          9709 => x"9f",
          9710 => x"56",
          9711 => x"7c",
          9712 => x"38",
          9713 => x"ff",
          9714 => x"dd",
          9715 => x"77",
          9716 => x"76",
          9717 => x"2e",
          9718 => x"80",
          9719 => x"83",
          9720 => x"72",
          9721 => x"56",
          9722 => x"82",
          9723 => x"83",
          9724 => x"53",
          9725 => x"82",
          9726 => x"80",
          9727 => x"77",
          9728 => x"70",
          9729 => x"78",
          9730 => x"38",
          9731 => x"fe",
          9732 => x"17",
          9733 => x"2e",
          9734 => x"14",
          9735 => x"54",
          9736 => x"09",
          9737 => x"38",
          9738 => x"1d",
          9739 => x"74",
          9740 => x"56",
          9741 => x"53",
          9742 => x"72",
          9743 => x"88",
          9744 => x"22",
          9745 => x"57",
          9746 => x"80",
          9747 => x"38",
          9748 => x"83",
          9749 => x"ae",
          9750 => x"70",
          9751 => x"5a",
          9752 => x"2e",
          9753 => x"72",
          9754 => x"72",
          9755 => x"26",
          9756 => x"59",
          9757 => x"70",
          9758 => x"07",
          9759 => x"7c",
          9760 => x"54",
          9761 => x"2e",
          9762 => x"7c",
          9763 => x"83",
          9764 => x"2e",
          9765 => x"83",
          9766 => x"77",
          9767 => x"76",
          9768 => x"8b",
          9769 => x"81",
          9770 => x"18",
          9771 => x"77",
          9772 => x"81",
          9773 => x"53",
          9774 => x"38",
          9775 => x"57",
          9776 => x"2e",
          9777 => x"7c",
          9778 => x"e3",
          9779 => x"06",
          9780 => x"2e",
          9781 => x"7d",
          9782 => x"74",
          9783 => x"e3",
          9784 => x"2a",
          9785 => x"75",
          9786 => x"81",
          9787 => x"80",
          9788 => x"79",
          9789 => x"7d",
          9790 => x"06",
          9791 => x"2e",
          9792 => x"88",
          9793 => x"ab",
          9794 => x"51",
          9795 => x"84",
          9796 => x"ab",
          9797 => x"54",
          9798 => x"08",
          9799 => x"ac",
          9800 => x"8c",
          9801 => x"09",
          9802 => x"f7",
          9803 => x"2a",
          9804 => x"79",
          9805 => x"f0",
          9806 => x"2a",
          9807 => x"78",
          9808 => x"7b",
          9809 => x"56",
          9810 => x"16",
          9811 => x"57",
          9812 => x"81",
          9813 => x"79",
          9814 => x"40",
          9815 => x"7c",
          9816 => x"38",
          9817 => x"fd",
          9818 => x"83",
          9819 => x"8a",
          9820 => x"22",
          9821 => x"2e",
          9822 => x"fc",
          9823 => x"22",
          9824 => x"2e",
          9825 => x"fc",
          9826 => x"10",
          9827 => x"7b",
          9828 => x"a0",
          9829 => x"ae",
          9830 => x"26",
          9831 => x"54",
          9832 => x"81",
          9833 => x"81",
          9834 => x"73",
          9835 => x"79",
          9836 => x"77",
          9837 => x"7b",
          9838 => x"3f",
          9839 => x"08",
          9840 => x"56",
          9841 => x"8c",
          9842 => x"38",
          9843 => x"81",
          9844 => x"fa",
          9845 => x"1c",
          9846 => x"2a",
          9847 => x"5d",
          9848 => x"83",
          9849 => x"1c",
          9850 => x"06",
          9851 => x"d3",
          9852 => x"d2",
          9853 => x"88",
          9854 => x"33",
          9855 => x"54",
          9856 => x"82",
          9857 => x"88",
          9858 => x"08",
          9859 => x"fe",
          9860 => x"22",
          9861 => x"2e",
          9862 => x"76",
          9863 => x"fb",
          9864 => x"ab",
          9865 => x"07",
          9866 => x"5a",
          9867 => x"7d",
          9868 => x"fc",
          9869 => x"06",
          9870 => x"8c",
          9871 => x"06",
          9872 => x"79",
          9873 => x"fd",
          9874 => x"0b",
          9875 => x"7c",
          9876 => x"81",
          9877 => x"38",
          9878 => x"80",
          9879 => x"34",
          9880 => x"ba",
          9881 => x"3d",
          9882 => x"80",
          9883 => x"38",
          9884 => x"27",
          9885 => x"ff",
          9886 => x"7b",
          9887 => x"38",
          9888 => x"7d",
          9889 => x"5c",
          9890 => x"39",
          9891 => x"5a",
          9892 => x"74",
          9893 => x"f6",
          9894 => x"8c",
          9895 => x"ff",
          9896 => x"2a",
          9897 => x"55",
          9898 => x"c4",
          9899 => x"ff",
          9900 => x"9c",
          9901 => x"54",
          9902 => x"26",
          9903 => x"74",
          9904 => x"85",
          9905 => x"b4",
          9906 => x"b4",
          9907 => x"ff",
          9908 => x"59",
          9909 => x"80",
          9910 => x"75",
          9911 => x"81",
          9912 => x"70",
          9913 => x"56",
          9914 => x"ee",
          9915 => x"ff",
          9916 => x"80",
          9917 => x"bf",
          9918 => x"99",
          9919 => x"7d",
          9920 => x"81",
          9921 => x"53",
          9922 => x"59",
          9923 => x"93",
          9924 => x"07",
          9925 => x"06",
          9926 => x"83",
          9927 => x"58",
          9928 => x"7b",
          9929 => x"59",
          9930 => x"81",
          9931 => x"16",
          9932 => x"39",
          9933 => x"b3",
          9934 => x"b4",
          9935 => x"ff",
          9936 => x"78",
          9937 => x"ae",
          9938 => x"7a",
          9939 => x"1d",
          9940 => x"5b",
          9941 => x"34",
          9942 => x"d2",
          9943 => x"14",
          9944 => x"15",
          9945 => x"2b",
          9946 => x"07",
          9947 => x"1f",
          9948 => x"fd",
          9949 => x"1b",
          9950 => x"88",
          9951 => x"72",
          9952 => x"1b",
          9953 => x"05",
          9954 => x"79",
          9955 => x"5b",
          9956 => x"79",
          9957 => x"1d",
          9958 => x"76",
          9959 => x"09",
          9960 => x"a3",
          9961 => x"39",
          9962 => x"81",
          9963 => x"f6",
          9964 => x"0b",
          9965 => x"0c",
          9966 => x"04",
          9967 => x"67",
          9968 => x"05",
          9969 => x"33",
          9970 => x"80",
          9971 => x"7e",
          9972 => x"5b",
          9973 => x"2e",
          9974 => x"79",
          9975 => x"5b",
          9976 => x"26",
          9977 => x"ba",
          9978 => x"38",
          9979 => x"75",
          9980 => x"c7",
          9981 => x"e8",
          9982 => x"76",
          9983 => x"38",
          9984 => x"84",
          9985 => x"70",
          9986 => x"8c",
          9987 => x"2e",
          9988 => x"76",
          9989 => x"81",
          9990 => x"33",
          9991 => x"80",
          9992 => x"81",
          9993 => x"ff",
          9994 => x"84",
          9995 => x"81",
          9996 => x"81",
          9997 => x"7c",
          9998 => x"96",
          9999 => x"34",
         10000 => x"84",
         10001 => x"33",
         10002 => x"81",
         10003 => x"33",
         10004 => x"a4",
         10005 => x"8c",
         10006 => x"06",
         10007 => x"41",
         10008 => x"7f",
         10009 => x"78",
         10010 => x"38",
         10011 => x"81",
         10012 => x"58",
         10013 => x"38",
         10014 => x"83",
         10015 => x"0b",
         10016 => x"7a",
         10017 => x"81",
         10018 => x"b8",
         10019 => x"81",
         10020 => x"58",
         10021 => x"3f",
         10022 => x"08",
         10023 => x"38",
         10024 => x"59",
         10025 => x"0c",
         10026 => x"99",
         10027 => x"17",
         10028 => x"18",
         10029 => x"2b",
         10030 => x"83",
         10031 => x"d4",
         10032 => x"a5",
         10033 => x"26",
         10034 => x"ba",
         10035 => x"42",
         10036 => x"38",
         10037 => x"84",
         10038 => x"38",
         10039 => x"81",
         10040 => x"38",
         10041 => x"33",
         10042 => x"33",
         10043 => x"07",
         10044 => x"84",
         10045 => x"81",
         10046 => x"38",
         10047 => x"33",
         10048 => x"33",
         10049 => x"07",
         10050 => x"a4",
         10051 => x"17",
         10052 => x"82",
         10053 => x"90",
         10054 => x"2b",
         10055 => x"33",
         10056 => x"88",
         10057 => x"71",
         10058 => x"45",
         10059 => x"56",
         10060 => x"0c",
         10061 => x"33",
         10062 => x"80",
         10063 => x"ff",
         10064 => x"ff",
         10065 => x"59",
         10066 => x"81",
         10067 => x"38",
         10068 => x"06",
         10069 => x"80",
         10070 => x"5a",
         10071 => x"8a",
         10072 => x"59",
         10073 => x"87",
         10074 => x"18",
         10075 => x"61",
         10076 => x"80",
         10077 => x"80",
         10078 => x"71",
         10079 => x"56",
         10080 => x"18",
         10081 => x"8f",
         10082 => x"8d",
         10083 => x"98",
         10084 => x"17",
         10085 => x"18",
         10086 => x"2b",
         10087 => x"74",
         10088 => x"d8",
         10089 => x"33",
         10090 => x"71",
         10091 => x"88",
         10092 => x"14",
         10093 => x"07",
         10094 => x"33",
         10095 => x"44",
         10096 => x"42",
         10097 => x"17",
         10098 => x"18",
         10099 => x"2b",
         10100 => x"8d",
         10101 => x"2e",
         10102 => x"7d",
         10103 => x"2a",
         10104 => x"75",
         10105 => x"38",
         10106 => x"7a",
         10107 => x"ed",
         10108 => x"ba",
         10109 => x"84",
         10110 => x"80",
         10111 => x"38",
         10112 => x"08",
         10113 => x"ff",
         10114 => x"38",
         10115 => x"83",
         10116 => x"83",
         10117 => x"75",
         10118 => x"85",
         10119 => x"5d",
         10120 => x"9c",
         10121 => x"a4",
         10122 => x"1d",
         10123 => x"0c",
         10124 => x"1a",
         10125 => x"7c",
         10126 => x"87",
         10127 => x"22",
         10128 => x"7b",
         10129 => x"e0",
         10130 => x"ac",
         10131 => x"19",
         10132 => x"2e",
         10133 => x"10",
         10134 => x"2a",
         10135 => x"05",
         10136 => x"ff",
         10137 => x"59",
         10138 => x"a0",
         10139 => x"b8",
         10140 => x"94",
         10141 => x"0b",
         10142 => x"ff",
         10143 => x"18",
         10144 => x"2e",
         10145 => x"7c",
         10146 => x"d1",
         10147 => x"05",
         10148 => x"d1",
         10149 => x"86",
         10150 => x"d1",
         10151 => x"18",
         10152 => x"98",
         10153 => x"58",
         10154 => x"8c",
         10155 => x"0d",
         10156 => x"84",
         10157 => x"97",
         10158 => x"76",
         10159 => x"70",
         10160 => x"57",
         10161 => x"89",
         10162 => x"82",
         10163 => x"ff",
         10164 => x"5d",
         10165 => x"2e",
         10166 => x"80",
         10167 => x"e5",
         10168 => x"5c",
         10169 => x"5a",
         10170 => x"81",
         10171 => x"79",
         10172 => x"5b",
         10173 => x"12",
         10174 => x"77",
         10175 => x"38",
         10176 => x"81",
         10177 => x"55",
         10178 => x"58",
         10179 => x"89",
         10180 => x"70",
         10181 => x"58",
         10182 => x"70",
         10183 => x"55",
         10184 => x"09",
         10185 => x"38",
         10186 => x"38",
         10187 => x"70",
         10188 => x"07",
         10189 => x"07",
         10190 => x"7a",
         10191 => x"98",
         10192 => x"84",
         10193 => x"83",
         10194 => x"98",
         10195 => x"f9",
         10196 => x"80",
         10197 => x"38",
         10198 => x"81",
         10199 => x"58",
         10200 => x"38",
         10201 => x"c0",
         10202 => x"33",
         10203 => x"81",
         10204 => x"81",
         10205 => x"81",
         10206 => x"eb",
         10207 => x"70",
         10208 => x"07",
         10209 => x"77",
         10210 => x"75",
         10211 => x"83",
         10212 => x"3d",
         10213 => x"83",
         10214 => x"16",
         10215 => x"5b",
         10216 => x"a5",
         10217 => x"16",
         10218 => x"17",
         10219 => x"2b",
         10220 => x"07",
         10221 => x"33",
         10222 => x"88",
         10223 => x"1b",
         10224 => x"52",
         10225 => x"40",
         10226 => x"70",
         10227 => x"0c",
         10228 => x"17",
         10229 => x"80",
         10230 => x"38",
         10231 => x"1d",
         10232 => x"70",
         10233 => x"71",
         10234 => x"71",
         10235 => x"f0",
         10236 => x"1c",
         10237 => x"43",
         10238 => x"08",
         10239 => x"7a",
         10240 => x"fb",
         10241 => x"83",
         10242 => x"0b",
         10243 => x"7a",
         10244 => x"7a",
         10245 => x"38",
         10246 => x"53",
         10247 => x"81",
         10248 => x"ff",
         10249 => x"84",
         10250 => x"76",
         10251 => x"ff",
         10252 => x"74",
         10253 => x"84",
         10254 => x"38",
         10255 => x"7f",
         10256 => x"2b",
         10257 => x"83",
         10258 => x"d4",
         10259 => x"81",
         10260 => x"80",
         10261 => x"33",
         10262 => x"81",
         10263 => x"b7",
         10264 => x"eb",
         10265 => x"70",
         10266 => x"07",
         10267 => x"7f",
         10268 => x"81",
         10269 => x"38",
         10270 => x"81",
         10271 => x"80",
         10272 => x"81",
         10273 => x"58",
         10274 => x"09",
         10275 => x"38",
         10276 => x"76",
         10277 => x"38",
         10278 => x"f8",
         10279 => x"1a",
         10280 => x"5a",
         10281 => x"fe",
         10282 => x"a8",
         10283 => x"80",
         10284 => x"e5",
         10285 => x"58",
         10286 => x"05",
         10287 => x"70",
         10288 => x"33",
         10289 => x"ff",
         10290 => x"56",
         10291 => x"2e",
         10292 => x"75",
         10293 => x"38",
         10294 => x"8a",
         10295 => x"c0",
         10296 => x"7b",
         10297 => x"5d",
         10298 => x"81",
         10299 => x"71",
         10300 => x"1b",
         10301 => x"40",
         10302 => x"85",
         10303 => x"80",
         10304 => x"82",
         10305 => x"39",
         10306 => x"fa",
         10307 => x"84",
         10308 => x"97",
         10309 => x"75",
         10310 => x"2e",
         10311 => x"85",
         10312 => x"18",
         10313 => x"40",
         10314 => x"b7",
         10315 => x"84",
         10316 => x"97",
         10317 => x"83",
         10318 => x"18",
         10319 => x"5c",
         10320 => x"70",
         10321 => x"33",
         10322 => x"05",
         10323 => x"71",
         10324 => x"5b",
         10325 => x"77",
         10326 => x"d1",
         10327 => x"2e",
         10328 => x"0b",
         10329 => x"83",
         10330 => x"5a",
         10331 => x"81",
         10332 => x"7a",
         10333 => x"5c",
         10334 => x"31",
         10335 => x"58",
         10336 => x"80",
         10337 => x"38",
         10338 => x"e1",
         10339 => x"77",
         10340 => x"59",
         10341 => x"81",
         10342 => x"39",
         10343 => x"33",
         10344 => x"33",
         10345 => x"07",
         10346 => x"81",
         10347 => x"06",
         10348 => x"81",
         10349 => x"5a",
         10350 => x"78",
         10351 => x"83",
         10352 => x"7a",
         10353 => x"81",
         10354 => x"38",
         10355 => x"53",
         10356 => x"81",
         10357 => x"ff",
         10358 => x"84",
         10359 => x"80",
         10360 => x"ff",
         10361 => x"77",
         10362 => x"79",
         10363 => x"79",
         10364 => x"84",
         10365 => x"84",
         10366 => x"71",
         10367 => x"57",
         10368 => x"d4",
         10369 => x"81",
         10370 => x"38",
         10371 => x"11",
         10372 => x"33",
         10373 => x"71",
         10374 => x"81",
         10375 => x"72",
         10376 => x"75",
         10377 => x"5e",
         10378 => x"42",
         10379 => x"84",
         10380 => x"d2",
         10381 => x"06",
         10382 => x"84",
         10383 => x"11",
         10384 => x"33",
         10385 => x"71",
         10386 => x"81",
         10387 => x"72",
         10388 => x"75",
         10389 => x"47",
         10390 => x"5c",
         10391 => x"86",
         10392 => x"f2",
         10393 => x"06",
         10394 => x"84",
         10395 => x"11",
         10396 => x"33",
         10397 => x"71",
         10398 => x"81",
         10399 => x"72",
         10400 => x"75",
         10401 => x"94",
         10402 => x"84",
         10403 => x"11",
         10404 => x"33",
         10405 => x"71",
         10406 => x"81",
         10407 => x"72",
         10408 => x"75",
         10409 => x"62",
         10410 => x"59",
         10411 => x"5c",
         10412 => x"5b",
         10413 => x"77",
         10414 => x"e4",
         10415 => x"5d",
         10416 => x"e4",
         10417 => x"18",
         10418 => x"ec",
         10419 => x"0c",
         10420 => x"18",
         10421 => x"39",
         10422 => x"f8",
         10423 => x"7a",
         10424 => x"f2",
         10425 => x"54",
         10426 => x"53",
         10427 => x"53",
         10428 => x"52",
         10429 => x"b3",
         10430 => x"8c",
         10431 => x"09",
         10432 => x"a4",
         10433 => x"8c",
         10434 => x"34",
         10435 => x"a8",
         10436 => x"40",
         10437 => x"08",
         10438 => x"82",
         10439 => x"60",
         10440 => x"8d",
         10441 => x"8c",
         10442 => x"a0",
         10443 => x"74",
         10444 => x"91",
         10445 => x"81",
         10446 => x"e5",
         10447 => x"58",
         10448 => x"80",
         10449 => x"80",
         10450 => x"71",
         10451 => x"5f",
         10452 => x"7d",
         10453 => x"88",
         10454 => x"61",
         10455 => x"80",
         10456 => x"11",
         10457 => x"33",
         10458 => x"71",
         10459 => x"81",
         10460 => x"72",
         10461 => x"75",
         10462 => x"ac",
         10463 => x"7d",
         10464 => x"43",
         10465 => x"40",
         10466 => x"75",
         10467 => x"2e",
         10468 => x"82",
         10469 => x"39",
         10470 => x"f2",
         10471 => x"3d",
         10472 => x"83",
         10473 => x"39",
         10474 => x"f5",
         10475 => x"bf",
         10476 => x"b4",
         10477 => x"18",
         10478 => x"78",
         10479 => x"33",
         10480 => x"e7",
         10481 => x"39",
         10482 => x"02",
         10483 => x"33",
         10484 => x"93",
         10485 => x"5d",
         10486 => x"40",
         10487 => x"80",
         10488 => x"70",
         10489 => x"33",
         10490 => x"55",
         10491 => x"2e",
         10492 => x"73",
         10493 => x"ba",
         10494 => x"38",
         10495 => x"33",
         10496 => x"24",
         10497 => x"73",
         10498 => x"d1",
         10499 => x"08",
         10500 => x"80",
         10501 => x"80",
         10502 => x"54",
         10503 => x"86",
         10504 => x"34",
         10505 => x"75",
         10506 => x"7c",
         10507 => x"38",
         10508 => x"3d",
         10509 => x"05",
         10510 => x"3f",
         10511 => x"08",
         10512 => x"ba",
         10513 => x"3d",
         10514 => x"0b",
         10515 => x"0c",
         10516 => x"04",
         10517 => x"11",
         10518 => x"06",
         10519 => x"73",
         10520 => x"38",
         10521 => x"81",
         10522 => x"05",
         10523 => x"79",
         10524 => x"38",
         10525 => x"83",
         10526 => x"5f",
         10527 => x"7e",
         10528 => x"70",
         10529 => x"33",
         10530 => x"05",
         10531 => x"9f",
         10532 => x"55",
         10533 => x"89",
         10534 => x"70",
         10535 => x"56",
         10536 => x"16",
         10537 => x"26",
         10538 => x"16",
         10539 => x"06",
         10540 => x"30",
         10541 => x"58",
         10542 => x"2e",
         10543 => x"85",
         10544 => x"be",
         10545 => x"32",
         10546 => x"72",
         10547 => x"79",
         10548 => x"54",
         10549 => x"92",
         10550 => x"84",
         10551 => x"83",
         10552 => x"99",
         10553 => x"fe",
         10554 => x"83",
         10555 => x"7a",
         10556 => x"54",
         10557 => x"e6",
         10558 => x"02",
         10559 => x"fb",
         10560 => x"59",
         10561 => x"80",
         10562 => x"74",
         10563 => x"54",
         10564 => x"05",
         10565 => x"84",
         10566 => x"ed",
         10567 => x"ba",
         10568 => x"84",
         10569 => x"80",
         10570 => x"80",
         10571 => x"56",
         10572 => x"8c",
         10573 => x"0d",
         10574 => x"6d",
         10575 => x"70",
         10576 => x"9a",
         10577 => x"8c",
         10578 => x"ba",
         10579 => x"2e",
         10580 => x"77",
         10581 => x"7c",
         10582 => x"ca",
         10583 => x"2e",
         10584 => x"76",
         10585 => x"ea",
         10586 => x"07",
         10587 => x"bb",
         10588 => x"2a",
         10589 => x"7a",
         10590 => x"d1",
         10591 => x"11",
         10592 => x"33",
         10593 => x"07",
         10594 => x"42",
         10595 => x"56",
         10596 => x"84",
         10597 => x"0b",
         10598 => x"80",
         10599 => x"34",
         10600 => x"17",
         10601 => x"0b",
         10602 => x"66",
         10603 => x"8b",
         10604 => x"67",
         10605 => x"0b",
         10606 => x"80",
         10607 => x"34",
         10608 => x"7c",
         10609 => x"a9",
         10610 => x"80",
         10611 => x"34",
         10612 => x"1c",
         10613 => x"9e",
         10614 => x"0b",
         10615 => x"7e",
         10616 => x"83",
         10617 => x"80",
         10618 => x"38",
         10619 => x"08",
         10620 => x"53",
         10621 => x"81",
         10622 => x"38",
         10623 => x"7c",
         10624 => x"38",
         10625 => x"79",
         10626 => x"39",
         10627 => x"05",
         10628 => x"2b",
         10629 => x"80",
         10630 => x"38",
         10631 => x"06",
         10632 => x"fe",
         10633 => x"fe",
         10634 => x"80",
         10635 => x"70",
         10636 => x"06",
         10637 => x"82",
         10638 => x"81",
         10639 => x"5e",
         10640 => x"89",
         10641 => x"06",
         10642 => x"f6",
         10643 => x"2a",
         10644 => x"75",
         10645 => x"38",
         10646 => x"07",
         10647 => x"11",
         10648 => x"0c",
         10649 => x"0c",
         10650 => x"33",
         10651 => x"71",
         10652 => x"73",
         10653 => x"40",
         10654 => x"83",
         10655 => x"38",
         10656 => x"0c",
         10657 => x"11",
         10658 => x"33",
         10659 => x"71",
         10660 => x"81",
         10661 => x"72",
         10662 => x"75",
         10663 => x"70",
         10664 => x"0c",
         10665 => x"51",
         10666 => x"57",
         10667 => x"1a",
         10668 => x"23",
         10669 => x"34",
         10670 => x"1a",
         10671 => x"9c",
         10672 => x"85",
         10673 => x"55",
         10674 => x"84",
         10675 => x"80",
         10676 => x"38",
         10677 => x"0c",
         10678 => x"70",
         10679 => x"52",
         10680 => x"30",
         10681 => x"80",
         10682 => x"79",
         10683 => x"92",
         10684 => x"76",
         10685 => x"7d",
         10686 => x"86",
         10687 => x"78",
         10688 => x"db",
         10689 => x"8c",
         10690 => x"ba",
         10691 => x"26",
         10692 => x"57",
         10693 => x"08",
         10694 => x"cb",
         10695 => x"31",
         10696 => x"02",
         10697 => x"33",
         10698 => x"7d",
         10699 => x"82",
         10700 => x"55",
         10701 => x"fc",
         10702 => x"57",
         10703 => x"fb",
         10704 => x"57",
         10705 => x"fb",
         10706 => x"57",
         10707 => x"fb",
         10708 => x"51",
         10709 => x"84",
         10710 => x"78",
         10711 => x"57",
         10712 => x"38",
         10713 => x"7a",
         10714 => x"57",
         10715 => x"39",
         10716 => x"94",
         10717 => x"98",
         10718 => x"2b",
         10719 => x"5d",
         10720 => x"fc",
         10721 => x"7c",
         10722 => x"bd",
         10723 => x"79",
         10724 => x"cb",
         10725 => x"8c",
         10726 => x"ba",
         10727 => x"2e",
         10728 => x"84",
         10729 => x"81",
         10730 => x"38",
         10731 => x"08",
         10732 => x"99",
         10733 => x"74",
         10734 => x"ff",
         10735 => x"84",
         10736 => x"83",
         10737 => x"17",
         10738 => x"94",
         10739 => x"56",
         10740 => x"27",
         10741 => x"81",
         10742 => x"0c",
         10743 => x"81",
         10744 => x"84",
         10745 => x"55",
         10746 => x"ff",
         10747 => x"d9",
         10748 => x"94",
         10749 => x"0b",
         10750 => x"fb",
         10751 => x"16",
         10752 => x"33",
         10753 => x"71",
         10754 => x"7e",
         10755 => x"5b",
         10756 => x"17",
         10757 => x"8f",
         10758 => x"0b",
         10759 => x"80",
         10760 => x"17",
         10761 => x"a0",
         10762 => x"34",
         10763 => x"5e",
         10764 => x"17",
         10765 => x"9b",
         10766 => x"33",
         10767 => x"2e",
         10768 => x"fb",
         10769 => x"a9",
         10770 => x"7f",
         10771 => x"57",
         10772 => x"08",
         10773 => x"38",
         10774 => x"5a",
         10775 => x"09",
         10776 => x"38",
         10777 => x"53",
         10778 => x"81",
         10779 => x"ff",
         10780 => x"84",
         10781 => x"80",
         10782 => x"ff",
         10783 => x"76",
         10784 => x"7e",
         10785 => x"1d",
         10786 => x"57",
         10787 => x"fb",
         10788 => x"79",
         10789 => x"39",
         10790 => x"16",
         10791 => x"16",
         10792 => x"17",
         10793 => x"ff",
         10794 => x"84",
         10795 => x"7d",
         10796 => x"06",
         10797 => x"84",
         10798 => x"83",
         10799 => x"16",
         10800 => x"08",
         10801 => x"8c",
         10802 => x"74",
         10803 => x"27",
         10804 => x"82",
         10805 => x"74",
         10806 => x"81",
         10807 => x"38",
         10808 => x"16",
         10809 => x"08",
         10810 => x"52",
         10811 => x"51",
         10812 => x"3f",
         10813 => x"ec",
         10814 => x"1a",
         10815 => x"f8",
         10816 => x"98",
         10817 => x"f8",
         10818 => x"83",
         10819 => x"79",
         10820 => x"9a",
         10821 => x"19",
         10822 => x"fe",
         10823 => x"5a",
         10824 => x"f9",
         10825 => x"1a",
         10826 => x"29",
         10827 => x"05",
         10828 => x"80",
         10829 => x"38",
         10830 => x"15",
         10831 => x"76",
         10832 => x"39",
         10833 => x"0c",
         10834 => x"e4",
         10835 => x"80",
         10836 => x"da",
         10837 => x"8c",
         10838 => x"79",
         10839 => x"39",
         10840 => x"5b",
         10841 => x"f0",
         10842 => x"65",
         10843 => x"40",
         10844 => x"7e",
         10845 => x"79",
         10846 => x"38",
         10847 => x"75",
         10848 => x"38",
         10849 => x"74",
         10850 => x"38",
         10851 => x"84",
         10852 => x"59",
         10853 => x"84",
         10854 => x"55",
         10855 => x"55",
         10856 => x"38",
         10857 => x"55",
         10858 => x"38",
         10859 => x"81",
         10860 => x"56",
         10861 => x"81",
         10862 => x"1a",
         10863 => x"08",
         10864 => x"56",
         10865 => x"81",
         10866 => x"80",
         10867 => x"38",
         10868 => x"83",
         10869 => x"7a",
         10870 => x"8a",
         10871 => x"05",
         10872 => x"06",
         10873 => x"38",
         10874 => x"38",
         10875 => x"55",
         10876 => x"84",
         10877 => x"ff",
         10878 => x"38",
         10879 => x"0c",
         10880 => x"1a",
         10881 => x"9c",
         10882 => x"05",
         10883 => x"60",
         10884 => x"38",
         10885 => x"70",
         10886 => x"1b",
         10887 => x"56",
         10888 => x"83",
         10889 => x"15",
         10890 => x"59",
         10891 => x"2e",
         10892 => x"77",
         10893 => x"75",
         10894 => x"75",
         10895 => x"77",
         10896 => x"7c",
         10897 => x"33",
         10898 => x"e0",
         10899 => x"8c",
         10900 => x"38",
         10901 => x"33",
         10902 => x"80",
         10903 => x"b4",
         10904 => x"31",
         10905 => x"27",
         10906 => x"80",
         10907 => x"1e",
         10908 => x"58",
         10909 => x"81",
         10910 => x"77",
         10911 => x"59",
         10912 => x"55",
         10913 => x"77",
         10914 => x"7b",
         10915 => x"08",
         10916 => x"78",
         10917 => x"08",
         10918 => x"94",
         10919 => x"5c",
         10920 => x"38",
         10921 => x"84",
         10922 => x"92",
         10923 => x"74",
         10924 => x"0c",
         10925 => x"04",
         10926 => x"8e",
         10927 => x"08",
         10928 => x"ff",
         10929 => x"71",
         10930 => x"7b",
         10931 => x"38",
         10932 => x"56",
         10933 => x"77",
         10934 => x"80",
         10935 => x"33",
         10936 => x"5f",
         10937 => x"09",
         10938 => x"e4",
         10939 => x"76",
         10940 => x"52",
         10941 => x"51",
         10942 => x"3f",
         10943 => x"08",
         10944 => x"38",
         10945 => x"5b",
         10946 => x"0c",
         10947 => x"38",
         10948 => x"08",
         10949 => x"11",
         10950 => x"58",
         10951 => x"59",
         10952 => x"fe",
         10953 => x"70",
         10954 => x"33",
         10955 => x"05",
         10956 => x"16",
         10957 => x"2e",
         10958 => x"74",
         10959 => x"56",
         10960 => x"81",
         10961 => x"ff",
         10962 => x"da",
         10963 => x"39",
         10964 => x"19",
         10965 => x"19",
         10966 => x"1a",
         10967 => x"ff",
         10968 => x"81",
         10969 => x"8c",
         10970 => x"09",
         10971 => x"9c",
         10972 => x"8c",
         10973 => x"34",
         10974 => x"a8",
         10975 => x"84",
         10976 => x"5c",
         10977 => x"1a",
         10978 => x"e1",
         10979 => x"33",
         10980 => x"2e",
         10981 => x"fe",
         10982 => x"54",
         10983 => x"a0",
         10984 => x"53",
         10985 => x"19",
         10986 => x"9d",
         10987 => x"5b",
         10988 => x"76",
         10989 => x"94",
         10990 => x"fe",
         10991 => x"1a",
         10992 => x"51",
         10993 => x"3f",
         10994 => x"08",
         10995 => x"39",
         10996 => x"51",
         10997 => x"3f",
         10998 => x"08",
         10999 => x"74",
         11000 => x"74",
         11001 => x"57",
         11002 => x"81",
         11003 => x"34",
         11004 => x"ba",
         11005 => x"3d",
         11006 => x"0b",
         11007 => x"82",
         11008 => x"8c",
         11009 => x"0d",
         11010 => x"0d",
         11011 => x"66",
         11012 => x"5a",
         11013 => x"89",
         11014 => x"2e",
         11015 => x"08",
         11016 => x"2e",
         11017 => x"33",
         11018 => x"2e",
         11019 => x"16",
         11020 => x"22",
         11021 => x"78",
         11022 => x"38",
         11023 => x"41",
         11024 => x"82",
         11025 => x"1a",
         11026 => x"82",
         11027 => x"1a",
         11028 => x"2a",
         11029 => x"58",
         11030 => x"80",
         11031 => x"38",
         11032 => x"7b",
         11033 => x"7b",
         11034 => x"38",
         11035 => x"7a",
         11036 => x"81",
         11037 => x"ff",
         11038 => x"82",
         11039 => x"8a",
         11040 => x"05",
         11041 => x"06",
         11042 => x"aa",
         11043 => x"9e",
         11044 => x"08",
         11045 => x"2e",
         11046 => x"74",
         11047 => x"a1",
         11048 => x"2e",
         11049 => x"74",
         11050 => x"88",
         11051 => x"38",
         11052 => x"0c",
         11053 => x"16",
         11054 => x"08",
         11055 => x"38",
         11056 => x"fe",
         11057 => x"08",
         11058 => x"58",
         11059 => x"85",
         11060 => x"16",
         11061 => x"29",
         11062 => x"05",
         11063 => x"80",
         11064 => x"38",
         11065 => x"89",
         11066 => x"77",
         11067 => x"98",
         11068 => x"5f",
         11069 => x"85",
         11070 => x"31",
         11071 => x"7b",
         11072 => x"81",
         11073 => x"ff",
         11074 => x"84",
         11075 => x"85",
         11076 => x"b4",
         11077 => x"31",
         11078 => x"78",
         11079 => x"84",
         11080 => x"18",
         11081 => x"1f",
         11082 => x"74",
         11083 => x"56",
         11084 => x"81",
         11085 => x"ff",
         11086 => x"ef",
         11087 => x"75",
         11088 => x"77",
         11089 => x"7a",
         11090 => x"08",
         11091 => x"79",
         11092 => x"08",
         11093 => x"94",
         11094 => x"1e",
         11095 => x"57",
         11096 => x"75",
         11097 => x"74",
         11098 => x"1b",
         11099 => x"85",
         11100 => x"33",
         11101 => x"c0",
         11102 => x"90",
         11103 => x"56",
         11104 => x"8c",
         11105 => x"0d",
         11106 => x"ba",
         11107 => x"3d",
         11108 => x"16",
         11109 => x"82",
         11110 => x"56",
         11111 => x"60",
         11112 => x"59",
         11113 => x"ff",
         11114 => x"71",
         11115 => x"7a",
         11116 => x"38",
         11117 => x"57",
         11118 => x"78",
         11119 => x"80",
         11120 => x"33",
         11121 => x"5f",
         11122 => x"09",
         11123 => x"d5",
         11124 => x"77",
         11125 => x"52",
         11126 => x"51",
         11127 => x"3f",
         11128 => x"08",
         11129 => x"38",
         11130 => x"5c",
         11131 => x"0c",
         11132 => x"38",
         11133 => x"08",
         11134 => x"11",
         11135 => x"05",
         11136 => x"58",
         11137 => x"95",
         11138 => x"81",
         11139 => x"75",
         11140 => x"57",
         11141 => x"56",
         11142 => x"60",
         11143 => x"83",
         11144 => x"a3",
         11145 => x"b4",
         11146 => x"b8",
         11147 => x"81",
         11148 => x"40",
         11149 => x"3f",
         11150 => x"ba",
         11151 => x"2e",
         11152 => x"ff",
         11153 => x"ba",
         11154 => x"17",
         11155 => x"08",
         11156 => x"31",
         11157 => x"08",
         11158 => x"a0",
         11159 => x"fe",
         11160 => x"16",
         11161 => x"82",
         11162 => x"06",
         11163 => x"81",
         11164 => x"08",
         11165 => x"05",
         11166 => x"81",
         11167 => x"ff",
         11168 => x"7e",
         11169 => x"39",
         11170 => x"57",
         11171 => x"77",
         11172 => x"83",
         11173 => x"7f",
         11174 => x"60",
         11175 => x"0c",
         11176 => x"58",
         11177 => x"9c",
         11178 => x"fd",
         11179 => x"1a",
         11180 => x"51",
         11181 => x"3f",
         11182 => x"08",
         11183 => x"8c",
         11184 => x"38",
         11185 => x"58",
         11186 => x"76",
         11187 => x"ff",
         11188 => x"84",
         11189 => x"55",
         11190 => x"08",
         11191 => x"e4",
         11192 => x"b4",
         11193 => x"b8",
         11194 => x"81",
         11195 => x"57",
         11196 => x"3f",
         11197 => x"08",
         11198 => x"84",
         11199 => x"83",
         11200 => x"16",
         11201 => x"08",
         11202 => x"a0",
         11203 => x"fd",
         11204 => x"16",
         11205 => x"82",
         11206 => x"06",
         11207 => x"81",
         11208 => x"08",
         11209 => x"05",
         11210 => x"81",
         11211 => x"ff",
         11212 => x"60",
         11213 => x"39",
         11214 => x"51",
         11215 => x"3f",
         11216 => x"08",
         11217 => x"74",
         11218 => x"74",
         11219 => x"57",
         11220 => x"81",
         11221 => x"08",
         11222 => x"70",
         11223 => x"33",
         11224 => x"96",
         11225 => x"ba",
         11226 => x"c6",
         11227 => x"8c",
         11228 => x"34",
         11229 => x"a8",
         11230 => x"55",
         11231 => x"08",
         11232 => x"38",
         11233 => x"58",
         11234 => x"09",
         11235 => x"8b",
         11236 => x"b4",
         11237 => x"17",
         11238 => x"76",
         11239 => x"33",
         11240 => x"87",
         11241 => x"b4",
         11242 => x"1b",
         11243 => x"fd",
         11244 => x"0b",
         11245 => x"81",
         11246 => x"8c",
         11247 => x"0d",
         11248 => x"91",
         11249 => x"0b",
         11250 => x"0c",
         11251 => x"04",
         11252 => x"7d",
         11253 => x"77",
         11254 => x"38",
         11255 => x"75",
         11256 => x"38",
         11257 => x"74",
         11258 => x"38",
         11259 => x"84",
         11260 => x"59",
         11261 => x"83",
         11262 => x"55",
         11263 => x"56",
         11264 => x"38",
         11265 => x"70",
         11266 => x"06",
         11267 => x"80",
         11268 => x"38",
         11269 => x"08",
         11270 => x"17",
         11271 => x"ac",
         11272 => x"33",
         11273 => x"bc",
         11274 => x"78",
         11275 => x"52",
         11276 => x"51",
         11277 => x"3f",
         11278 => x"08",
         11279 => x"38",
         11280 => x"56",
         11281 => x"0c",
         11282 => x"38",
         11283 => x"8b",
         11284 => x"07",
         11285 => x"8b",
         11286 => x"08",
         11287 => x"70",
         11288 => x"06",
         11289 => x"7a",
         11290 => x"7a",
         11291 => x"79",
         11292 => x"9c",
         11293 => x"96",
         11294 => x"5b",
         11295 => x"81",
         11296 => x"18",
         11297 => x"7b",
         11298 => x"2a",
         11299 => x"18",
         11300 => x"2a",
         11301 => x"18",
         11302 => x"2a",
         11303 => x"18",
         11304 => x"34",
         11305 => x"18",
         11306 => x"98",
         11307 => x"cc",
         11308 => x"34",
         11309 => x"18",
         11310 => x"93",
         11311 => x"5b",
         11312 => x"1c",
         11313 => x"ff",
         11314 => x"84",
         11315 => x"90",
         11316 => x"bf",
         11317 => x"79",
         11318 => x"75",
         11319 => x"0c",
         11320 => x"04",
         11321 => x"17",
         11322 => x"17",
         11323 => x"18",
         11324 => x"ff",
         11325 => x"81",
         11326 => x"8c",
         11327 => x"38",
         11328 => x"08",
         11329 => x"b4",
         11330 => x"18",
         11331 => x"ba",
         11332 => x"55",
         11333 => x"08",
         11334 => x"38",
         11335 => x"55",
         11336 => x"09",
         11337 => x"81",
         11338 => x"b4",
         11339 => x"18",
         11340 => x"7a",
         11341 => x"33",
         11342 => x"ef",
         11343 => x"fd",
         11344 => x"90",
         11345 => x"94",
         11346 => x"88",
         11347 => x"95",
         11348 => x"18",
         11349 => x"7b",
         11350 => x"2a",
         11351 => x"18",
         11352 => x"2a",
         11353 => x"18",
         11354 => x"2a",
         11355 => x"18",
         11356 => x"34",
         11357 => x"18",
         11358 => x"98",
         11359 => x"cc",
         11360 => x"34",
         11361 => x"18",
         11362 => x"93",
         11363 => x"5b",
         11364 => x"1c",
         11365 => x"ff",
         11366 => x"84",
         11367 => x"90",
         11368 => x"bf",
         11369 => x"79",
         11370 => x"fe",
         11371 => x"16",
         11372 => x"90",
         11373 => x"ba",
         11374 => x"06",
         11375 => x"ba",
         11376 => x"08",
         11377 => x"b4",
         11378 => x"0d",
         11379 => x"55",
         11380 => x"84",
         11381 => x"54",
         11382 => x"08",
         11383 => x"56",
         11384 => x"9e",
         11385 => x"53",
         11386 => x"96",
         11387 => x"52",
         11388 => x"8e",
         11389 => x"22",
         11390 => x"58",
         11391 => x"2e",
         11392 => x"52",
         11393 => x"54",
         11394 => x"75",
         11395 => x"84",
         11396 => x"89",
         11397 => x"81",
         11398 => x"ff",
         11399 => x"84",
         11400 => x"81",
         11401 => x"da",
         11402 => x"08",
         11403 => x"39",
         11404 => x"ff",
         11405 => x"57",
         11406 => x"2e",
         11407 => x"70",
         11408 => x"33",
         11409 => x"52",
         11410 => x"2e",
         11411 => x"ee",
         11412 => x"2e",
         11413 => x"d1",
         11414 => x"80",
         11415 => x"38",
         11416 => x"e8",
         11417 => x"84",
         11418 => x"8c",
         11419 => x"8b",
         11420 => x"8c",
         11421 => x"0d",
         11422 => x"d0",
         11423 => x"ff",
         11424 => x"53",
         11425 => x"91",
         11426 => x"73",
         11427 => x"d0",
         11428 => x"73",
         11429 => x"f5",
         11430 => x"83",
         11431 => x"58",
         11432 => x"56",
         11433 => x"81",
         11434 => x"75",
         11435 => x"57",
         11436 => x"12",
         11437 => x"70",
         11438 => x"38",
         11439 => x"81",
         11440 => x"54",
         11441 => x"51",
         11442 => x"89",
         11443 => x"70",
         11444 => x"54",
         11445 => x"70",
         11446 => x"51",
         11447 => x"09",
         11448 => x"38",
         11449 => x"38",
         11450 => x"70",
         11451 => x"07",
         11452 => x"07",
         11453 => x"76",
         11454 => x"38",
         11455 => x"1b",
         11456 => x"78",
         11457 => x"38",
         11458 => x"cf",
         11459 => x"24",
         11460 => x"76",
         11461 => x"c3",
         11462 => x"0d",
         11463 => x"3d",
         11464 => x"99",
         11465 => x"94",
         11466 => x"8c",
         11467 => x"ba",
         11468 => x"2e",
         11469 => x"84",
         11470 => x"98",
         11471 => x"7a",
         11472 => x"98",
         11473 => x"51",
         11474 => x"84",
         11475 => x"55",
         11476 => x"08",
         11477 => x"02",
         11478 => x"33",
         11479 => x"58",
         11480 => x"24",
         11481 => x"02",
         11482 => x"70",
         11483 => x"06",
         11484 => x"80",
         11485 => x"7a",
         11486 => x"33",
         11487 => x"71",
         11488 => x"73",
         11489 => x"5b",
         11490 => x"83",
         11491 => x"76",
         11492 => x"74",
         11493 => x"0c",
         11494 => x"04",
         11495 => x"08",
         11496 => x"81",
         11497 => x"38",
         11498 => x"ba",
         11499 => x"3d",
         11500 => x"16",
         11501 => x"33",
         11502 => x"71",
         11503 => x"79",
         11504 => x"0c",
         11505 => x"39",
         11506 => x"12",
         11507 => x"84",
         11508 => x"98",
         11509 => x"ff",
         11510 => x"80",
         11511 => x"80",
         11512 => x"5d",
         11513 => x"34",
         11514 => x"e4",
         11515 => x"05",
         11516 => x"3d",
         11517 => x"3f",
         11518 => x"08",
         11519 => x"8c",
         11520 => x"38",
         11521 => x"3d",
         11522 => x"98",
         11523 => x"dd",
         11524 => x"80",
         11525 => x"5b",
         11526 => x"2e",
         11527 => x"80",
         11528 => x"3d",
         11529 => x"52",
         11530 => x"a4",
         11531 => x"ba",
         11532 => x"84",
         11533 => x"83",
         11534 => x"80",
         11535 => x"58",
         11536 => x"08",
         11537 => x"38",
         11538 => x"08",
         11539 => x"5f",
         11540 => x"c7",
         11541 => x"76",
         11542 => x"52",
         11543 => x"51",
         11544 => x"3f",
         11545 => x"08",
         11546 => x"38",
         11547 => x"59",
         11548 => x"0c",
         11549 => x"38",
         11550 => x"08",
         11551 => x"9a",
         11552 => x"88",
         11553 => x"70",
         11554 => x"59",
         11555 => x"83",
         11556 => x"38",
         11557 => x"3d",
         11558 => x"7a",
         11559 => x"b7",
         11560 => x"8c",
         11561 => x"ba",
         11562 => x"9f",
         11563 => x"7a",
         11564 => x"f5",
         11565 => x"8c",
         11566 => x"ba",
         11567 => x"38",
         11568 => x"08",
         11569 => x"9a",
         11570 => x"88",
         11571 => x"70",
         11572 => x"59",
         11573 => x"83",
         11574 => x"38",
         11575 => x"a4",
         11576 => x"8c",
         11577 => x"51",
         11578 => x"3f",
         11579 => x"08",
         11580 => x"8c",
         11581 => x"ff",
         11582 => x"84",
         11583 => x"38",
         11584 => x"38",
         11585 => x"fd",
         11586 => x"7a",
         11587 => x"89",
         11588 => x"82",
         11589 => x"57",
         11590 => x"90",
         11591 => x"56",
         11592 => x"17",
         11593 => x"57",
         11594 => x"38",
         11595 => x"75",
         11596 => x"95",
         11597 => x"2e",
         11598 => x"17",
         11599 => x"ff",
         11600 => x"3d",
         11601 => x"19",
         11602 => x"59",
         11603 => x"33",
         11604 => x"eb",
         11605 => x"80",
         11606 => x"11",
         11607 => x"7e",
         11608 => x"3d",
         11609 => x"fd",
         11610 => x"60",
         11611 => x"38",
         11612 => x"d1",
         11613 => x"10",
         11614 => x"fc",
         11615 => x"70",
         11616 => x"59",
         11617 => x"7a",
         11618 => x"81",
         11619 => x"70",
         11620 => x"5a",
         11621 => x"82",
         11622 => x"78",
         11623 => x"80",
         11624 => x"27",
         11625 => x"16",
         11626 => x"7c",
         11627 => x"5e",
         11628 => x"57",
         11629 => x"ee",
         11630 => x"70",
         11631 => x"34",
         11632 => x"09",
         11633 => x"df",
         11634 => x"80",
         11635 => x"84",
         11636 => x"80",
         11637 => x"04",
         11638 => x"94",
         11639 => x"98",
         11640 => x"2b",
         11641 => x"59",
         11642 => x"f0",
         11643 => x"33",
         11644 => x"71",
         11645 => x"90",
         11646 => x"07",
         11647 => x"0c",
         11648 => x"52",
         11649 => x"a0",
         11650 => x"ba",
         11651 => x"84",
         11652 => x"80",
         11653 => x"38",
         11654 => x"81",
         11655 => x"08",
         11656 => x"70",
         11657 => x"33",
         11658 => x"88",
         11659 => x"59",
         11660 => x"08",
         11661 => x"84",
         11662 => x"83",
         11663 => x"16",
         11664 => x"08",
         11665 => x"8c",
         11666 => x"74",
         11667 => x"27",
         11668 => x"82",
         11669 => x"74",
         11670 => x"81",
         11671 => x"38",
         11672 => x"16",
         11673 => x"08",
         11674 => x"52",
         11675 => x"51",
         11676 => x"3f",
         11677 => x"dd",
         11678 => x"80",
         11679 => x"11",
         11680 => x"7b",
         11681 => x"84",
         11682 => x"70",
         11683 => x"e5",
         11684 => x"08",
         11685 => x"59",
         11686 => x"7e",
         11687 => x"81",
         11688 => x"38",
         11689 => x"80",
         11690 => x"18",
         11691 => x"5a",
         11692 => x"70",
         11693 => x"34",
         11694 => x"fe",
         11695 => x"e5",
         11696 => x"81",
         11697 => x"79",
         11698 => x"81",
         11699 => x"7f",
         11700 => x"38",
         11701 => x"82",
         11702 => x"34",
         11703 => x"8c",
         11704 => x"3d",
         11705 => x"3d",
         11706 => x"58",
         11707 => x"74",
         11708 => x"38",
         11709 => x"73",
         11710 => x"38",
         11711 => x"72",
         11712 => x"38",
         11713 => x"84",
         11714 => x"59",
         11715 => x"83",
         11716 => x"53",
         11717 => x"53",
         11718 => x"38",
         11719 => x"53",
         11720 => x"38",
         11721 => x"56",
         11722 => x"81",
         11723 => x"15",
         11724 => x"58",
         11725 => x"81",
         11726 => x"8a",
         11727 => x"89",
         11728 => x"56",
         11729 => x"81",
         11730 => x"52",
         11731 => x"fd",
         11732 => x"84",
         11733 => x"ff",
         11734 => x"70",
         11735 => x"fd",
         11736 => x"84",
         11737 => x"73",
         11738 => x"38",
         11739 => x"06",
         11740 => x"0c",
         11741 => x"98",
         11742 => x"58",
         11743 => x"2e",
         11744 => x"75",
         11745 => x"d9",
         11746 => x"31",
         11747 => x"17",
         11748 => x"90",
         11749 => x"81",
         11750 => x"51",
         11751 => x"80",
         11752 => x"38",
         11753 => x"51",
         11754 => x"3f",
         11755 => x"08",
         11756 => x"8c",
         11757 => x"81",
         11758 => x"ff",
         11759 => x"81",
         11760 => x"b4",
         11761 => x"73",
         11762 => x"27",
         11763 => x"73",
         11764 => x"ff",
         11765 => x"0b",
         11766 => x"81",
         11767 => x"ba",
         11768 => x"3d",
         11769 => x"15",
         11770 => x"2a",
         11771 => x"58",
         11772 => x"38",
         11773 => x"08",
         11774 => x"58",
         11775 => x"09",
         11776 => x"b6",
         11777 => x"16",
         11778 => x"08",
         11779 => x"27",
         11780 => x"8c",
         11781 => x"15",
         11782 => x"07",
         11783 => x"16",
         11784 => x"ff",
         11785 => x"80",
         11786 => x"9c",
         11787 => x"2e",
         11788 => x"9c",
         11789 => x"0b",
         11790 => x"0c",
         11791 => x"04",
         11792 => x"16",
         11793 => x"08",
         11794 => x"2e",
         11795 => x"73",
         11796 => x"73",
         11797 => x"c2",
         11798 => x"39",
         11799 => x"08",
         11800 => x"08",
         11801 => x"0c",
         11802 => x"06",
         11803 => x"2e",
         11804 => x"fe",
         11805 => x"08",
         11806 => x"55",
         11807 => x"27",
         11808 => x"8a",
         11809 => x"71",
         11810 => x"08",
         11811 => x"2a",
         11812 => x"53",
         11813 => x"80",
         11814 => x"15",
         11815 => x"e9",
         11816 => x"74",
         11817 => x"b7",
         11818 => x"8c",
         11819 => x"8a",
         11820 => x"33",
         11821 => x"a2",
         11822 => x"8c",
         11823 => x"53",
         11824 => x"38",
         11825 => x"54",
         11826 => x"39",
         11827 => x"51",
         11828 => x"3f",
         11829 => x"08",
         11830 => x"8c",
         11831 => x"98",
         11832 => x"8c",
         11833 => x"fd",
         11834 => x"ba",
         11835 => x"16",
         11836 => x"16",
         11837 => x"39",
         11838 => x"16",
         11839 => x"84",
         11840 => x"8b",
         11841 => x"f6",
         11842 => x"56",
         11843 => x"80",
         11844 => x"80",
         11845 => x"fc",
         11846 => x"3d",
         11847 => x"c5",
         11848 => x"ba",
         11849 => x"84",
         11850 => x"80",
         11851 => x"80",
         11852 => x"54",
         11853 => x"8c",
         11854 => x"0d",
         11855 => x"0c",
         11856 => x"51",
         11857 => x"3f",
         11858 => x"08",
         11859 => x"8c",
         11860 => x"38",
         11861 => x"70",
         11862 => x"59",
         11863 => x"af",
         11864 => x"33",
         11865 => x"81",
         11866 => x"79",
         11867 => x"c5",
         11868 => x"08",
         11869 => x"9a",
         11870 => x"88",
         11871 => x"70",
         11872 => x"5a",
         11873 => x"83",
         11874 => x"77",
         11875 => x"7a",
         11876 => x"22",
         11877 => x"74",
         11878 => x"ff",
         11879 => x"84",
         11880 => x"55",
         11881 => x"8d",
         11882 => x"2e",
         11883 => x"80",
         11884 => x"fe",
         11885 => x"80",
         11886 => x"f6",
         11887 => x"33",
         11888 => x"71",
         11889 => x"90",
         11890 => x"07",
         11891 => x"5a",
         11892 => x"39",
         11893 => x"78",
         11894 => x"74",
         11895 => x"38",
         11896 => x"72",
         11897 => x"38",
         11898 => x"71",
         11899 => x"38",
         11900 => x"84",
         11901 => x"52",
         11902 => x"94",
         11903 => x"71",
         11904 => x"38",
         11905 => x"73",
         11906 => x"0c",
         11907 => x"04",
         11908 => x"51",
         11909 => x"3f",
         11910 => x"08",
         11911 => x"71",
         11912 => x"75",
         11913 => x"d7",
         11914 => x"0d",
         11915 => x"55",
         11916 => x"80",
         11917 => x"74",
         11918 => x"80",
         11919 => x"73",
         11920 => x"80",
         11921 => x"86",
         11922 => x"16",
         11923 => x"72",
         11924 => x"97",
         11925 => x"72",
         11926 => x"75",
         11927 => x"76",
         11928 => x"f3",
         11929 => x"74",
         11930 => x"bd",
         11931 => x"8c",
         11932 => x"ba",
         11933 => x"2e",
         11934 => x"ba",
         11935 => x"38",
         11936 => x"51",
         11937 => x"3f",
         11938 => x"51",
         11939 => x"3f",
         11940 => x"08",
         11941 => x"30",
         11942 => x"9f",
         11943 => x"8c",
         11944 => x"57",
         11945 => x"ba",
         11946 => x"3d",
         11947 => x"77",
         11948 => x"53",
         11949 => x"3f",
         11950 => x"51",
         11951 => x"3f",
         11952 => x"08",
         11953 => x"30",
         11954 => x"9f",
         11955 => x"8c",
         11956 => x"57",
         11957 => x"75",
         11958 => x"ff",
         11959 => x"84",
         11960 => x"84",
         11961 => x"8a",
         11962 => x"81",
         11963 => x"fe",
         11964 => x"84",
         11965 => x"81",
         11966 => x"fe",
         11967 => x"75",
         11968 => x"fe",
         11969 => x"3d",
         11970 => x"80",
         11971 => x"70",
         11972 => x"52",
         11973 => x"3f",
         11974 => x"08",
         11975 => x"8c",
         11976 => x"8a",
         11977 => x"ba",
         11978 => x"3d",
         11979 => x"52",
         11980 => x"b5",
         11981 => x"ba",
         11982 => x"84",
         11983 => x"e5",
         11984 => x"cb",
         11985 => x"98",
         11986 => x"80",
         11987 => x"38",
         11988 => x"d1",
         11989 => x"75",
         11990 => x"bd",
         11991 => x"ba",
         11992 => x"3d",
         11993 => x"0b",
         11994 => x"0c",
         11995 => x"04",
         11996 => x"66",
         11997 => x"80",
         11998 => x"ec",
         11999 => x"3d",
         12000 => x"3f",
         12001 => x"08",
         12002 => x"8c",
         12003 => x"7f",
         12004 => x"08",
         12005 => x"fe",
         12006 => x"08",
         12007 => x"57",
         12008 => x"8d",
         12009 => x"0c",
         12010 => x"8c",
         12011 => x"0d",
         12012 => x"8c",
         12013 => x"5a",
         12014 => x"2e",
         12015 => x"77",
         12016 => x"84",
         12017 => x"5a",
         12018 => x"80",
         12019 => x"81",
         12020 => x"5d",
         12021 => x"08",
         12022 => x"ef",
         12023 => x"33",
         12024 => x"7c",
         12025 => x"81",
         12026 => x"b8",
         12027 => x"17",
         12028 => x"fc",
         12029 => x"ba",
         12030 => x"2e",
         12031 => x"5a",
         12032 => x"b4",
         12033 => x"7e",
         12034 => x"80",
         12035 => x"33",
         12036 => x"2e",
         12037 => x"77",
         12038 => x"83",
         12039 => x"12",
         12040 => x"2b",
         12041 => x"07",
         12042 => x"70",
         12043 => x"2b",
         12044 => x"80",
         12045 => x"80",
         12046 => x"30",
         12047 => x"63",
         12048 => x"05",
         12049 => x"62",
         12050 => x"41",
         12051 => x"52",
         12052 => x"5e",
         12053 => x"f2",
         12054 => x"0c",
         12055 => x"0c",
         12056 => x"81",
         12057 => x"84",
         12058 => x"84",
         12059 => x"95",
         12060 => x"81",
         12061 => x"08",
         12062 => x"70",
         12063 => x"33",
         12064 => x"fc",
         12065 => x"5e",
         12066 => x"08",
         12067 => x"84",
         12068 => x"83",
         12069 => x"17",
         12070 => x"08",
         12071 => x"8c",
         12072 => x"74",
         12073 => x"27",
         12074 => x"82",
         12075 => x"74",
         12076 => x"81",
         12077 => x"38",
         12078 => x"17",
         12079 => x"08",
         12080 => x"52",
         12081 => x"51",
         12082 => x"3f",
         12083 => x"97",
         12084 => x"42",
         12085 => x"56",
         12086 => x"51",
         12087 => x"3f",
         12088 => x"08",
         12089 => x"e8",
         12090 => x"8c",
         12091 => x"80",
         12092 => x"ba",
         12093 => x"70",
         12094 => x"08",
         12095 => x"7c",
         12096 => x"62",
         12097 => x"5c",
         12098 => x"76",
         12099 => x"7a",
         12100 => x"94",
         12101 => x"17",
         12102 => x"58",
         12103 => x"34",
         12104 => x"77",
         12105 => x"81",
         12106 => x"33",
         12107 => x"07",
         12108 => x"80",
         12109 => x"1d",
         12110 => x"ff",
         12111 => x"5f",
         12112 => x"55",
         12113 => x"38",
         12114 => x"77",
         12115 => x"39",
         12116 => x"5a",
         12117 => x"7a",
         12118 => x"84",
         12119 => x"07",
         12120 => x"18",
         12121 => x"39",
         12122 => x"5a",
         12123 => x"3d",
         12124 => x"89",
         12125 => x"2e",
         12126 => x"08",
         12127 => x"2e",
         12128 => x"33",
         12129 => x"2e",
         12130 => x"15",
         12131 => x"22",
         12132 => x"78",
         12133 => x"38",
         12134 => x"5a",
         12135 => x"38",
         12136 => x"56",
         12137 => x"38",
         12138 => x"70",
         12139 => x"06",
         12140 => x"55",
         12141 => x"80",
         12142 => x"17",
         12143 => x"8c",
         12144 => x"b7",
         12145 => x"d5",
         12146 => x"08",
         12147 => x"54",
         12148 => x"88",
         12149 => x"08",
         12150 => x"38",
         12151 => x"0b",
         12152 => x"94",
         12153 => x"18",
         12154 => x"c0",
         12155 => x"90",
         12156 => x"80",
         12157 => x"75",
         12158 => x"75",
         12159 => x"ba",
         12160 => x"3d",
         12161 => x"54",
         12162 => x"80",
         12163 => x"52",
         12164 => x"fe",
         12165 => x"ba",
         12166 => x"84",
         12167 => x"80",
         12168 => x"38",
         12169 => x"08",
         12170 => x"d8",
         12171 => x"8c",
         12172 => x"82",
         12173 => x"53",
         12174 => x"51",
         12175 => x"3f",
         12176 => x"08",
         12177 => x"9c",
         12178 => x"11",
         12179 => x"57",
         12180 => x"74",
         12181 => x"38",
         12182 => x"17",
         12183 => x"33",
         12184 => x"73",
         12185 => x"78",
         12186 => x"26",
         12187 => x"9c",
         12188 => x"33",
         12189 => x"e2",
         12190 => x"8c",
         12191 => x"54",
         12192 => x"38",
         12193 => x"55",
         12194 => x"39",
         12195 => x"18",
         12196 => x"73",
         12197 => x"88",
         12198 => x"c7",
         12199 => x"08",
         12200 => x"fe",
         12201 => x"84",
         12202 => x"ff",
         12203 => x"38",
         12204 => x"08",
         12205 => x"be",
         12206 => x"ae",
         12207 => x"84",
         12208 => x"9c",
         12209 => x"81",
         12210 => x"ba",
         12211 => x"18",
         12212 => x"58",
         12213 => x"0b",
         12214 => x"08",
         12215 => x"38",
         12216 => x"08",
         12217 => x"27",
         12218 => x"74",
         12219 => x"38",
         12220 => x"52",
         12221 => x"83",
         12222 => x"ba",
         12223 => x"84",
         12224 => x"80",
         12225 => x"52",
         12226 => x"fc",
         12227 => x"ba",
         12228 => x"84",
         12229 => x"80",
         12230 => x"38",
         12231 => x"08",
         12232 => x"dc",
         12233 => x"8c",
         12234 => x"80",
         12235 => x"53",
         12236 => x"51",
         12237 => x"3f",
         12238 => x"08",
         12239 => x"9c",
         12240 => x"11",
         12241 => x"57",
         12242 => x"74",
         12243 => x"81",
         12244 => x"0c",
         12245 => x"81",
         12246 => x"84",
         12247 => x"54",
         12248 => x"ff",
         12249 => x"55",
         12250 => x"17",
         12251 => x"f3",
         12252 => x"fe",
         12253 => x"0b",
         12254 => x"59",
         12255 => x"39",
         12256 => x"39",
         12257 => x"18",
         12258 => x"fe",
         12259 => x"ba",
         12260 => x"18",
         12261 => x"fd",
         12262 => x"0b",
         12263 => x"59",
         12264 => x"39",
         12265 => x"08",
         12266 => x"81",
         12267 => x"39",
         12268 => x"82",
         12269 => x"ff",
         12270 => x"a8",
         12271 => x"b7",
         12272 => x"ba",
         12273 => x"84",
         12274 => x"80",
         12275 => x"75",
         12276 => x"0c",
         12277 => x"04",
         12278 => x"3d",
         12279 => x"3d",
         12280 => x"ff",
         12281 => x"84",
         12282 => x"56",
         12283 => x"08",
         12284 => x"81",
         12285 => x"70",
         12286 => x"06",
         12287 => x"56",
         12288 => x"76",
         12289 => x"80",
         12290 => x"38",
         12291 => x"05",
         12292 => x"06",
         12293 => x"56",
         12294 => x"38",
         12295 => x"08",
         12296 => x"9a",
         12297 => x"88",
         12298 => x"33",
         12299 => x"57",
         12300 => x"2e",
         12301 => x"76",
         12302 => x"06",
         12303 => x"2e",
         12304 => x"87",
         12305 => x"08",
         12306 => x"83",
         12307 => x"7a",
         12308 => x"8c",
         12309 => x"3d",
         12310 => x"ff",
         12311 => x"84",
         12312 => x"56",
         12313 => x"08",
         12314 => x"84",
         12315 => x"52",
         12316 => x"91",
         12317 => x"ba",
         12318 => x"84",
         12319 => x"a0",
         12320 => x"84",
         12321 => x"a7",
         12322 => x"95",
         12323 => x"17",
         12324 => x"2b",
         12325 => x"07",
         12326 => x"5d",
         12327 => x"39",
         12328 => x"08",
         12329 => x"38",
         12330 => x"08",
         12331 => x"78",
         12332 => x"3d",
         12333 => x"57",
         12334 => x"80",
         12335 => x"52",
         12336 => x"8b",
         12337 => x"ba",
         12338 => x"84",
         12339 => x"80",
         12340 => x"75",
         12341 => x"07",
         12342 => x"5a",
         12343 => x"9a",
         12344 => x"2e",
         12345 => x"79",
         12346 => x"81",
         12347 => x"38",
         12348 => x"7b",
         12349 => x"38",
         12350 => x"fd",
         12351 => x"51",
         12352 => x"3f",
         12353 => x"08",
         12354 => x"0c",
         12355 => x"04",
         12356 => x"98",
         12357 => x"80",
         12358 => x"08",
         12359 => x"b9",
         12360 => x"33",
         12361 => x"74",
         12362 => x"81",
         12363 => x"38",
         12364 => x"53",
         12365 => x"81",
         12366 => x"fe",
         12367 => x"84",
         12368 => x"80",
         12369 => x"ff",
         12370 => x"75",
         12371 => x"77",
         12372 => x"38",
         12373 => x"58",
         12374 => x"81",
         12375 => x"34",
         12376 => x"7c",
         12377 => x"38",
         12378 => x"51",
         12379 => x"3f",
         12380 => x"08",
         12381 => x"8c",
         12382 => x"ff",
         12383 => x"84",
         12384 => x"06",
         12385 => x"82",
         12386 => x"39",
         12387 => x"17",
         12388 => x"52",
         12389 => x"51",
         12390 => x"3f",
         12391 => x"ba",
         12392 => x"2e",
         12393 => x"ff",
         12394 => x"ba",
         12395 => x"18",
         12396 => x"08",
         12397 => x"31",
         12398 => x"08",
         12399 => x"a0",
         12400 => x"fe",
         12401 => x"17",
         12402 => x"82",
         12403 => x"06",
         12404 => x"81",
         12405 => x"08",
         12406 => x"05",
         12407 => x"81",
         12408 => x"fe",
         12409 => x"79",
         12410 => x"39",
         12411 => x"78",
         12412 => x"38",
         12413 => x"51",
         12414 => x"3f",
         12415 => x"08",
         12416 => x"8c",
         12417 => x"80",
         12418 => x"ba",
         12419 => x"2e",
         12420 => x"84",
         12421 => x"ff",
         12422 => x"38",
         12423 => x"52",
         12424 => x"fd",
         12425 => x"ba",
         12426 => x"38",
         12427 => x"fe",
         12428 => x"08",
         12429 => x"75",
         12430 => x"b0",
         12431 => x"94",
         12432 => x"17",
         12433 => x"5c",
         12434 => x"34",
         12435 => x"7a",
         12436 => x"38",
         12437 => x"a2",
         12438 => x"fd",
         12439 => x"ba",
         12440 => x"fd",
         12441 => x"56",
         12442 => x"e3",
         12443 => x"53",
         12444 => x"bc",
         12445 => x"3d",
         12446 => x"c0",
         12447 => x"8c",
         12448 => x"ba",
         12449 => x"2e",
         12450 => x"84",
         12451 => x"9f",
         12452 => x"7d",
         12453 => x"93",
         12454 => x"5a",
         12455 => x"3f",
         12456 => x"08",
         12457 => x"8c",
         12458 => x"88",
         12459 => x"8c",
         12460 => x"0d",
         12461 => x"8c",
         12462 => x"09",
         12463 => x"38",
         12464 => x"05",
         12465 => x"2a",
         12466 => x"58",
         12467 => x"ff",
         12468 => x"5f",
         12469 => x"3d",
         12470 => x"ff",
         12471 => x"84",
         12472 => x"75",
         12473 => x"ba",
         12474 => x"38",
         12475 => x"ba",
         12476 => x"2e",
         12477 => x"84",
         12478 => x"ff",
         12479 => x"38",
         12480 => x"38",
         12481 => x"8c",
         12482 => x"33",
         12483 => x"7a",
         12484 => x"fe",
         12485 => x"08",
         12486 => x"56",
         12487 => x"79",
         12488 => x"8a",
         12489 => x"71",
         12490 => x"08",
         12491 => x"7a",
         12492 => x"b8",
         12493 => x"80",
         12494 => x"80",
         12495 => x"05",
         12496 => x"15",
         12497 => x"38",
         12498 => x"17",
         12499 => x"75",
         12500 => x"38",
         12501 => x"1b",
         12502 => x"81",
         12503 => x"fe",
         12504 => x"84",
         12505 => x"81",
         12506 => x"18",
         12507 => x"82",
         12508 => x"39",
         12509 => x"17",
         12510 => x"17",
         12511 => x"18",
         12512 => x"fe",
         12513 => x"81",
         12514 => x"8c",
         12515 => x"84",
         12516 => x"83",
         12517 => x"17",
         12518 => x"08",
         12519 => x"a0",
         12520 => x"fe",
         12521 => x"17",
         12522 => x"82",
         12523 => x"06",
         12524 => x"75",
         12525 => x"08",
         12526 => x"05",
         12527 => x"81",
         12528 => x"fe",
         12529 => x"fe",
         12530 => x"56",
         12531 => x"58",
         12532 => x"27",
         12533 => x"7b",
         12534 => x"27",
         12535 => x"74",
         12536 => x"fe",
         12537 => x"84",
         12538 => x"5a",
         12539 => x"08",
         12540 => x"96",
         12541 => x"8c",
         12542 => x"fd",
         12543 => x"ba",
         12544 => x"2e",
         12545 => x"80",
         12546 => x"76",
         12547 => x"b0",
         12548 => x"8c",
         12549 => x"38",
         12550 => x"fe",
         12551 => x"08",
         12552 => x"77",
         12553 => x"38",
         12554 => x"18",
         12555 => x"33",
         12556 => x"7b",
         12557 => x"79",
         12558 => x"26",
         12559 => x"75",
         12560 => x"0c",
         12561 => x"04",
         12562 => x"55",
         12563 => x"ff",
         12564 => x"56",
         12565 => x"09",
         12566 => x"f0",
         12567 => x"b8",
         12568 => x"a0",
         12569 => x"05",
         12570 => x"16",
         12571 => x"38",
         12572 => x"0b",
         12573 => x"7d",
         12574 => x"80",
         12575 => x"7d",
         12576 => x"ce",
         12577 => x"80",
         12578 => x"a1",
         12579 => x"1a",
         12580 => x"0b",
         12581 => x"34",
         12582 => x"ff",
         12583 => x"56",
         12584 => x"17",
         12585 => x"2a",
         12586 => x"d3",
         12587 => x"33",
         12588 => x"2e",
         12589 => x"7d",
         12590 => x"80",
         12591 => x"1b",
         12592 => x"74",
         12593 => x"56",
         12594 => x"81",
         12595 => x"ff",
         12596 => x"ef",
         12597 => x"ae",
         12598 => x"17",
         12599 => x"71",
         12600 => x"06",
         12601 => x"78",
         12602 => x"34",
         12603 => x"5b",
         12604 => x"17",
         12605 => x"55",
         12606 => x"80",
         12607 => x"5b",
         12608 => x"1c",
         12609 => x"ff",
         12610 => x"84",
         12611 => x"56",
         12612 => x"08",
         12613 => x"69",
         12614 => x"8c",
         12615 => x"34",
         12616 => x"08",
         12617 => x"a1",
         12618 => x"34",
         12619 => x"99",
         12620 => x"6a",
         12621 => x"9a",
         12622 => x"88",
         12623 => x"9b",
         12624 => x"33",
         12625 => x"2e",
         12626 => x"69",
         12627 => x"8b",
         12628 => x"57",
         12629 => x"18",
         12630 => x"fe",
         12631 => x"84",
         12632 => x"56",
         12633 => x"8c",
         12634 => x"0d",
         12635 => x"2a",
         12636 => x"ec",
         12637 => x"88",
         12638 => x"80",
         12639 => x"fe",
         12640 => x"90",
         12641 => x"80",
         12642 => x"7a",
         12643 => x"74",
         12644 => x"34",
         12645 => x"0b",
         12646 => x"b8",
         12647 => x"56",
         12648 => x"7b",
         12649 => x"77",
         12650 => x"77",
         12651 => x"7b",
         12652 => x"69",
         12653 => x"8b",
         12654 => x"57",
         12655 => x"18",
         12656 => x"fe",
         12657 => x"84",
         12658 => x"56",
         12659 => x"d1",
         12660 => x"3d",
         12661 => x"70",
         12662 => x"79",
         12663 => x"38",
         12664 => x"05",
         12665 => x"9f",
         12666 => x"75",
         12667 => x"b8",
         12668 => x"38",
         12669 => x"81",
         12670 => x"53",
         12671 => x"fc",
         12672 => x"3d",
         12673 => x"b4",
         12674 => x"8c",
         12675 => x"ba",
         12676 => x"2e",
         12677 => x"84",
         12678 => x"b1",
         12679 => x"7f",
         12680 => x"b2",
         12681 => x"a5",
         12682 => x"59",
         12683 => x"3f",
         12684 => x"08",
         12685 => x"8c",
         12686 => x"02",
         12687 => x"33",
         12688 => x"5d",
         12689 => x"ce",
         12690 => x"92",
         12691 => x"08",
         12692 => x"75",
         12693 => x"57",
         12694 => x"81",
         12695 => x"ff",
         12696 => x"ef",
         12697 => x"58",
         12698 => x"58",
         12699 => x"70",
         12700 => x"33",
         12701 => x"05",
         12702 => x"15",
         12703 => x"38",
         12704 => x"52",
         12705 => x"9e",
         12706 => x"ba",
         12707 => x"84",
         12708 => x"85",
         12709 => x"a8",
         12710 => x"81",
         12711 => x"0b",
         12712 => x"0c",
         12713 => x"04",
         12714 => x"11",
         12715 => x"06",
         12716 => x"74",
         12717 => x"38",
         12718 => x"81",
         12719 => x"05",
         12720 => x"7a",
         12721 => x"38",
         12722 => x"83",
         12723 => x"08",
         12724 => x"5f",
         12725 => x"70",
         12726 => x"33",
         12727 => x"05",
         12728 => x"9f",
         12729 => x"56",
         12730 => x"89",
         12731 => x"70",
         12732 => x"57",
         12733 => x"17",
         12734 => x"26",
         12735 => x"17",
         12736 => x"06",
         12737 => x"30",
         12738 => x"59",
         12739 => x"2e",
         12740 => x"85",
         12741 => x"be",
         12742 => x"32",
         12743 => x"72",
         12744 => x"7a",
         12745 => x"55",
         12746 => x"95",
         12747 => x"84",
         12748 => x"7b",
         12749 => x"c2",
         12750 => x"7e",
         12751 => x"96",
         12752 => x"24",
         12753 => x"79",
         12754 => x"53",
         12755 => x"fc",
         12756 => x"3d",
         12757 => x"e4",
         12758 => x"8c",
         12759 => x"ba",
         12760 => x"b2",
         12761 => x"39",
         12762 => x"08",
         12763 => x"06",
         12764 => x"77",
         12765 => x"a8",
         12766 => x"8c",
         12767 => x"ba",
         12768 => x"92",
         12769 => x"93",
         12770 => x"02",
         12771 => x"cd",
         12772 => x"5a",
         12773 => x"05",
         12774 => x"70",
         12775 => x"34",
         12776 => x"79",
         12777 => x"80",
         12778 => x"8b",
         12779 => x"18",
         12780 => x"2a",
         12781 => x"56",
         12782 => x"75",
         12783 => x"76",
         12784 => x"7f",
         12785 => x"83",
         12786 => x"18",
         12787 => x"2a",
         12788 => x"5c",
         12789 => x"81",
         12790 => x"3d",
         12791 => x"81",
         12792 => x"9b",
         12793 => x"1a",
         12794 => x"2b",
         12795 => x"41",
         12796 => x"7d",
         12797 => x"e0",
         12798 => x"9c",
         12799 => x"05",
         12800 => x"7d",
         12801 => x"38",
         12802 => x"76",
         12803 => x"19",
         12804 => x"5e",
         12805 => x"82",
         12806 => x"7a",
         12807 => x"17",
         12808 => x"aa",
         12809 => x"33",
         12810 => x"bc",
         12811 => x"75",
         12812 => x"52",
         12813 => x"51",
         12814 => x"3f",
         12815 => x"08",
         12816 => x"38",
         12817 => x"5c",
         12818 => x"0c",
         12819 => x"80",
         12820 => x"56",
         12821 => x"38",
         12822 => x"5a",
         12823 => x"09",
         12824 => x"38",
         12825 => x"ff",
         12826 => x"56",
         12827 => x"18",
         12828 => x"2a",
         12829 => x"f3",
         12830 => x"33",
         12831 => x"2e",
         12832 => x"93",
         12833 => x"2a",
         12834 => x"ec",
         12835 => x"88",
         12836 => x"80",
         12837 => x"7f",
         12838 => x"83",
         12839 => x"08",
         12840 => x"b2",
         12841 => x"5c",
         12842 => x"2e",
         12843 => x"52",
         12844 => x"fb",
         12845 => x"ba",
         12846 => x"84",
         12847 => x"80",
         12848 => x"16",
         12849 => x"08",
         12850 => x"b4",
         12851 => x"2e",
         12852 => x"16",
         12853 => x"5f",
         12854 => x"09",
         12855 => x"a8",
         12856 => x"76",
         12857 => x"52",
         12858 => x"51",
         12859 => x"3f",
         12860 => x"08",
         12861 => x"38",
         12862 => x"58",
         12863 => x"0c",
         12864 => x"aa",
         12865 => x"08",
         12866 => x"34",
         12867 => x"17",
         12868 => x"08",
         12869 => x"38",
         12870 => x"51",
         12871 => x"3f",
         12872 => x"08",
         12873 => x"8c",
         12874 => x"ff",
         12875 => x"56",
         12876 => x"f9",
         12877 => x"56",
         12878 => x"38",
         12879 => x"e5",
         12880 => x"ba",
         12881 => x"ba",
         12882 => x"3d",
         12883 => x"0b",
         12884 => x"0c",
         12885 => x"04",
         12886 => x"94",
         12887 => x"98",
         12888 => x"2b",
         12889 => x"58",
         12890 => x"8d",
         12891 => x"8c",
         12892 => x"fb",
         12893 => x"ba",
         12894 => x"2e",
         12895 => x"75",
         12896 => x"0c",
         12897 => x"04",
         12898 => x"16",
         12899 => x"52",
         12900 => x"51",
         12901 => x"3f",
         12902 => x"ba",
         12903 => x"2e",
         12904 => x"fe",
         12905 => x"ba",
         12906 => x"17",
         12907 => x"08",
         12908 => x"31",
         12909 => x"08",
         12910 => x"a0",
         12911 => x"fe",
         12912 => x"16",
         12913 => x"82",
         12914 => x"06",
         12915 => x"81",
         12916 => x"08",
         12917 => x"05",
         12918 => x"81",
         12919 => x"fe",
         12920 => x"79",
         12921 => x"39",
         12922 => x"17",
         12923 => x"17",
         12924 => x"18",
         12925 => x"fe",
         12926 => x"81",
         12927 => x"8c",
         12928 => x"38",
         12929 => x"08",
         12930 => x"b4",
         12931 => x"18",
         12932 => x"ba",
         12933 => x"55",
         12934 => x"08",
         12935 => x"38",
         12936 => x"5d",
         12937 => x"09",
         12938 => x"81",
         12939 => x"b4",
         12940 => x"18",
         12941 => x"7a",
         12942 => x"33",
         12943 => x"eb",
         12944 => x"fb",
         12945 => x"3d",
         12946 => x"df",
         12947 => x"84",
         12948 => x"05",
         12949 => x"82",
         12950 => x"cc",
         12951 => x"3d",
         12952 => x"d8",
         12953 => x"8c",
         12954 => x"ba",
         12955 => x"2e",
         12956 => x"84",
         12957 => x"96",
         12958 => x"78",
         12959 => x"96",
         12960 => x"51",
         12961 => x"3f",
         12962 => x"08",
         12963 => x"8c",
         12964 => x"02",
         12965 => x"33",
         12966 => x"54",
         12967 => x"d2",
         12968 => x"06",
         12969 => x"8b",
         12970 => x"06",
         12971 => x"07",
         12972 => x"55",
         12973 => x"34",
         12974 => x"0b",
         12975 => x"78",
         12976 => x"9a",
         12977 => x"8c",
         12978 => x"8c",
         12979 => x"0d",
         12980 => x"0d",
         12981 => x"53",
         12982 => x"05",
         12983 => x"51",
         12984 => x"3f",
         12985 => x"08",
         12986 => x"8c",
         12987 => x"8a",
         12988 => x"ba",
         12989 => x"3d",
         12990 => x"5a",
         12991 => x"3d",
         12992 => x"ff",
         12993 => x"84",
         12994 => x"55",
         12995 => x"08",
         12996 => x"80",
         12997 => x"81",
         12998 => x"86",
         12999 => x"38",
         13000 => x"22",
         13001 => x"71",
         13002 => x"59",
         13003 => x"96",
         13004 => x"88",
         13005 => x"97",
         13006 => x"90",
         13007 => x"98",
         13008 => x"98",
         13009 => x"99",
         13010 => x"57",
         13011 => x"18",
         13012 => x"fe",
         13013 => x"84",
         13014 => x"84",
         13015 => x"96",
         13016 => x"e8",
         13017 => x"6d",
         13018 => x"53",
         13019 => x"05",
         13020 => x"51",
         13021 => x"3f",
         13022 => x"08",
         13023 => x"08",
         13024 => x"ba",
         13025 => x"80",
         13026 => x"57",
         13027 => x"8b",
         13028 => x"76",
         13029 => x"78",
         13030 => x"76",
         13031 => x"07",
         13032 => x"5b",
         13033 => x"81",
         13034 => x"70",
         13035 => x"58",
         13036 => x"81",
         13037 => x"a4",
         13038 => x"56",
         13039 => x"16",
         13040 => x"82",
         13041 => x"16",
         13042 => x"55",
         13043 => x"09",
         13044 => x"98",
         13045 => x"76",
         13046 => x"52",
         13047 => x"51",
         13048 => x"3f",
         13049 => x"08",
         13050 => x"38",
         13051 => x"59",
         13052 => x"0c",
         13053 => x"bd",
         13054 => x"33",
         13055 => x"c3",
         13056 => x"2e",
         13057 => x"e4",
         13058 => x"2e",
         13059 => x"56",
         13060 => x"05",
         13061 => x"82",
         13062 => x"90",
         13063 => x"2b",
         13064 => x"33",
         13065 => x"88",
         13066 => x"71",
         13067 => x"5f",
         13068 => x"59",
         13069 => x"ba",
         13070 => x"3d",
         13071 => x"5e",
         13072 => x"52",
         13073 => x"52",
         13074 => x"8b",
         13075 => x"8c",
         13076 => x"ba",
         13077 => x"2e",
         13078 => x"76",
         13079 => x"81",
         13080 => x"38",
         13081 => x"80",
         13082 => x"39",
         13083 => x"16",
         13084 => x"16",
         13085 => x"17",
         13086 => x"fe",
         13087 => x"77",
         13088 => x"8c",
         13089 => x"09",
         13090 => x"e8",
         13091 => x"8c",
         13092 => x"34",
         13093 => x"a8",
         13094 => x"84",
         13095 => x"5a",
         13096 => x"17",
         13097 => x"ad",
         13098 => x"33",
         13099 => x"2e",
         13100 => x"fe",
         13101 => x"54",
         13102 => x"a0",
         13103 => x"53",
         13104 => x"16",
         13105 => x"db",
         13106 => x"59",
         13107 => x"53",
         13108 => x"81",
         13109 => x"fe",
         13110 => x"84",
         13111 => x"80",
         13112 => x"38",
         13113 => x"75",
         13114 => x"fe",
         13115 => x"84",
         13116 => x"57",
         13117 => x"08",
         13118 => x"84",
         13119 => x"84",
         13120 => x"66",
         13121 => x"79",
         13122 => x"7c",
         13123 => x"56",
         13124 => x"34",
         13125 => x"8a",
         13126 => x"38",
         13127 => x"57",
         13128 => x"34",
         13129 => x"fc",
         13130 => x"18",
         13131 => x"33",
         13132 => x"79",
         13133 => x"38",
         13134 => x"79",
         13135 => x"39",
         13136 => x"82",
         13137 => x"ff",
         13138 => x"a2",
         13139 => x"9c",
         13140 => x"ba",
         13141 => x"84",
         13142 => x"82",
         13143 => x"3d",
         13144 => x"57",
         13145 => x"70",
         13146 => x"34",
         13147 => x"74",
         13148 => x"a3",
         13149 => x"33",
         13150 => x"06",
         13151 => x"5a",
         13152 => x"81",
         13153 => x"3d",
         13154 => x"5c",
         13155 => x"06",
         13156 => x"55",
         13157 => x"38",
         13158 => x"74",
         13159 => x"26",
         13160 => x"74",
         13161 => x"3f",
         13162 => x"84",
         13163 => x"51",
         13164 => x"84",
         13165 => x"83",
         13166 => x"57",
         13167 => x"81",
         13168 => x"e7",
         13169 => x"e7",
         13170 => x"81",
         13171 => x"56",
         13172 => x"2e",
         13173 => x"74",
         13174 => x"2e",
         13175 => x"18",
         13176 => x"81",
         13177 => x"57",
         13178 => x"2e",
         13179 => x"77",
         13180 => x"06",
         13181 => x"81",
         13182 => x"78",
         13183 => x"81",
         13184 => x"81",
         13185 => x"89",
         13186 => x"38",
         13187 => x"27",
         13188 => x"88",
         13189 => x"7b",
         13190 => x"5d",
         13191 => x"5a",
         13192 => x"81",
         13193 => x"81",
         13194 => x"08",
         13195 => x"81",
         13196 => x"58",
         13197 => x"9f",
         13198 => x"38",
         13199 => x"57",
         13200 => x"81",
         13201 => x"38",
         13202 => x"99",
         13203 => x"05",
         13204 => x"70",
         13205 => x"7a",
         13206 => x"81",
         13207 => x"ff",
         13208 => x"ed",
         13209 => x"80",
         13210 => x"95",
         13211 => x"56",
         13212 => x"3f",
         13213 => x"08",
         13214 => x"8c",
         13215 => x"b4",
         13216 => x"75",
         13217 => x"0c",
         13218 => x"04",
         13219 => x"74",
         13220 => x"3f",
         13221 => x"08",
         13222 => x"06",
         13223 => x"f8",
         13224 => x"75",
         13225 => x"0c",
         13226 => x"04",
         13227 => x"33",
         13228 => x"39",
         13229 => x"51",
         13230 => x"3f",
         13231 => x"08",
         13232 => x"8c",
         13233 => x"38",
         13234 => x"82",
         13235 => x"6c",
         13236 => x"55",
         13237 => x"05",
         13238 => x"70",
         13239 => x"34",
         13240 => x"74",
         13241 => x"5d",
         13242 => x"1e",
         13243 => x"fe",
         13244 => x"84",
         13245 => x"55",
         13246 => x"87",
         13247 => x"27",
         13248 => x"86",
         13249 => x"39",
         13250 => x"08",
         13251 => x"81",
         13252 => x"38",
         13253 => x"75",
         13254 => x"38",
         13255 => x"53",
         13256 => x"fe",
         13257 => x"84",
         13258 => x"57",
         13259 => x"08",
         13260 => x"81",
         13261 => x"38",
         13262 => x"08",
         13263 => x"5a",
         13264 => x"57",
         13265 => x"18",
         13266 => x"b2",
         13267 => x"33",
         13268 => x"2e",
         13269 => x"81",
         13270 => x"54",
         13271 => x"18",
         13272 => x"33",
         13273 => x"c4",
         13274 => x"8c",
         13275 => x"85",
         13276 => x"81",
         13277 => x"19",
         13278 => x"78",
         13279 => x"9c",
         13280 => x"33",
         13281 => x"74",
         13282 => x"81",
         13283 => x"30",
         13284 => x"78",
         13285 => x"74",
         13286 => x"d7",
         13287 => x"5a",
         13288 => x"a5",
         13289 => x"75",
         13290 => x"a1",
         13291 => x"8c",
         13292 => x"ba",
         13293 => x"2e",
         13294 => x"87",
         13295 => x"2e",
         13296 => x"76",
         13297 => x"b9",
         13298 => x"57",
         13299 => x"70",
         13300 => x"34",
         13301 => x"74",
         13302 => x"56",
         13303 => x"17",
         13304 => x"7e",
         13305 => x"76",
         13306 => x"58",
         13307 => x"81",
         13308 => x"ff",
         13309 => x"80",
         13310 => x"38",
         13311 => x"05",
         13312 => x"70",
         13313 => x"34",
         13314 => x"74",
         13315 => x"d6",
         13316 => x"e5",
         13317 => x"5d",
         13318 => x"1e",
         13319 => x"fe",
         13320 => x"84",
         13321 => x"55",
         13322 => x"81",
         13323 => x"39",
         13324 => x"18",
         13325 => x"52",
         13326 => x"51",
         13327 => x"3f",
         13328 => x"08",
         13329 => x"81",
         13330 => x"38",
         13331 => x"08",
         13332 => x"b4",
         13333 => x"19",
         13334 => x"7b",
         13335 => x"27",
         13336 => x"18",
         13337 => x"82",
         13338 => x"84",
         13339 => x"59",
         13340 => x"74",
         13341 => x"75",
         13342 => x"d1",
         13343 => x"8c",
         13344 => x"ba",
         13345 => x"2e",
         13346 => x"fe",
         13347 => x"70",
         13348 => x"80",
         13349 => x"38",
         13350 => x"81",
         13351 => x"08",
         13352 => x"05",
         13353 => x"81",
         13354 => x"fe",
         13355 => x"fd",
         13356 => x"3d",
         13357 => x"02",
         13358 => x"cb",
         13359 => x"5b",
         13360 => x"76",
         13361 => x"38",
         13362 => x"74",
         13363 => x"38",
         13364 => x"73",
         13365 => x"38",
         13366 => x"84",
         13367 => x"59",
         13368 => x"81",
         13369 => x"54",
         13370 => x"81",
         13371 => x"17",
         13372 => x"81",
         13373 => x"80",
         13374 => x"38",
         13375 => x"81",
         13376 => x"17",
         13377 => x"2a",
         13378 => x"5d",
         13379 => x"81",
         13380 => x"8a",
         13381 => x"89",
         13382 => x"7c",
         13383 => x"59",
         13384 => x"3f",
         13385 => x"06",
         13386 => x"72",
         13387 => x"84",
         13388 => x"05",
         13389 => x"79",
         13390 => x"55",
         13391 => x"27",
         13392 => x"19",
         13393 => x"83",
         13394 => x"77",
         13395 => x"80",
         13396 => x"76",
         13397 => x"87",
         13398 => x"7f",
         13399 => x"14",
         13400 => x"83",
         13401 => x"84",
         13402 => x"81",
         13403 => x"38",
         13404 => x"08",
         13405 => x"d8",
         13406 => x"8c",
         13407 => x"38",
         13408 => x"78",
         13409 => x"38",
         13410 => x"09",
         13411 => x"38",
         13412 => x"54",
         13413 => x"8c",
         13414 => x"0d",
         13415 => x"84",
         13416 => x"90",
         13417 => x"81",
         13418 => x"fe",
         13419 => x"84",
         13420 => x"81",
         13421 => x"fe",
         13422 => x"77",
         13423 => x"fe",
         13424 => x"80",
         13425 => x"38",
         13426 => x"58",
         13427 => x"ab",
         13428 => x"54",
         13429 => x"80",
         13430 => x"53",
         13431 => x"51",
         13432 => x"3f",
         13433 => x"08",
         13434 => x"8c",
         13435 => x"38",
         13436 => x"ff",
         13437 => x"5e",
         13438 => x"7e",
         13439 => x"0c",
         13440 => x"2e",
         13441 => x"7a",
         13442 => x"79",
         13443 => x"90",
         13444 => x"c0",
         13445 => x"90",
         13446 => x"15",
         13447 => x"94",
         13448 => x"5a",
         13449 => x"fe",
         13450 => x"7d",
         13451 => x"0c",
         13452 => x"81",
         13453 => x"84",
         13454 => x"54",
         13455 => x"ff",
         13456 => x"39",
         13457 => x"59",
         13458 => x"82",
         13459 => x"39",
         13460 => x"c0",
         13461 => x"5e",
         13462 => x"84",
         13463 => x"e3",
         13464 => x"3d",
         13465 => x"08",
         13466 => x"81",
         13467 => x"44",
         13468 => x"0b",
         13469 => x"70",
         13470 => x"79",
         13471 => x"8a",
         13472 => x"81",
         13473 => x"70",
         13474 => x"56",
         13475 => x"85",
         13476 => x"ed",
         13477 => x"2e",
         13478 => x"84",
         13479 => x"56",
         13480 => x"84",
         13481 => x"10",
         13482 => x"d4",
         13483 => x"56",
         13484 => x"2e",
         13485 => x"75",
         13486 => x"84",
         13487 => x"33",
         13488 => x"12",
         13489 => x"5d",
         13490 => x"51",
         13491 => x"3f",
         13492 => x"08",
         13493 => x"70",
         13494 => x"56",
         13495 => x"84",
         13496 => x"82",
         13497 => x"40",
         13498 => x"84",
         13499 => x"3d",
         13500 => x"83",
         13501 => x"fe",
         13502 => x"84",
         13503 => x"84",
         13504 => x"55",
         13505 => x"84",
         13506 => x"82",
         13507 => x"84",
         13508 => x"15",
         13509 => x"74",
         13510 => x"7e",
         13511 => x"38",
         13512 => x"26",
         13513 => x"7e",
         13514 => x"26",
         13515 => x"ff",
         13516 => x"55",
         13517 => x"38",
         13518 => x"a6",
         13519 => x"2a",
         13520 => x"77",
         13521 => x"5b",
         13522 => x"85",
         13523 => x"30",
         13524 => x"77",
         13525 => x"91",
         13526 => x"b0",
         13527 => x"2e",
         13528 => x"81",
         13529 => x"60",
         13530 => x"fe",
         13531 => x"81",
         13532 => x"8c",
         13533 => x"38",
         13534 => x"05",
         13535 => x"fe",
         13536 => x"88",
         13537 => x"56",
         13538 => x"82",
         13539 => x"09",
         13540 => x"f8",
         13541 => x"29",
         13542 => x"b2",
         13543 => x"58",
         13544 => x"82",
         13545 => x"b6",
         13546 => x"33",
         13547 => x"71",
         13548 => x"88",
         13549 => x"14",
         13550 => x"07",
         13551 => x"33",
         13552 => x"ba",
         13553 => x"33",
         13554 => x"71",
         13555 => x"88",
         13556 => x"14",
         13557 => x"07",
         13558 => x"33",
         13559 => x"a2",
         13560 => x"a3",
         13561 => x"3d",
         13562 => x"54",
         13563 => x"41",
         13564 => x"4d",
         13565 => x"ff",
         13566 => x"90",
         13567 => x"7a",
         13568 => x"82",
         13569 => x"81",
         13570 => x"06",
         13571 => x"80",
         13572 => x"38",
         13573 => x"45",
         13574 => x"89",
         13575 => x"06",
         13576 => x"f4",
         13577 => x"70",
         13578 => x"43",
         13579 => x"83",
         13580 => x"38",
         13581 => x"78",
         13582 => x"81",
         13583 => x"b0",
         13584 => x"74",
         13585 => x"38",
         13586 => x"98",
         13587 => x"b0",
         13588 => x"82",
         13589 => x"57",
         13590 => x"80",
         13591 => x"76",
         13592 => x"38",
         13593 => x"51",
         13594 => x"3f",
         13595 => x"08",
         13596 => x"55",
         13597 => x"08",
         13598 => x"96",
         13599 => x"84",
         13600 => x"10",
         13601 => x"08",
         13602 => x"72",
         13603 => x"57",
         13604 => x"ff",
         13605 => x"5d",
         13606 => x"47",
         13607 => x"11",
         13608 => x"11",
         13609 => x"6b",
         13610 => x"58",
         13611 => x"62",
         13612 => x"b8",
         13613 => x"5d",
         13614 => x"16",
         13615 => x"56",
         13616 => x"26",
         13617 => x"78",
         13618 => x"31",
         13619 => x"68",
         13620 => x"fc",
         13621 => x"84",
         13622 => x"40",
         13623 => x"89",
         13624 => x"82",
         13625 => x"06",
         13626 => x"83",
         13627 => x"84",
         13628 => x"27",
         13629 => x"7a",
         13630 => x"77",
         13631 => x"80",
         13632 => x"ef",
         13633 => x"fe",
         13634 => x"57",
         13635 => x"8c",
         13636 => x"0d",
         13637 => x"0c",
         13638 => x"fb",
         13639 => x"0b",
         13640 => x"0c",
         13641 => x"84",
         13642 => x"04",
         13643 => x"11",
         13644 => x"06",
         13645 => x"74",
         13646 => x"38",
         13647 => x"81",
         13648 => x"05",
         13649 => x"7a",
         13650 => x"38",
         13651 => x"e5",
         13652 => x"7d",
         13653 => x"5b",
         13654 => x"05",
         13655 => x"70",
         13656 => x"33",
         13657 => x"45",
         13658 => x"99",
         13659 => x"e0",
         13660 => x"ff",
         13661 => x"ff",
         13662 => x"64",
         13663 => x"38",
         13664 => x"81",
         13665 => x"46",
         13666 => x"9f",
         13667 => x"76",
         13668 => x"81",
         13669 => x"78",
         13670 => x"75",
         13671 => x"30",
         13672 => x"9f",
         13673 => x"5d",
         13674 => x"80",
         13675 => x"38",
         13676 => x"1f",
         13677 => x"7c",
         13678 => x"38",
         13679 => x"e0",
         13680 => x"f8",
         13681 => x"52",
         13682 => x"ca",
         13683 => x"57",
         13684 => x"08",
         13685 => x"61",
         13686 => x"06",
         13687 => x"08",
         13688 => x"83",
         13689 => x"6c",
         13690 => x"7e",
         13691 => x"9c",
         13692 => x"31",
         13693 => x"39",
         13694 => x"d2",
         13695 => x"24",
         13696 => x"7b",
         13697 => x"0c",
         13698 => x"39",
         13699 => x"48",
         13700 => x"80",
         13701 => x"38",
         13702 => x"30",
         13703 => x"fc",
         13704 => x"ba",
         13705 => x"f5",
         13706 => x"7a",
         13707 => x"18",
         13708 => x"7b",
         13709 => x"38",
         13710 => x"84",
         13711 => x"9f",
         13712 => x"ba",
         13713 => x"80",
         13714 => x"2e",
         13715 => x"9f",
         13716 => x"8b",
         13717 => x"06",
         13718 => x"7a",
         13719 => x"84",
         13720 => x"55",
         13721 => x"81",
         13722 => x"ff",
         13723 => x"f4",
         13724 => x"83",
         13725 => x"57",
         13726 => x"81",
         13727 => x"76",
         13728 => x"58",
         13729 => x"55",
         13730 => x"60",
         13731 => x"74",
         13732 => x"61",
         13733 => x"77",
         13734 => x"34",
         13735 => x"ff",
         13736 => x"61",
         13737 => x"6a",
         13738 => x"7b",
         13739 => x"34",
         13740 => x"05",
         13741 => x"32",
         13742 => x"48",
         13743 => x"05",
         13744 => x"2a",
         13745 => x"68",
         13746 => x"34",
         13747 => x"83",
         13748 => x"86",
         13749 => x"83",
         13750 => x"55",
         13751 => x"05",
         13752 => x"2a",
         13753 => x"94",
         13754 => x"61",
         13755 => x"bf",
         13756 => x"34",
         13757 => x"05",
         13758 => x"9a",
         13759 => x"61",
         13760 => x"7e",
         13761 => x"34",
         13762 => x"48",
         13763 => x"05",
         13764 => x"2a",
         13765 => x"9e",
         13766 => x"98",
         13767 => x"98",
         13768 => x"98",
         13769 => x"05",
         13770 => x"2e",
         13771 => x"80",
         13772 => x"34",
         13773 => x"05",
         13774 => x"a9",
         13775 => x"cc",
         13776 => x"34",
         13777 => x"ff",
         13778 => x"61",
         13779 => x"74",
         13780 => x"6a",
         13781 => x"34",
         13782 => x"a4",
         13783 => x"61",
         13784 => x"93",
         13785 => x"83",
         13786 => x"57",
         13787 => x"81",
         13788 => x"76",
         13789 => x"58",
         13790 => x"55",
         13791 => x"60",
         13792 => x"49",
         13793 => x"34",
         13794 => x"05",
         13795 => x"6b",
         13796 => x"7e",
         13797 => x"79",
         13798 => x"8f",
         13799 => x"84",
         13800 => x"fa",
         13801 => x"17",
         13802 => x"2e",
         13803 => x"69",
         13804 => x"80",
         13805 => x"05",
         13806 => x"15",
         13807 => x"38",
         13808 => x"5b",
         13809 => x"86",
         13810 => x"ff",
         13811 => x"62",
         13812 => x"38",
         13813 => x"61",
         13814 => x"2a",
         13815 => x"74",
         13816 => x"05",
         13817 => x"90",
         13818 => x"64",
         13819 => x"46",
         13820 => x"2a",
         13821 => x"34",
         13822 => x"59",
         13823 => x"83",
         13824 => x"78",
         13825 => x"60",
         13826 => x"fe",
         13827 => x"84",
         13828 => x"85",
         13829 => x"80",
         13830 => x"80",
         13831 => x"05",
         13832 => x"15",
         13833 => x"38",
         13834 => x"7a",
         13835 => x"76",
         13836 => x"81",
         13837 => x"80",
         13838 => x"38",
         13839 => x"83",
         13840 => x"66",
         13841 => x"75",
         13842 => x"38",
         13843 => x"54",
         13844 => x"52",
         13845 => x"c4",
         13846 => x"ba",
         13847 => x"9b",
         13848 => x"76",
         13849 => x"5b",
         13850 => x"8c",
         13851 => x"2e",
         13852 => x"58",
         13853 => x"ff",
         13854 => x"84",
         13855 => x"2e",
         13856 => x"58",
         13857 => x"38",
         13858 => x"81",
         13859 => x"81",
         13860 => x"80",
         13861 => x"80",
         13862 => x"05",
         13863 => x"19",
         13864 => x"38",
         13865 => x"34",
         13866 => x"34",
         13867 => x"05",
         13868 => x"34",
         13869 => x"05",
         13870 => x"82",
         13871 => x"67",
         13872 => x"77",
         13873 => x"34",
         13874 => x"fd",
         13875 => x"1f",
         13876 => x"d1",
         13877 => x"85",
         13878 => x"ba",
         13879 => x"2a",
         13880 => x"76",
         13881 => x"34",
         13882 => x"08",
         13883 => x"34",
         13884 => x"c6",
         13885 => x"61",
         13886 => x"34",
         13887 => x"c8",
         13888 => x"ba",
         13889 => x"83",
         13890 => x"62",
         13891 => x"05",
         13892 => x"2a",
         13893 => x"83",
         13894 => x"62",
         13895 => x"77",
         13896 => x"05",
         13897 => x"2a",
         13898 => x"83",
         13899 => x"81",
         13900 => x"60",
         13901 => x"fe",
         13902 => x"81",
         13903 => x"8c",
         13904 => x"38",
         13905 => x"52",
         13906 => x"c3",
         13907 => x"57",
         13908 => x"08",
         13909 => x"84",
         13910 => x"84",
         13911 => x"9f",
         13912 => x"ba",
         13913 => x"62",
         13914 => x"39",
         13915 => x"16",
         13916 => x"c4",
         13917 => x"38",
         13918 => x"57",
         13919 => x"e7",
         13920 => x"58",
         13921 => x"9d",
         13922 => x"26",
         13923 => x"e7",
         13924 => x"10",
         13925 => x"22",
         13926 => x"74",
         13927 => x"38",
         13928 => x"ee",
         13929 => x"78",
         13930 => x"f9",
         13931 => x"8c",
         13932 => x"84",
         13933 => x"89",
         13934 => x"a0",
         13935 => x"84",
         13936 => x"fc",
         13937 => x"58",
         13938 => x"f0",
         13939 => x"f5",
         13940 => x"57",
         13941 => x"84",
         13942 => x"83",
         13943 => x"f8",
         13944 => x"f8",
         13945 => x"81",
         13946 => x"f4",
         13947 => x"57",
         13948 => x"68",
         13949 => x"63",
         13950 => x"af",
         13951 => x"f4",
         13952 => x"61",
         13953 => x"75",
         13954 => x"68",
         13955 => x"34",
         13956 => x"5b",
         13957 => x"05",
         13958 => x"2a",
         13959 => x"a3",
         13960 => x"c6",
         13961 => x"80",
         13962 => x"80",
         13963 => x"05",
         13964 => x"80",
         13965 => x"80",
         13966 => x"c6",
         13967 => x"61",
         13968 => x"7c",
         13969 => x"7b",
         13970 => x"34",
         13971 => x"59",
         13972 => x"05",
         13973 => x"2a",
         13974 => x"a7",
         13975 => x"61",
         13976 => x"80",
         13977 => x"34",
         13978 => x"05",
         13979 => x"af",
         13980 => x"61",
         13981 => x"80",
         13982 => x"34",
         13983 => x"05",
         13984 => x"b3",
         13985 => x"80",
         13986 => x"05",
         13987 => x"80",
         13988 => x"93",
         13989 => x"05",
         13990 => x"59",
         13991 => x"70",
         13992 => x"33",
         13993 => x"05",
         13994 => x"15",
         13995 => x"2e",
         13996 => x"76",
         13997 => x"58",
         13998 => x"81",
         13999 => x"ff",
         14000 => x"da",
         14001 => x"39",
         14002 => x"53",
         14003 => x"51",
         14004 => x"3f",
         14005 => x"ba",
         14006 => x"b0",
         14007 => x"29",
         14008 => x"77",
         14009 => x"05",
         14010 => x"84",
         14011 => x"53",
         14012 => x"51",
         14013 => x"3f",
         14014 => x"81",
         14015 => x"8c",
         14016 => x"0d",
         14017 => x"0c",
         14018 => x"34",
         14019 => x"6a",
         14020 => x"4c",
         14021 => x"70",
         14022 => x"34",
         14023 => x"ff",
         14024 => x"34",
         14025 => x"05",
         14026 => x"86",
         14027 => x"61",
         14028 => x"ff",
         14029 => x"34",
         14030 => x"05",
         14031 => x"8a",
         14032 => x"65",
         14033 => x"f9",
         14034 => x"54",
         14035 => x"60",
         14036 => x"fe",
         14037 => x"84",
         14038 => x"57",
         14039 => x"81",
         14040 => x"ff",
         14041 => x"f4",
         14042 => x"80",
         14043 => x"81",
         14044 => x"7b",
         14045 => x"75",
         14046 => x"57",
         14047 => x"75",
         14048 => x"57",
         14049 => x"75",
         14050 => x"61",
         14051 => x"34",
         14052 => x"83",
         14053 => x"80",
         14054 => x"e6",
         14055 => x"e1",
         14056 => x"05",
         14057 => x"05",
         14058 => x"83",
         14059 => x"7a",
         14060 => x"78",
         14061 => x"05",
         14062 => x"2a",
         14063 => x"83",
         14064 => x"7a",
         14065 => x"7f",
         14066 => x"05",
         14067 => x"83",
         14068 => x"76",
         14069 => x"05",
         14070 => x"83",
         14071 => x"76",
         14072 => x"05",
         14073 => x"69",
         14074 => x"6b",
         14075 => x"87",
         14076 => x"52",
         14077 => x"bd",
         14078 => x"54",
         14079 => x"60",
         14080 => x"fe",
         14081 => x"69",
         14082 => x"f7",
         14083 => x"3d",
         14084 => x"5b",
         14085 => x"61",
         14086 => x"57",
         14087 => x"25",
         14088 => x"3d",
         14089 => x"f8",
         14090 => x"53",
         14091 => x"51",
         14092 => x"3f",
         14093 => x"09",
         14094 => x"38",
         14095 => x"55",
         14096 => x"90",
         14097 => x"70",
         14098 => x"34",
         14099 => x"74",
         14100 => x"38",
         14101 => x"cd",
         14102 => x"34",
         14103 => x"83",
         14104 => x"74",
         14105 => x"0c",
         14106 => x"04",
         14107 => x"7b",
         14108 => x"b3",
         14109 => x"57",
         14110 => x"80",
         14111 => x"17",
         14112 => x"76",
         14113 => x"88",
         14114 => x"17",
         14115 => x"59",
         14116 => x"81",
         14117 => x"bb",
         14118 => x"74",
         14119 => x"81",
         14120 => x"0c",
         14121 => x"04",
         14122 => x"05",
         14123 => x"8c",
         14124 => x"08",
         14125 => x"d1",
         14126 => x"32",
         14127 => x"72",
         14128 => x"70",
         14129 => x"0c",
         14130 => x"1b",
         14131 => x"56",
         14132 => x"52",
         14133 => x"94",
         14134 => x"39",
         14135 => x"02",
         14136 => x"33",
         14137 => x"58",
         14138 => x"57",
         14139 => x"70",
         14140 => x"34",
         14141 => x"74",
         14142 => x"3d",
         14143 => x"77",
         14144 => x"f7",
         14145 => x"80",
         14146 => x"c0",
         14147 => x"17",
         14148 => x"59",
         14149 => x"81",
         14150 => x"bb",
         14151 => x"74",
         14152 => x"81",
         14153 => x"0c",
         14154 => x"75",
         14155 => x"9f",
         14156 => x"11",
         14157 => x"c0",
         14158 => x"08",
         14159 => x"c9",
         14160 => x"8c",
         14161 => x"7c",
         14162 => x"38",
         14163 => x"ba",
         14164 => x"3d",
         14165 => x"3d",
         14166 => x"55",
         14167 => x"05",
         14168 => x"51",
         14169 => x"3f",
         14170 => x"70",
         14171 => x"07",
         14172 => x"30",
         14173 => x"56",
         14174 => x"8d",
         14175 => x"fd",
         14176 => x"81",
         14177 => x"ba",
         14178 => x"3d",
         14179 => x"3d",
         14180 => x"84",
         14181 => x"22",
         14182 => x"52",
         14183 => x"26",
         14184 => x"83",
         14185 => x"52",
         14186 => x"8c",
         14187 => x"0d",
         14188 => x"ff",
         14189 => x"70",
         14190 => x"09",
         14191 => x"38",
         14192 => x"e4",
         14193 => x"d0",
         14194 => x"71",
         14195 => x"81",
         14196 => x"ff",
         14197 => x"54",
         14198 => x"26",
         14199 => x"10",
         14200 => x"05",
         14201 => x"51",
         14202 => x"80",
         14203 => x"ff",
         14204 => x"8c",
         14205 => x"3d",
         14206 => x"3d",
         14207 => x"05",
         14208 => x"05",
         14209 => x"53",
         14210 => x"70",
         14211 => x"8c",
         14212 => x"72",
         14213 => x"0c",
         14214 => x"04",
         14215 => x"2e",
         14216 => x"ef",
         14217 => x"ff",
         14218 => x"70",
         14219 => x"d0",
         14220 => x"84",
         14221 => x"51",
         14222 => x"04",
         14223 => x"77",
         14224 => x"ff",
         14225 => x"e1",
         14226 => x"ff",
         14227 => x"e9",
         14228 => x"75",
         14229 => x"80",
         14230 => x"70",
         14231 => x"22",
         14232 => x"70",
         14233 => x"7a",
         14234 => x"56",
         14235 => x"b7",
         14236 => x"82",
         14237 => x"72",
         14238 => x"54",
         14239 => x"06",
         14240 => x"54",
         14241 => x"b1",
         14242 => x"38",
         14243 => x"70",
         14244 => x"52",
         14245 => x"30",
         14246 => x"75",
         14247 => x"53",
         14248 => x"80",
         14249 => x"75",
         14250 => x"ba",
         14251 => x"3d",
         14252 => x"ed",
         14253 => x"a2",
         14254 => x"26",
         14255 => x"10",
         14256 => x"a8",
         14257 => x"08",
         14258 => x"16",
         14259 => x"ff",
         14260 => x"75",
         14261 => x"ff",
         14262 => x"83",
         14263 => x"57",
         14264 => x"88",
         14265 => x"ff",
         14266 => x"51",
         14267 => x"16",
         14268 => x"ff",
         14269 => x"db",
         14270 => x"70",
         14271 => x"06",
         14272 => x"39",
         14273 => x"83",
         14274 => x"57",
         14275 => x"f0",
         14276 => x"ff",
         14277 => x"51",
         14278 => x"75",
         14279 => x"06",
         14280 => x"70",
         14281 => x"06",
         14282 => x"ff",
         14283 => x"73",
         14284 => x"05",
         14285 => x"52",
         14286 => x"00",
         14287 => x"ff",
         14288 => x"ff",
         14289 => x"ff",
         14290 => x"00",
         14291 => x"8b",
         14292 => x"80",
         14293 => x"75",
         14294 => x"6a",
         14295 => x"5f",
         14296 => x"54",
         14297 => x"49",
         14298 => x"3e",
         14299 => x"33",
         14300 => x"28",
         14301 => x"1d",
         14302 => x"12",
         14303 => x"07",
         14304 => x"fc",
         14305 => x"f1",
         14306 => x"e6",
         14307 => x"db",
         14308 => x"d0",
         14309 => x"c5",
         14310 => x"ba",
         14311 => x"bf",
         14312 => x"59",
         14313 => x"59",
         14314 => x"59",
         14315 => x"59",
         14316 => x"59",
         14317 => x"59",
         14318 => x"59",
         14319 => x"59",
         14320 => x"59",
         14321 => x"59",
         14322 => x"59",
         14323 => x"59",
         14324 => x"59",
         14325 => x"59",
         14326 => x"59",
         14327 => x"59",
         14328 => x"59",
         14329 => x"59",
         14330 => x"59",
         14331 => x"59",
         14332 => x"59",
         14333 => x"59",
         14334 => x"59",
         14335 => x"59",
         14336 => x"59",
         14337 => x"59",
         14338 => x"59",
         14339 => x"59",
         14340 => x"59",
         14341 => x"59",
         14342 => x"59",
         14343 => x"59",
         14344 => x"59",
         14345 => x"59",
         14346 => x"59",
         14347 => x"59",
         14348 => x"59",
         14349 => x"59",
         14350 => x"59",
         14351 => x"59",
         14352 => x"59",
         14353 => x"59",
         14354 => x"7b",
         14355 => x"59",
         14356 => x"59",
         14357 => x"59",
         14358 => x"59",
         14359 => x"59",
         14360 => x"59",
         14361 => x"59",
         14362 => x"59",
         14363 => x"59",
         14364 => x"59",
         14365 => x"59",
         14366 => x"59",
         14367 => x"59",
         14368 => x"59",
         14369 => x"59",
         14370 => x"59",
         14371 => x"11",
         14372 => x"10",
         14373 => x"59",
         14374 => x"94",
         14375 => x"b2",
         14376 => x"71",
         14377 => x"36",
         14378 => x"d8",
         14379 => x"59",
         14380 => x"59",
         14381 => x"59",
         14382 => x"59",
         14383 => x"59",
         14384 => x"59",
         14385 => x"59",
         14386 => x"59",
         14387 => x"59",
         14388 => x"59",
         14389 => x"59",
         14390 => x"59",
         14391 => x"59",
         14392 => x"59",
         14393 => x"59",
         14394 => x"59",
         14395 => x"59",
         14396 => x"59",
         14397 => x"59",
         14398 => x"59",
         14399 => x"59",
         14400 => x"59",
         14401 => x"59",
         14402 => x"59",
         14403 => x"59",
         14404 => x"59",
         14405 => x"59",
         14406 => x"59",
         14407 => x"59",
         14408 => x"59",
         14409 => x"59",
         14410 => x"59",
         14411 => x"59",
         14412 => x"59",
         14413 => x"59",
         14414 => x"59",
         14415 => x"59",
         14416 => x"59",
         14417 => x"59",
         14418 => x"59",
         14419 => x"59",
         14420 => x"59",
         14421 => x"59",
         14422 => x"59",
         14423 => x"59",
         14424 => x"59",
         14425 => x"59",
         14426 => x"59",
         14427 => x"59",
         14428 => x"59",
         14429 => x"59",
         14430 => x"59",
         14431 => x"b5",
         14432 => x"7a",
         14433 => x"59",
         14434 => x"59",
         14435 => x"59",
         14436 => x"59",
         14437 => x"59",
         14438 => x"59",
         14439 => x"59",
         14440 => x"59",
         14441 => x"6d",
         14442 => x"62",
         14443 => x"59",
         14444 => x"4b",
         14445 => x"59",
         14446 => x"5b",
         14447 => x"51",
         14448 => x"44",
         14449 => x"1c",
         14450 => x"34",
         14451 => x"40",
         14452 => x"4c",
         14453 => x"58",
         14454 => x"28",
         14455 => x"91",
         14456 => x"7f",
         14457 => x"fb",
         14458 => x"49",
         14459 => x"1b",
         14460 => x"d8",
         14461 => x"95",
         14462 => x"6e",
         14463 => x"c5",
         14464 => x"9d",
         14465 => x"0c",
         14466 => x"24",
         14467 => x"d8",
         14468 => x"fb",
         14469 => x"05",
         14470 => x"95",
         14471 => x"d8",
         14472 => x"d8",
         14473 => x"0c",
         14474 => x"9d",
         14475 => x"6e",
         14476 => x"49",
         14477 => x"76",
         14478 => x"8f",
         14479 => x"b4",
         14480 => x"d5",
         14481 => x"36",
         14482 => x"fa",
         14483 => x"4f",
         14484 => x"9f",
         14485 => x"5c",
         14486 => x"5c",
         14487 => x"5c",
         14488 => x"5c",
         14489 => x"5c",
         14490 => x"5c",
         14491 => x"35",
         14492 => x"5c",
         14493 => x"5c",
         14494 => x"5c",
         14495 => x"5c",
         14496 => x"5c",
         14497 => x"5c",
         14498 => x"5c",
         14499 => x"5c",
         14500 => x"5c",
         14501 => x"5c",
         14502 => x"5c",
         14503 => x"5c",
         14504 => x"5c",
         14505 => x"5c",
         14506 => x"5c",
         14507 => x"5c",
         14508 => x"5c",
         14509 => x"5c",
         14510 => x"5c",
         14511 => x"5c",
         14512 => x"5c",
         14513 => x"5c",
         14514 => x"74",
         14515 => x"62",
         14516 => x"4f",
         14517 => x"3c",
         14518 => x"66",
         14519 => x"2a",
         14520 => x"17",
         14521 => x"7f",
         14522 => x"5c",
         14523 => x"7f",
         14524 => x"07",
         14525 => x"84",
         14526 => x"b0",
         14527 => x"8e",
         14528 => x"f5",
         14529 => x"e3",
         14530 => x"d1",
         14531 => x"c2",
         14532 => x"5c",
         14533 => x"66",
         14534 => x"02",
         14535 => x"71",
         14536 => x"43",
         14537 => x"9a",
         14538 => x"77",
         14539 => x"56",
         14540 => x"2c",
         14541 => x"fc",
         14542 => x"83",
         14543 => x"d6",
         14544 => x"c5",
         14545 => x"83",
         14546 => x"83",
         14547 => x"83",
         14548 => x"83",
         14549 => x"83",
         14550 => x"83",
         14551 => x"9f",
         14552 => x"ad",
         14553 => x"64",
         14554 => x"83",
         14555 => x"83",
         14556 => x"83",
         14557 => x"83",
         14558 => x"83",
         14559 => x"83",
         14560 => x"83",
         14561 => x"83",
         14562 => x"83",
         14563 => x"83",
         14564 => x"83",
         14565 => x"83",
         14566 => x"83",
         14567 => x"83",
         14568 => x"83",
         14569 => x"83",
         14570 => x"83",
         14571 => x"83",
         14572 => x"83",
         14573 => x"21",
         14574 => x"83",
         14575 => x"83",
         14576 => x"83",
         14577 => x"c4",
         14578 => x"d3",
         14579 => x"75",
         14580 => x"83",
         14581 => x"83",
         14582 => x"83",
         14583 => x"83",
         14584 => x"5a",
         14585 => x"83",
         14586 => x"3d",
         14587 => x"a6",
         14588 => x"1b",
         14589 => x"1b",
         14590 => x"1b",
         14591 => x"1b",
         14592 => x"1b",
         14593 => x"1b",
         14594 => x"f6",
         14595 => x"1b",
         14596 => x"1b",
         14597 => x"1b",
         14598 => x"1b",
         14599 => x"1b",
         14600 => x"1b",
         14601 => x"1b",
         14602 => x"1b",
         14603 => x"1b",
         14604 => x"1b",
         14605 => x"1b",
         14606 => x"1b",
         14607 => x"1b",
         14608 => x"1b",
         14609 => x"1b",
         14610 => x"1b",
         14611 => x"1b",
         14612 => x"1b",
         14613 => x"1b",
         14614 => x"1b",
         14615 => x"1b",
         14616 => x"1b",
         14617 => x"b8",
         14618 => x"00",
         14619 => x"ed",
         14620 => x"da",
         14621 => x"c8",
         14622 => x"8b",
         14623 => x"78",
         14624 => x"68",
         14625 => x"1b",
         14626 => x"58",
         14627 => x"48",
         14628 => x"36",
         14629 => x"24",
         14630 => x"12",
         14631 => x"83",
         14632 => x"72",
         14633 => x"61",
         14634 => x"4a",
         14635 => x"1b",
         14636 => x"94",
         14637 => x"75",
         14638 => x"d1",
         14639 => x"d1",
         14640 => x"d1",
         14641 => x"d1",
         14642 => x"d1",
         14643 => x"d1",
         14644 => x"d1",
         14645 => x"d1",
         14646 => x"d1",
         14647 => x"d1",
         14648 => x"d1",
         14649 => x"d1",
         14650 => x"d1",
         14651 => x"f3",
         14652 => x"d1",
         14653 => x"d1",
         14654 => x"d1",
         14655 => x"d1",
         14656 => x"d1",
         14657 => x"d1",
         14658 => x"bf",
         14659 => x"d1",
         14660 => x"d1",
         14661 => x"4a",
         14662 => x"d1",
         14663 => x"61",
         14664 => x"d2",
         14665 => x"33",
         14666 => x"2e",
         14667 => x"1b",
         14668 => x"0f",
         14669 => x"04",
         14670 => x"f9",
         14671 => x"ee",
         14672 => x"e3",
         14673 => x"d7",
         14674 => x"c9",
         14675 => x"01",
         14676 => x"fd",
         14677 => x"fd",
         14678 => x"49",
         14679 => x"fd",
         14680 => x"fd",
         14681 => x"fd",
         14682 => x"fd",
         14683 => x"fd",
         14684 => x"fd",
         14685 => x"fd",
         14686 => x"fd",
         14687 => x"fd",
         14688 => x"7f",
         14689 => x"0d",
         14690 => x"fd",
         14691 => x"fd",
         14692 => x"fd",
         14693 => x"fd",
         14694 => x"fd",
         14695 => x"fd",
         14696 => x"fd",
         14697 => x"fd",
         14698 => x"fd",
         14699 => x"fd",
         14700 => x"fd",
         14701 => x"fd",
         14702 => x"fd",
         14703 => x"fd",
         14704 => x"fd",
         14705 => x"fd",
         14706 => x"fd",
         14707 => x"fd",
         14708 => x"fd",
         14709 => x"fd",
         14710 => x"fd",
         14711 => x"fd",
         14712 => x"fd",
         14713 => x"fd",
         14714 => x"fd",
         14715 => x"fd",
         14716 => x"fd",
         14717 => x"fd",
         14718 => x"fd",
         14719 => x"fd",
         14720 => x"fd",
         14721 => x"fd",
         14722 => x"fd",
         14723 => x"fd",
         14724 => x"fd",
         14725 => x"fd",
         14726 => x"1d",
         14727 => x"fd",
         14728 => x"fd",
         14729 => x"fd",
         14730 => x"fd",
         14731 => x"17",
         14732 => x"fd",
         14733 => x"fd",
         14734 => x"fd",
         14735 => x"fd",
         14736 => x"fd",
         14737 => x"fd",
         14738 => x"fd",
         14739 => x"fd",
         14740 => x"fd",
         14741 => x"fd",
         14742 => x"2b",
         14743 => x"e1",
         14744 => x"b8",
         14745 => x"b8",
         14746 => x"b8",
         14747 => x"fd",
         14748 => x"e1",
         14749 => x"fd",
         14750 => x"fd",
         14751 => x"ff",
         14752 => x"fd",
         14753 => x"fd",
         14754 => x"16",
         14755 => x"0f",
         14756 => x"fd",
         14757 => x"fd",
         14758 => x"58",
         14759 => x"fd",
         14760 => x"18",
         14761 => x"fd",
         14762 => x"fd",
         14763 => x"17",
         14764 => x"69",
         14765 => x"00",
         14766 => x"63",
         14767 => x"00",
         14768 => x"69",
         14769 => x"00",
         14770 => x"61",
         14771 => x"00",
         14772 => x"65",
         14773 => x"00",
         14774 => x"65",
         14775 => x"00",
         14776 => x"70",
         14777 => x"00",
         14778 => x"66",
         14779 => x"00",
         14780 => x"6d",
         14781 => x"00",
         14782 => x"00",
         14783 => x"00",
         14784 => x"00",
         14785 => x"00",
         14786 => x"00",
         14787 => x"00",
         14788 => x"00",
         14789 => x"6c",
         14790 => x"00",
         14791 => x"00",
         14792 => x"74",
         14793 => x"00",
         14794 => x"65",
         14795 => x"00",
         14796 => x"6f",
         14797 => x"00",
         14798 => x"74",
         14799 => x"00",
         14800 => x"00",
         14801 => x"00",
         14802 => x"73",
         14803 => x"00",
         14804 => x"73",
         14805 => x"00",
         14806 => x"6f",
         14807 => x"00",
         14808 => x"00",
         14809 => x"6e",
         14810 => x"20",
         14811 => x"6f",
         14812 => x"00",
         14813 => x"61",
         14814 => x"65",
         14815 => x"69",
         14816 => x"72",
         14817 => x"74",
         14818 => x"00",
         14819 => x"20",
         14820 => x"79",
         14821 => x"65",
         14822 => x"69",
         14823 => x"2e",
         14824 => x"00",
         14825 => x"75",
         14826 => x"63",
         14827 => x"74",
         14828 => x"6d",
         14829 => x"2e",
         14830 => x"00",
         14831 => x"65",
         14832 => x"20",
         14833 => x"6b",
         14834 => x"00",
         14835 => x"65",
         14836 => x"2c",
         14837 => x"65",
         14838 => x"69",
         14839 => x"63",
         14840 => x"65",
         14841 => x"64",
         14842 => x"00",
         14843 => x"6d",
         14844 => x"61",
         14845 => x"74",
         14846 => x"00",
         14847 => x"63",
         14848 => x"61",
         14849 => x"6c",
         14850 => x"69",
         14851 => x"79",
         14852 => x"6d",
         14853 => x"75",
         14854 => x"6f",
         14855 => x"69",
         14856 => x"00",
         14857 => x"6b",
         14858 => x"74",
         14859 => x"61",
         14860 => x"64",
         14861 => x"00",
         14862 => x"76",
         14863 => x"75",
         14864 => x"72",
         14865 => x"20",
         14866 => x"61",
         14867 => x"2e",
         14868 => x"00",
         14869 => x"69",
         14870 => x"72",
         14871 => x"20",
         14872 => x"74",
         14873 => x"65",
         14874 => x"00",
         14875 => x"65",
         14876 => x"6e",
         14877 => x"20",
         14878 => x"61",
         14879 => x"2e",
         14880 => x"00",
         14881 => x"65",
         14882 => x"72",
         14883 => x"79",
         14884 => x"69",
         14885 => x"2e",
         14886 => x"00",
         14887 => x"65",
         14888 => x"64",
         14889 => x"65",
         14890 => x"00",
         14891 => x"61",
         14892 => x"20",
         14893 => x"65",
         14894 => x"65",
         14895 => x"00",
         14896 => x"70",
         14897 => x"20",
         14898 => x"6e",
         14899 => x"00",
         14900 => x"66",
         14901 => x"20",
         14902 => x"6e",
         14903 => x"00",
         14904 => x"6b",
         14905 => x"74",
         14906 => x"61",
         14907 => x"00",
         14908 => x"65",
         14909 => x"6c",
         14910 => x"72",
         14911 => x"00",
         14912 => x"6b",
         14913 => x"72",
         14914 => x"00",
         14915 => x"63",
         14916 => x"2e",
         14917 => x"00",
         14918 => x"75",
         14919 => x"74",
         14920 => x"25",
         14921 => x"74",
         14922 => x"75",
         14923 => x"74",
         14924 => x"73",
         14925 => x"0a",
         14926 => x"00",
         14927 => x"64",
         14928 => x"00",
         14929 => x"6c",
         14930 => x"00",
         14931 => x"00",
         14932 => x"58",
         14933 => x"00",
         14934 => x"00",
         14935 => x"00",
         14936 => x"00",
         14937 => x"58",
         14938 => x"00",
         14939 => x"20",
         14940 => x"20",
         14941 => x"00",
         14942 => x"00",
         14943 => x"25",
         14944 => x"00",
         14945 => x"31",
         14946 => x"30",
         14947 => x"00",
         14948 => x"31",
         14949 => x"00",
         14950 => x"55",
         14951 => x"65",
         14952 => x"30",
         14953 => x"20",
         14954 => x"25",
         14955 => x"2a",
         14956 => x"00",
         14957 => x"20",
         14958 => x"65",
         14959 => x"70",
         14960 => x"61",
         14961 => x"65",
         14962 => x"00",
         14963 => x"54",
         14964 => x"58",
         14965 => x"74",
         14966 => x"75",
         14967 => x"00",
         14968 => x"54",
         14969 => x"58",
         14970 => x"74",
         14971 => x"75",
         14972 => x"00",
         14973 => x"54",
         14974 => x"58",
         14975 => x"74",
         14976 => x"75",
         14977 => x"00",
         14978 => x"54",
         14979 => x"58",
         14980 => x"74",
         14981 => x"75",
         14982 => x"00",
         14983 => x"54",
         14984 => x"52",
         14985 => x"74",
         14986 => x"75",
         14987 => x"00",
         14988 => x"54",
         14989 => x"44",
         14990 => x"74",
         14991 => x"75",
         14992 => x"00",
         14993 => x"20",
         14994 => x"65",
         14995 => x"70",
         14996 => x"00",
         14997 => x"65",
         14998 => x"6e",
         14999 => x"72",
         15000 => x"00",
         15001 => x"74",
         15002 => x"20",
         15003 => x"74",
         15004 => x"72",
         15005 => x"00",
         15006 => x"62",
         15007 => x"67",
         15008 => x"6d",
         15009 => x"2e",
         15010 => x"00",
         15011 => x"6f",
         15012 => x"63",
         15013 => x"74",
         15014 => x"00",
         15015 => x"5f",
         15016 => x"2e",
         15017 => x"00",
         15018 => x"6c",
         15019 => x"74",
         15020 => x"6e",
         15021 => x"61",
         15022 => x"65",
         15023 => x"20",
         15024 => x"64",
         15025 => x"20",
         15026 => x"61",
         15027 => x"69",
         15028 => x"20",
         15029 => x"75",
         15030 => x"79",
         15031 => x"00",
         15032 => x"00",
         15033 => x"5c",
         15034 => x"00",
         15035 => x"6b",
         15036 => x"69",
         15037 => x"6c",
         15038 => x"64",
         15039 => x"00",
         15040 => x"00",
         15041 => x"20",
         15042 => x"6d",
         15043 => x"2e",
         15044 => x"00",
         15045 => x"00",
         15046 => x"00",
         15047 => x"5c",
         15048 => x"25",
         15049 => x"73",
         15050 => x"00",
         15051 => x"64",
         15052 => x"62",
         15053 => x"69",
         15054 => x"2e",
         15055 => x"00",
         15056 => x"74",
         15057 => x"69",
         15058 => x"61",
         15059 => x"69",
         15060 => x"69",
         15061 => x"2e",
         15062 => x"00",
         15063 => x"6c",
         15064 => x"20",
         15065 => x"65",
         15066 => x"25",
         15067 => x"78",
         15068 => x"2e",
         15069 => x"00",
         15070 => x"6c",
         15071 => x"74",
         15072 => x"65",
         15073 => x"6f",
         15074 => x"28",
         15075 => x"2e",
         15076 => x"00",
         15077 => x"63",
         15078 => x"6e",
         15079 => x"6f",
         15080 => x"40",
         15081 => x"38",
         15082 => x"2e",
         15083 => x"00",
         15084 => x"6c",
         15085 => x"30",
         15086 => x"2d",
         15087 => x"00",
         15088 => x"6c",
         15089 => x"30",
         15090 => x"00",
         15091 => x"70",
         15092 => x"6e",
         15093 => x"2e",
         15094 => x"00",
         15095 => x"6c",
         15096 => x"30",
         15097 => x"2d",
         15098 => x"38",
         15099 => x"25",
         15100 => x"29",
         15101 => x"00",
         15102 => x"79",
         15103 => x"2e",
         15104 => x"00",
         15105 => x"6c",
         15106 => x"30",
         15107 => x"00",
         15108 => x"61",
         15109 => x"67",
         15110 => x"2e",
         15111 => x"00",
         15112 => x"70",
         15113 => x"6d",
         15114 => x"00",
         15115 => x"6d",
         15116 => x"74",
         15117 => x"00",
         15118 => x"5c",
         15119 => x"25",
         15120 => x"00",
         15121 => x"6f",
         15122 => x"65",
         15123 => x"75",
         15124 => x"64",
         15125 => x"61",
         15126 => x"74",
         15127 => x"6f",
         15128 => x"73",
         15129 => x"6d",
         15130 => x"64",
         15131 => x"00",
         15132 => x"00",
         15133 => x"25",
         15134 => x"64",
         15135 => x"3a",
         15136 => x"25",
         15137 => x"64",
         15138 => x"00",
         15139 => x"20",
         15140 => x"66",
         15141 => x"72",
         15142 => x"6f",
         15143 => x"00",
         15144 => x"65",
         15145 => x"65",
         15146 => x"6d",
         15147 => x"6d",
         15148 => x"65",
         15149 => x"00",
         15150 => x"72",
         15151 => x"65",
         15152 => x"00",
         15153 => x"20",
         15154 => x"20",
         15155 => x"65",
         15156 => x"65",
         15157 => x"72",
         15158 => x"64",
         15159 => x"73",
         15160 => x"25",
         15161 => x"0a",
         15162 => x"00",
         15163 => x"20",
         15164 => x"20",
         15165 => x"6f",
         15166 => x"53",
         15167 => x"74",
         15168 => x"64",
         15169 => x"73",
         15170 => x"25",
         15171 => x"0a",
         15172 => x"00",
         15173 => x"20",
         15174 => x"63",
         15175 => x"74",
         15176 => x"20",
         15177 => x"72",
         15178 => x"20",
         15179 => x"20",
         15180 => x"25",
         15181 => x"0a",
         15182 => x"00",
         15183 => x"63",
         15184 => x"00",
         15185 => x"20",
         15186 => x"20",
         15187 => x"20",
         15188 => x"20",
         15189 => x"20",
         15190 => x"20",
         15191 => x"20",
         15192 => x"25",
         15193 => x"0a",
         15194 => x"00",
         15195 => x"20",
         15196 => x"74",
         15197 => x"43",
         15198 => x"6b",
         15199 => x"65",
         15200 => x"20",
         15201 => x"20",
         15202 => x"25",
         15203 => x"30",
         15204 => x"48",
         15205 => x"00",
         15206 => x"20",
         15207 => x"68",
         15208 => x"65",
         15209 => x"52",
         15210 => x"43",
         15211 => x"6b",
         15212 => x"65",
         15213 => x"25",
         15214 => x"30",
         15215 => x"48",
         15216 => x"00",
         15217 => x"20",
         15218 => x"41",
         15219 => x"6c",
         15220 => x"20",
         15221 => x"71",
         15222 => x"20",
         15223 => x"20",
         15224 => x"25",
         15225 => x"30",
         15226 => x"48",
         15227 => x"00",
         15228 => x"20",
         15229 => x"00",
         15230 => x"20",
         15231 => x"00",
         15232 => x"20",
         15233 => x"54",
         15234 => x"00",
         15235 => x"20",
         15236 => x"49",
         15237 => x"00",
         15238 => x"20",
         15239 => x"48",
         15240 => x"45",
         15241 => x"53",
         15242 => x"00",
         15243 => x"20",
         15244 => x"52",
         15245 => x"52",
         15246 => x"43",
         15247 => x"6e",
         15248 => x"3d",
         15249 => x"64",
         15250 => x"00",
         15251 => x"20",
         15252 => x"45",
         15253 => x"20",
         15254 => x"54",
         15255 => x"72",
         15256 => x"3d",
         15257 => x"64",
         15258 => x"00",
         15259 => x"20",
         15260 => x"43",
         15261 => x"20",
         15262 => x"44",
         15263 => x"63",
         15264 => x"3d",
         15265 => x"64",
         15266 => x"00",
         15267 => x"20",
         15268 => x"20",
         15269 => x"20",
         15270 => x"25",
         15271 => x"3a",
         15272 => x"58",
         15273 => x"00",
         15274 => x"20",
         15275 => x"4d",
         15276 => x"20",
         15277 => x"25",
         15278 => x"3a",
         15279 => x"58",
         15280 => x"00",
         15281 => x"20",
         15282 => x"4e",
         15283 => x"41",
         15284 => x"25",
         15285 => x"3a",
         15286 => x"58",
         15287 => x"00",
         15288 => x"20",
         15289 => x"41",
         15290 => x"20",
         15291 => x"25",
         15292 => x"3a",
         15293 => x"58",
         15294 => x"00",
         15295 => x"20",
         15296 => x"53",
         15297 => x"4d",
         15298 => x"25",
         15299 => x"3a",
         15300 => x"58",
         15301 => x"00",
         15302 => x"72",
         15303 => x"53",
         15304 => x"63",
         15305 => x"69",
         15306 => x"00",
         15307 => x"6e",
         15308 => x"00",
         15309 => x"6d",
         15310 => x"00",
         15311 => x"6c",
         15312 => x"00",
         15313 => x"69",
         15314 => x"00",
         15315 => x"78",
         15316 => x"00",
         15317 => x"00",
         15318 => x"b4",
         15319 => x"00",
         15320 => x"02",
         15321 => x"b0",
         15322 => x"00",
         15323 => x"03",
         15324 => x"ac",
         15325 => x"00",
         15326 => x"04",
         15327 => x"a8",
         15328 => x"00",
         15329 => x"05",
         15330 => x"a4",
         15331 => x"00",
         15332 => x"06",
         15333 => x"a0",
         15334 => x"00",
         15335 => x"07",
         15336 => x"9c",
         15337 => x"00",
         15338 => x"01",
         15339 => x"98",
         15340 => x"00",
         15341 => x"08",
         15342 => x"94",
         15343 => x"00",
         15344 => x"0b",
         15345 => x"90",
         15346 => x"00",
         15347 => x"09",
         15348 => x"8c",
         15349 => x"00",
         15350 => x"0a",
         15351 => x"88",
         15352 => x"00",
         15353 => x"0d",
         15354 => x"84",
         15355 => x"00",
         15356 => x"0c",
         15357 => x"80",
         15358 => x"00",
         15359 => x"0e",
         15360 => x"7c",
         15361 => x"00",
         15362 => x"0f",
         15363 => x"78",
         15364 => x"00",
         15365 => x"0f",
         15366 => x"74",
         15367 => x"00",
         15368 => x"10",
         15369 => x"70",
         15370 => x"00",
         15371 => x"11",
         15372 => x"6c",
         15373 => x"00",
         15374 => x"12",
         15375 => x"68",
         15376 => x"00",
         15377 => x"13",
         15378 => x"64",
         15379 => x"00",
         15380 => x"14",
         15381 => x"60",
         15382 => x"00",
         15383 => x"15",
         15384 => x"00",
         15385 => x"00",
         15386 => x"00",
         15387 => x"00",
         15388 => x"7e",
         15389 => x"7e",
         15390 => x"7e",
         15391 => x"00",
         15392 => x"7e",
         15393 => x"7e",
         15394 => x"7e",
         15395 => x"00",
         15396 => x"00",
         15397 => x"00",
         15398 => x"00",
         15399 => x"00",
         15400 => x"00",
         15401 => x"00",
         15402 => x"00",
         15403 => x"00",
         15404 => x"00",
         15405 => x"00",
         15406 => x"6e",
         15407 => x"6f",
         15408 => x"2f",
         15409 => x"61",
         15410 => x"68",
         15411 => x"6f",
         15412 => x"66",
         15413 => x"2c",
         15414 => x"73",
         15415 => x"69",
         15416 => x"00",
         15417 => x"74",
         15418 => x"00",
         15419 => x"74",
         15420 => x"00",
         15421 => x"00",
         15422 => x"6c",
         15423 => x"25",
         15424 => x"00",
         15425 => x"6c",
         15426 => x"74",
         15427 => x"65",
         15428 => x"20",
         15429 => x"20",
         15430 => x"74",
         15431 => x"20",
         15432 => x"65",
         15433 => x"20",
         15434 => x"2e",
         15435 => x"00",
         15436 => x"0a",
         15437 => x"00",
         15438 => x"7e",
         15439 => x"00",
         15440 => x"00",
         15441 => x"00",
         15442 => x"00",
         15443 => x"00",
         15444 => x"30",
         15445 => x"00",
         15446 => x"31",
         15447 => x"00",
         15448 => x"32",
         15449 => x"00",
         15450 => x"33",
         15451 => x"00",
         15452 => x"34",
         15453 => x"00",
         15454 => x"35",
         15455 => x"00",
         15456 => x"37",
         15457 => x"00",
         15458 => x"38",
         15459 => x"00",
         15460 => x"39",
         15461 => x"00",
         15462 => x"30",
         15463 => x"00",
         15464 => x"7e",
         15465 => x"00",
         15466 => x"7e",
         15467 => x"00",
         15468 => x"00",
         15469 => x"7e",
         15470 => x"00",
         15471 => x"7e",
         15472 => x"00",
         15473 => x"64",
         15474 => x"2c",
         15475 => x"25",
         15476 => x"64",
         15477 => x"3a",
         15478 => x"78",
         15479 => x"00",
         15480 => x"64",
         15481 => x"2d",
         15482 => x"25",
         15483 => x"64",
         15484 => x"2c",
         15485 => x"00",
         15486 => x"00",
         15487 => x"64",
         15488 => x"00",
         15489 => x"78",
         15490 => x"00",
         15491 => x"25",
         15492 => x"64",
         15493 => x"00",
         15494 => x"6f",
         15495 => x"43",
         15496 => x"6f",
         15497 => x"00",
         15498 => x"25",
         15499 => x"20",
         15500 => x"78",
         15501 => x"00",
         15502 => x"25",
         15503 => x"20",
         15504 => x"78",
         15505 => x"00",
         15506 => x"25",
         15507 => x"20",
         15508 => x"00",
         15509 => x"20",
         15510 => x"74",
         15511 => x"44",
         15512 => x"69",
         15513 => x"00",
         15514 => x"20",
         15515 => x"74",
         15516 => x"44",
         15517 => x"61",
         15518 => x"00",
         15519 => x"20",
         15520 => x"74",
         15521 => x"44",
         15522 => x"69",
         15523 => x"00",
         15524 => x"74",
         15525 => x"20",
         15526 => x"69",
         15527 => x"2e",
         15528 => x"00",
         15529 => x"00",
         15530 => x"3c",
         15531 => x"7f",
         15532 => x"00",
         15533 => x"3d",
         15534 => x"00",
         15535 => x"00",
         15536 => x"33",
         15537 => x"00",
         15538 => x"4d",
         15539 => x"53",
         15540 => x"00",
         15541 => x"4e",
         15542 => x"20",
         15543 => x"46",
         15544 => x"20",
         15545 => x"00",
         15546 => x"4e",
         15547 => x"20",
         15548 => x"46",
         15549 => x"32",
         15550 => x"00",
         15551 => x"a4",
         15552 => x"00",
         15553 => x"00",
         15554 => x"00",
         15555 => x"07",
         15556 => x"12",
         15557 => x"1c",
         15558 => x"00",
         15559 => x"41",
         15560 => x"80",
         15561 => x"49",
         15562 => x"8f",
         15563 => x"4f",
         15564 => x"55",
         15565 => x"9b",
         15566 => x"9f",
         15567 => x"55",
         15568 => x"a7",
         15569 => x"ab",
         15570 => x"af",
         15571 => x"b3",
         15572 => x"b7",
         15573 => x"bb",
         15574 => x"bf",
         15575 => x"c3",
         15576 => x"c7",
         15577 => x"cb",
         15578 => x"cf",
         15579 => x"d3",
         15580 => x"d7",
         15581 => x"db",
         15582 => x"df",
         15583 => x"e3",
         15584 => x"e7",
         15585 => x"eb",
         15586 => x"ef",
         15587 => x"f3",
         15588 => x"f7",
         15589 => x"fb",
         15590 => x"ff",
         15591 => x"3b",
         15592 => x"2f",
         15593 => x"3a",
         15594 => x"7c",
         15595 => x"00",
         15596 => x"04",
         15597 => x"40",
         15598 => x"00",
         15599 => x"00",
         15600 => x"02",
         15601 => x"08",
         15602 => x"20",
         15603 => x"00",
         15604 => x"fc",
         15605 => x"e2",
         15606 => x"e0",
         15607 => x"e7",
         15608 => x"eb",
         15609 => x"ef",
         15610 => x"ec",
         15611 => x"c5",
         15612 => x"e6",
         15613 => x"f4",
         15614 => x"f2",
         15615 => x"f9",
         15616 => x"d6",
         15617 => x"a2",
         15618 => x"a5",
         15619 => x"92",
         15620 => x"ed",
         15621 => x"fa",
         15622 => x"d1",
         15623 => x"ba",
         15624 => x"10",
         15625 => x"bd",
         15626 => x"a1",
         15627 => x"bb",
         15628 => x"92",
         15629 => x"02",
         15630 => x"61",
         15631 => x"56",
         15632 => x"63",
         15633 => x"57",
         15634 => x"5c",
         15635 => x"10",
         15636 => x"34",
         15637 => x"1c",
         15638 => x"3c",
         15639 => x"5f",
         15640 => x"54",
         15641 => x"66",
         15642 => x"50",
         15643 => x"67",
         15644 => x"64",
         15645 => x"59",
         15646 => x"52",
         15647 => x"6b",
         15648 => x"18",
         15649 => x"88",
         15650 => x"8c",
         15651 => x"80",
         15652 => x"df",
         15653 => x"c0",
         15654 => x"c3",
         15655 => x"c4",
         15656 => x"98",
         15657 => x"b4",
         15658 => x"c6",
         15659 => x"29",
         15660 => x"b1",
         15661 => x"64",
         15662 => x"21",
         15663 => x"48",
         15664 => x"19",
         15665 => x"1a",
         15666 => x"b2",
         15667 => x"a0",
         15668 => x"1a",
         15669 => x"17",
         15670 => x"07",
         15671 => x"01",
         15672 => x"00",
         15673 => x"32",
         15674 => x"39",
         15675 => x"4a",
         15676 => x"79",
         15677 => x"80",
         15678 => x"43",
         15679 => x"82",
         15680 => x"84",
         15681 => x"86",
         15682 => x"87",
         15683 => x"8a",
         15684 => x"8b",
         15685 => x"8e",
         15686 => x"90",
         15687 => x"91",
         15688 => x"94",
         15689 => x"96",
         15690 => x"98",
         15691 => x"3d",
         15692 => x"9c",
         15693 => x"20",
         15694 => x"a0",
         15695 => x"a2",
         15696 => x"a4",
         15697 => x"a6",
         15698 => x"a7",
         15699 => x"aa",
         15700 => x"ac",
         15701 => x"ae",
         15702 => x"af",
         15703 => x"b2",
         15704 => x"b3",
         15705 => x"b5",
         15706 => x"b8",
         15707 => x"ba",
         15708 => x"bc",
         15709 => x"be",
         15710 => x"c0",
         15711 => x"c2",
         15712 => x"c4",
         15713 => x"c4",
         15714 => x"c8",
         15715 => x"ca",
         15716 => x"ca",
         15717 => x"10",
         15718 => x"01",
         15719 => x"de",
         15720 => x"f3",
         15721 => x"f1",
         15722 => x"f4",
         15723 => x"28",
         15724 => x"12",
         15725 => x"09",
         15726 => x"3b",
         15727 => x"3d",
         15728 => x"3f",
         15729 => x"41",
         15730 => x"46",
         15731 => x"53",
         15732 => x"81",
         15733 => x"55",
         15734 => x"8a",
         15735 => x"8f",
         15736 => x"90",
         15737 => x"5d",
         15738 => x"5f",
         15739 => x"61",
         15740 => x"94",
         15741 => x"65",
         15742 => x"67",
         15743 => x"96",
         15744 => x"62",
         15745 => x"6d",
         15746 => x"9c",
         15747 => x"71",
         15748 => x"73",
         15749 => x"9f",
         15750 => x"77",
         15751 => x"79",
         15752 => x"7b",
         15753 => x"64",
         15754 => x"7f",
         15755 => x"81",
         15756 => x"a9",
         15757 => x"85",
         15758 => x"87",
         15759 => x"44",
         15760 => x"b2",
         15761 => x"8d",
         15762 => x"8f",
         15763 => x"91",
         15764 => x"7b",
         15765 => x"fd",
         15766 => x"ff",
         15767 => x"04",
         15768 => x"88",
         15769 => x"8a",
         15770 => x"11",
         15771 => x"02",
         15772 => x"a3",
         15773 => x"08",
         15774 => x"03",
         15775 => x"8e",
         15776 => x"d8",
         15777 => x"f2",
         15778 => x"f9",
         15779 => x"f4",
         15780 => x"f6",
         15781 => x"f7",
         15782 => x"fa",
         15783 => x"30",
         15784 => x"50",
         15785 => x"60",
         15786 => x"8a",
         15787 => x"c1",
         15788 => x"cf",
         15789 => x"c0",
         15790 => x"44",
         15791 => x"26",
         15792 => x"00",
         15793 => x"01",
         15794 => x"00",
         15795 => x"a0",
         15796 => x"00",
         15797 => x"10",
         15798 => x"20",
         15799 => x"30",
         15800 => x"40",
         15801 => x"51",
         15802 => x"59",
         15803 => x"5b",
         15804 => x"5d",
         15805 => x"5f",
         15806 => x"08",
         15807 => x"0e",
         15808 => x"bb",
         15809 => x"c9",
         15810 => x"cb",
         15811 => x"db",
         15812 => x"f9",
         15813 => x"eb",
         15814 => x"fb",
         15815 => x"08",
         15816 => x"08",
         15817 => x"08",
         15818 => x"04",
         15819 => x"b9",
         15820 => x"bc",
         15821 => x"01",
         15822 => x"d0",
         15823 => x"e0",
         15824 => x"e5",
         15825 => x"ec",
         15826 => x"01",
         15827 => x"4e",
         15828 => x"32",
         15829 => x"10",
         15830 => x"01",
         15831 => x"d0",
         15832 => x"30",
         15833 => x"60",
         15834 => x"67",
         15835 => x"75",
         15836 => x"80",
         15837 => x"00",
         15838 => x"41",
         15839 => x"00",
         15840 => x"00",
         15841 => x"b0",
         15842 => x"00",
         15843 => x"00",
         15844 => x"00",
         15845 => x"b8",
         15846 => x"00",
         15847 => x"00",
         15848 => x"00",
         15849 => x"c0",
         15850 => x"00",
         15851 => x"00",
         15852 => x"00",
         15853 => x"c8",
         15854 => x"00",
         15855 => x"00",
         15856 => x"00",
         15857 => x"d0",
         15858 => x"00",
         15859 => x"00",
         15860 => x"00",
         15861 => x"d8",
         15862 => x"00",
         15863 => x"00",
         15864 => x"00",
         15865 => x"e0",
         15866 => x"00",
         15867 => x"00",
         15868 => x"00",
         15869 => x"e8",
         15870 => x"00",
         15871 => x"00",
         15872 => x"00",
         15873 => x"f0",
         15874 => x"00",
         15875 => x"00",
         15876 => x"00",
         15877 => x"f8",
         15878 => x"00",
         15879 => x"00",
         15880 => x"00",
         15881 => x"fc",
         15882 => x"00",
         15883 => x"00",
         15884 => x"00",
         15885 => x"00",
         15886 => x"00",
         15887 => x"00",
         15888 => x"00",
         15889 => x"04",
         15890 => x"00",
         15891 => x"00",
         15892 => x"00",
         15893 => x"08",
         15894 => x"00",
         15895 => x"00",
         15896 => x"00",
         15897 => x"0c",
         15898 => x"00",
         15899 => x"00",
         15900 => x"00",
         15901 => x"10",
         15902 => x"00",
         15903 => x"00",
         15904 => x"00",
         15905 => x"14",
         15906 => x"00",
         15907 => x"00",
         15908 => x"00",
         15909 => x"1c",
         15910 => x"00",
         15911 => x"00",
         15912 => x"00",
         15913 => x"20",
         15914 => x"00",
         15915 => x"00",
         15916 => x"00",
         15917 => x"28",
         15918 => x"00",
         15919 => x"00",
         15920 => x"00",
         15921 => x"30",
         15922 => x"00",
         15923 => x"00",
         15924 => x"00",
         15925 => x"38",
         15926 => x"00",
         15927 => x"00",
         15928 => x"00",
         15929 => x"40",
         15930 => x"00",
         15931 => x"00",
         15932 => x"00",
         15933 => x"44",
         15934 => x"00",
         15935 => x"00",
         15936 => x"00",
         15937 => x"48",
         15938 => x"00",
         15939 => x"00",
         15940 => x"00",
         15941 => x"50",
         15942 => x"00",
         15943 => x"00",
         15944 => x"00",
         15945 => x"58",
         15946 => x"00",
         15947 => x"00",
         15948 => x"00",
         15949 => x"60",
         15950 => x"00",
         15951 => x"00",
         15952 => x"00",
         15953 => x"00",
         15954 => x"00",
         15955 => x"ff",
         15956 => x"00",
         15957 => x"ff",
         15958 => x"00",
         15959 => x"ff",
         15960 => x"00",
         15961 => x"00",
         15962 => x"00",
         15963 => x"ff",
         15964 => x"00",
         15965 => x"00",
         15966 => x"00",
         15967 => x"00",
         15968 => x"00",
         15969 => x"00",
         15970 => x"00",
         15971 => x"00",
         15972 => x"01",
         15973 => x"01",
         15974 => x"01",
         15975 => x"00",
         15976 => x"00",
         15977 => x"00",
         15978 => x"00",
         15979 => x"00",
         15980 => x"00",
         15981 => x"00",
         15982 => x"00",
         15983 => x"00",
         15984 => x"00",
         15985 => x"00",
         15986 => x"00",
         15987 => x"00",
         15988 => x"00",
         15989 => x"00",
         15990 => x"00",
         15991 => x"00",
         15992 => x"00",
         15993 => x"00",
         15994 => x"00",
         15995 => x"00",
         15996 => x"00",
         15997 => x"00",
         15998 => x"00",
         15999 => x"00",
         16000 => x"e4",
         16001 => x"00",
         16002 => x"ec",
         16003 => x"00",
         16004 => x"f4",
         16005 => x"00",
         16006 => x"80",
         16007 => x"fd",
         16008 => x"0d",
         16009 => x"5b",
         16010 => x"f0",
         16011 => x"74",
         16012 => x"78",
         16013 => x"6c",
         16014 => x"70",
         16015 => x"64",
         16016 => x"68",
         16017 => x"34",
         16018 => x"38",
         16019 => x"20",
         16020 => x"2e",
         16021 => x"f4",
         16022 => x"2f",
         16023 => x"f0",
         16024 => x"f0",
         16025 => x"83",
         16026 => x"f0",
         16027 => x"fd",
         16028 => x"0d",
         16029 => x"5b",
         16030 => x"f0",
         16031 => x"54",
         16032 => x"58",
         16033 => x"4c",
         16034 => x"50",
         16035 => x"44",
         16036 => x"48",
         16037 => x"34",
         16038 => x"38",
         16039 => x"20",
         16040 => x"2e",
         16041 => x"f4",
         16042 => x"2f",
         16043 => x"f0",
         16044 => x"f0",
         16045 => x"83",
         16046 => x"f0",
         16047 => x"fd",
         16048 => x"0d",
         16049 => x"7b",
         16050 => x"f0",
         16051 => x"54",
         16052 => x"58",
         16053 => x"4c",
         16054 => x"50",
         16055 => x"44",
         16056 => x"48",
         16057 => x"24",
         16058 => x"28",
         16059 => x"20",
         16060 => x"3e",
         16061 => x"e1",
         16062 => x"2f",
         16063 => x"f0",
         16064 => x"f0",
         16065 => x"88",
         16066 => x"f0",
         16067 => x"fa",
         16068 => x"f0",
         16069 => x"1b",
         16070 => x"f0",
         16071 => x"14",
         16072 => x"18",
         16073 => x"0c",
         16074 => x"10",
         16075 => x"04",
         16076 => x"08",
         16077 => x"f0",
         16078 => x"f0",
         16079 => x"f0",
         16080 => x"f0",
         16081 => x"f0",
         16082 => x"1c",
         16083 => x"f0",
         16084 => x"f0",
         16085 => x"83",
         16086 => x"f0",
         16087 => x"c9",
         16088 => x"cd",
         16089 => x"b3",
         16090 => x"f0",
         16091 => x"31",
         16092 => x"dd",
         16093 => x"56",
         16094 => x"b1",
         16095 => x"48",
         16096 => x"73",
         16097 => x"3b",
         16098 => x"a2",
         16099 => x"00",
         16100 => x"b9",
         16101 => x"c1",
         16102 => x"be",
         16103 => x"f0",
         16104 => x"f0",
         16105 => x"83",
         16106 => x"f0",
         16107 => x"00",
         16108 => x"00",
         16109 => x"00",
         16110 => x"00",
         16111 => x"00",
         16112 => x"00",
         16113 => x"00",
         16114 => x"00",
         16115 => x"00",
         16116 => x"00",
         16117 => x"00",
         16118 => x"00",
         16119 => x"00",
         16120 => x"00",
         16121 => x"00",
         16122 => x"00",
         16123 => x"00",
         16124 => x"00",
         16125 => x"00",
         16126 => x"00",
         16127 => x"00",
         16128 => x"00",
         16129 => x"00",
         16130 => x"00",
         16131 => x"00",
         16132 => x"00",
         16133 => x"00",
         16134 => x"00",
         16135 => x"38",
         16136 => x"00",
         16137 => x"40",
         16138 => x"00",
         16139 => x"44",
         16140 => x"00",
         16141 => x"48",
         16142 => x"00",
         16143 => x"4c",
         16144 => x"00",
         16145 => x"50",
         16146 => x"00",
         16147 => x"58",
         16148 => x"00",
         16149 => x"60",
         16150 => x"00",
         16151 => x"68",
         16152 => x"00",
         16153 => x"70",
         16154 => x"00",
         16155 => x"78",
         16156 => x"00",
         16157 => x"80",
         16158 => x"00",
         16159 => x"88",
         16160 => x"00",
         16161 => x"90",
         16162 => x"00",
         16163 => x"98",
         16164 => x"00",
         16165 => x"a0",
         16166 => x"00",
         16167 => x"a8",
         16168 => x"00",
         16169 => x"b0",
         16170 => x"00",
         16171 => x"b4",
         16172 => x"00",
         16173 => x"bc",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"00",
         18159 => x"00",
         18160 => x"00",
         18161 => x"00",
         18162 => x"00",
         18163 => x"00",
         18164 => x"00",
         18165 => x"00",
         18166 => x"00",
         18167 => x"00",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"19",
         18176 => x"01",
         18177 => x"00",
         18178 => x"f3",
         18179 => x"f7",
         18180 => x"fb",
         18181 => x"ff",
         18182 => x"c3",
         18183 => x"e2",
         18184 => x"e6",
         18185 => x"f4",
         18186 => x"63",
         18187 => x"67",
         18188 => x"6a",
         18189 => x"2d",
         18190 => x"23",
         18191 => x"27",
         18192 => x"2c",
         18193 => x"49",
         18194 => x"03",
         18195 => x"07",
         18196 => x"0b",
         18197 => x"0f",
         18198 => x"13",
         18199 => x"17",
         18200 => x"52",
         18201 => x"3c",
         18202 => x"83",
         18203 => x"87",
         18204 => x"8b",
         18205 => x"8f",
         18206 => x"93",
         18207 => x"97",
         18208 => x"bc",
         18209 => x"c0",
         18210 => x"00",
         18211 => x"00",
         18212 => x"00",
         18213 => x"00",
         18214 => x"00",
         18215 => x"00",
         18216 => x"00",
         18217 => x"00",
         18218 => x"00",
         18219 => x"00",
         18220 => x"00",
         18221 => x"00",
         18222 => x"00",
         18223 => x"00",
         18224 => x"00",
         18225 => x"00",
         18226 => x"00",
         18227 => x"00",
         18228 => x"00",
         18229 => x"00",
         18230 => x"00",
         18231 => x"00",
         18232 => x"00",
         18233 => x"00",
         18234 => x"00",
         18235 => x"00",
         18236 => x"00",
         18237 => x"00",
         18238 => x"00",
         18239 => x"00",
         18240 => x"03",
         18241 => x"01",
         18242 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"0b",
             2 => x"e9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"83",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a6",
           270 => x"0b",
           271 => x"0b",
           272 => x"c6",
           273 => x"0b",
           274 => x"0b",
           275 => x"e6",
           276 => x"0b",
           277 => x"0b",
           278 => x"86",
           279 => x"0b",
           280 => x"0b",
           281 => x"a6",
           282 => x"0b",
           283 => x"0b",
           284 => x"c6",
           285 => x"0b",
           286 => x"0b",
           287 => x"e8",
           288 => x"0b",
           289 => x"0b",
           290 => x"8a",
           291 => x"0b",
           292 => x"0b",
           293 => x"ac",
           294 => x"0b",
           295 => x"0b",
           296 => x"ce",
           297 => x"0b",
           298 => x"0b",
           299 => x"f0",
           300 => x"0b",
           301 => x"0b",
           302 => x"92",
           303 => x"0b",
           304 => x"0b",
           305 => x"b4",
           306 => x"0b",
           307 => x"0b",
           308 => x"d6",
           309 => x"0b",
           310 => x"0b",
           311 => x"f8",
           312 => x"0b",
           313 => x"0b",
           314 => x"9a",
           315 => x"0b",
           316 => x"0b",
           317 => x"bc",
           318 => x"0b",
           319 => x"0b",
           320 => x"de",
           321 => x"0b",
           322 => x"0b",
           323 => x"80",
           324 => x"0b",
           325 => x"0b",
           326 => x"a2",
           327 => x"0b",
           328 => x"0b",
           329 => x"c4",
           330 => x"0b",
           331 => x"0b",
           332 => x"e6",
           333 => x"0b",
           334 => x"0b",
           335 => x"88",
           336 => x"0b",
           337 => x"0b",
           338 => x"aa",
           339 => x"0b",
           340 => x"0b",
           341 => x"cb",
           342 => x"0b",
           343 => x"0b",
           344 => x"ed",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"ba",
           386 => x"d5",
           387 => x"ba",
           388 => x"c0",
           389 => x"84",
           390 => x"a2",
           391 => x"ba",
           392 => x"c0",
           393 => x"84",
           394 => x"a0",
           395 => x"ba",
           396 => x"c0",
           397 => x"84",
           398 => x"a0",
           399 => x"ba",
           400 => x"c0",
           401 => x"84",
           402 => x"94",
           403 => x"ba",
           404 => x"c0",
           405 => x"84",
           406 => x"a1",
           407 => x"ba",
           408 => x"c0",
           409 => x"84",
           410 => x"af",
           411 => x"ba",
           412 => x"c0",
           413 => x"84",
           414 => x"ad",
           415 => x"ba",
           416 => x"c0",
           417 => x"84",
           418 => x"94",
           419 => x"ba",
           420 => x"c0",
           421 => x"84",
           422 => x"95",
           423 => x"ba",
           424 => x"c0",
           425 => x"84",
           426 => x"95",
           427 => x"ba",
           428 => x"c0",
           429 => x"84",
           430 => x"b1",
           431 => x"ba",
           432 => x"c0",
           433 => x"84",
           434 => x"80",
           435 => x"84",
           436 => x"80",
           437 => x"04",
           438 => x"0c",
           439 => x"2d",
           440 => x"08",
           441 => x"90",
           442 => x"98",
           443 => x"97",
           444 => x"98",
           445 => x"80",
           446 => x"ba",
           447 => x"d3",
           448 => x"ba",
           449 => x"c0",
           450 => x"84",
           451 => x"82",
           452 => x"84",
           453 => x"80",
           454 => x"04",
           455 => x"0c",
           456 => x"2d",
           457 => x"08",
           458 => x"90",
           459 => x"98",
           460 => x"e7",
           461 => x"98",
           462 => x"80",
           463 => x"ba",
           464 => x"d8",
           465 => x"ba",
           466 => x"c0",
           467 => x"84",
           468 => x"82",
           469 => x"84",
           470 => x"80",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"90",
           476 => x"98",
           477 => x"d0",
           478 => x"98",
           479 => x"80",
           480 => x"ba",
           481 => x"f2",
           482 => x"ba",
           483 => x"c0",
           484 => x"84",
           485 => x"82",
           486 => x"84",
           487 => x"80",
           488 => x"04",
           489 => x"0c",
           490 => x"2d",
           491 => x"08",
           492 => x"90",
           493 => x"98",
           494 => x"eb",
           495 => x"98",
           496 => x"80",
           497 => x"ba",
           498 => x"ff",
           499 => x"ba",
           500 => x"c0",
           501 => x"84",
           502 => x"83",
           503 => x"84",
           504 => x"80",
           505 => x"04",
           506 => x"0c",
           507 => x"2d",
           508 => x"08",
           509 => x"90",
           510 => x"98",
           511 => x"c6",
           512 => x"98",
           513 => x"80",
           514 => x"ba",
           515 => x"95",
           516 => x"ba",
           517 => x"c0",
           518 => x"84",
           519 => x"82",
           520 => x"84",
           521 => x"80",
           522 => x"04",
           523 => x"0c",
           524 => x"2d",
           525 => x"08",
           526 => x"90",
           527 => x"98",
           528 => x"d7",
           529 => x"98",
           530 => x"80",
           531 => x"ba",
           532 => x"f6",
           533 => x"ba",
           534 => x"c0",
           535 => x"84",
           536 => x"83",
           537 => x"84",
           538 => x"80",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"90",
           544 => x"98",
           545 => x"b2",
           546 => x"98",
           547 => x"80",
           548 => x"ba",
           549 => x"c7",
           550 => x"ba",
           551 => x"c0",
           552 => x"84",
           553 => x"83",
           554 => x"84",
           555 => x"80",
           556 => x"04",
           557 => x"0c",
           558 => x"2d",
           559 => x"08",
           560 => x"90",
           561 => x"98",
           562 => x"8e",
           563 => x"98",
           564 => x"80",
           565 => x"ba",
           566 => x"f4",
           567 => x"ba",
           568 => x"c0",
           569 => x"84",
           570 => x"81",
           571 => x"84",
           572 => x"80",
           573 => x"04",
           574 => x"0c",
           575 => x"2d",
           576 => x"08",
           577 => x"90",
           578 => x"98",
           579 => x"99",
           580 => x"98",
           581 => x"80",
           582 => x"ba",
           583 => x"d1",
           584 => x"ba",
           585 => x"c0",
           586 => x"84",
           587 => x"80",
           588 => x"84",
           589 => x"80",
           590 => x"04",
           591 => x"0c",
           592 => x"84",
           593 => x"80",
           594 => x"04",
           595 => x"0c",
           596 => x"2d",
           597 => x"08",
           598 => x"90",
           599 => x"98",
           600 => x"85",
           601 => x"98",
           602 => x"80",
           603 => x"ba",
           604 => x"f2",
           605 => x"ba",
           606 => x"c0",
           607 => x"84",
           608 => x"81",
           609 => x"84",
           610 => x"80",
           611 => x"04",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"04",
           621 => x"81",
           622 => x"83",
           623 => x"05",
           624 => x"10",
           625 => x"72",
           626 => x"51",
           627 => x"72",
           628 => x"06",
           629 => x"72",
           630 => x"10",
           631 => x"10",
           632 => x"ed",
           633 => x"53",
           634 => x"ba",
           635 => x"d5",
           636 => x"38",
           637 => x"84",
           638 => x"0b",
           639 => x"ec",
           640 => x"51",
           641 => x"04",
           642 => x"0d",
           643 => x"70",
           644 => x"08",
           645 => x"52",
           646 => x"08",
           647 => x"3f",
           648 => x"04",
           649 => x"78",
           650 => x"11",
           651 => x"81",
           652 => x"25",
           653 => x"55",
           654 => x"72",
           655 => x"81",
           656 => x"38",
           657 => x"74",
           658 => x"30",
           659 => x"9f",
           660 => x"55",
           661 => x"74",
           662 => x"71",
           663 => x"38",
           664 => x"fa",
           665 => x"8c",
           666 => x"ba",
           667 => x"2e",
           668 => x"ba",
           669 => x"70",
           670 => x"34",
           671 => x"8a",
           672 => x"70",
           673 => x"2a",
           674 => x"54",
           675 => x"cb",
           676 => x"34",
           677 => x"84",
           678 => x"88",
           679 => x"80",
           680 => x"8c",
           681 => x"0d",
           682 => x"0d",
           683 => x"02",
           684 => x"05",
           685 => x"fe",
           686 => x"3d",
           687 => x"7e",
           688 => x"e4",
           689 => x"3f",
           690 => x"80",
           691 => x"3d",
           692 => x"3d",
           693 => x"88",
           694 => x"52",
           695 => x"3f",
           696 => x"04",
           697 => x"61",
           698 => x"5d",
           699 => x"8c",
           700 => x"1e",
           701 => x"2a",
           702 => x"06",
           703 => x"ff",
           704 => x"2e",
           705 => x"80",
           706 => x"33",
           707 => x"2e",
           708 => x"81",
           709 => x"06",
           710 => x"80",
           711 => x"38",
           712 => x"7e",
           713 => x"a3",
           714 => x"32",
           715 => x"80",
           716 => x"55",
           717 => x"72",
           718 => x"38",
           719 => x"70",
           720 => x"06",
           721 => x"80",
           722 => x"7a",
           723 => x"5b",
           724 => x"76",
           725 => x"8c",
           726 => x"73",
           727 => x"0c",
           728 => x"04",
           729 => x"54",
           730 => x"10",
           731 => x"70",
           732 => x"98",
           733 => x"81",
           734 => x"8b",
           735 => x"98",
           736 => x"5b",
           737 => x"79",
           738 => x"38",
           739 => x"53",
           740 => x"38",
           741 => x"58",
           742 => x"f7",
           743 => x"39",
           744 => x"09",
           745 => x"38",
           746 => x"5a",
           747 => x"7c",
           748 => x"76",
           749 => x"ff",
           750 => x"52",
           751 => x"af",
           752 => x"57",
           753 => x"38",
           754 => x"7a",
           755 => x"81",
           756 => x"78",
           757 => x"70",
           758 => x"54",
           759 => x"e0",
           760 => x"80",
           761 => x"38",
           762 => x"83",
           763 => x"54",
           764 => x"73",
           765 => x"59",
           766 => x"27",
           767 => x"52",
           768 => x"eb",
           769 => x"33",
           770 => x"fe",
           771 => x"c7",
           772 => x"59",
           773 => x"88",
           774 => x"84",
           775 => x"7d",
           776 => x"06",
           777 => x"54",
           778 => x"5e",
           779 => x"51",
           780 => x"84",
           781 => x"81",
           782 => x"ba",
           783 => x"df",
           784 => x"72",
           785 => x"38",
           786 => x"08",
           787 => x"74",
           788 => x"05",
           789 => x"52",
           790 => x"ca",
           791 => x"8c",
           792 => x"ba",
           793 => x"38",
           794 => x"9c",
           795 => x"7b",
           796 => x"56",
           797 => x"8f",
           798 => x"80",
           799 => x"80",
           800 => x"90",
           801 => x"7a",
           802 => x"81",
           803 => x"73",
           804 => x"38",
           805 => x"80",
           806 => x"80",
           807 => x"90",
           808 => x"77",
           809 => x"29",
           810 => x"05",
           811 => x"2c",
           812 => x"2a",
           813 => x"54",
           814 => x"2e",
           815 => x"98",
           816 => x"ff",
           817 => x"78",
           818 => x"cc",
           819 => x"ff",
           820 => x"83",
           821 => x"2a",
           822 => x"74",
           823 => x"73",
           824 => x"f0",
           825 => x"31",
           826 => x"90",
           827 => x"80",
           828 => x"53",
           829 => x"85",
           830 => x"81",
           831 => x"54",
           832 => x"38",
           833 => x"81",
           834 => x"86",
           835 => x"85",
           836 => x"54",
           837 => x"38",
           838 => x"54",
           839 => x"38",
           840 => x"81",
           841 => x"80",
           842 => x"77",
           843 => x"80",
           844 => x"80",
           845 => x"2c",
           846 => x"80",
           847 => x"38",
           848 => x"51",
           849 => x"77",
           850 => x"80",
           851 => x"80",
           852 => x"2c",
           853 => x"73",
           854 => x"38",
           855 => x"53",
           856 => x"b2",
           857 => x"81",
           858 => x"81",
           859 => x"70",
           860 => x"55",
           861 => x"25",
           862 => x"52",
           863 => x"ef",
           864 => x"81",
           865 => x"81",
           866 => x"70",
           867 => x"55",
           868 => x"24",
           869 => x"87",
           870 => x"06",
           871 => x"80",
           872 => x"38",
           873 => x"2e",
           874 => x"76",
           875 => x"81",
           876 => x"80",
           877 => x"e2",
           878 => x"ba",
           879 => x"38",
           880 => x"1e",
           881 => x"5e",
           882 => x"7d",
           883 => x"2e",
           884 => x"ec",
           885 => x"06",
           886 => x"2e",
           887 => x"77",
           888 => x"80",
           889 => x"80",
           890 => x"2c",
           891 => x"80",
           892 => x"91",
           893 => x"a0",
           894 => x"3f",
           895 => x"90",
           896 => x"a0",
           897 => x"58",
           898 => x"87",
           899 => x"39",
           900 => x"07",
           901 => x"57",
           902 => x"84",
           903 => x"7e",
           904 => x"06",
           905 => x"55",
           906 => x"39",
           907 => x"05",
           908 => x"0a",
           909 => x"33",
           910 => x"72",
           911 => x"80",
           912 => x"80",
           913 => x"90",
           914 => x"5a",
           915 => x"5f",
           916 => x"70",
           917 => x"55",
           918 => x"38",
           919 => x"80",
           920 => x"80",
           921 => x"90",
           922 => x"5f",
           923 => x"fe",
           924 => x"52",
           925 => x"f7",
           926 => x"ff",
           927 => x"ff",
           928 => x"57",
           929 => x"ff",
           930 => x"38",
           931 => x"70",
           932 => x"33",
           933 => x"3f",
           934 => x"1a",
           935 => x"ff",
           936 => x"79",
           937 => x"2e",
           938 => x"7c",
           939 => x"81",
           940 => x"51",
           941 => x"e2",
           942 => x"0a",
           943 => x"0a",
           944 => x"80",
           945 => x"80",
           946 => x"90",
           947 => x"56",
           948 => x"87",
           949 => x"06",
           950 => x"7a",
           951 => x"fe",
           952 => x"60",
           953 => x"08",
           954 => x"41",
           955 => x"24",
           956 => x"7a",
           957 => x"06",
           958 => x"9c",
           959 => x"39",
           960 => x"7c",
           961 => x"76",
           962 => x"f8",
           963 => x"88",
           964 => x"7c",
           965 => x"76",
           966 => x"f8",
           967 => x"60",
           968 => x"08",
           969 => x"56",
           970 => x"72",
           971 => x"75",
           972 => x"3f",
           973 => x"08",
           974 => x"06",
           975 => x"90",
           976 => x"72",
           977 => x"fe",
           978 => x"80",
           979 => x"33",
           980 => x"f7",
           981 => x"ff",
           982 => x"84",
           983 => x"77",
           984 => x"58",
           985 => x"81",
           986 => x"51",
           987 => x"84",
           988 => x"83",
           989 => x"78",
           990 => x"2b",
           991 => x"39",
           992 => x"07",
           993 => x"5b",
           994 => x"38",
           995 => x"77",
           996 => x"80",
           997 => x"80",
           998 => x"2c",
           999 => x"80",
          1000 => x"d6",
          1001 => x"a0",
          1002 => x"3f",
          1003 => x"52",
          1004 => x"bb",
          1005 => x"2e",
          1006 => x"fa",
          1007 => x"52",
          1008 => x"ab",
          1009 => x"2a",
          1010 => x"7e",
          1011 => x"8c",
          1012 => x"39",
          1013 => x"78",
          1014 => x"2b",
          1015 => x"7d",
          1016 => x"57",
          1017 => x"73",
          1018 => x"ff",
          1019 => x"52",
          1020 => x"fb",
          1021 => x"06",
          1022 => x"2e",
          1023 => x"ff",
          1024 => x"52",
          1025 => x"51",
          1026 => x"74",
          1027 => x"7a",
          1028 => x"f1",
          1029 => x"39",
          1030 => x"98",
          1031 => x"2c",
          1032 => x"b7",
          1033 => x"ab",
          1034 => x"3f",
          1035 => x"52",
          1036 => x"bb",
          1037 => x"39",
          1038 => x"51",
          1039 => x"84",
          1040 => x"83",
          1041 => x"78",
          1042 => x"2b",
          1043 => x"f3",
          1044 => x"07",
          1045 => x"83",
          1046 => x"52",
          1047 => x"99",
          1048 => x"0d",
          1049 => x"08",
          1050 => x"74",
          1051 => x"3f",
          1052 => x"04",
          1053 => x"78",
          1054 => x"84",
          1055 => x"85",
          1056 => x"81",
          1057 => x"70",
          1058 => x"56",
          1059 => x"ff",
          1060 => x"2e",
          1061 => x"80",
          1062 => x"70",
          1063 => x"33",
          1064 => x"2e",
          1065 => x"d5",
          1066 => x"72",
          1067 => x"08",
          1068 => x"84",
          1069 => x"80",
          1070 => x"ff",
          1071 => x"81",
          1072 => x"53",
          1073 => x"88",
          1074 => x"f0",
          1075 => x"39",
          1076 => x"08",
          1077 => x"f0",
          1078 => x"51",
          1079 => x"55",
          1080 => x"ba",
          1081 => x"2e",
          1082 => x"57",
          1083 => x"84",
          1084 => x"88",
          1085 => x"fa",
          1086 => x"7a",
          1087 => x"0b",
          1088 => x"70",
          1089 => x"32",
          1090 => x"51",
          1091 => x"ff",
          1092 => x"2e",
          1093 => x"92",
          1094 => x"81",
          1095 => x"53",
          1096 => x"09",
          1097 => x"38",
          1098 => x"84",
          1099 => x"88",
          1100 => x"73",
          1101 => x"55",
          1102 => x"80",
          1103 => x"74",
          1104 => x"90",
          1105 => x"72",
          1106 => x"8c",
          1107 => x"e3",
          1108 => x"70",
          1109 => x"33",
          1110 => x"e3",
          1111 => x"ff",
          1112 => x"d5",
          1113 => x"73",
          1114 => x"83",
          1115 => x"fa",
          1116 => x"7a",
          1117 => x"70",
          1118 => x"32",
          1119 => x"56",
          1120 => x"56",
          1121 => x"73",
          1122 => x"06",
          1123 => x"2e",
          1124 => x"15",
          1125 => x"88",
          1126 => x"91",
          1127 => x"56",
          1128 => x"74",
          1129 => x"75",
          1130 => x"08",
          1131 => x"8c",
          1132 => x"56",
          1133 => x"8c",
          1134 => x"0d",
          1135 => x"76",
          1136 => x"51",
          1137 => x"54",
          1138 => x"56",
          1139 => x"08",
          1140 => x"15",
          1141 => x"8c",
          1142 => x"56",
          1143 => x"3d",
          1144 => x"11",
          1145 => x"ff",
          1146 => x"32",
          1147 => x"55",
          1148 => x"54",
          1149 => x"72",
          1150 => x"06",
          1151 => x"38",
          1152 => x"81",
          1153 => x"80",
          1154 => x"38",
          1155 => x"33",
          1156 => x"80",
          1157 => x"38",
          1158 => x"0c",
          1159 => x"81",
          1160 => x"0c",
          1161 => x"06",
          1162 => x"ba",
          1163 => x"3d",
          1164 => x"ff",
          1165 => x"72",
          1166 => x"8c",
          1167 => x"05",
          1168 => x"84",
          1169 => x"ba",
          1170 => x"3d",
          1171 => x"51",
          1172 => x"55",
          1173 => x"ba",
          1174 => x"84",
          1175 => x"80",
          1176 => x"38",
          1177 => x"70",
          1178 => x"52",
          1179 => x"08",
          1180 => x"38",
          1181 => x"53",
          1182 => x"34",
          1183 => x"84",
          1184 => x"87",
          1185 => x"74",
          1186 => x"72",
          1187 => x"ff",
          1188 => x"fd",
          1189 => x"77",
          1190 => x"54",
          1191 => x"05",
          1192 => x"70",
          1193 => x"12",
          1194 => x"81",
          1195 => x"51",
          1196 => x"81",
          1197 => x"70",
          1198 => x"84",
          1199 => x"85",
          1200 => x"fc",
          1201 => x"79",
          1202 => x"55",
          1203 => x"80",
          1204 => x"73",
          1205 => x"38",
          1206 => x"93",
          1207 => x"81",
          1208 => x"73",
          1209 => x"55",
          1210 => x"51",
          1211 => x"73",
          1212 => x"0c",
          1213 => x"04",
          1214 => x"73",
          1215 => x"38",
          1216 => x"53",
          1217 => x"ff",
          1218 => x"71",
          1219 => x"ff",
          1220 => x"80",
          1221 => x"ff",
          1222 => x"53",
          1223 => x"73",
          1224 => x"51",
          1225 => x"c7",
          1226 => x"0d",
          1227 => x"53",
          1228 => x"05",
          1229 => x"70",
          1230 => x"12",
          1231 => x"84",
          1232 => x"51",
          1233 => x"04",
          1234 => x"75",
          1235 => x"54",
          1236 => x"81",
          1237 => x"51",
          1238 => x"81",
          1239 => x"70",
          1240 => x"84",
          1241 => x"85",
          1242 => x"fd",
          1243 => x"78",
          1244 => x"55",
          1245 => x"80",
          1246 => x"71",
          1247 => x"53",
          1248 => x"81",
          1249 => x"ff",
          1250 => x"ef",
          1251 => x"ba",
          1252 => x"3d",
          1253 => x"3d",
          1254 => x"7a",
          1255 => x"72",
          1256 => x"38",
          1257 => x"70",
          1258 => x"33",
          1259 => x"71",
          1260 => x"06",
          1261 => x"14",
          1262 => x"2e",
          1263 => x"13",
          1264 => x"38",
          1265 => x"84",
          1266 => x"86",
          1267 => x"72",
          1268 => x"38",
          1269 => x"ff",
          1270 => x"2e",
          1271 => x"15",
          1272 => x"51",
          1273 => x"de",
          1274 => x"31",
          1275 => x"0c",
          1276 => x"04",
          1277 => x"8c",
          1278 => x"0d",
          1279 => x"0d",
          1280 => x"70",
          1281 => x"c1",
          1282 => x"8c",
          1283 => x"8c",
          1284 => x"52",
          1285 => x"b3",
          1286 => x"8c",
          1287 => x"ba",
          1288 => x"2e",
          1289 => x"ba",
          1290 => x"54",
          1291 => x"74",
          1292 => x"84",
          1293 => x"51",
          1294 => x"84",
          1295 => x"54",
          1296 => x"8c",
          1297 => x"0d",
          1298 => x"0d",
          1299 => x"71",
          1300 => x"54",
          1301 => x"9f",
          1302 => x"81",
          1303 => x"51",
          1304 => x"8c",
          1305 => x"52",
          1306 => x"09",
          1307 => x"38",
          1308 => x"75",
          1309 => x"70",
          1310 => x"0c",
          1311 => x"04",
          1312 => x"75",
          1313 => x"55",
          1314 => x"70",
          1315 => x"38",
          1316 => x"81",
          1317 => x"ff",
          1318 => x"f4",
          1319 => x"ba",
          1320 => x"3d",
          1321 => x"3d",
          1322 => x"58",
          1323 => x"76",
          1324 => x"38",
          1325 => x"f5",
          1326 => x"8c",
          1327 => x"12",
          1328 => x"2e",
          1329 => x"51",
          1330 => x"71",
          1331 => x"08",
          1332 => x"52",
          1333 => x"80",
          1334 => x"52",
          1335 => x"80",
          1336 => x"13",
          1337 => x"a0",
          1338 => x"71",
          1339 => x"54",
          1340 => x"74",
          1341 => x"38",
          1342 => x"9f",
          1343 => x"10",
          1344 => x"72",
          1345 => x"9f",
          1346 => x"06",
          1347 => x"75",
          1348 => x"1c",
          1349 => x"52",
          1350 => x"53",
          1351 => x"73",
          1352 => x"52",
          1353 => x"8c",
          1354 => x"0d",
          1355 => x"0d",
          1356 => x"80",
          1357 => x"30",
          1358 => x"80",
          1359 => x"2b",
          1360 => x"75",
          1361 => x"83",
          1362 => x"70",
          1363 => x"25",
          1364 => x"71",
          1365 => x"2a",
          1366 => x"06",
          1367 => x"80",
          1368 => x"84",
          1369 => x"71",
          1370 => x"75",
          1371 => x"8c",
          1372 => x"70",
          1373 => x"82",
          1374 => x"71",
          1375 => x"2a",
          1376 => x"81",
          1377 => x"82",
          1378 => x"75",
          1379 => x"ba",
          1380 => x"52",
          1381 => x"54",
          1382 => x"55",
          1383 => x"56",
          1384 => x"51",
          1385 => x"52",
          1386 => x"04",
          1387 => x"75",
          1388 => x"71",
          1389 => x"81",
          1390 => x"ba",
          1391 => x"29",
          1392 => x"84",
          1393 => x"53",
          1394 => x"04",
          1395 => x"78",
          1396 => x"a0",
          1397 => x"2e",
          1398 => x"51",
          1399 => x"84",
          1400 => x"53",
          1401 => x"73",
          1402 => x"38",
          1403 => x"bd",
          1404 => x"ba",
          1405 => x"52",
          1406 => x"9f",
          1407 => x"38",
          1408 => x"9f",
          1409 => x"81",
          1410 => x"2a",
          1411 => x"76",
          1412 => x"54",
          1413 => x"56",
          1414 => x"a8",
          1415 => x"74",
          1416 => x"74",
          1417 => x"78",
          1418 => x"11",
          1419 => x"81",
          1420 => x"06",
          1421 => x"ff",
          1422 => x"52",
          1423 => x"55",
          1424 => x"38",
          1425 => x"8c",
          1426 => x"0d",
          1427 => x"0d",
          1428 => x"7a",
          1429 => x"9f",
          1430 => x"7c",
          1431 => x"32",
          1432 => x"71",
          1433 => x"72",
          1434 => x"59",
          1435 => x"56",
          1436 => x"84",
          1437 => x"75",
          1438 => x"84",
          1439 => x"88",
          1440 => x"f7",
          1441 => x"7d",
          1442 => x"70",
          1443 => x"08",
          1444 => x"56",
          1445 => x"2e",
          1446 => x"8f",
          1447 => x"70",
          1448 => x"33",
          1449 => x"a0",
          1450 => x"73",
          1451 => x"f5",
          1452 => x"2e",
          1453 => x"d0",
          1454 => x"56",
          1455 => x"80",
          1456 => x"58",
          1457 => x"74",
          1458 => x"38",
          1459 => x"27",
          1460 => x"14",
          1461 => x"06",
          1462 => x"14",
          1463 => x"06",
          1464 => x"73",
          1465 => x"f9",
          1466 => x"ff",
          1467 => x"89",
          1468 => x"89",
          1469 => x"27",
          1470 => x"77",
          1471 => x"81",
          1472 => x"0c",
          1473 => x"56",
          1474 => x"26",
          1475 => x"78",
          1476 => x"38",
          1477 => x"75",
          1478 => x"56",
          1479 => x"8c",
          1480 => x"0d",
          1481 => x"16",
          1482 => x"70",
          1483 => x"59",
          1484 => x"09",
          1485 => x"ff",
          1486 => x"70",
          1487 => x"33",
          1488 => x"80",
          1489 => x"38",
          1490 => x"80",
          1491 => x"38",
          1492 => x"74",
          1493 => x"d0",
          1494 => x"56",
          1495 => x"73",
          1496 => x"38",
          1497 => x"8c",
          1498 => x"0d",
          1499 => x"81",
          1500 => x"0c",
          1501 => x"55",
          1502 => x"ca",
          1503 => x"84",
          1504 => x"8b",
          1505 => x"f7",
          1506 => x"7d",
          1507 => x"70",
          1508 => x"08",
          1509 => x"56",
          1510 => x"2e",
          1511 => x"8f",
          1512 => x"70",
          1513 => x"33",
          1514 => x"a0",
          1515 => x"73",
          1516 => x"f5",
          1517 => x"2e",
          1518 => x"d0",
          1519 => x"56",
          1520 => x"80",
          1521 => x"58",
          1522 => x"74",
          1523 => x"38",
          1524 => x"27",
          1525 => x"14",
          1526 => x"06",
          1527 => x"14",
          1528 => x"06",
          1529 => x"73",
          1530 => x"f9",
          1531 => x"ff",
          1532 => x"89",
          1533 => x"89",
          1534 => x"27",
          1535 => x"77",
          1536 => x"81",
          1537 => x"0c",
          1538 => x"56",
          1539 => x"26",
          1540 => x"78",
          1541 => x"38",
          1542 => x"75",
          1543 => x"56",
          1544 => x"8c",
          1545 => x"0d",
          1546 => x"16",
          1547 => x"70",
          1548 => x"59",
          1549 => x"09",
          1550 => x"ff",
          1551 => x"70",
          1552 => x"33",
          1553 => x"80",
          1554 => x"38",
          1555 => x"80",
          1556 => x"38",
          1557 => x"74",
          1558 => x"d0",
          1559 => x"56",
          1560 => x"73",
          1561 => x"38",
          1562 => x"8c",
          1563 => x"0d",
          1564 => x"81",
          1565 => x"0c",
          1566 => x"55",
          1567 => x"ca",
          1568 => x"84",
          1569 => x"8b",
          1570 => x"80",
          1571 => x"84",
          1572 => x"81",
          1573 => x"ba",
          1574 => x"ff",
          1575 => x"52",
          1576 => x"8c",
          1577 => x"10",
          1578 => x"05",
          1579 => x"04",
          1580 => x"51",
          1581 => x"83",
          1582 => x"83",
          1583 => x"ef",
          1584 => x"3d",
          1585 => x"cf",
          1586 => x"a8",
          1587 => x"0d",
          1588 => x"a4",
          1589 => x"3f",
          1590 => x"04",
          1591 => x"51",
          1592 => x"83",
          1593 => x"83",
          1594 => x"ef",
          1595 => x"3d",
          1596 => x"cf",
          1597 => x"fc",
          1598 => x"0d",
          1599 => x"fc",
          1600 => x"3f",
          1601 => x"04",
          1602 => x"51",
          1603 => x"83",
          1604 => x"83",
          1605 => x"ee",
          1606 => x"3d",
          1607 => x"d0",
          1608 => x"d0",
          1609 => x"0d",
          1610 => x"ec",
          1611 => x"3f",
          1612 => x"04",
          1613 => x"51",
          1614 => x"83",
          1615 => x"83",
          1616 => x"ee",
          1617 => x"3d",
          1618 => x"d1",
          1619 => x"a4",
          1620 => x"0d",
          1621 => x"c0",
          1622 => x"3f",
          1623 => x"04",
          1624 => x"51",
          1625 => x"83",
          1626 => x"83",
          1627 => x"ee",
          1628 => x"3d",
          1629 => x"d1",
          1630 => x"f8",
          1631 => x"0d",
          1632 => x"80",
          1633 => x"3f",
          1634 => x"04",
          1635 => x"51",
          1636 => x"83",
          1637 => x"ec",
          1638 => x"02",
          1639 => x"e3",
          1640 => x"58",
          1641 => x"30",
          1642 => x"73",
          1643 => x"57",
          1644 => x"75",
          1645 => x"83",
          1646 => x"74",
          1647 => x"81",
          1648 => x"55",
          1649 => x"80",
          1650 => x"53",
          1651 => x"3d",
          1652 => x"82",
          1653 => x"84",
          1654 => x"57",
          1655 => x"08",
          1656 => x"d0",
          1657 => x"82",
          1658 => x"76",
          1659 => x"07",
          1660 => x"30",
          1661 => x"72",
          1662 => x"57",
          1663 => x"2e",
          1664 => x"c0",
          1665 => x"55",
          1666 => x"26",
          1667 => x"74",
          1668 => x"e8",
          1669 => x"8e",
          1670 => x"8c",
          1671 => x"d2",
          1672 => x"52",
          1673 => x"51",
          1674 => x"76",
          1675 => x"0c",
          1676 => x"04",
          1677 => x"08",
          1678 => x"88",
          1679 => x"8c",
          1680 => x"3d",
          1681 => x"84",
          1682 => x"52",
          1683 => x"9e",
          1684 => x"ba",
          1685 => x"84",
          1686 => x"ff",
          1687 => x"55",
          1688 => x"ff",
          1689 => x"19",
          1690 => x"59",
          1691 => x"e8",
          1692 => x"f4",
          1693 => x"ba",
          1694 => x"78",
          1695 => x"3f",
          1696 => x"08",
          1697 => x"bc",
          1698 => x"83",
          1699 => x"de",
          1700 => x"97",
          1701 => x"0d",
          1702 => x"05",
          1703 => x"58",
          1704 => x"80",
          1705 => x"7a",
          1706 => x"3f",
          1707 => x"08",
          1708 => x"80",
          1709 => x"76",
          1710 => x"38",
          1711 => x"8c",
          1712 => x"0d",
          1713 => x"84",
          1714 => x"61",
          1715 => x"84",
          1716 => x"7f",
          1717 => x"78",
          1718 => x"8c",
          1719 => x"8c",
          1720 => x"0d",
          1721 => x"0d",
          1722 => x"02",
          1723 => x"cf",
          1724 => x"73",
          1725 => x"5f",
          1726 => x"5d",
          1727 => x"2e",
          1728 => x"7a",
          1729 => x"c4",
          1730 => x"3f",
          1731 => x"51",
          1732 => x"80",
          1733 => x"27",
          1734 => x"90",
          1735 => x"38",
          1736 => x"82",
          1737 => x"18",
          1738 => x"27",
          1739 => x"72",
          1740 => x"d2",
          1741 => x"d1",
          1742 => x"84",
          1743 => x"53",
          1744 => x"ec",
          1745 => x"74",
          1746 => x"83",
          1747 => x"dd",
          1748 => x"56",
          1749 => x"80",
          1750 => x"18",
          1751 => x"53",
          1752 => x"7a",
          1753 => x"81",
          1754 => x"9f",
          1755 => x"38",
          1756 => x"73",
          1757 => x"ff",
          1758 => x"74",
          1759 => x"38",
          1760 => x"27",
          1761 => x"84",
          1762 => x"52",
          1763 => x"df",
          1764 => x"56",
          1765 => x"c2",
          1766 => x"dc",
          1767 => x"3f",
          1768 => x"1c",
          1769 => x"51",
          1770 => x"84",
          1771 => x"98",
          1772 => x"2c",
          1773 => x"a0",
          1774 => x"38",
          1775 => x"82",
          1776 => x"1e",
          1777 => x"26",
          1778 => x"ff",
          1779 => x"8c",
          1780 => x"0d",
          1781 => x"e0",
          1782 => x"3f",
          1783 => x"d5",
          1784 => x"54",
          1785 => x"87",
          1786 => x"26",
          1787 => x"fe",
          1788 => x"d2",
          1789 => x"91",
          1790 => x"84",
          1791 => x"53",
          1792 => x"ea",
          1793 => x"79",
          1794 => x"38",
          1795 => x"72",
          1796 => x"38",
          1797 => x"83",
          1798 => x"db",
          1799 => x"14",
          1800 => x"08",
          1801 => x"51",
          1802 => x"78",
          1803 => x"38",
          1804 => x"83",
          1805 => x"db",
          1806 => x"14",
          1807 => x"08",
          1808 => x"51",
          1809 => x"73",
          1810 => x"ff",
          1811 => x"53",
          1812 => x"df",
          1813 => x"52",
          1814 => x"51",
          1815 => x"84",
          1816 => x"f0",
          1817 => x"a0",
          1818 => x"3f",
          1819 => x"dd",
          1820 => x"39",
          1821 => x"08",
          1822 => x"e9",
          1823 => x"16",
          1824 => x"39",
          1825 => x"3f",
          1826 => x"08",
          1827 => x"53",
          1828 => x"a8",
          1829 => x"38",
          1830 => x"80",
          1831 => x"81",
          1832 => x"38",
          1833 => x"db",
          1834 => x"9b",
          1835 => x"ba",
          1836 => x"2b",
          1837 => x"70",
          1838 => x"30",
          1839 => x"70",
          1840 => x"07",
          1841 => x"06",
          1842 => x"59",
          1843 => x"72",
          1844 => x"e8",
          1845 => x"9b",
          1846 => x"ba",
          1847 => x"2b",
          1848 => x"70",
          1849 => x"30",
          1850 => x"70",
          1851 => x"07",
          1852 => x"06",
          1853 => x"59",
          1854 => x"80",
          1855 => x"a9",
          1856 => x"39",
          1857 => x"ba",
          1858 => x"3d",
          1859 => x"3d",
          1860 => x"96",
          1861 => x"aa",
          1862 => x"51",
          1863 => x"83",
          1864 => x"9d",
          1865 => x"51",
          1866 => x"72",
          1867 => x"81",
          1868 => x"71",
          1869 => x"72",
          1870 => x"81",
          1871 => x"71",
          1872 => x"72",
          1873 => x"81",
          1874 => x"71",
          1875 => x"72",
          1876 => x"81",
          1877 => x"71",
          1878 => x"72",
          1879 => x"81",
          1880 => x"71",
          1881 => x"72",
          1882 => x"81",
          1883 => x"71",
          1884 => x"72",
          1885 => x"81",
          1886 => x"71",
          1887 => x"88",
          1888 => x"53",
          1889 => x"a9",
          1890 => x"3d",
          1891 => x"51",
          1892 => x"83",
          1893 => x"9c",
          1894 => x"51",
          1895 => x"a9",
          1896 => x"3d",
          1897 => x"51",
          1898 => x"83",
          1899 => x"9b",
          1900 => x"51",
          1901 => x"72",
          1902 => x"06",
          1903 => x"2e",
          1904 => x"39",
          1905 => x"cd",
          1906 => x"f4",
          1907 => x"3f",
          1908 => x"c1",
          1909 => x"2a",
          1910 => x"51",
          1911 => x"2e",
          1912 => x"c2",
          1913 => x"9b",
          1914 => x"d4",
          1915 => x"bd",
          1916 => x"9b",
          1917 => x"86",
          1918 => x"06",
          1919 => x"80",
          1920 => x"38",
          1921 => x"81",
          1922 => x"3f",
          1923 => x"51",
          1924 => x"80",
          1925 => x"3f",
          1926 => x"70",
          1927 => x"52",
          1928 => x"fe",
          1929 => x"bd",
          1930 => x"9a",
          1931 => x"d4",
          1932 => x"f9",
          1933 => x"9a",
          1934 => x"84",
          1935 => x"06",
          1936 => x"80",
          1937 => x"38",
          1938 => x"81",
          1939 => x"3f",
          1940 => x"51",
          1941 => x"80",
          1942 => x"3f",
          1943 => x"70",
          1944 => x"52",
          1945 => x"fd",
          1946 => x"bd",
          1947 => x"9a",
          1948 => x"d4",
          1949 => x"b5",
          1950 => x"9a",
          1951 => x"82",
          1952 => x"06",
          1953 => x"80",
          1954 => x"38",
          1955 => x"ca",
          1956 => x"70",
          1957 => x"61",
          1958 => x"0c",
          1959 => x"60",
          1960 => x"d5",
          1961 => x"8c",
          1962 => x"06",
          1963 => x"59",
          1964 => x"84",
          1965 => x"d5",
          1966 => x"b8",
          1967 => x"43",
          1968 => x"51",
          1969 => x"7e",
          1970 => x"53",
          1971 => x"51",
          1972 => x"0b",
          1973 => x"80",
          1974 => x"ff",
          1975 => x"79",
          1976 => x"f1",
          1977 => x"2e",
          1978 => x"78",
          1979 => x"5e",
          1980 => x"83",
          1981 => x"70",
          1982 => x"80",
          1983 => x"38",
          1984 => x"7b",
          1985 => x"81",
          1986 => x"81",
          1987 => x"5d",
          1988 => x"2e",
          1989 => x"5c",
          1990 => x"be",
          1991 => x"29",
          1992 => x"05",
          1993 => x"5b",
          1994 => x"84",
          1995 => x"84",
          1996 => x"54",
          1997 => x"08",
          1998 => x"da",
          1999 => x"8c",
          2000 => x"84",
          2001 => x"7d",
          2002 => x"80",
          2003 => x"70",
          2004 => x"5d",
          2005 => x"27",
          2006 => x"3d",
          2007 => x"80",
          2008 => x"38",
          2009 => x"7e",
          2010 => x"3f",
          2011 => x"08",
          2012 => x"8c",
          2013 => x"8d",
          2014 => x"ba",
          2015 => x"b8",
          2016 => x"05",
          2017 => x"3f",
          2018 => x"08",
          2019 => x"5c",
          2020 => x"2e",
          2021 => x"84",
          2022 => x"51",
          2023 => x"84",
          2024 => x"8f",
          2025 => x"38",
          2026 => x"3d",
          2027 => x"82",
          2028 => x"38",
          2029 => x"8c",
          2030 => x"81",
          2031 => x"38",
          2032 => x"53",
          2033 => x"52",
          2034 => x"dd",
          2035 => x"c8",
          2036 => x"bc",
          2037 => x"67",
          2038 => x"90",
          2039 => x"90",
          2040 => x"7c",
          2041 => x"3f",
          2042 => x"08",
          2043 => x"08",
          2044 => x"70",
          2045 => x"25",
          2046 => x"42",
          2047 => x"83",
          2048 => x"81",
          2049 => x"06",
          2050 => x"2e",
          2051 => x"1b",
          2052 => x"06",
          2053 => x"ff",
          2054 => x"81",
          2055 => x"32",
          2056 => x"81",
          2057 => x"ff",
          2058 => x"38",
          2059 => x"95",
          2060 => x"d5",
          2061 => x"d1",
          2062 => x"80",
          2063 => x"52",
          2064 => x"bc",
          2065 => x"83",
          2066 => x"70",
          2067 => x"5b",
          2068 => x"91",
          2069 => x"83",
          2070 => x"84",
          2071 => x"82",
          2072 => x"84",
          2073 => x"80",
          2074 => x"0b",
          2075 => x"ef",
          2076 => x"d1",
          2077 => x"f8",
          2078 => x"82",
          2079 => x"84",
          2080 => x"80",
          2081 => x"84",
          2082 => x"51",
          2083 => x"0b",
          2084 => x"80",
          2085 => x"ff",
          2086 => x"7d",
          2087 => x"81",
          2088 => x"38",
          2089 => x"d1",
          2090 => x"a2",
          2091 => x"0b",
          2092 => x"ef",
          2093 => x"d5",
          2094 => x"f8",
          2095 => x"a7",
          2096 => x"70",
          2097 => x"fc",
          2098 => x"39",
          2099 => x"0c",
          2100 => x"59",
          2101 => x"26",
          2102 => x"78",
          2103 => x"bf",
          2104 => x"79",
          2105 => x"d5",
          2106 => x"88",
          2107 => x"5f",
          2108 => x"d6",
          2109 => x"51",
          2110 => x"60",
          2111 => x"84",
          2112 => x"82",
          2113 => x"84",
          2114 => x"61",
          2115 => x"06",
          2116 => x"81",
          2117 => x"45",
          2118 => x"a4",
          2119 => x"84",
          2120 => x"3f",
          2121 => x"93",
          2122 => x"86",
          2123 => x"94",
          2124 => x"83",
          2125 => x"80",
          2126 => x"9c",
          2127 => x"d2",
          2128 => x"89",
          2129 => x"e3",
          2130 => x"39",
          2131 => x"fa",
          2132 => x"52",
          2133 => x"94",
          2134 => x"39",
          2135 => x"3f",
          2136 => x"83",
          2137 => x"de",
          2138 => x"59",
          2139 => x"d6",
          2140 => x"80",
          2141 => x"3f",
          2142 => x"b8",
          2143 => x"11",
          2144 => x"05",
          2145 => x"3f",
          2146 => x"08",
          2147 => x"b0",
          2148 => x"83",
          2149 => x"d0",
          2150 => x"5a",
          2151 => x"ba",
          2152 => x"2e",
          2153 => x"84",
          2154 => x"52",
          2155 => x"51",
          2156 => x"fa",
          2157 => x"3d",
          2158 => x"53",
          2159 => x"51",
          2160 => x"84",
          2161 => x"80",
          2162 => x"38",
          2163 => x"d7",
          2164 => x"b5",
          2165 => x"78",
          2166 => x"fe",
          2167 => x"ff",
          2168 => x"e9",
          2169 => x"ba",
          2170 => x"2e",
          2171 => x"b8",
          2172 => x"11",
          2173 => x"05",
          2174 => x"3f",
          2175 => x"08",
          2176 => x"64",
          2177 => x"53",
          2178 => x"d7",
          2179 => x"f9",
          2180 => x"ec",
          2181 => x"f8",
          2182 => x"d0",
          2183 => x"48",
          2184 => x"78",
          2185 => x"98",
          2186 => x"26",
          2187 => x"64",
          2188 => x"46",
          2189 => x"b8",
          2190 => x"11",
          2191 => x"05",
          2192 => x"3f",
          2193 => x"08",
          2194 => x"f4",
          2195 => x"fe",
          2196 => x"ff",
          2197 => x"e8",
          2198 => x"ba",
          2199 => x"b0",
          2200 => x"78",
          2201 => x"52",
          2202 => x"51",
          2203 => x"84",
          2204 => x"53",
          2205 => x"7e",
          2206 => x"3f",
          2207 => x"33",
          2208 => x"2e",
          2209 => x"78",
          2210 => x"ca",
          2211 => x"05",
          2212 => x"cf",
          2213 => x"ff",
          2214 => x"ff",
          2215 => x"e9",
          2216 => x"ba",
          2217 => x"2e",
          2218 => x"b8",
          2219 => x"11",
          2220 => x"05",
          2221 => x"3f",
          2222 => x"08",
          2223 => x"80",
          2224 => x"fe",
          2225 => x"ff",
          2226 => x"e9",
          2227 => x"ba",
          2228 => x"2e",
          2229 => x"83",
          2230 => x"ce",
          2231 => x"67",
          2232 => x"7c",
          2233 => x"38",
          2234 => x"7a",
          2235 => x"5a",
          2236 => x"95",
          2237 => x"79",
          2238 => x"53",
          2239 => x"d7",
          2240 => x"85",
          2241 => x"5b",
          2242 => x"81",
          2243 => x"d2",
          2244 => x"ff",
          2245 => x"ff",
          2246 => x"e8",
          2247 => x"ba",
          2248 => x"2e",
          2249 => x"b8",
          2250 => x"11",
          2251 => x"05",
          2252 => x"3f",
          2253 => x"08",
          2254 => x"84",
          2255 => x"fe",
          2256 => x"ff",
          2257 => x"e8",
          2258 => x"ba",
          2259 => x"2e",
          2260 => x"83",
          2261 => x"cd",
          2262 => x"5a",
          2263 => x"82",
          2264 => x"5c",
          2265 => x"05",
          2266 => x"34",
          2267 => x"46",
          2268 => x"3d",
          2269 => x"53",
          2270 => x"51",
          2271 => x"84",
          2272 => x"80",
          2273 => x"38",
          2274 => x"fc",
          2275 => x"80",
          2276 => x"f3",
          2277 => x"8c",
          2278 => x"68",
          2279 => x"52",
          2280 => x"51",
          2281 => x"84",
          2282 => x"53",
          2283 => x"7e",
          2284 => x"3f",
          2285 => x"33",
          2286 => x"2e",
          2287 => x"78",
          2288 => x"97",
          2289 => x"05",
          2290 => x"68",
          2291 => x"db",
          2292 => x"34",
          2293 => x"49",
          2294 => x"fc",
          2295 => x"80",
          2296 => x"a3",
          2297 => x"8c",
          2298 => x"f5",
          2299 => x"59",
          2300 => x"05",
          2301 => x"68",
          2302 => x"b8",
          2303 => x"11",
          2304 => x"05",
          2305 => x"3f",
          2306 => x"08",
          2307 => x"f5",
          2308 => x"3d",
          2309 => x"53",
          2310 => x"51",
          2311 => x"84",
          2312 => x"80",
          2313 => x"38",
          2314 => x"fc",
          2315 => x"80",
          2316 => x"d3",
          2317 => x"8c",
          2318 => x"f5",
          2319 => x"3d",
          2320 => x"53",
          2321 => x"51",
          2322 => x"84",
          2323 => x"86",
          2324 => x"8c",
          2325 => x"d8",
          2326 => x"ad",
          2327 => x"5b",
          2328 => x"27",
          2329 => x"5b",
          2330 => x"84",
          2331 => x"79",
          2332 => x"38",
          2333 => x"e7",
          2334 => x"39",
          2335 => x"80",
          2336 => x"96",
          2337 => x"8c",
          2338 => x"ff",
          2339 => x"59",
          2340 => x"81",
          2341 => x"8c",
          2342 => x"51",
          2343 => x"84",
          2344 => x"80",
          2345 => x"38",
          2346 => x"08",
          2347 => x"3f",
          2348 => x"b8",
          2349 => x"11",
          2350 => x"05",
          2351 => x"3f",
          2352 => x"08",
          2353 => x"f3",
          2354 => x"79",
          2355 => x"c0",
          2356 => x"c8",
          2357 => x"3d",
          2358 => x"53",
          2359 => x"51",
          2360 => x"84",
          2361 => x"91",
          2362 => x"90",
          2363 => x"80",
          2364 => x"38",
          2365 => x"08",
          2366 => x"fe",
          2367 => x"ff",
          2368 => x"e5",
          2369 => x"ba",
          2370 => x"2e",
          2371 => x"66",
          2372 => x"88",
          2373 => x"81",
          2374 => x"32",
          2375 => x"72",
          2376 => x"7e",
          2377 => x"5d",
          2378 => x"88",
          2379 => x"2e",
          2380 => x"46",
          2381 => x"51",
          2382 => x"80",
          2383 => x"65",
          2384 => x"68",
          2385 => x"3f",
          2386 => x"51",
          2387 => x"f2",
          2388 => x"64",
          2389 => x"64",
          2390 => x"b8",
          2391 => x"11",
          2392 => x"05",
          2393 => x"3f",
          2394 => x"08",
          2395 => x"d0",
          2396 => x"71",
          2397 => x"84",
          2398 => x"3d",
          2399 => x"53",
          2400 => x"51",
          2401 => x"84",
          2402 => x"c6",
          2403 => x"39",
          2404 => x"80",
          2405 => x"7e",
          2406 => x"40",
          2407 => x"b8",
          2408 => x"11",
          2409 => x"05",
          2410 => x"3f",
          2411 => x"08",
          2412 => x"8c",
          2413 => x"02",
          2414 => x"22",
          2415 => x"05",
          2416 => x"45",
          2417 => x"f0",
          2418 => x"80",
          2419 => x"b3",
          2420 => x"8c",
          2421 => x"38",
          2422 => x"b8",
          2423 => x"11",
          2424 => x"05",
          2425 => x"3f",
          2426 => x"08",
          2427 => x"dc",
          2428 => x"02",
          2429 => x"33",
          2430 => x"81",
          2431 => x"9b",
          2432 => x"fe",
          2433 => x"ff",
          2434 => x"e0",
          2435 => x"ba",
          2436 => x"2e",
          2437 => x"64",
          2438 => x"5d",
          2439 => x"70",
          2440 => x"e1",
          2441 => x"2e",
          2442 => x"f3",
          2443 => x"55",
          2444 => x"54",
          2445 => x"d8",
          2446 => x"51",
          2447 => x"f3",
          2448 => x"52",
          2449 => x"80",
          2450 => x"39",
          2451 => x"51",
          2452 => x"f0",
          2453 => x"3d",
          2454 => x"53",
          2455 => x"51",
          2456 => x"84",
          2457 => x"80",
          2458 => x"64",
          2459 => x"ce",
          2460 => x"70",
          2461 => x"23",
          2462 => x"e7",
          2463 => x"91",
          2464 => x"80",
          2465 => x"38",
          2466 => x"08",
          2467 => x"39",
          2468 => x"33",
          2469 => x"2e",
          2470 => x"f2",
          2471 => x"fc",
          2472 => x"d8",
          2473 => x"cc",
          2474 => x"f7",
          2475 => x"d8",
          2476 => x"c0",
          2477 => x"f6",
          2478 => x"f3",
          2479 => x"78",
          2480 => x"38",
          2481 => x"08",
          2482 => x"39",
          2483 => x"51",
          2484 => x"f9",
          2485 => x"f3",
          2486 => x"78",
          2487 => x"38",
          2488 => x"08",
          2489 => x"39",
          2490 => x"33",
          2491 => x"2e",
          2492 => x"f2",
          2493 => x"fb",
          2494 => x"f3",
          2495 => x"7d",
          2496 => x"38",
          2497 => x"08",
          2498 => x"39",
          2499 => x"33",
          2500 => x"2e",
          2501 => x"f2",
          2502 => x"fb",
          2503 => x"f3",
          2504 => x"7c",
          2505 => x"38",
          2506 => x"08",
          2507 => x"39",
          2508 => x"08",
          2509 => x"49",
          2510 => x"83",
          2511 => x"88",
          2512 => x"b5",
          2513 => x"0d",
          2514 => x"ba",
          2515 => x"c0",
          2516 => x"08",
          2517 => x"84",
          2518 => x"51",
          2519 => x"84",
          2520 => x"90",
          2521 => x"57",
          2522 => x"80",
          2523 => x"da",
          2524 => x"84",
          2525 => x"07",
          2526 => x"c0",
          2527 => x"08",
          2528 => x"84",
          2529 => x"51",
          2530 => x"84",
          2531 => x"90",
          2532 => x"57",
          2533 => x"80",
          2534 => x"da",
          2535 => x"84",
          2536 => x"07",
          2537 => x"80",
          2538 => x"c0",
          2539 => x"8c",
          2540 => x"87",
          2541 => x"0c",
          2542 => x"5c",
          2543 => x"5d",
          2544 => x"05",
          2545 => x"80",
          2546 => x"ec",
          2547 => x"70",
          2548 => x"70",
          2549 => x"d5",
          2550 => x"b6",
          2551 => x"83",
          2552 => x"3f",
          2553 => x"94",
          2554 => x"d2",
          2555 => x"d2",
          2556 => x"95",
          2557 => x"fc",
          2558 => x"55",
          2559 => x"83",
          2560 => x"83",
          2561 => x"81",
          2562 => x"83",
          2563 => x"c3",
          2564 => x"97",
          2565 => x"3f",
          2566 => x"3d",
          2567 => x"08",
          2568 => x"75",
          2569 => x"73",
          2570 => x"38",
          2571 => x"81",
          2572 => x"52",
          2573 => x"09",
          2574 => x"38",
          2575 => x"33",
          2576 => x"06",
          2577 => x"70",
          2578 => x"38",
          2579 => x"06",
          2580 => x"2e",
          2581 => x"74",
          2582 => x"2e",
          2583 => x"80",
          2584 => x"81",
          2585 => x"54",
          2586 => x"2e",
          2587 => x"54",
          2588 => x"8b",
          2589 => x"2e",
          2590 => x"12",
          2591 => x"80",
          2592 => x"06",
          2593 => x"a0",
          2594 => x"06",
          2595 => x"54",
          2596 => x"70",
          2597 => x"25",
          2598 => x"52",
          2599 => x"2e",
          2600 => x"72",
          2601 => x"54",
          2602 => x"0c",
          2603 => x"84",
          2604 => x"87",
          2605 => x"70",
          2606 => x"38",
          2607 => x"ff",
          2608 => x"12",
          2609 => x"33",
          2610 => x"06",
          2611 => x"70",
          2612 => x"38",
          2613 => x"39",
          2614 => x"81",
          2615 => x"72",
          2616 => x"81",
          2617 => x"38",
          2618 => x"3d",
          2619 => x"72",
          2620 => x"80",
          2621 => x"8c",
          2622 => x"0d",
          2623 => x"fc",
          2624 => x"51",
          2625 => x"84",
          2626 => x"80",
          2627 => x"74",
          2628 => x"0c",
          2629 => x"04",
          2630 => x"76",
          2631 => x"ff",
          2632 => x"81",
          2633 => x"26",
          2634 => x"83",
          2635 => x"05",
          2636 => x"73",
          2637 => x"8a",
          2638 => x"33",
          2639 => x"70",
          2640 => x"fe",
          2641 => x"33",
          2642 => x"73",
          2643 => x"f2",
          2644 => x"33",
          2645 => x"74",
          2646 => x"e6",
          2647 => x"22",
          2648 => x"74",
          2649 => x"80",
          2650 => x"13",
          2651 => x"52",
          2652 => x"26",
          2653 => x"81",
          2654 => x"98",
          2655 => x"22",
          2656 => x"bc",
          2657 => x"33",
          2658 => x"b8",
          2659 => x"33",
          2660 => x"b4",
          2661 => x"33",
          2662 => x"b0",
          2663 => x"33",
          2664 => x"ac",
          2665 => x"33",
          2666 => x"a8",
          2667 => x"c0",
          2668 => x"73",
          2669 => x"a0",
          2670 => x"87",
          2671 => x"0c",
          2672 => x"84",
          2673 => x"86",
          2674 => x"f3",
          2675 => x"5b",
          2676 => x"9c",
          2677 => x"0c",
          2678 => x"bc",
          2679 => x"7b",
          2680 => x"98",
          2681 => x"7b",
          2682 => x"87",
          2683 => x"08",
          2684 => x"1c",
          2685 => x"98",
          2686 => x"7b",
          2687 => x"87",
          2688 => x"08",
          2689 => x"1c",
          2690 => x"98",
          2691 => x"7b",
          2692 => x"87",
          2693 => x"08",
          2694 => x"1c",
          2695 => x"98",
          2696 => x"79",
          2697 => x"80",
          2698 => x"83",
          2699 => x"59",
          2700 => x"ff",
          2701 => x"1b",
          2702 => x"1b",
          2703 => x"1b",
          2704 => x"1b",
          2705 => x"1b",
          2706 => x"83",
          2707 => x"52",
          2708 => x"51",
          2709 => x"3f",
          2710 => x"04",
          2711 => x"02",
          2712 => x"53",
          2713 => x"a8",
          2714 => x"80",
          2715 => x"84",
          2716 => x"98",
          2717 => x"2c",
          2718 => x"ff",
          2719 => x"06",
          2720 => x"83",
          2721 => x"71",
          2722 => x"0c",
          2723 => x"04",
          2724 => x"e8",
          2725 => x"ba",
          2726 => x"2b",
          2727 => x"51",
          2728 => x"2e",
          2729 => x"df",
          2730 => x"80",
          2731 => x"84",
          2732 => x"98",
          2733 => x"2c",
          2734 => x"ff",
          2735 => x"c7",
          2736 => x"0d",
          2737 => x"52",
          2738 => x"54",
          2739 => x"e7",
          2740 => x"ba",
          2741 => x"2b",
          2742 => x"51",
          2743 => x"2e",
          2744 => x"72",
          2745 => x"54",
          2746 => x"25",
          2747 => x"84",
          2748 => x"85",
          2749 => x"fc",
          2750 => x"9b",
          2751 => x"f2",
          2752 => x"81",
          2753 => x"55",
          2754 => x"2e",
          2755 => x"87",
          2756 => x"08",
          2757 => x"70",
          2758 => x"54",
          2759 => x"2e",
          2760 => x"91",
          2761 => x"06",
          2762 => x"e3",
          2763 => x"32",
          2764 => x"72",
          2765 => x"38",
          2766 => x"81",
          2767 => x"cf",
          2768 => x"ff",
          2769 => x"c0",
          2770 => x"70",
          2771 => x"38",
          2772 => x"90",
          2773 => x"0c",
          2774 => x"8c",
          2775 => x"0d",
          2776 => x"2a",
          2777 => x"51",
          2778 => x"38",
          2779 => x"81",
          2780 => x"80",
          2781 => x"71",
          2782 => x"06",
          2783 => x"2e",
          2784 => x"c0",
          2785 => x"70",
          2786 => x"81",
          2787 => x"52",
          2788 => x"d8",
          2789 => x"0d",
          2790 => x"33",
          2791 => x"9f",
          2792 => x"52",
          2793 => x"c4",
          2794 => x"0d",
          2795 => x"0d",
          2796 => x"75",
          2797 => x"52",
          2798 => x"2e",
          2799 => x"81",
          2800 => x"c4",
          2801 => x"ff",
          2802 => x"55",
          2803 => x"80",
          2804 => x"c0",
          2805 => x"70",
          2806 => x"81",
          2807 => x"52",
          2808 => x"8c",
          2809 => x"2a",
          2810 => x"51",
          2811 => x"38",
          2812 => x"81",
          2813 => x"80",
          2814 => x"71",
          2815 => x"06",
          2816 => x"38",
          2817 => x"06",
          2818 => x"94",
          2819 => x"80",
          2820 => x"87",
          2821 => x"52",
          2822 => x"81",
          2823 => x"55",
          2824 => x"9b",
          2825 => x"ba",
          2826 => x"3d",
          2827 => x"91",
          2828 => x"06",
          2829 => x"98",
          2830 => x"32",
          2831 => x"72",
          2832 => x"38",
          2833 => x"81",
          2834 => x"80",
          2835 => x"38",
          2836 => x"84",
          2837 => x"2a",
          2838 => x"53",
          2839 => x"ce",
          2840 => x"ff",
          2841 => x"c0",
          2842 => x"70",
          2843 => x"06",
          2844 => x"80",
          2845 => x"38",
          2846 => x"a4",
          2847 => x"c8",
          2848 => x"9e",
          2849 => x"f2",
          2850 => x"c0",
          2851 => x"83",
          2852 => x"87",
          2853 => x"08",
          2854 => x"0c",
          2855 => x"9c",
          2856 => x"d8",
          2857 => x"9e",
          2858 => x"f2",
          2859 => x"c0",
          2860 => x"83",
          2861 => x"87",
          2862 => x"08",
          2863 => x"0c",
          2864 => x"b4",
          2865 => x"e8",
          2866 => x"9e",
          2867 => x"f2",
          2868 => x"c0",
          2869 => x"83",
          2870 => x"87",
          2871 => x"08",
          2872 => x"0c",
          2873 => x"c4",
          2874 => x"f8",
          2875 => x"9e",
          2876 => x"71",
          2877 => x"23",
          2878 => x"84",
          2879 => x"80",
          2880 => x"9e",
          2881 => x"f3",
          2882 => x"c0",
          2883 => x"83",
          2884 => x"81",
          2885 => x"8c",
          2886 => x"87",
          2887 => x"08",
          2888 => x"0a",
          2889 => x"52",
          2890 => x"38",
          2891 => x"8d",
          2892 => x"87",
          2893 => x"08",
          2894 => x"0a",
          2895 => x"52",
          2896 => x"83",
          2897 => x"71",
          2898 => x"34",
          2899 => x"c0",
          2900 => x"70",
          2901 => x"06",
          2902 => x"70",
          2903 => x"38",
          2904 => x"83",
          2905 => x"80",
          2906 => x"9e",
          2907 => x"88",
          2908 => x"51",
          2909 => x"80",
          2910 => x"81",
          2911 => x"f3",
          2912 => x"0b",
          2913 => x"90",
          2914 => x"80",
          2915 => x"52",
          2916 => x"2e",
          2917 => x"52",
          2918 => x"91",
          2919 => x"87",
          2920 => x"08",
          2921 => x"80",
          2922 => x"52",
          2923 => x"83",
          2924 => x"71",
          2925 => x"34",
          2926 => x"c0",
          2927 => x"70",
          2928 => x"06",
          2929 => x"70",
          2930 => x"38",
          2931 => x"83",
          2932 => x"80",
          2933 => x"9e",
          2934 => x"82",
          2935 => x"51",
          2936 => x"80",
          2937 => x"81",
          2938 => x"f3",
          2939 => x"0b",
          2940 => x"90",
          2941 => x"80",
          2942 => x"52",
          2943 => x"2e",
          2944 => x"52",
          2945 => x"95",
          2946 => x"87",
          2947 => x"08",
          2948 => x"80",
          2949 => x"52",
          2950 => x"83",
          2951 => x"71",
          2952 => x"34",
          2953 => x"c0",
          2954 => x"70",
          2955 => x"51",
          2956 => x"80",
          2957 => x"81",
          2958 => x"f3",
          2959 => x"c0",
          2960 => x"98",
          2961 => x"8a",
          2962 => x"71",
          2963 => x"34",
          2964 => x"c0",
          2965 => x"70",
          2966 => x"51",
          2967 => x"80",
          2968 => x"81",
          2969 => x"f3",
          2970 => x"c0",
          2971 => x"83",
          2972 => x"84",
          2973 => x"71",
          2974 => x"34",
          2975 => x"c0",
          2976 => x"70",
          2977 => x"52",
          2978 => x"2e",
          2979 => x"52",
          2980 => x"9b",
          2981 => x"9e",
          2982 => x"06",
          2983 => x"f3",
          2984 => x"3d",
          2985 => x"52",
          2986 => x"fb",
          2987 => x"d9",
          2988 => x"b6",
          2989 => x"f3",
          2990 => x"73",
          2991 => x"83",
          2992 => x"c3",
          2993 => x"f3",
          2994 => x"74",
          2995 => x"83",
          2996 => x"54",
          2997 => x"38",
          2998 => x"33",
          2999 => x"a8",
          3000 => x"91",
          3001 => x"84",
          3002 => x"f3",
          3003 => x"73",
          3004 => x"83",
          3005 => x"56",
          3006 => x"38",
          3007 => x"33",
          3008 => x"90",
          3009 => x"99",
          3010 => x"83",
          3011 => x"f3",
          3012 => x"75",
          3013 => x"83",
          3014 => x"54",
          3015 => x"38",
          3016 => x"33",
          3017 => x"93",
          3018 => x"95",
          3019 => x"82",
          3020 => x"f3",
          3021 => x"73",
          3022 => x"83",
          3023 => x"c2",
          3024 => x"f2",
          3025 => x"83",
          3026 => x"ff",
          3027 => x"83",
          3028 => x"52",
          3029 => x"51",
          3030 => x"3f",
          3031 => x"08",
          3032 => x"94",
          3033 => x"a1",
          3034 => x"bc",
          3035 => x"3f",
          3036 => x"22",
          3037 => x"c4",
          3038 => x"8d",
          3039 => x"80",
          3040 => x"84",
          3041 => x"51",
          3042 => x"84",
          3043 => x"bd",
          3044 => x"76",
          3045 => x"54",
          3046 => x"08",
          3047 => x"ec",
          3048 => x"e5",
          3049 => x"93",
          3050 => x"80",
          3051 => x"f3",
          3052 => x"74",
          3053 => x"51",
          3054 => x"87",
          3055 => x"83",
          3056 => x"56",
          3057 => x"52",
          3058 => x"da",
          3059 => x"8c",
          3060 => x"c0",
          3061 => x"31",
          3062 => x"ba",
          3063 => x"83",
          3064 => x"ff",
          3065 => x"8a",
          3066 => x"3f",
          3067 => x"04",
          3068 => x"08",
          3069 => x"c0",
          3070 => x"c9",
          3071 => x"ba",
          3072 => x"84",
          3073 => x"71",
          3074 => x"84",
          3075 => x"52",
          3076 => x"51",
          3077 => x"3f",
          3078 => x"33",
          3079 => x"2e",
          3080 => x"ff",
          3081 => x"db",
          3082 => x"c8",
          3083 => x"b8",
          3084 => x"3f",
          3085 => x"08",
          3086 => x"c4",
          3087 => x"c9",
          3088 => x"f4",
          3089 => x"d9",
          3090 => x"b3",
          3091 => x"f2",
          3092 => x"83",
          3093 => x"ff",
          3094 => x"83",
          3095 => x"c0",
          3096 => x"f2",
          3097 => x"83",
          3098 => x"ff",
          3099 => x"83",
          3100 => x"56",
          3101 => x"52",
          3102 => x"aa",
          3103 => x"8c",
          3104 => x"c0",
          3105 => x"31",
          3106 => x"ba",
          3107 => x"83",
          3108 => x"ff",
          3109 => x"83",
          3110 => x"55",
          3111 => x"fe",
          3112 => x"cc",
          3113 => x"f8",
          3114 => x"c8",
          3115 => x"96",
          3116 => x"80",
          3117 => x"38",
          3118 => x"83",
          3119 => x"ff",
          3120 => x"83",
          3121 => x"56",
          3122 => x"fc",
          3123 => x"39",
          3124 => x"51",
          3125 => x"3f",
          3126 => x"33",
          3127 => x"2e",
          3128 => x"d7",
          3129 => x"98",
          3130 => x"88",
          3131 => x"8f",
          3132 => x"80",
          3133 => x"38",
          3134 => x"f3",
          3135 => x"83",
          3136 => x"ff",
          3137 => x"83",
          3138 => x"56",
          3139 => x"fc",
          3140 => x"39",
          3141 => x"33",
          3142 => x"cc",
          3143 => x"e9",
          3144 => x"99",
          3145 => x"80",
          3146 => x"38",
          3147 => x"f3",
          3148 => x"83",
          3149 => x"ff",
          3150 => x"83",
          3151 => x"54",
          3152 => x"fb",
          3153 => x"39",
          3154 => x"08",
          3155 => x"08",
          3156 => x"83",
          3157 => x"ff",
          3158 => x"83",
          3159 => x"56",
          3160 => x"fb",
          3161 => x"39",
          3162 => x"08",
          3163 => x"08",
          3164 => x"83",
          3165 => x"ff",
          3166 => x"83",
          3167 => x"54",
          3168 => x"fa",
          3169 => x"39",
          3170 => x"08",
          3171 => x"08",
          3172 => x"83",
          3173 => x"ff",
          3174 => x"83",
          3175 => x"55",
          3176 => x"fa",
          3177 => x"39",
          3178 => x"08",
          3179 => x"08",
          3180 => x"83",
          3181 => x"ff",
          3182 => x"83",
          3183 => x"56",
          3184 => x"fa",
          3185 => x"39",
          3186 => x"08",
          3187 => x"08",
          3188 => x"83",
          3189 => x"ff",
          3190 => x"83",
          3191 => x"54",
          3192 => x"f9",
          3193 => x"39",
          3194 => x"51",
          3195 => x"3f",
          3196 => x"51",
          3197 => x"3f",
          3198 => x"33",
          3199 => x"2e",
          3200 => x"c4",
          3201 => x"0d",
          3202 => x"33",
          3203 => x"26",
          3204 => x"10",
          3205 => x"c4",
          3206 => x"08",
          3207 => x"ac",
          3208 => x"e5",
          3209 => x"0d",
          3210 => x"b4",
          3211 => x"d9",
          3212 => x"0d",
          3213 => x"bc",
          3214 => x"cd",
          3215 => x"0d",
          3216 => x"c4",
          3217 => x"c1",
          3218 => x"0d",
          3219 => x"cc",
          3220 => x"b5",
          3221 => x"0d",
          3222 => x"d4",
          3223 => x"a9",
          3224 => x"0d",
          3225 => x"80",
          3226 => x"0b",
          3227 => x"84",
          3228 => x"f3",
          3229 => x"c0",
          3230 => x"04",
          3231 => x"aa",
          3232 => x"3d",
          3233 => x"81",
          3234 => x"80",
          3235 => x"f8",
          3236 => x"88",
          3237 => x"ba",
          3238 => x"ed",
          3239 => x"57",
          3240 => x"f3",
          3241 => x"55",
          3242 => x"76",
          3243 => x"df",
          3244 => x"8c",
          3245 => x"a4",
          3246 => x"c0",
          3247 => x"ba",
          3248 => x"17",
          3249 => x"0b",
          3250 => x"08",
          3251 => x"84",
          3252 => x"ff",
          3253 => x"55",
          3254 => x"34",
          3255 => x"30",
          3256 => x"9f",
          3257 => x"55",
          3258 => x"85",
          3259 => x"b0",
          3260 => x"f8",
          3261 => x"08",
          3262 => x"87",
          3263 => x"ba",
          3264 => x"38",
          3265 => x"9a",
          3266 => x"ba",
          3267 => x"3d",
          3268 => x"e2",
          3269 => x"ad",
          3270 => x"76",
          3271 => x"06",
          3272 => x"52",
          3273 => x"a0",
          3274 => x"ff",
          3275 => x"ab",
          3276 => x"84",
          3277 => x"76",
          3278 => x"83",
          3279 => x"ff",
          3280 => x"80",
          3281 => x"8c",
          3282 => x"0d",
          3283 => x"0d",
          3284 => x"ad",
          3285 => x"72",
          3286 => x"57",
          3287 => x"73",
          3288 => x"91",
          3289 => x"8d",
          3290 => x"75",
          3291 => x"83",
          3292 => x"70",
          3293 => x"ff",
          3294 => x"84",
          3295 => x"53",
          3296 => x"08",
          3297 => x"3f",
          3298 => x"08",
          3299 => x"14",
          3300 => x"81",
          3301 => x"38",
          3302 => x"99",
          3303 => x"70",
          3304 => x"57",
          3305 => x"27",
          3306 => x"54",
          3307 => x"8c",
          3308 => x"0d",
          3309 => x"5a",
          3310 => x"84",
          3311 => x"80",
          3312 => x"c3",
          3313 => x"8c",
          3314 => x"d1",
          3315 => x"53",
          3316 => x"51",
          3317 => x"84",
          3318 => x"81",
          3319 => x"73",
          3320 => x"38",
          3321 => x"81",
          3322 => x"54",
          3323 => x"fe",
          3324 => x"b6",
          3325 => x"77",
          3326 => x"76",
          3327 => x"38",
          3328 => x"5b",
          3329 => x"55",
          3330 => x"09",
          3331 => x"d5",
          3332 => x"26",
          3333 => x"0b",
          3334 => x"56",
          3335 => x"73",
          3336 => x"08",
          3337 => x"f8",
          3338 => x"82",
          3339 => x"84",
          3340 => x"80",
          3341 => x"f3",
          3342 => x"80",
          3343 => x"51",
          3344 => x"3f",
          3345 => x"08",
          3346 => x"38",
          3347 => x"bd",
          3348 => x"ba",
          3349 => x"80",
          3350 => x"8c",
          3351 => x"38",
          3352 => x"08",
          3353 => x"19",
          3354 => x"77",
          3355 => x"75",
          3356 => x"83",
          3357 => x"56",
          3358 => x"3f",
          3359 => x"09",
          3360 => x"b2",
          3361 => x"84",
          3362 => x"aa",
          3363 => x"ce",
          3364 => x"3d",
          3365 => x"08",
          3366 => x"5a",
          3367 => x"0b",
          3368 => x"83",
          3369 => x"83",
          3370 => x"56",
          3371 => x"38",
          3372 => x"f4",
          3373 => x"74",
          3374 => x"cb",
          3375 => x"2e",
          3376 => x"81",
          3377 => x"5a",
          3378 => x"a0",
          3379 => x"2e",
          3380 => x"93",
          3381 => x"5f",
          3382 => x"ea",
          3383 => x"ba",
          3384 => x"2b",
          3385 => x"5b",
          3386 => x"2e",
          3387 => x"81",
          3388 => x"d1",
          3389 => x"98",
          3390 => x"2c",
          3391 => x"33",
          3392 => x"70",
          3393 => x"98",
          3394 => x"10",
          3395 => x"d8",
          3396 => x"15",
          3397 => x"53",
          3398 => x"52",
          3399 => x"59",
          3400 => x"79",
          3401 => x"38",
          3402 => x"81",
          3403 => x"81",
          3404 => x"81",
          3405 => x"70",
          3406 => x"55",
          3407 => x"81",
          3408 => x"10",
          3409 => x"2b",
          3410 => x"0b",
          3411 => x"16",
          3412 => x"77",
          3413 => x"38",
          3414 => x"15",
          3415 => x"33",
          3416 => x"75",
          3417 => x"38",
          3418 => x"c2",
          3419 => x"d1",
          3420 => x"57",
          3421 => x"81",
          3422 => x"1b",
          3423 => x"70",
          3424 => x"d1",
          3425 => x"98",
          3426 => x"2c",
          3427 => x"05",
          3428 => x"83",
          3429 => x"33",
          3430 => x"5d",
          3431 => x"57",
          3432 => x"81",
          3433 => x"84",
          3434 => x"fe",
          3435 => x"57",
          3436 => x"38",
          3437 => x"0a",
          3438 => x"0a",
          3439 => x"2c",
          3440 => x"06",
          3441 => x"76",
          3442 => x"c0",
          3443 => x"16",
          3444 => x"51",
          3445 => x"83",
          3446 => x"33",
          3447 => x"61",
          3448 => x"83",
          3449 => x"08",
          3450 => x"42",
          3451 => x"2e",
          3452 => x"76",
          3453 => x"bc",
          3454 => x"39",
          3455 => x"80",
          3456 => x"38",
          3457 => x"81",
          3458 => x"39",
          3459 => x"fe",
          3460 => x"84",
          3461 => x"76",
          3462 => x"34",
          3463 => x"76",
          3464 => x"55",
          3465 => x"fd",
          3466 => x"10",
          3467 => x"dc",
          3468 => x"08",
          3469 => x"e0",
          3470 => x"0c",
          3471 => x"d1",
          3472 => x"0b",
          3473 => x"34",
          3474 => x"d1",
          3475 => x"75",
          3476 => x"85",
          3477 => x"f0",
          3478 => x"51",
          3479 => x"3f",
          3480 => x"33",
          3481 => x"76",
          3482 => x"34",
          3483 => x"84",
          3484 => x"70",
          3485 => x"84",
          3486 => x"5b",
          3487 => x"79",
          3488 => x"38",
          3489 => x"08",
          3490 => x"58",
          3491 => x"d0",
          3492 => x"70",
          3493 => x"ff",
          3494 => x"fc",
          3495 => x"93",
          3496 => x"38",
          3497 => x"83",
          3498 => x"70",
          3499 => x"75",
          3500 => x"75",
          3501 => x"34",
          3502 => x"84",
          3503 => x"84",
          3504 => x"56",
          3505 => x"2e",
          3506 => x"d5",
          3507 => x"88",
          3508 => x"9b",
          3509 => x"f0",
          3510 => x"51",
          3511 => x"3f",
          3512 => x"08",
          3513 => x"ff",
          3514 => x"84",
          3515 => x"ff",
          3516 => x"84",
          3517 => x"7a",
          3518 => x"55",
          3519 => x"7b",
          3520 => x"85",
          3521 => x"d1",
          3522 => x"cd",
          3523 => x"38",
          3524 => x"08",
          3525 => x"9e",
          3526 => x"10",
          3527 => x"05",
          3528 => x"57",
          3529 => x"f9",
          3530 => x"56",
          3531 => x"fb",
          3532 => x"51",
          3533 => x"3f",
          3534 => x"08",
          3535 => x"34",
          3536 => x"08",
          3537 => x"81",
          3538 => x"52",
          3539 => x"b8",
          3540 => x"d1",
          3541 => x"d1",
          3542 => x"56",
          3543 => x"ff",
          3544 => x"d5",
          3545 => x"88",
          3546 => x"83",
          3547 => x"f0",
          3548 => x"51",
          3549 => x"3f",
          3550 => x"08",
          3551 => x"ff",
          3552 => x"84",
          3553 => x"ff",
          3554 => x"84",
          3555 => x"74",
          3556 => x"55",
          3557 => x"d1",
          3558 => x"81",
          3559 => x"d1",
          3560 => x"57",
          3561 => x"27",
          3562 => x"84",
          3563 => x"52",
          3564 => x"76",
          3565 => x"34",
          3566 => x"33",
          3567 => x"b3",
          3568 => x"d1",
          3569 => x"81",
          3570 => x"d1",
          3571 => x"57",
          3572 => x"27",
          3573 => x"84",
          3574 => x"52",
          3575 => x"76",
          3576 => x"34",
          3577 => x"33",
          3578 => x"b3",
          3579 => x"d1",
          3580 => x"81",
          3581 => x"d1",
          3582 => x"57",
          3583 => x"26",
          3584 => x"f9",
          3585 => x"d1",
          3586 => x"d1",
          3587 => x"56",
          3588 => x"f9",
          3589 => x"15",
          3590 => x"d1",
          3591 => x"98",
          3592 => x"2c",
          3593 => x"06",
          3594 => x"60",
          3595 => x"ef",
          3596 => x"f0",
          3597 => x"51",
          3598 => x"3f",
          3599 => x"33",
          3600 => x"70",
          3601 => x"d1",
          3602 => x"57",
          3603 => x"77",
          3604 => x"38",
          3605 => x"08",
          3606 => x"ff",
          3607 => x"74",
          3608 => x"29",
          3609 => x"05",
          3610 => x"84",
          3611 => x"5d",
          3612 => x"7b",
          3613 => x"38",
          3614 => x"08",
          3615 => x"ff",
          3616 => x"74",
          3617 => x"29",
          3618 => x"05",
          3619 => x"84",
          3620 => x"5d",
          3621 => x"75",
          3622 => x"38",
          3623 => x"7b",
          3624 => x"18",
          3625 => x"84",
          3626 => x"52",
          3627 => x"ff",
          3628 => x"75",
          3629 => x"29",
          3630 => x"05",
          3631 => x"84",
          3632 => x"5b",
          3633 => x"79",
          3634 => x"38",
          3635 => x"81",
          3636 => x"34",
          3637 => x"08",
          3638 => x"51",
          3639 => x"3f",
          3640 => x"0a",
          3641 => x"0a",
          3642 => x"2c",
          3643 => x"33",
          3644 => x"78",
          3645 => x"a7",
          3646 => x"39",
          3647 => x"33",
          3648 => x"2e",
          3649 => x"84",
          3650 => x"52",
          3651 => x"b0",
          3652 => x"d1",
          3653 => x"05",
          3654 => x"d1",
          3655 => x"81",
          3656 => x"dd",
          3657 => x"cc",
          3658 => x"5f",
          3659 => x"84",
          3660 => x"52",
          3661 => x"b0",
          3662 => x"d1",
          3663 => x"51",
          3664 => x"84",
          3665 => x"81",
          3666 => x"77",
          3667 => x"84",
          3668 => x"57",
          3669 => x"80",
          3670 => x"f3",
          3671 => x"10",
          3672 => x"a4",
          3673 => x"57",
          3674 => x"8b",
          3675 => x"82",
          3676 => x"06",
          3677 => x"05",
          3678 => x"53",
          3679 => x"e8",
          3680 => x"ba",
          3681 => x"0c",
          3682 => x"33",
          3683 => x"83",
          3684 => x"70",
          3685 => x"41",
          3686 => x"38",
          3687 => x"08",
          3688 => x"2e",
          3689 => x"f3",
          3690 => x"77",
          3691 => x"bc",
          3692 => x"84",
          3693 => x"80",
          3694 => x"cc",
          3695 => x"ba",
          3696 => x"3d",
          3697 => x"d1",
          3698 => x"74",
          3699 => x"38",
          3700 => x"08",
          3701 => x"ff",
          3702 => x"84",
          3703 => x"52",
          3704 => x"af",
          3705 => x"d5",
          3706 => x"88",
          3707 => x"ff",
          3708 => x"d0",
          3709 => x"56",
          3710 => x"d0",
          3711 => x"ff",
          3712 => x"cc",
          3713 => x"b8",
          3714 => x"fd",
          3715 => x"84",
          3716 => x"80",
          3717 => x"cc",
          3718 => x"39",
          3719 => x"80",
          3720 => x"34",
          3721 => x"33",
          3722 => x"2e",
          3723 => x"d5",
          3724 => x"88",
          3725 => x"b7",
          3726 => x"f0",
          3727 => x"51",
          3728 => x"3f",
          3729 => x"08",
          3730 => x"ff",
          3731 => x"84",
          3732 => x"ff",
          3733 => x"84",
          3734 => x"7c",
          3735 => x"55",
          3736 => x"83",
          3737 => x"ff",
          3738 => x"80",
          3739 => x"d0",
          3740 => x"84",
          3741 => x"7b",
          3742 => x"0c",
          3743 => x"04",
          3744 => x"33",
          3745 => x"06",
          3746 => x"80",
          3747 => x"38",
          3748 => x"33",
          3749 => x"78",
          3750 => x"34",
          3751 => x"77",
          3752 => x"34",
          3753 => x"08",
          3754 => x"ff",
          3755 => x"84",
          3756 => x"70",
          3757 => x"98",
          3758 => x"cc",
          3759 => x"5b",
          3760 => x"24",
          3761 => x"84",
          3762 => x"52",
          3763 => x"ad",
          3764 => x"d1",
          3765 => x"98",
          3766 => x"2c",
          3767 => x"33",
          3768 => x"56",
          3769 => x"f3",
          3770 => x"d5",
          3771 => x"88",
          3772 => x"fb",
          3773 => x"80",
          3774 => x"80",
          3775 => x"98",
          3776 => x"cc",
          3777 => x"55",
          3778 => x"f3",
          3779 => x"d5",
          3780 => x"88",
          3781 => x"d7",
          3782 => x"80",
          3783 => x"80",
          3784 => x"98",
          3785 => x"cc",
          3786 => x"55",
          3787 => x"ff",
          3788 => x"a5",
          3789 => x"57",
          3790 => x"77",
          3791 => x"f0",
          3792 => x"33",
          3793 => x"a7",
          3794 => x"80",
          3795 => x"80",
          3796 => x"98",
          3797 => x"cc",
          3798 => x"5b",
          3799 => x"fe",
          3800 => x"16",
          3801 => x"33",
          3802 => x"d5",
          3803 => x"76",
          3804 => x"ab",
          3805 => x"81",
          3806 => x"81",
          3807 => x"70",
          3808 => x"d1",
          3809 => x"57",
          3810 => x"24",
          3811 => x"fe",
          3812 => x"d1",
          3813 => x"81",
          3814 => x"58",
          3815 => x"f2",
          3816 => x"d1",
          3817 => x"76",
          3818 => x"38",
          3819 => x"70",
          3820 => x"41",
          3821 => x"a1",
          3822 => x"5b",
          3823 => x"1c",
          3824 => x"80",
          3825 => x"ff",
          3826 => x"98",
          3827 => x"d0",
          3828 => x"58",
          3829 => x"e1",
          3830 => x"55",
          3831 => x"d0",
          3832 => x"ff",
          3833 => x"5a",
          3834 => x"7a",
          3835 => x"cc",
          3836 => x"60",
          3837 => x"81",
          3838 => x"84",
          3839 => x"75",
          3840 => x"d0",
          3841 => x"80",
          3842 => x"ff",
          3843 => x"98",
          3844 => x"ff",
          3845 => x"5c",
          3846 => x"24",
          3847 => x"77",
          3848 => x"98",
          3849 => x"ff",
          3850 => x"59",
          3851 => x"f1",
          3852 => x"d5",
          3853 => x"88",
          3854 => x"b3",
          3855 => x"80",
          3856 => x"80",
          3857 => x"98",
          3858 => x"cc",
          3859 => x"41",
          3860 => x"f1",
          3861 => x"d5",
          3862 => x"88",
          3863 => x"8f",
          3864 => x"80",
          3865 => x"80",
          3866 => x"98",
          3867 => x"cc",
          3868 => x"41",
          3869 => x"ff",
          3870 => x"dd",
          3871 => x"a4",
          3872 => x"80",
          3873 => x"38",
          3874 => x"ad",
          3875 => x"ba",
          3876 => x"d1",
          3877 => x"ba",
          3878 => x"ff",
          3879 => x"53",
          3880 => x"51",
          3881 => x"3f",
          3882 => x"33",
          3883 => x"33",
          3884 => x"80",
          3885 => x"38",
          3886 => x"08",
          3887 => x"ff",
          3888 => x"84",
          3889 => x"52",
          3890 => x"a9",
          3891 => x"d5",
          3892 => x"88",
          3893 => x"97",
          3894 => x"d0",
          3895 => x"5b",
          3896 => x"d0",
          3897 => x"ff",
          3898 => x"39",
          3899 => x"e1",
          3900 => x"ba",
          3901 => x"f3",
          3902 => x"ba",
          3903 => x"a5",
          3904 => x"f3",
          3905 => x"ef",
          3906 => x"c3",
          3907 => x"f0",
          3908 => x"16",
          3909 => x"58",
          3910 => x"3f",
          3911 => x"0a",
          3912 => x"0a",
          3913 => x"2c",
          3914 => x"33",
          3915 => x"76",
          3916 => x"38",
          3917 => x"33",
          3918 => x"70",
          3919 => x"81",
          3920 => x"58",
          3921 => x"7a",
          3922 => x"38",
          3923 => x"83",
          3924 => x"80",
          3925 => x"38",
          3926 => x"57",
          3927 => x"08",
          3928 => x"38",
          3929 => x"18",
          3930 => x"80",
          3931 => x"80",
          3932 => x"fc",
          3933 => x"f8",
          3934 => x"80",
          3935 => x"38",
          3936 => x"e8",
          3937 => x"f3",
          3938 => x"80",
          3939 => x"80",
          3940 => x"f8",
          3941 => x"b4",
          3942 => x"ee",
          3943 => x"51",
          3944 => x"3f",
          3945 => x"ff",
          3946 => x"58",
          3947 => x"25",
          3948 => x"ff",
          3949 => x"51",
          3950 => x"3f",
          3951 => x"08",
          3952 => x"34",
          3953 => x"08",
          3954 => x"81",
          3955 => x"52",
          3956 => x"ab",
          3957 => x"0b",
          3958 => x"33",
          3959 => x"33",
          3960 => x"74",
          3961 => x"97",
          3962 => x"f0",
          3963 => x"51",
          3964 => x"3f",
          3965 => x"08",
          3966 => x"ff",
          3967 => x"84",
          3968 => x"52",
          3969 => x"a6",
          3970 => x"d1",
          3971 => x"05",
          3972 => x"d1",
          3973 => x"81",
          3974 => x"c7",
          3975 => x"34",
          3976 => x"d1",
          3977 => x"0b",
          3978 => x"34",
          3979 => x"8c",
          3980 => x"0d",
          3981 => x"ff",
          3982 => x"84",
          3983 => x"84",
          3984 => x"84",
          3985 => x"81",
          3986 => x"05",
          3987 => x"7b",
          3988 => x"97",
          3989 => x"70",
          3990 => x"84",
          3991 => x"84",
          3992 => x"58",
          3993 => x"74",
          3994 => x"93",
          3995 => x"f0",
          3996 => x"51",
          3997 => x"3f",
          3998 => x"08",
          3999 => x"ff",
          4000 => x"84",
          4001 => x"52",
          4002 => x"a5",
          4003 => x"d1",
          4004 => x"05",
          4005 => x"d1",
          4006 => x"81",
          4007 => x"c7",
          4008 => x"ff",
          4009 => x"84",
          4010 => x"84",
          4011 => x"84",
          4012 => x"81",
          4013 => x"05",
          4014 => x"7b",
          4015 => x"ab",
          4016 => x"70",
          4017 => x"84",
          4018 => x"84",
          4019 => x"58",
          4020 => x"74",
          4021 => x"a7",
          4022 => x"f0",
          4023 => x"51",
          4024 => x"3f",
          4025 => x"08",
          4026 => x"ff",
          4027 => x"84",
          4028 => x"52",
          4029 => x"a4",
          4030 => x"d1",
          4031 => x"05",
          4032 => x"d1",
          4033 => x"81",
          4034 => x"c7",
          4035 => x"80",
          4036 => x"83",
          4037 => x"70",
          4038 => x"fc",
          4039 => x"a4",
          4040 => x"70",
          4041 => x"56",
          4042 => x"3f",
          4043 => x"08",
          4044 => x"f3",
          4045 => x"10",
          4046 => x"a4",
          4047 => x"57",
          4048 => x"80",
          4049 => x"38",
          4050 => x"52",
          4051 => x"a8",
          4052 => x"f3",
          4053 => x"05",
          4054 => x"06",
          4055 => x"79",
          4056 => x"38",
          4057 => x"fc",
          4058 => x"39",
          4059 => x"f8",
          4060 => x"53",
          4061 => x"51",
          4062 => x"3f",
          4063 => x"08",
          4064 => x"82",
          4065 => x"83",
          4066 => x"51",
          4067 => x"3f",
          4068 => x"d1",
          4069 => x"0b",
          4070 => x"34",
          4071 => x"8c",
          4072 => x"0d",
          4073 => x"77",
          4074 => x"8c",
          4075 => x"ca",
          4076 => x"ba",
          4077 => x"a5",
          4078 => x"8c",
          4079 => x"5c",
          4080 => x"f8",
          4081 => x"f8",
          4082 => x"82",
          4083 => x"84",
          4084 => x"5a",
          4085 => x"08",
          4086 => x"81",
          4087 => x"38",
          4088 => x"08",
          4089 => x"c1",
          4090 => x"8c",
          4091 => x"0b",
          4092 => x"08",
          4093 => x"38",
          4094 => x"08",
          4095 => x"1b",
          4096 => x"77",
          4097 => x"ff",
          4098 => x"fc",
          4099 => x"10",
          4100 => x"05",
          4101 => x"40",
          4102 => x"80",
          4103 => x"82",
          4104 => x"06",
          4105 => x"05",
          4106 => x"53",
          4107 => x"db",
          4108 => x"ba",
          4109 => x"0c",
          4110 => x"33",
          4111 => x"83",
          4112 => x"70",
          4113 => x"41",
          4114 => x"81",
          4115 => x"ff",
          4116 => x"93",
          4117 => x"38",
          4118 => x"ff",
          4119 => x"06",
          4120 => x"77",
          4121 => x"f9",
          4122 => x"53",
          4123 => x"51",
          4124 => x"3f",
          4125 => x"33",
          4126 => x"81",
          4127 => x"57",
          4128 => x"80",
          4129 => x"0b",
          4130 => x"34",
          4131 => x"74",
          4132 => x"c7",
          4133 => x"fc",
          4134 => x"2b",
          4135 => x"83",
          4136 => x"81",
          4137 => x"52",
          4138 => x"da",
          4139 => x"ba",
          4140 => x"0c",
          4141 => x"33",
          4142 => x"83",
          4143 => x"70",
          4144 => x"41",
          4145 => x"ff",
          4146 => x"9e",
          4147 => x"f3",
          4148 => x"f7",
          4149 => x"f3",
          4150 => x"c0",
          4151 => x"b8",
          4152 => x"90",
          4153 => x"eb",
          4154 => x"39",
          4155 => x"02",
          4156 => x"33",
          4157 => x"80",
          4158 => x"5b",
          4159 => x"26",
          4160 => x"72",
          4161 => x"8b",
          4162 => x"25",
          4163 => x"72",
          4164 => x"a8",
          4165 => x"a0",
          4166 => x"a3",
          4167 => x"5e",
          4168 => x"9f",
          4169 => x"76",
          4170 => x"75",
          4171 => x"34",
          4172 => x"bd",
          4173 => x"f9",
          4174 => x"f9",
          4175 => x"98",
          4176 => x"2b",
          4177 => x"2b",
          4178 => x"7a",
          4179 => x"56",
          4180 => x"27",
          4181 => x"74",
          4182 => x"56",
          4183 => x"70",
          4184 => x"0c",
          4185 => x"ee",
          4186 => x"27",
          4187 => x"f9",
          4188 => x"98",
          4189 => x"78",
          4190 => x"55",
          4191 => x"e0",
          4192 => x"74",
          4193 => x"56",
          4194 => x"53",
          4195 => x"90",
          4196 => x"87",
          4197 => x"0b",
          4198 => x"33",
          4199 => x"11",
          4200 => x"33",
          4201 => x"11",
          4202 => x"41",
          4203 => x"87",
          4204 => x"0b",
          4205 => x"33",
          4206 => x"06",
          4207 => x"33",
          4208 => x"06",
          4209 => x"22",
          4210 => x"ff",
          4211 => x"29",
          4212 => x"58",
          4213 => x"5d",
          4214 => x"87",
          4215 => x"31",
          4216 => x"79",
          4217 => x"7e",
          4218 => x"7c",
          4219 => x"7a",
          4220 => x"06",
          4221 => x"06",
          4222 => x"14",
          4223 => x"57",
          4224 => x"74",
          4225 => x"83",
          4226 => x"74",
          4227 => x"70",
          4228 => x"59",
          4229 => x"06",
          4230 => x"2e",
          4231 => x"78",
          4232 => x"72",
          4233 => x"c1",
          4234 => x"70",
          4235 => x"34",
          4236 => x"33",
          4237 => x"05",
          4238 => x"39",
          4239 => x"80",
          4240 => x"b0",
          4241 => x"b8",
          4242 => x"81",
          4243 => x"b7",
          4244 => x"81",
          4245 => x"f9",
          4246 => x"74",
          4247 => x"5d",
          4248 => x"5e",
          4249 => x"27",
          4250 => x"73",
          4251 => x"73",
          4252 => x"71",
          4253 => x"5a",
          4254 => x"80",
          4255 => x"38",
          4256 => x"f9",
          4257 => x"0b",
          4258 => x"34",
          4259 => x"33",
          4260 => x"71",
          4261 => x"71",
          4262 => x"71",
          4263 => x"56",
          4264 => x"76",
          4265 => x"ae",
          4266 => x"39",
          4267 => x"38",
          4268 => x"33",
          4269 => x"06",
          4270 => x"11",
          4271 => x"33",
          4272 => x"11",
          4273 => x"80",
          4274 => x"5b",
          4275 => x"87",
          4276 => x"70",
          4277 => x"80",
          4278 => x"ff",
          4279 => x"ff",
          4280 => x"ff",
          4281 => x"ba",
          4282 => x"ff",
          4283 => x"75",
          4284 => x"5e",
          4285 => x"58",
          4286 => x"57",
          4287 => x"8b",
          4288 => x"31",
          4289 => x"29",
          4290 => x"7d",
          4291 => x"74",
          4292 => x"71",
          4293 => x"83",
          4294 => x"62",
          4295 => x"70",
          4296 => x"5f",
          4297 => x"55",
          4298 => x"85",
          4299 => x"29",
          4300 => x"31",
          4301 => x"06",
          4302 => x"fd",
          4303 => x"83",
          4304 => x"fd",
          4305 => x"f2",
          4306 => x"31",
          4307 => x"fe",
          4308 => x"3d",
          4309 => x"80",
          4310 => x"f4",
          4311 => x"b0",
          4312 => x"ee",
          4313 => x"80",
          4314 => x"73",
          4315 => x"80",
          4316 => x"76",
          4317 => x"34",
          4318 => x"34",
          4319 => x"8c",
          4320 => x"75",
          4321 => x"34",
          4322 => x"81",
          4323 => x"52",
          4324 => x"d8",
          4325 => x"87",
          4326 => x"54",
          4327 => x"56",
          4328 => x"f8",
          4329 => x"84",
          4330 => x"72",
          4331 => x"08",
          4332 => x"06",
          4333 => x"51",
          4334 => x"34",
          4335 => x"cc",
          4336 => x"06",
          4337 => x"53",
          4338 => x"81",
          4339 => x"08",
          4340 => x"88",
          4341 => x"75",
          4342 => x"0b",
          4343 => x"34",
          4344 => x"ba",
          4345 => x"3d",
          4346 => x"b8",
          4347 => x"ba",
          4348 => x"f7",
          4349 => x"af",
          4350 => x"84",
          4351 => x"33",
          4352 => x"33",
          4353 => x"81",
          4354 => x"26",
          4355 => x"84",
          4356 => x"83",
          4357 => x"83",
          4358 => x"72",
          4359 => x"87",
          4360 => x"11",
          4361 => x"22",
          4362 => x"59",
          4363 => x"05",
          4364 => x"ff",
          4365 => x"92",
          4366 => x"58",
          4367 => x"2e",
          4368 => x"83",
          4369 => x"76",
          4370 => x"83",
          4371 => x"83",
          4372 => x"76",
          4373 => x"ff",
          4374 => x"ff",
          4375 => x"55",
          4376 => x"82",
          4377 => x"19",
          4378 => x"f9",
          4379 => x"f9",
          4380 => x"83",
          4381 => x"84",
          4382 => x"5c",
          4383 => x"74",
          4384 => x"38",
          4385 => x"33",
          4386 => x"54",
          4387 => x"72",
          4388 => x"ac",
          4389 => x"de",
          4390 => x"55",
          4391 => x"33",
          4392 => x"34",
          4393 => x"05",
          4394 => x"70",
          4395 => x"34",
          4396 => x"84",
          4397 => x"27",
          4398 => x"9f",
          4399 => x"38",
          4400 => x"33",
          4401 => x"15",
          4402 => x"0b",
          4403 => x"34",
          4404 => x"81",
          4405 => x"81",
          4406 => x"9f",
          4407 => x"38",
          4408 => x"33",
          4409 => x"75",
          4410 => x"23",
          4411 => x"81",
          4412 => x"83",
          4413 => x"54",
          4414 => x"26",
          4415 => x"72",
          4416 => x"05",
          4417 => x"33",
          4418 => x"58",
          4419 => x"55",
          4420 => x"80",
          4421 => x"b0",
          4422 => x"ff",
          4423 => x"ff",
          4424 => x"29",
          4425 => x"54",
          4426 => x"27",
          4427 => x"98",
          4428 => x"e0",
          4429 => x"53",
          4430 => x"13",
          4431 => x"81",
          4432 => x"73",
          4433 => x"55",
          4434 => x"81",
          4435 => x"81",
          4436 => x"80",
          4437 => x"ff",
          4438 => x"29",
          4439 => x"5a",
          4440 => x"26",
          4441 => x"53",
          4442 => x"8c",
          4443 => x"0d",
          4444 => x"f9",
          4445 => x"f9",
          4446 => x"83",
          4447 => x"84",
          4448 => x"5c",
          4449 => x"7a",
          4450 => x"38",
          4451 => x"fe",
          4452 => x"81",
          4453 => x"05",
          4454 => x"33",
          4455 => x"75",
          4456 => x"06",
          4457 => x"73",
          4458 => x"05",
          4459 => x"33",
          4460 => x"78",
          4461 => x"56",
          4462 => x"73",
          4463 => x"ae",
          4464 => x"b8",
          4465 => x"de",
          4466 => x"31",
          4467 => x"a0",
          4468 => x"16",
          4469 => x"70",
          4470 => x"34",
          4471 => x"72",
          4472 => x"8a",
          4473 => x"e0",
          4474 => x"75",
          4475 => x"05",
          4476 => x"13",
          4477 => x"38",
          4478 => x"80",
          4479 => x"80",
          4480 => x"fe",
          4481 => x"f9",
          4482 => x"59",
          4483 => x"19",
          4484 => x"84",
          4485 => x"59",
          4486 => x"fc",
          4487 => x"02",
          4488 => x"05",
          4489 => x"70",
          4490 => x"38",
          4491 => x"83",
          4492 => x"51",
          4493 => x"84",
          4494 => x"51",
          4495 => x"86",
          4496 => x"f9",
          4497 => x"0b",
          4498 => x"0c",
          4499 => x"04",
          4500 => x"f9",
          4501 => x"f9",
          4502 => x"81",
          4503 => x"52",
          4504 => x"e2",
          4505 => x"51",
          4506 => x"bc",
          4507 => x"84",
          4508 => x"86",
          4509 => x"83",
          4510 => x"70",
          4511 => x"09",
          4512 => x"72",
          4513 => x"53",
          4514 => x"f9",
          4515 => x"39",
          4516 => x"33",
          4517 => x"b7",
          4518 => x"11",
          4519 => x"70",
          4520 => x"38",
          4521 => x"83",
          4522 => x"80",
          4523 => x"8c",
          4524 => x"0d",
          4525 => x"bd",
          4526 => x"31",
          4527 => x"9f",
          4528 => x"54",
          4529 => x"70",
          4530 => x"34",
          4531 => x"ba",
          4532 => x"3d",
          4533 => x"f9",
          4534 => x"05",
          4535 => x"33",
          4536 => x"55",
          4537 => x"25",
          4538 => x"53",
          4539 => x"bd",
          4540 => x"84",
          4541 => x"86",
          4542 => x"80",
          4543 => x"bd",
          4544 => x"bc",
          4545 => x"ff",
          4546 => x"56",
          4547 => x"25",
          4548 => x"81",
          4549 => x"83",
          4550 => x"fe",
          4551 => x"3d",
          4552 => x"05",
          4553 => x"b1",
          4554 => x"70",
          4555 => x"c4",
          4556 => x"70",
          4557 => x"f9",
          4558 => x"80",
          4559 => x"84",
          4560 => x"06",
          4561 => x"2a",
          4562 => x"53",
          4563 => x"f0",
          4564 => x"06",
          4565 => x"f2",
          4566 => x"b8",
          4567 => x"84",
          4568 => x"83",
          4569 => x"83",
          4570 => x"81",
          4571 => x"07",
          4572 => x"f9",
          4573 => x"0b",
          4574 => x"0c",
          4575 => x"04",
          4576 => x"33",
          4577 => x"51",
          4578 => x"b8",
          4579 => x"83",
          4580 => x"81",
          4581 => x"07",
          4582 => x"f9",
          4583 => x"39",
          4584 => x"83",
          4585 => x"80",
          4586 => x"8c",
          4587 => x"0d",
          4588 => x"b8",
          4589 => x"06",
          4590 => x"70",
          4591 => x"34",
          4592 => x"83",
          4593 => x"87",
          4594 => x"83",
          4595 => x"ff",
          4596 => x"f9",
          4597 => x"fd",
          4598 => x"51",
          4599 => x"b8",
          4600 => x"39",
          4601 => x"33",
          4602 => x"83",
          4603 => x"83",
          4604 => x"ff",
          4605 => x"f9",
          4606 => x"f9",
          4607 => x"51",
          4608 => x"b8",
          4609 => x"39",
          4610 => x"33",
          4611 => x"51",
          4612 => x"b8",
          4613 => x"39",
          4614 => x"33",
          4615 => x"80",
          4616 => x"70",
          4617 => x"34",
          4618 => x"83",
          4619 => x"81",
          4620 => x"07",
          4621 => x"f9",
          4622 => x"ba",
          4623 => x"b8",
          4624 => x"06",
          4625 => x"51",
          4626 => x"b8",
          4627 => x"39",
          4628 => x"33",
          4629 => x"80",
          4630 => x"70",
          4631 => x"34",
          4632 => x"83",
          4633 => x"81",
          4634 => x"07",
          4635 => x"f9",
          4636 => x"82",
          4637 => x"b8",
          4638 => x"06",
          4639 => x"f9",
          4640 => x"f2",
          4641 => x"b8",
          4642 => x"06",
          4643 => x"70",
          4644 => x"34",
          4645 => x"f3",
          4646 => x"bf",
          4647 => x"84",
          4648 => x"05",
          4649 => x"bc",
          4650 => x"bb",
          4651 => x"bd",
          4652 => x"82",
          4653 => x"5f",
          4654 => x"78",
          4655 => x"a1",
          4656 => x"24",
          4657 => x"81",
          4658 => x"38",
          4659 => x"82",
          4660 => x"84",
          4661 => x"7a",
          4662 => x"34",
          4663 => x"ba",
          4664 => x"f9",
          4665 => x"3d",
          4666 => x"83",
          4667 => x"06",
          4668 => x"0b",
          4669 => x"34",
          4670 => x"b8",
          4671 => x"0b",
          4672 => x"34",
          4673 => x"f9",
          4674 => x"0b",
          4675 => x"23",
          4676 => x"b8",
          4677 => x"84",
          4678 => x"56",
          4679 => x"33",
          4680 => x"7c",
          4681 => x"83",
          4682 => x"ff",
          4683 => x"7d",
          4684 => x"34",
          4685 => x"b8",
          4686 => x"83",
          4687 => x"7b",
          4688 => x"23",
          4689 => x"bd",
          4690 => x"0d",
          4691 => x"84",
          4692 => x"81",
          4693 => x"84",
          4694 => x"83",
          4695 => x"a8",
          4696 => x"bd",
          4697 => x"83",
          4698 => x"84",
          4699 => x"58",
          4700 => x"33",
          4701 => x"8d",
          4702 => x"55",
          4703 => x"53",
          4704 => x"e3",
          4705 => x"81",
          4706 => x"0b",
          4707 => x"33",
          4708 => x"79",
          4709 => x"79",
          4710 => x"e0",
          4711 => x"53",
          4712 => x"f8",
          4713 => x"e1",
          4714 => x"70",
          4715 => x"84",
          4716 => x"52",
          4717 => x"7a",
          4718 => x"83",
          4719 => x"ff",
          4720 => x"7d",
          4721 => x"34",
          4722 => x"b8",
          4723 => x"83",
          4724 => x"7b",
          4725 => x"23",
          4726 => x"bd",
          4727 => x"0d",
          4728 => x"84",
          4729 => x"81",
          4730 => x"84",
          4731 => x"83",
          4732 => x"a8",
          4733 => x"bd",
          4734 => x"83",
          4735 => x"83",
          4736 => x"ff",
          4737 => x"84",
          4738 => x"52",
          4739 => x"51",
          4740 => x"3f",
          4741 => x"f7",
          4742 => x"92",
          4743 => x"84",
          4744 => x"27",
          4745 => x"83",
          4746 => x"33",
          4747 => x"84",
          4748 => x"d5",
          4749 => x"70",
          4750 => x"5a",
          4751 => x"f9",
          4752 => x"02",
          4753 => x"05",
          4754 => x"80",
          4755 => x"bd",
          4756 => x"bc",
          4757 => x"29",
          4758 => x"a0",
          4759 => x"f9",
          4760 => x"51",
          4761 => x"7c",
          4762 => x"83",
          4763 => x"83",
          4764 => x"52",
          4765 => x"57",
          4766 => x"2e",
          4767 => x"75",
          4768 => x"f9",
          4769 => x"24",
          4770 => x"75",
          4771 => x"85",
          4772 => x"2e",
          4773 => x"84",
          4774 => x"83",
          4775 => x"83",
          4776 => x"72",
          4777 => x"55",
          4778 => x"b8",
          4779 => x"87",
          4780 => x"14",
          4781 => x"80",
          4782 => x"bd",
          4783 => x"ba",
          4784 => x"29",
          4785 => x"56",
          4786 => x"f9",
          4787 => x"83",
          4788 => x"73",
          4789 => x"58",
          4790 => x"b8",
          4791 => x"b0",
          4792 => x"84",
          4793 => x"70",
          4794 => x"83",
          4795 => x"83",
          4796 => x"72",
          4797 => x"57",
          4798 => x"57",
          4799 => x"33",
          4800 => x"14",
          4801 => x"70",
          4802 => x"59",
          4803 => x"26",
          4804 => x"84",
          4805 => x"58",
          4806 => x"38",
          4807 => x"72",
          4808 => x"34",
          4809 => x"33",
          4810 => x"2e",
          4811 => x"b8",
          4812 => x"76",
          4813 => x"fb",
          4814 => x"84",
          4815 => x"89",
          4816 => x"75",
          4817 => x"38",
          4818 => x"80",
          4819 => x"8a",
          4820 => x"06",
          4821 => x"81",
          4822 => x"f1",
          4823 => x"0b",
          4824 => x"34",
          4825 => x"83",
          4826 => x"33",
          4827 => x"88",
          4828 => x"34",
          4829 => x"09",
          4830 => x"89",
          4831 => x"76",
          4832 => x"fd",
          4833 => x"13",
          4834 => x"06",
          4835 => x"83",
          4836 => x"38",
          4837 => x"51",
          4838 => x"81",
          4839 => x"ff",
          4840 => x"83",
          4841 => x"38",
          4842 => x"74",
          4843 => x"34",
          4844 => x"75",
          4845 => x"f9",
          4846 => x"0b",
          4847 => x"0c",
          4848 => x"04",
          4849 => x"2e",
          4850 => x"fd",
          4851 => x"f9",
          4852 => x"81",
          4853 => x"ff",
          4854 => x"83",
          4855 => x"72",
          4856 => x"34",
          4857 => x"51",
          4858 => x"83",
          4859 => x"70",
          4860 => x"55",
          4861 => x"73",
          4862 => x"73",
          4863 => x"f9",
          4864 => x"a0",
          4865 => x"83",
          4866 => x"81",
          4867 => x"ef",
          4868 => x"90",
          4869 => x"75",
          4870 => x"3f",
          4871 => x"e6",
          4872 => x"80",
          4873 => x"84",
          4874 => x"57",
          4875 => x"2e",
          4876 => x"75",
          4877 => x"82",
          4878 => x"2e",
          4879 => x"78",
          4880 => x"d1",
          4881 => x"2e",
          4882 => x"78",
          4883 => x"8f",
          4884 => x"80",
          4885 => x"bc",
          4886 => x"bd",
          4887 => x"29",
          4888 => x"5c",
          4889 => x"19",
          4890 => x"a0",
          4891 => x"84",
          4892 => x"83",
          4893 => x"83",
          4894 => x"72",
          4895 => x"5a",
          4896 => x"78",
          4897 => x"18",
          4898 => x"bc",
          4899 => x"29",
          4900 => x"5a",
          4901 => x"33",
          4902 => x"b0",
          4903 => x"84",
          4904 => x"70",
          4905 => x"83",
          4906 => x"83",
          4907 => x"72",
          4908 => x"42",
          4909 => x"59",
          4910 => x"33",
          4911 => x"1f",
          4912 => x"70",
          4913 => x"42",
          4914 => x"26",
          4915 => x"84",
          4916 => x"5a",
          4917 => x"38",
          4918 => x"75",
          4919 => x"34",
          4920 => x"ba",
          4921 => x"3d",
          4922 => x"b7",
          4923 => x"38",
          4924 => x"81",
          4925 => x"b8",
          4926 => x"38",
          4927 => x"2e",
          4928 => x"80",
          4929 => x"88",
          4930 => x"80",
          4931 => x"bc",
          4932 => x"bd",
          4933 => x"29",
          4934 => x"40",
          4935 => x"19",
          4936 => x"a0",
          4937 => x"84",
          4938 => x"83",
          4939 => x"83",
          4940 => x"72",
          4941 => x"41",
          4942 => x"78",
          4943 => x"1f",
          4944 => x"bc",
          4945 => x"29",
          4946 => x"83",
          4947 => x"87",
          4948 => x"1b",
          4949 => x"80",
          4950 => x"ff",
          4951 => x"ba",
          4952 => x"bd",
          4953 => x"29",
          4954 => x"43",
          4955 => x"f9",
          4956 => x"84",
          4957 => x"34",
          4958 => x"77",
          4959 => x"41",
          4960 => x"fe",
          4961 => x"83",
          4962 => x"80",
          4963 => x"8c",
          4964 => x"0d",
          4965 => x"2e",
          4966 => x"78",
          4967 => x"81",
          4968 => x"2e",
          4969 => x"fd",
          4970 => x"0b",
          4971 => x"34",
          4972 => x"ba",
          4973 => x"3d",
          4974 => x"9b",
          4975 => x"38",
          4976 => x"75",
          4977 => x"d0",
          4978 => x"8c",
          4979 => x"59",
          4980 => x"b9",
          4981 => x"84",
          4982 => x"34",
          4983 => x"06",
          4984 => x"84",
          4985 => x"34",
          4986 => x"ba",
          4987 => x"3d",
          4988 => x"9b",
          4989 => x"38",
          4990 => x"b9",
          4991 => x"b8",
          4992 => x"f9",
          4993 => x"f9",
          4994 => x"72",
          4995 => x"40",
          4996 => x"88",
          4997 => x"a3",
          4998 => x"34",
          4999 => x"33",
          5000 => x"33",
          5001 => x"22",
          5002 => x"12",
          5003 => x"56",
          5004 => x"be",
          5005 => x"f9",
          5006 => x"71",
          5007 => x"57",
          5008 => x"33",
          5009 => x"80",
          5010 => x"b8",
          5011 => x"81",
          5012 => x"f9",
          5013 => x"f9",
          5014 => x"72",
          5015 => x"42",
          5016 => x"83",
          5017 => x"60",
          5018 => x"05",
          5019 => x"58",
          5020 => x"81",
          5021 => x"ea",
          5022 => x"0b",
          5023 => x"34",
          5024 => x"84",
          5025 => x"83",
          5026 => x"70",
          5027 => x"83",
          5028 => x"73",
          5029 => x"87",
          5030 => x"05",
          5031 => x"22",
          5032 => x"72",
          5033 => x"70",
          5034 => x"06",
          5035 => x"33",
          5036 => x"5a",
          5037 => x"2e",
          5038 => x"78",
          5039 => x"ff",
          5040 => x"76",
          5041 => x"76",
          5042 => x"f9",
          5043 => x"90",
          5044 => x"84",
          5045 => x"80",
          5046 => x"8d",
          5047 => x"84",
          5048 => x"80",
          5049 => x"8f",
          5050 => x"84",
          5051 => x"80",
          5052 => x"8c",
          5053 => x"0d",
          5054 => x"bc",
          5055 => x"f4",
          5056 => x"bd",
          5057 => x"f5",
          5058 => x"bb",
          5059 => x"f6",
          5060 => x"84",
          5061 => x"80",
          5062 => x"8c",
          5063 => x"0d",
          5064 => x"ff",
          5065 => x"06",
          5066 => x"83",
          5067 => x"84",
          5068 => x"70",
          5069 => x"83",
          5070 => x"70",
          5071 => x"72",
          5072 => x"87",
          5073 => x"05",
          5074 => x"22",
          5075 => x"7b",
          5076 => x"83",
          5077 => x"83",
          5078 => x"44",
          5079 => x"42",
          5080 => x"81",
          5081 => x"38",
          5082 => x"06",
          5083 => x"56",
          5084 => x"75",
          5085 => x"f9",
          5086 => x"81",
          5087 => x"81",
          5088 => x"81",
          5089 => x"72",
          5090 => x"40",
          5091 => x"a8",
          5092 => x"a0",
          5093 => x"84",
          5094 => x"83",
          5095 => x"83",
          5096 => x"72",
          5097 => x"5a",
          5098 => x"a0",
          5099 => x"be",
          5100 => x"f9",
          5101 => x"71",
          5102 => x"5a",
          5103 => x"b8",
          5104 => x"b0",
          5105 => x"84",
          5106 => x"70",
          5107 => x"83",
          5108 => x"83",
          5109 => x"72",
          5110 => x"43",
          5111 => x"59",
          5112 => x"33",
          5113 => x"de",
          5114 => x"1a",
          5115 => x"06",
          5116 => x"7b",
          5117 => x"38",
          5118 => x"33",
          5119 => x"d0",
          5120 => x"58",
          5121 => x"bd",
          5122 => x"bd",
          5123 => x"ff",
          5124 => x"05",
          5125 => x"39",
          5126 => x"95",
          5127 => x"bd",
          5128 => x"38",
          5129 => x"95",
          5130 => x"b9",
          5131 => x"7e",
          5132 => x"ff",
          5133 => x"75",
          5134 => x"c8",
          5135 => x"10",
          5136 => x"05",
          5137 => x"04",
          5138 => x"f9",
          5139 => x"52",
          5140 => x"9f",
          5141 => x"84",
          5142 => x"9c",
          5143 => x"83",
          5144 => x"84",
          5145 => x"70",
          5146 => x"83",
          5147 => x"70",
          5148 => x"72",
          5149 => x"87",
          5150 => x"05",
          5151 => x"22",
          5152 => x"7b",
          5153 => x"83",
          5154 => x"83",
          5155 => x"46",
          5156 => x"59",
          5157 => x"81",
          5158 => x"38",
          5159 => x"81",
          5160 => x"81",
          5161 => x"81",
          5162 => x"72",
          5163 => x"58",
          5164 => x"a8",
          5165 => x"a0",
          5166 => x"84",
          5167 => x"83",
          5168 => x"83",
          5169 => x"72",
          5170 => x"5e",
          5171 => x"a0",
          5172 => x"be",
          5173 => x"f9",
          5174 => x"71",
          5175 => x"5e",
          5176 => x"33",
          5177 => x"80",
          5178 => x"b8",
          5179 => x"81",
          5180 => x"f9",
          5181 => x"f9",
          5182 => x"72",
          5183 => x"44",
          5184 => x"83",
          5185 => x"84",
          5186 => x"34",
          5187 => x"70",
          5188 => x"5b",
          5189 => x"26",
          5190 => x"84",
          5191 => x"58",
          5192 => x"38",
          5193 => x"75",
          5194 => x"34",
          5195 => x"81",
          5196 => x"59",
          5197 => x"f7",
          5198 => x"f9",
          5199 => x"b8",
          5200 => x"f9",
          5201 => x"81",
          5202 => x"81",
          5203 => x"81",
          5204 => x"72",
          5205 => x"5b",
          5206 => x"5b",
          5207 => x"33",
          5208 => x"80",
          5209 => x"b8",
          5210 => x"f9",
          5211 => x"f9",
          5212 => x"71",
          5213 => x"41",
          5214 => x"0b",
          5215 => x"1c",
          5216 => x"bc",
          5217 => x"29",
          5218 => x"83",
          5219 => x"87",
          5220 => x"1a",
          5221 => x"80",
          5222 => x"ff",
          5223 => x"ba",
          5224 => x"bd",
          5225 => x"29",
          5226 => x"5a",
          5227 => x"f9",
          5228 => x"98",
          5229 => x"60",
          5230 => x"81",
          5231 => x"58",
          5232 => x"fe",
          5233 => x"83",
          5234 => x"fe",
          5235 => x"0b",
          5236 => x"0c",
          5237 => x"ba",
          5238 => x"3d",
          5239 => x"f9",
          5240 => x"59",
          5241 => x"19",
          5242 => x"83",
          5243 => x"70",
          5244 => x"58",
          5245 => x"f9",
          5246 => x"0b",
          5247 => x"34",
          5248 => x"ba",
          5249 => x"3d",
          5250 => x"f9",
          5251 => x"5b",
          5252 => x"1b",
          5253 => x"83",
          5254 => x"84",
          5255 => x"83",
          5256 => x"5b",
          5257 => x"5c",
          5258 => x"84",
          5259 => x"9c",
          5260 => x"53",
          5261 => x"ff",
          5262 => x"84",
          5263 => x"80",
          5264 => x"38",
          5265 => x"33",
          5266 => x"5a",
          5267 => x"8d",
          5268 => x"83",
          5269 => x"02",
          5270 => x"22",
          5271 => x"e0",
          5272 => x"cf",
          5273 => x"be",
          5274 => x"84",
          5275 => x"33",
          5276 => x"f9",
          5277 => x"b8",
          5278 => x"f9",
          5279 => x"5b",
          5280 => x"39",
          5281 => x"33",
          5282 => x"33",
          5283 => x"33",
          5284 => x"05",
          5285 => x"84",
          5286 => x"33",
          5287 => x"a0",
          5288 => x"84",
          5289 => x"83",
          5290 => x"83",
          5291 => x"72",
          5292 => x"5a",
          5293 => x"78",
          5294 => x"18",
          5295 => x"bc",
          5296 => x"29",
          5297 => x"83",
          5298 => x"60",
          5299 => x"80",
          5300 => x"b8",
          5301 => x"81",
          5302 => x"f9",
          5303 => x"f9",
          5304 => x"72",
          5305 => x"5f",
          5306 => x"83",
          5307 => x"84",
          5308 => x"34",
          5309 => x"81",
          5310 => x"58",
          5311 => x"90",
          5312 => x"b8",
          5313 => x"77",
          5314 => x"ff",
          5315 => x"83",
          5316 => x"80",
          5317 => x"88",
          5318 => x"83",
          5319 => x"80",
          5320 => x"38",
          5321 => x"33",
          5322 => x"b4",
          5323 => x"81",
          5324 => x"3f",
          5325 => x"ba",
          5326 => x"3d",
          5327 => x"b9",
          5328 => x"f9",
          5329 => x"b9",
          5330 => x"f9",
          5331 => x"b9",
          5332 => x"76",
          5333 => x"23",
          5334 => x"83",
          5335 => x"84",
          5336 => x"83",
          5337 => x"84",
          5338 => x"83",
          5339 => x"84",
          5340 => x"ff",
          5341 => x"b9",
          5342 => x"7a",
          5343 => x"93",
          5344 => x"e0",
          5345 => x"86",
          5346 => x"06",
          5347 => x"83",
          5348 => x"81",
          5349 => x"f9",
          5350 => x"05",
          5351 => x"83",
          5352 => x"94",
          5353 => x"57",
          5354 => x"3f",
          5355 => x"fe",
          5356 => x"ba",
          5357 => x"ff",
          5358 => x"90",
          5359 => x"05",
          5360 => x"24",
          5361 => x"76",
          5362 => x"f0",
          5363 => x"c3",
          5364 => x"39",
          5365 => x"b9",
          5366 => x"58",
          5367 => x"06",
          5368 => x"27",
          5369 => x"77",
          5370 => x"e0",
          5371 => x"33",
          5372 => x"b1",
          5373 => x"38",
          5374 => x"83",
          5375 => x"5f",
          5376 => x"84",
          5377 => x"5e",
          5378 => x"8f",
          5379 => x"f9",
          5380 => x"b9",
          5381 => x"71",
          5382 => x"70",
          5383 => x"06",
          5384 => x"5e",
          5385 => x"f9",
          5386 => x"e7",
          5387 => x"8d",
          5388 => x"80",
          5389 => x"38",
          5390 => x"33",
          5391 => x"81",
          5392 => x"b8",
          5393 => x"57",
          5394 => x"27",
          5395 => x"75",
          5396 => x"34",
          5397 => x"80",
          5398 => x"bd",
          5399 => x"bc",
          5400 => x"ff",
          5401 => x"7b",
          5402 => x"a7",
          5403 => x"56",
          5404 => x"bc",
          5405 => x"39",
          5406 => x"f9",
          5407 => x"f9",
          5408 => x"b7",
          5409 => x"05",
          5410 => x"76",
          5411 => x"38",
          5412 => x"75",
          5413 => x"34",
          5414 => x"84",
          5415 => x"40",
          5416 => x"8d",
          5417 => x"f9",
          5418 => x"b9",
          5419 => x"71",
          5420 => x"70",
          5421 => x"06",
          5422 => x"42",
          5423 => x"f9",
          5424 => x"cf",
          5425 => x"8d",
          5426 => x"80",
          5427 => x"38",
          5428 => x"22",
          5429 => x"2e",
          5430 => x"fc",
          5431 => x"b8",
          5432 => x"f9",
          5433 => x"f9",
          5434 => x"71",
          5435 => x"a3",
          5436 => x"83",
          5437 => x"43",
          5438 => x"71",
          5439 => x"70",
          5440 => x"06",
          5441 => x"08",
          5442 => x"80",
          5443 => x"5d",
          5444 => x"82",
          5445 => x"bf",
          5446 => x"83",
          5447 => x"fb",
          5448 => x"b9",
          5449 => x"79",
          5450 => x"e7",
          5451 => x"e0",
          5452 => x"99",
          5453 => x"06",
          5454 => x"81",
          5455 => x"91",
          5456 => x"39",
          5457 => x"33",
          5458 => x"2e",
          5459 => x"84",
          5460 => x"83",
          5461 => x"5d",
          5462 => x"b8",
          5463 => x"11",
          5464 => x"75",
          5465 => x"38",
          5466 => x"83",
          5467 => x"fb",
          5468 => x"b9",
          5469 => x"76",
          5470 => x"c8",
          5471 => x"e1",
          5472 => x"bc",
          5473 => x"05",
          5474 => x"33",
          5475 => x"41",
          5476 => x"25",
          5477 => x"57",
          5478 => x"bc",
          5479 => x"39",
          5480 => x"51",
          5481 => x"3f",
          5482 => x"b9",
          5483 => x"57",
          5484 => x"8b",
          5485 => x"10",
          5486 => x"05",
          5487 => x"5a",
          5488 => x"51",
          5489 => x"3f",
          5490 => x"81",
          5491 => x"b9",
          5492 => x"58",
          5493 => x"82",
          5494 => x"8d",
          5495 => x"7d",
          5496 => x"38",
          5497 => x"22",
          5498 => x"26",
          5499 => x"57",
          5500 => x"81",
          5501 => x"d5",
          5502 => x"97",
          5503 => x"8d",
          5504 => x"77",
          5505 => x"38",
          5506 => x"33",
          5507 => x"81",
          5508 => x"b9",
          5509 => x"05",
          5510 => x"06",
          5511 => x"33",
          5512 => x"06",
          5513 => x"43",
          5514 => x"5c",
          5515 => x"27",
          5516 => x"5a",
          5517 => x"ba",
          5518 => x"ff",
          5519 => x"58",
          5520 => x"27",
          5521 => x"57",
          5522 => x"bc",
          5523 => x"80",
          5524 => x"57",
          5525 => x"27",
          5526 => x"7a",
          5527 => x"f9",
          5528 => x"af",
          5529 => x"8d",
          5530 => x"80",
          5531 => x"38",
          5532 => x"33",
          5533 => x"33",
          5534 => x"7f",
          5535 => x"38",
          5536 => x"33",
          5537 => x"33",
          5538 => x"06",
          5539 => x"33",
          5540 => x"11",
          5541 => x"80",
          5542 => x"ba",
          5543 => x"71",
          5544 => x"70",
          5545 => x"06",
          5546 => x"33",
          5547 => x"59",
          5548 => x"81",
          5549 => x"38",
          5550 => x"ff",
          5551 => x"31",
          5552 => x"7c",
          5553 => x"38",
          5554 => x"33",
          5555 => x"27",
          5556 => x"ff",
          5557 => x"83",
          5558 => x"7c",
          5559 => x"70",
          5560 => x"57",
          5561 => x"8e",
          5562 => x"b7",
          5563 => x"76",
          5564 => x"ee",
          5565 => x"56",
          5566 => x"bc",
          5567 => x"ff",
          5568 => x"ba",
          5569 => x"80",
          5570 => x"26",
          5571 => x"77",
          5572 => x"7e",
          5573 => x"71",
          5574 => x"5e",
          5575 => x"87",
          5576 => x"5b",
          5577 => x"80",
          5578 => x"06",
          5579 => x"06",
          5580 => x"1d",
          5581 => x"5c",
          5582 => x"f7",
          5583 => x"98",
          5584 => x"e0",
          5585 => x"5f",
          5586 => x"1f",
          5587 => x"81",
          5588 => x"76",
          5589 => x"58",
          5590 => x"81",
          5591 => x"81",
          5592 => x"80",
          5593 => x"ff",
          5594 => x"29",
          5595 => x"5e",
          5596 => x"27",
          5597 => x"e0",
          5598 => x"5f",
          5599 => x"1f",
          5600 => x"81",
          5601 => x"76",
          5602 => x"58",
          5603 => x"81",
          5604 => x"81",
          5605 => x"80",
          5606 => x"ff",
          5607 => x"29",
          5608 => x"5e",
          5609 => x"26",
          5610 => x"f6",
          5611 => x"b9",
          5612 => x"75",
          5613 => x"e0",
          5614 => x"84",
          5615 => x"51",
          5616 => x"f6",
          5617 => x"0b",
          5618 => x"33",
          5619 => x"b9",
          5620 => x"59",
          5621 => x"78",
          5622 => x"84",
          5623 => x"56",
          5624 => x"09",
          5625 => x"be",
          5626 => x"bd",
          5627 => x"81",
          5628 => x"f9",
          5629 => x"43",
          5630 => x"ff",
          5631 => x"38",
          5632 => x"33",
          5633 => x"26",
          5634 => x"7e",
          5635 => x"56",
          5636 => x"f5",
          5637 => x"76",
          5638 => x"27",
          5639 => x"f5",
          5640 => x"10",
          5641 => x"90",
          5642 => x"87",
          5643 => x"11",
          5644 => x"5a",
          5645 => x"80",
          5646 => x"06",
          5647 => x"75",
          5648 => x"79",
          5649 => x"76",
          5650 => x"83",
          5651 => x"70",
          5652 => x"90",
          5653 => x"88",
          5654 => x"07",
          5655 => x"52",
          5656 => x"7a",
          5657 => x"80",
          5658 => x"05",
          5659 => x"76",
          5660 => x"58",
          5661 => x"26",
          5662 => x"b8",
          5663 => x"b7",
          5664 => x"5f",
          5665 => x"06",
          5666 => x"06",
          5667 => x"22",
          5668 => x"64",
          5669 => x"59",
          5670 => x"26",
          5671 => x"78",
          5672 => x"7b",
          5673 => x"57",
          5674 => x"1d",
          5675 => x"76",
          5676 => x"38",
          5677 => x"33",
          5678 => x"18",
          5679 => x"0b",
          5680 => x"34",
          5681 => x"81",
          5682 => x"81",
          5683 => x"76",
          5684 => x"38",
          5685 => x"e0",
          5686 => x"78",
          5687 => x"5a",
          5688 => x"57",
          5689 => x"d6",
          5690 => x"39",
          5691 => x"81",
          5692 => x"58",
          5693 => x"83",
          5694 => x"70",
          5695 => x"71",
          5696 => x"f0",
          5697 => x"2a",
          5698 => x"57",
          5699 => x"2e",
          5700 => x"be",
          5701 => x"0b",
          5702 => x"34",
          5703 => x"81",
          5704 => x"56",
          5705 => x"83",
          5706 => x"33",
          5707 => x"88",
          5708 => x"34",
          5709 => x"33",
          5710 => x"33",
          5711 => x"22",
          5712 => x"33",
          5713 => x"5d",
          5714 => x"83",
          5715 => x"87",
          5716 => x"83",
          5717 => x"81",
          5718 => x"ff",
          5719 => x"f4",
          5720 => x"f9",
          5721 => x"fd",
          5722 => x"56",
          5723 => x"b8",
          5724 => x"83",
          5725 => x"81",
          5726 => x"07",
          5727 => x"f9",
          5728 => x"39",
          5729 => x"33",
          5730 => x"81",
          5731 => x"83",
          5732 => x"c3",
          5733 => x"b8",
          5734 => x"06",
          5735 => x"75",
          5736 => x"34",
          5737 => x"80",
          5738 => x"f9",
          5739 => x"18",
          5740 => x"06",
          5741 => x"a4",
          5742 => x"b8",
          5743 => x"06",
          5744 => x"f9",
          5745 => x"8f",
          5746 => x"b8",
          5747 => x"06",
          5748 => x"75",
          5749 => x"34",
          5750 => x"83",
          5751 => x"81",
          5752 => x"e0",
          5753 => x"83",
          5754 => x"fe",
          5755 => x"f9",
          5756 => x"cf",
          5757 => x"07",
          5758 => x"f9",
          5759 => x"d7",
          5760 => x"b8",
          5761 => x"06",
          5762 => x"75",
          5763 => x"34",
          5764 => x"83",
          5765 => x"81",
          5766 => x"07",
          5767 => x"f9",
          5768 => x"b3",
          5769 => x"b8",
          5770 => x"06",
          5771 => x"75",
          5772 => x"34",
          5773 => x"83",
          5774 => x"81",
          5775 => x"07",
          5776 => x"f9",
          5777 => x"8f",
          5778 => x"b8",
          5779 => x"06",
          5780 => x"f9",
          5781 => x"ff",
          5782 => x"b8",
          5783 => x"07",
          5784 => x"f9",
          5785 => x"ef",
          5786 => x"b8",
          5787 => x"07",
          5788 => x"f9",
          5789 => x"df",
          5790 => x"b8",
          5791 => x"06",
          5792 => x"56",
          5793 => x"b8",
          5794 => x"39",
          5795 => x"33",
          5796 => x"b0",
          5797 => x"83",
          5798 => x"fd",
          5799 => x"0b",
          5800 => x"34",
          5801 => x"51",
          5802 => x"ec",
          5803 => x"b9",
          5804 => x"f9",
          5805 => x"b9",
          5806 => x"f9",
          5807 => x"b9",
          5808 => x"78",
          5809 => x"23",
          5810 => x"b9",
          5811 => x"c7",
          5812 => x"84",
          5813 => x"80",
          5814 => x"8c",
          5815 => x"0d",
          5816 => x"f9",
          5817 => x"f9",
          5818 => x"81",
          5819 => x"ff",
          5820 => x"cf",
          5821 => x"90",
          5822 => x"dc",
          5823 => x"05",
          5824 => x"83",
          5825 => x"8c",
          5826 => x"84",
          5827 => x"84",
          5828 => x"80",
          5829 => x"8c",
          5830 => x"84",
          5831 => x"9c",
          5832 => x"77",
          5833 => x"34",
          5834 => x"84",
          5835 => x"81",
          5836 => x"7a",
          5837 => x"34",
          5838 => x"fe",
          5839 => x"80",
          5840 => x"84",
          5841 => x"23",
          5842 => x"b9",
          5843 => x"39",
          5844 => x"f9",
          5845 => x"52",
          5846 => x"97",
          5847 => x"bd",
          5848 => x"ff",
          5849 => x"05",
          5850 => x"39",
          5851 => x"f9",
          5852 => x"52",
          5853 => x"fb",
          5854 => x"39",
          5855 => x"eb",
          5856 => x"8f",
          5857 => x"bd",
          5858 => x"70",
          5859 => x"2c",
          5860 => x"5f",
          5861 => x"39",
          5862 => x"51",
          5863 => x"b8",
          5864 => x"75",
          5865 => x"eb",
          5866 => x"f9",
          5867 => x"e3",
          5868 => x"bc",
          5869 => x"70",
          5870 => x"2c",
          5871 => x"40",
          5872 => x"39",
          5873 => x"33",
          5874 => x"b7",
          5875 => x"11",
          5876 => x"75",
          5877 => x"c0",
          5878 => x"f3",
          5879 => x"b7",
          5880 => x"81",
          5881 => x"5c",
          5882 => x"ee",
          5883 => x"f9",
          5884 => x"b8",
          5885 => x"81",
          5886 => x"f9",
          5887 => x"74",
          5888 => x"a3",
          5889 => x"83",
          5890 => x"5f",
          5891 => x"29",
          5892 => x"ff",
          5893 => x"f8",
          5894 => x"5b",
          5895 => x"5d",
          5896 => x"81",
          5897 => x"83",
          5898 => x"ff",
          5899 => x"80",
          5900 => x"89",
          5901 => x"ff",
          5902 => x"76",
          5903 => x"38",
          5904 => x"75",
          5905 => x"23",
          5906 => x"06",
          5907 => x"57",
          5908 => x"83",
          5909 => x"b7",
          5910 => x"76",
          5911 => x"ec",
          5912 => x"56",
          5913 => x"bc",
          5914 => x"ff",
          5915 => x"ba",
          5916 => x"80",
          5917 => x"26",
          5918 => x"77",
          5919 => x"7e",
          5920 => x"71",
          5921 => x"5e",
          5922 => x"87",
          5923 => x"5b",
          5924 => x"80",
          5925 => x"06",
          5926 => x"06",
          5927 => x"1d",
          5928 => x"5d",
          5929 => x"ec",
          5930 => x"98",
          5931 => x"e0",
          5932 => x"5e",
          5933 => x"1e",
          5934 => x"81",
          5935 => x"76",
          5936 => x"58",
          5937 => x"81",
          5938 => x"81",
          5939 => x"80",
          5940 => x"ff",
          5941 => x"29",
          5942 => x"5d",
          5943 => x"27",
          5944 => x"e0",
          5945 => x"5e",
          5946 => x"1e",
          5947 => x"81",
          5948 => x"76",
          5949 => x"58",
          5950 => x"81",
          5951 => x"81",
          5952 => x"80",
          5953 => x"ff",
          5954 => x"29",
          5955 => x"5d",
          5956 => x"26",
          5957 => x"eb",
          5958 => x"f9",
          5959 => x"5c",
          5960 => x"1c",
          5961 => x"83",
          5962 => x"84",
          5963 => x"83",
          5964 => x"84",
          5965 => x"5f",
          5966 => x"fd",
          5967 => x"eb",
          5968 => x"b7",
          5969 => x"81",
          5970 => x"11",
          5971 => x"76",
          5972 => x"38",
          5973 => x"83",
          5974 => x"77",
          5975 => x"ff",
          5976 => x"80",
          5977 => x"38",
          5978 => x"83",
          5979 => x"84",
          5980 => x"70",
          5981 => x"ff",
          5982 => x"56",
          5983 => x"eb",
          5984 => x"56",
          5985 => x"bd",
          5986 => x"39",
          5987 => x"33",
          5988 => x"b8",
          5989 => x"11",
          5990 => x"75",
          5991 => x"ca",
          5992 => x"ef",
          5993 => x"81",
          5994 => x"06",
          5995 => x"83",
          5996 => x"70",
          5997 => x"83",
          5998 => x"7a",
          5999 => x"57",
          6000 => x"09",
          6001 => x"b8",
          6002 => x"39",
          6003 => x"75",
          6004 => x"34",
          6005 => x"ff",
          6006 => x"83",
          6007 => x"fc",
          6008 => x"7b",
          6009 => x"83",
          6010 => x"f2",
          6011 => x"7d",
          6012 => x"7a",
          6013 => x"38",
          6014 => x"81",
          6015 => x"83",
          6016 => x"77",
          6017 => x"59",
          6018 => x"26",
          6019 => x"80",
          6020 => x"05",
          6021 => x"f9",
          6022 => x"70",
          6023 => x"34",
          6024 => x"d4",
          6025 => x"39",
          6026 => x"56",
          6027 => x"ba",
          6028 => x"39",
          6029 => x"f9",
          6030 => x"ad",
          6031 => x"f9",
          6032 => x"84",
          6033 => x"83",
          6034 => x"f1",
          6035 => x"0b",
          6036 => x"34",
          6037 => x"83",
          6038 => x"33",
          6039 => x"88",
          6040 => x"34",
          6041 => x"f8",
          6042 => x"a7",
          6043 => x"0d",
          6044 => x"33",
          6045 => x"33",
          6046 => x"80",
          6047 => x"73",
          6048 => x"3f",
          6049 => x"ba",
          6050 => x"3d",
          6051 => x"52",
          6052 => x"ab",
          6053 => x"84",
          6054 => x"85",
          6055 => x"f3",
          6056 => x"bf",
          6057 => x"ff",
          6058 => x"90",
          6059 => x"ff",
          6060 => x"f0",
          6061 => x"55",
          6062 => x"80",
          6063 => x"38",
          6064 => x"75",
          6065 => x"34",
          6066 => x"84",
          6067 => x"8f",
          6068 => x"83",
          6069 => x"54",
          6070 => x"80",
          6071 => x"73",
          6072 => x"30",
          6073 => x"09",
          6074 => x"56",
          6075 => x"72",
          6076 => x"0c",
          6077 => x"54",
          6078 => x"09",
          6079 => x"38",
          6080 => x"83",
          6081 => x"70",
          6082 => x"07",
          6083 => x"79",
          6084 => x"c4",
          6085 => x"80",
          6086 => x"bd",
          6087 => x"bc",
          6088 => x"29",
          6089 => x"a0",
          6090 => x"f9",
          6091 => x"59",
          6092 => x"29",
          6093 => x"ff",
          6094 => x"f8",
          6095 => x"59",
          6096 => x"81",
          6097 => x"38",
          6098 => x"73",
          6099 => x"80",
          6100 => x"87",
          6101 => x"0c",
          6102 => x"88",
          6103 => x"80",
          6104 => x"86",
          6105 => x"08",
          6106 => x"f5",
          6107 => x"81",
          6108 => x"ff",
          6109 => x"81",
          6110 => x"cf",
          6111 => x"83",
          6112 => x"33",
          6113 => x"06",
          6114 => x"16",
          6115 => x"55",
          6116 => x"85",
          6117 => x"81",
          6118 => x"b4",
          6119 => x"f7",
          6120 => x"75",
          6121 => x"5a",
          6122 => x"2e",
          6123 => x"75",
          6124 => x"15",
          6125 => x"ac",
          6126 => x"f7",
          6127 => x"81",
          6128 => x"ff",
          6129 => x"89",
          6130 => x"b3",
          6131 => x"b4",
          6132 => x"2b",
          6133 => x"58",
          6134 => x"83",
          6135 => x"73",
          6136 => x"70",
          6137 => x"32",
          6138 => x"51",
          6139 => x"80",
          6140 => x"38",
          6141 => x"f7",
          6142 => x"09",
          6143 => x"72",
          6144 => x"e4",
          6145 => x"83",
          6146 => x"80",
          6147 => x"e5",
          6148 => x"ec",
          6149 => x"e6",
          6150 => x"f7",
          6151 => x"f7",
          6152 => x"5d",
          6153 => x"5e",
          6154 => x"c0",
          6155 => x"74",
          6156 => x"8d",
          6157 => x"d4",
          6158 => x"73",
          6159 => x"82",
          6160 => x"ca",
          6161 => x"72",
          6162 => x"8b",
          6163 => x"d4",
          6164 => x"73",
          6165 => x"74",
          6166 => x"54",
          6167 => x"2e",
          6168 => x"f7",
          6169 => x"53",
          6170 => x"81",
          6171 => x"81",
          6172 => x"72",
          6173 => x"84",
          6174 => x"f7",
          6175 => x"54",
          6176 => x"84",
          6177 => x"f7",
          6178 => x"e8",
          6179 => x"98",
          6180 => x"54",
          6181 => x"83",
          6182 => x"0b",
          6183 => x"9c",
          6184 => x"e0",
          6185 => x"16",
          6186 => x"06",
          6187 => x"76",
          6188 => x"38",
          6189 => x"e7",
          6190 => x"f7",
          6191 => x"9e",
          6192 => x"9c",
          6193 => x"38",
          6194 => x"83",
          6195 => x"5a",
          6196 => x"83",
          6197 => x"54",
          6198 => x"91",
          6199 => x"14",
          6200 => x"9c",
          6201 => x"7d",
          6202 => x"dc",
          6203 => x"83",
          6204 => x"54",
          6205 => x"2e",
          6206 => x"54",
          6207 => x"92",
          6208 => x"98",
          6209 => x"f8",
          6210 => x"81",
          6211 => x"77",
          6212 => x"38",
          6213 => x"17",
          6214 => x"b8",
          6215 => x"76",
          6216 => x"54",
          6217 => x"83",
          6218 => x"53",
          6219 => x"82",
          6220 => x"81",
          6221 => x"38",
          6222 => x"34",
          6223 => x"fc",
          6224 => x"58",
          6225 => x"80",
          6226 => x"83",
          6227 => x"2e",
          6228 => x"77",
          6229 => x"06",
          6230 => x"7d",
          6231 => x"ed",
          6232 => x"2e",
          6233 => x"79",
          6234 => x"59",
          6235 => x"75",
          6236 => x"54",
          6237 => x"a1",
          6238 => x"2e",
          6239 => x"17",
          6240 => x"06",
          6241 => x"fe",
          6242 => x"27",
          6243 => x"57",
          6244 => x"54",
          6245 => x"e1",
          6246 => x"10",
          6247 => x"05",
          6248 => x"2b",
          6249 => x"f4",
          6250 => x"33",
          6251 => x"78",
          6252 => x"9c",
          6253 => x"e0",
          6254 => x"ea",
          6255 => x"7d",
          6256 => x"a8",
          6257 => x"ff",
          6258 => x"a0",
          6259 => x"ff",
          6260 => x"ff",
          6261 => x"38",
          6262 => x"b8",
          6263 => x"54",
          6264 => x"83",
          6265 => x"82",
          6266 => x"70",
          6267 => x"07",
          6268 => x"7d",
          6269 => x"83",
          6270 => x"06",
          6271 => x"78",
          6272 => x"c6",
          6273 => x"72",
          6274 => x"83",
          6275 => x"70",
          6276 => x"78",
          6277 => x"ba",
          6278 => x"70",
          6279 => x"54",
          6280 => x"27",
          6281 => x"b8",
          6282 => x"72",
          6283 => x"9a",
          6284 => x"84",
          6285 => x"f9",
          6286 => x"81",
          6287 => x"82",
          6288 => x"3f",
          6289 => x"8c",
          6290 => x"0d",
          6291 => x"34",
          6292 => x"f9",
          6293 => x"81",
          6294 => x"38",
          6295 => x"14",
          6296 => x"5b",
          6297 => x"d4",
          6298 => x"c9",
          6299 => x"83",
          6300 => x"34",
          6301 => x"f7",
          6302 => x"ff",
          6303 => x"ca",
          6304 => x"b1",
          6305 => x"ff",
          6306 => x"81",
          6307 => x"96",
          6308 => x"d4",
          6309 => x"81",
          6310 => x"8a",
          6311 => x"ff",
          6312 => x"81",
          6313 => x"06",
          6314 => x"83",
          6315 => x"81",
          6316 => x"c0",
          6317 => x"54",
          6318 => x"27",
          6319 => x"87",
          6320 => x"08",
          6321 => x"0c",
          6322 => x"06",
          6323 => x"39",
          6324 => x"f7",
          6325 => x"f9",
          6326 => x"83",
          6327 => x"73",
          6328 => x"53",
          6329 => x"38",
          6330 => x"e6",
          6331 => x"83",
          6332 => x"83",
          6333 => x"83",
          6334 => x"70",
          6335 => x"33",
          6336 => x"33",
          6337 => x"5e",
          6338 => x"fa",
          6339 => x"82",
          6340 => x"06",
          6341 => x"7a",
          6342 => x"2e",
          6343 => x"79",
          6344 => x"81",
          6345 => x"38",
          6346 => x"ef",
          6347 => x"f0",
          6348 => x"39",
          6349 => x"b8",
          6350 => x"54",
          6351 => x"81",
          6352 => x"b8",
          6353 => x"59",
          6354 => x"80",
          6355 => x"82",
          6356 => x"76",
          6357 => x"54",
          6358 => x"82",
          6359 => x"f7",
          6360 => x"53",
          6361 => x"08",
          6362 => x"83",
          6363 => x"83",
          6364 => x"f6",
          6365 => x"b7",
          6366 => x"81",
          6367 => x"11",
          6368 => x"80",
          6369 => x"38",
          6370 => x"83",
          6371 => x"73",
          6372 => x"ff",
          6373 => x"80",
          6374 => x"38",
          6375 => x"83",
          6376 => x"84",
          6377 => x"70",
          6378 => x"56",
          6379 => x"80",
          6380 => x"38",
          6381 => x"83",
          6382 => x"ff",
          6383 => x"39",
          6384 => x"51",
          6385 => x"3f",
          6386 => x"aa",
          6387 => x"fc",
          6388 => x"14",
          6389 => x"f7",
          6390 => x"de",
          6391 => x"0b",
          6392 => x"34",
          6393 => x"33",
          6394 => x"39",
          6395 => x"81",
          6396 => x"3f",
          6397 => x"04",
          6398 => x"80",
          6399 => x"98",
          6400 => x"02",
          6401 => x"82",
          6402 => x"f4",
          6403 => x"80",
          6404 => x"85",
          6405 => x"98",
          6406 => x"fe",
          6407 => x"34",
          6408 => x"f0",
          6409 => x"87",
          6410 => x"08",
          6411 => x"08",
          6412 => x"90",
          6413 => x"c0",
          6414 => x"53",
          6415 => x"9c",
          6416 => x"73",
          6417 => x"81",
          6418 => x"c0",
          6419 => x"57",
          6420 => x"27",
          6421 => x"81",
          6422 => x"38",
          6423 => x"a4",
          6424 => x"56",
          6425 => x"80",
          6426 => x"56",
          6427 => x"80",
          6428 => x"c0",
          6429 => x"80",
          6430 => x"54",
          6431 => x"9c",
          6432 => x"c0",
          6433 => x"56",
          6434 => x"f6",
          6435 => x"33",
          6436 => x"9c",
          6437 => x"71",
          6438 => x"38",
          6439 => x"2e",
          6440 => x"c0",
          6441 => x"52",
          6442 => x"74",
          6443 => x"72",
          6444 => x"2e",
          6445 => x"80",
          6446 => x"75",
          6447 => x"53",
          6448 => x"38",
          6449 => x"95",
          6450 => x"ba",
          6451 => x"3d",
          6452 => x"17",
          6453 => x"06",
          6454 => x"df",
          6455 => x"83",
          6456 => x"58",
          6457 => x"3f",
          6458 => x"8c",
          6459 => x"0d",
          6460 => x"0d",
          6461 => x"05",
          6462 => x"57",
          6463 => x"83",
          6464 => x"74",
          6465 => x"fc",
          6466 => x"70",
          6467 => x"07",
          6468 => x"58",
          6469 => x"34",
          6470 => x"52",
          6471 => x"34",
          6472 => x"57",
          6473 => x"34",
          6474 => x"34",
          6475 => x"08",
          6476 => x"14",
          6477 => x"98",
          6478 => x"e1",
          6479 => x"0b",
          6480 => x"08",
          6481 => x"0b",
          6482 => x"80",
          6483 => x"80",
          6484 => x"c0",
          6485 => x"83",
          6486 => x"56",
          6487 => x"05",
          6488 => x"98",
          6489 => x"87",
          6490 => x"08",
          6491 => x"2e",
          6492 => x"15",
          6493 => x"98",
          6494 => x"53",
          6495 => x"87",
          6496 => x"fe",
          6497 => x"87",
          6498 => x"08",
          6499 => x"71",
          6500 => x"cf",
          6501 => x"72",
          6502 => x"c7",
          6503 => x"98",
          6504 => x"ce",
          6505 => x"87",
          6506 => x"08",
          6507 => x"98",
          6508 => x"75",
          6509 => x"38",
          6510 => x"87",
          6511 => x"08",
          6512 => x"74",
          6513 => x"72",
          6514 => x"db",
          6515 => x"98",
          6516 => x"ff",
          6517 => x"27",
          6518 => x"72",
          6519 => x"2e",
          6520 => x"76",
          6521 => x"dd",
          6522 => x"ff",
          6523 => x"fe",
          6524 => x"52",
          6525 => x"06",
          6526 => x"38",
          6527 => x"7c",
          6528 => x"56",
          6529 => x"74",
          6530 => x"72",
          6531 => x"54",
          6532 => x"81",
          6533 => x"73",
          6534 => x"38",
          6535 => x"8c",
          6536 => x"0d",
          6537 => x"83",
          6538 => x"58",
          6539 => x"3f",
          6540 => x"8c",
          6541 => x"0d",
          6542 => x"70",
          6543 => x"58",
          6544 => x"a5",
          6545 => x"ff",
          6546 => x"3d",
          6547 => x"84",
          6548 => x"33",
          6549 => x"0b",
          6550 => x"08",
          6551 => x"87",
          6552 => x"06",
          6553 => x"2a",
          6554 => x"56",
          6555 => x"16",
          6556 => x"2a",
          6557 => x"16",
          6558 => x"2a",
          6559 => x"16",
          6560 => x"16",
          6561 => x"f4",
          6562 => x"c6",
          6563 => x"13",
          6564 => x"52",
          6565 => x"97",
          6566 => x"81",
          6567 => x"73",
          6568 => x"55",
          6569 => x"26",
          6570 => x"f4",
          6571 => x"75",
          6572 => x"83",
          6573 => x"56",
          6574 => x"34",
          6575 => x"f4",
          6576 => x"57",
          6577 => x"16",
          6578 => x"86",
          6579 => x"34",
          6580 => x"9c",
          6581 => x"98",
          6582 => x"ce",
          6583 => x"87",
          6584 => x"08",
          6585 => x"98",
          6586 => x"71",
          6587 => x"38",
          6588 => x"87",
          6589 => x"08",
          6590 => x"74",
          6591 => x"72",
          6592 => x"db",
          6593 => x"98",
          6594 => x"ff",
          6595 => x"27",
          6596 => x"72",
          6597 => x"2e",
          6598 => x"87",
          6599 => x"08",
          6600 => x"05",
          6601 => x"98",
          6602 => x"87",
          6603 => x"08",
          6604 => x"2e",
          6605 => x"15",
          6606 => x"98",
          6607 => x"53",
          6608 => x"87",
          6609 => x"ff",
          6610 => x"87",
          6611 => x"08",
          6612 => x"71",
          6613 => x"38",
          6614 => x"ff",
          6615 => x"76",
          6616 => x"38",
          6617 => x"06",
          6618 => x"d8",
          6619 => x"81",
          6620 => x"52",
          6621 => x"77",
          6622 => x"0c",
          6623 => x"04",
          6624 => x"81",
          6625 => x"54",
          6626 => x"ff",
          6627 => x"06",
          6628 => x"80",
          6629 => x"81",
          6630 => x"fc",
          6631 => x"d1",
          6632 => x"84",
          6633 => x"89",
          6634 => x"fb",
          6635 => x"f4",
          6636 => x"80",
          6637 => x"85",
          6638 => x"98",
          6639 => x"fe",
          6640 => x"34",
          6641 => x"f0",
          6642 => x"87",
          6643 => x"08",
          6644 => x"08",
          6645 => x"90",
          6646 => x"c0",
          6647 => x"52",
          6648 => x"9c",
          6649 => x"72",
          6650 => x"81",
          6651 => x"c0",
          6652 => x"52",
          6653 => x"27",
          6654 => x"81",
          6655 => x"38",
          6656 => x"a4",
          6657 => x"53",
          6658 => x"80",
          6659 => x"53",
          6660 => x"80",
          6661 => x"c0",
          6662 => x"80",
          6663 => x"54",
          6664 => x"9c",
          6665 => x"c0",
          6666 => x"53",
          6667 => x"f6",
          6668 => x"33",
          6669 => x"9c",
          6670 => x"70",
          6671 => x"38",
          6672 => x"2e",
          6673 => x"c0",
          6674 => x"51",
          6675 => x"74",
          6676 => x"71",
          6677 => x"2e",
          6678 => x"80",
          6679 => x"72",
          6680 => x"52",
          6681 => x"38",
          6682 => x"16",
          6683 => x"06",
          6684 => x"39",
          6685 => x"83",
          6686 => x"fe",
          6687 => x"82",
          6688 => x"f9",
          6689 => x"b9",
          6690 => x"71",
          6691 => x"70",
          6692 => x"06",
          6693 => x"73",
          6694 => x"81",
          6695 => x"8b",
          6696 => x"2b",
          6697 => x"70",
          6698 => x"33",
          6699 => x"71",
          6700 => x"5c",
          6701 => x"53",
          6702 => x"52",
          6703 => x"80",
          6704 => x"af",
          6705 => x"82",
          6706 => x"12",
          6707 => x"2b",
          6708 => x"07",
          6709 => x"33",
          6710 => x"71",
          6711 => x"90",
          6712 => x"53",
          6713 => x"56",
          6714 => x"24",
          6715 => x"84",
          6716 => x"14",
          6717 => x"2b",
          6718 => x"07",
          6719 => x"88",
          6720 => x"56",
          6721 => x"13",
          6722 => x"ff",
          6723 => x"87",
          6724 => x"b9",
          6725 => x"17",
          6726 => x"85",
          6727 => x"88",
          6728 => x"88",
          6729 => x"59",
          6730 => x"84",
          6731 => x"85",
          6732 => x"b9",
          6733 => x"52",
          6734 => x"13",
          6735 => x"87",
          6736 => x"b9",
          6737 => x"74",
          6738 => x"73",
          6739 => x"84",
          6740 => x"16",
          6741 => x"12",
          6742 => x"2b",
          6743 => x"80",
          6744 => x"2a",
          6745 => x"52",
          6746 => x"75",
          6747 => x"89",
          6748 => x"86",
          6749 => x"13",
          6750 => x"2b",
          6751 => x"07",
          6752 => x"16",
          6753 => x"33",
          6754 => x"07",
          6755 => x"58",
          6756 => x"53",
          6757 => x"84",
          6758 => x"85",
          6759 => x"b9",
          6760 => x"16",
          6761 => x"85",
          6762 => x"8b",
          6763 => x"2b",
          6764 => x"5a",
          6765 => x"86",
          6766 => x"13",
          6767 => x"2b",
          6768 => x"2a",
          6769 => x"52",
          6770 => x"34",
          6771 => x"34",
          6772 => x"08",
          6773 => x"81",
          6774 => x"88",
          6775 => x"ff",
          6776 => x"88",
          6777 => x"54",
          6778 => x"34",
          6779 => x"34",
          6780 => x"08",
          6781 => x"33",
          6782 => x"71",
          6783 => x"83",
          6784 => x"05",
          6785 => x"12",
          6786 => x"2b",
          6787 => x"2b",
          6788 => x"06",
          6789 => x"88",
          6790 => x"53",
          6791 => x"57",
          6792 => x"82",
          6793 => x"83",
          6794 => x"b9",
          6795 => x"17",
          6796 => x"12",
          6797 => x"2b",
          6798 => x"07",
          6799 => x"33",
          6800 => x"71",
          6801 => x"81",
          6802 => x"70",
          6803 => x"52",
          6804 => x"57",
          6805 => x"73",
          6806 => x"14",
          6807 => x"fc",
          6808 => x"82",
          6809 => x"12",
          6810 => x"2b",
          6811 => x"07",
          6812 => x"33",
          6813 => x"71",
          6814 => x"90",
          6815 => x"53",
          6816 => x"57",
          6817 => x"80",
          6818 => x"38",
          6819 => x"13",
          6820 => x"2b",
          6821 => x"80",
          6822 => x"2a",
          6823 => x"76",
          6824 => x"81",
          6825 => x"b9",
          6826 => x"17",
          6827 => x"12",
          6828 => x"2b",
          6829 => x"07",
          6830 => x"14",
          6831 => x"33",
          6832 => x"07",
          6833 => x"57",
          6834 => x"58",
          6835 => x"72",
          6836 => x"75",
          6837 => x"89",
          6838 => x"f9",
          6839 => x"84",
          6840 => x"58",
          6841 => x"2e",
          6842 => x"80",
          6843 => x"77",
          6844 => x"3f",
          6845 => x"04",
          6846 => x"0b",
          6847 => x"0c",
          6848 => x"84",
          6849 => x"82",
          6850 => x"76",
          6851 => x"f4",
          6852 => x"ec",
          6853 => x"fc",
          6854 => x"75",
          6855 => x"81",
          6856 => x"b9",
          6857 => x"76",
          6858 => x"81",
          6859 => x"34",
          6860 => x"08",
          6861 => x"17",
          6862 => x"87",
          6863 => x"b9",
          6864 => x"b9",
          6865 => x"05",
          6866 => x"07",
          6867 => x"ff",
          6868 => x"2a",
          6869 => x"56",
          6870 => x"34",
          6871 => x"34",
          6872 => x"22",
          6873 => x"10",
          6874 => x"08",
          6875 => x"55",
          6876 => x"15",
          6877 => x"83",
          6878 => x"ee",
          6879 => x"0d",
          6880 => x"53",
          6881 => x"72",
          6882 => x"fb",
          6883 => x"82",
          6884 => x"ff",
          6885 => x"51",
          6886 => x"ff",
          6887 => x"fc",
          6888 => x"33",
          6889 => x"71",
          6890 => x"70",
          6891 => x"58",
          6892 => x"ff",
          6893 => x"2e",
          6894 => x"75",
          6895 => x"17",
          6896 => x"12",
          6897 => x"2b",
          6898 => x"ff",
          6899 => x"31",
          6900 => x"ff",
          6901 => x"27",
          6902 => x"5c",
          6903 => x"74",
          6904 => x"70",
          6905 => x"38",
          6906 => x"58",
          6907 => x"85",
          6908 => x"88",
          6909 => x"5a",
          6910 => x"73",
          6911 => x"2e",
          6912 => x"74",
          6913 => x"76",
          6914 => x"11",
          6915 => x"12",
          6916 => x"2b",
          6917 => x"ff",
          6918 => x"56",
          6919 => x"59",
          6920 => x"83",
          6921 => x"80",
          6922 => x"26",
          6923 => x"78",
          6924 => x"2e",
          6925 => x"72",
          6926 => x"88",
          6927 => x"70",
          6928 => x"11",
          6929 => x"80",
          6930 => x"2a",
          6931 => x"56",
          6932 => x"34",
          6933 => x"34",
          6934 => x"08",
          6935 => x"2a",
          6936 => x"82",
          6937 => x"83",
          6938 => x"b9",
          6939 => x"19",
          6940 => x"12",
          6941 => x"2b",
          6942 => x"2b",
          6943 => x"06",
          6944 => x"83",
          6945 => x"70",
          6946 => x"58",
          6947 => x"52",
          6948 => x"12",
          6949 => x"ff",
          6950 => x"83",
          6951 => x"b9",
          6952 => x"54",
          6953 => x"72",
          6954 => x"84",
          6955 => x"70",
          6956 => x"33",
          6957 => x"71",
          6958 => x"83",
          6959 => x"05",
          6960 => x"53",
          6961 => x"15",
          6962 => x"15",
          6963 => x"fc",
          6964 => x"55",
          6965 => x"11",
          6966 => x"33",
          6967 => x"07",
          6968 => x"54",
          6969 => x"70",
          6970 => x"71",
          6971 => x"84",
          6972 => x"70",
          6973 => x"33",
          6974 => x"71",
          6975 => x"83",
          6976 => x"05",
          6977 => x"5a",
          6978 => x"15",
          6979 => x"15",
          6980 => x"fc",
          6981 => x"55",
          6982 => x"11",
          6983 => x"33",
          6984 => x"07",
          6985 => x"54",
          6986 => x"70",
          6987 => x"79",
          6988 => x"84",
          6989 => x"18",
          6990 => x"70",
          6991 => x"0c",
          6992 => x"04",
          6993 => x"87",
          6994 => x"8b",
          6995 => x"2b",
          6996 => x"84",
          6997 => x"18",
          6998 => x"2b",
          6999 => x"2a",
          7000 => x"53",
          7001 => x"84",
          7002 => x"85",
          7003 => x"b9",
          7004 => x"19",
          7005 => x"85",
          7006 => x"8b",
          7007 => x"2b",
          7008 => x"86",
          7009 => x"15",
          7010 => x"2b",
          7011 => x"2a",
          7012 => x"52",
          7013 => x"52",
          7014 => x"34",
          7015 => x"34",
          7016 => x"08",
          7017 => x"81",
          7018 => x"88",
          7019 => x"ff",
          7020 => x"88",
          7021 => x"54",
          7022 => x"34",
          7023 => x"34",
          7024 => x"08",
          7025 => x"51",
          7026 => x"f9",
          7027 => x"84",
          7028 => x"58",
          7029 => x"2e",
          7030 => x"54",
          7031 => x"73",
          7032 => x"0c",
          7033 => x"04",
          7034 => x"91",
          7035 => x"8c",
          7036 => x"8c",
          7037 => x"0d",
          7038 => x"f4",
          7039 => x"fc",
          7040 => x"0b",
          7041 => x"23",
          7042 => x"53",
          7043 => x"ff",
          7044 => x"cc",
          7045 => x"b9",
          7046 => x"76",
          7047 => x"0b",
          7048 => x"84",
          7049 => x"54",
          7050 => x"34",
          7051 => x"15",
          7052 => x"fc",
          7053 => x"86",
          7054 => x"0b",
          7055 => x"84",
          7056 => x"84",
          7057 => x"ff",
          7058 => x"80",
          7059 => x"ff",
          7060 => x"88",
          7061 => x"55",
          7062 => x"17",
          7063 => x"17",
          7064 => x"f8",
          7065 => x"10",
          7066 => x"fc",
          7067 => x"05",
          7068 => x"82",
          7069 => x"0b",
          7070 => x"77",
          7071 => x"2e",
          7072 => x"fe",
          7073 => x"3d",
          7074 => x"41",
          7075 => x"84",
          7076 => x"59",
          7077 => x"61",
          7078 => x"38",
          7079 => x"85",
          7080 => x"80",
          7081 => x"38",
          7082 => x"60",
          7083 => x"7f",
          7084 => x"2a",
          7085 => x"83",
          7086 => x"55",
          7087 => x"ff",
          7088 => x"78",
          7089 => x"70",
          7090 => x"06",
          7091 => x"7a",
          7092 => x"81",
          7093 => x"88",
          7094 => x"75",
          7095 => x"ff",
          7096 => x"10",
          7097 => x"05",
          7098 => x"61",
          7099 => x"81",
          7100 => x"88",
          7101 => x"90",
          7102 => x"2c",
          7103 => x"46",
          7104 => x"43",
          7105 => x"59",
          7106 => x"42",
          7107 => x"85",
          7108 => x"15",
          7109 => x"33",
          7110 => x"07",
          7111 => x"10",
          7112 => x"81",
          7113 => x"98",
          7114 => x"2b",
          7115 => x"53",
          7116 => x"80",
          7117 => x"c9",
          7118 => x"27",
          7119 => x"63",
          7120 => x"62",
          7121 => x"38",
          7122 => x"85",
          7123 => x"1b",
          7124 => x"25",
          7125 => x"63",
          7126 => x"79",
          7127 => x"38",
          7128 => x"33",
          7129 => x"71",
          7130 => x"83",
          7131 => x"11",
          7132 => x"12",
          7133 => x"2b",
          7134 => x"07",
          7135 => x"52",
          7136 => x"58",
          7137 => x"8c",
          7138 => x"1e",
          7139 => x"83",
          7140 => x"8b",
          7141 => x"2b",
          7142 => x"86",
          7143 => x"12",
          7144 => x"2b",
          7145 => x"07",
          7146 => x"14",
          7147 => x"33",
          7148 => x"07",
          7149 => x"59",
          7150 => x"5b",
          7151 => x"5c",
          7152 => x"84",
          7153 => x"85",
          7154 => x"b9",
          7155 => x"17",
          7156 => x"85",
          7157 => x"8b",
          7158 => x"2b",
          7159 => x"86",
          7160 => x"15",
          7161 => x"2b",
          7162 => x"2a",
          7163 => x"52",
          7164 => x"57",
          7165 => x"34",
          7166 => x"34",
          7167 => x"08",
          7168 => x"81",
          7169 => x"88",
          7170 => x"ff",
          7171 => x"88",
          7172 => x"5e",
          7173 => x"34",
          7174 => x"34",
          7175 => x"08",
          7176 => x"11",
          7177 => x"33",
          7178 => x"71",
          7179 => x"74",
          7180 => x"81",
          7181 => x"88",
          7182 => x"88",
          7183 => x"45",
          7184 => x"55",
          7185 => x"34",
          7186 => x"34",
          7187 => x"08",
          7188 => x"33",
          7189 => x"71",
          7190 => x"83",
          7191 => x"05",
          7192 => x"83",
          7193 => x"88",
          7194 => x"88",
          7195 => x"45",
          7196 => x"55",
          7197 => x"1a",
          7198 => x"1a",
          7199 => x"fc",
          7200 => x"82",
          7201 => x"12",
          7202 => x"2b",
          7203 => x"62",
          7204 => x"2b",
          7205 => x"5d",
          7206 => x"05",
          7207 => x"a3",
          7208 => x"fc",
          7209 => x"05",
          7210 => x"1c",
          7211 => x"ff",
          7212 => x"5f",
          7213 => x"81",
          7214 => x"54",
          7215 => x"8c",
          7216 => x"0d",
          7217 => x"f4",
          7218 => x"fc",
          7219 => x"0b",
          7220 => x"23",
          7221 => x"53",
          7222 => x"ff",
          7223 => x"c7",
          7224 => x"b9",
          7225 => x"60",
          7226 => x"0b",
          7227 => x"84",
          7228 => x"5d",
          7229 => x"34",
          7230 => x"1e",
          7231 => x"fc",
          7232 => x"86",
          7233 => x"0b",
          7234 => x"84",
          7235 => x"84",
          7236 => x"ff",
          7237 => x"80",
          7238 => x"ff",
          7239 => x"88",
          7240 => x"5b",
          7241 => x"18",
          7242 => x"18",
          7243 => x"f8",
          7244 => x"10",
          7245 => x"fc",
          7246 => x"05",
          7247 => x"82",
          7248 => x"0b",
          7249 => x"84",
          7250 => x"57",
          7251 => x"38",
          7252 => x"82",
          7253 => x"54",
          7254 => x"fe",
          7255 => x"51",
          7256 => x"84",
          7257 => x"84",
          7258 => x"95",
          7259 => x"61",
          7260 => x"fc",
          7261 => x"2b",
          7262 => x"44",
          7263 => x"33",
          7264 => x"71",
          7265 => x"81",
          7266 => x"70",
          7267 => x"44",
          7268 => x"63",
          7269 => x"81",
          7270 => x"84",
          7271 => x"05",
          7272 => x"57",
          7273 => x"19",
          7274 => x"19",
          7275 => x"fc",
          7276 => x"70",
          7277 => x"33",
          7278 => x"07",
          7279 => x"8f",
          7280 => x"74",
          7281 => x"ff",
          7282 => x"88",
          7283 => x"47",
          7284 => x"5d",
          7285 => x"05",
          7286 => x"ff",
          7287 => x"63",
          7288 => x"84",
          7289 => x"1e",
          7290 => x"34",
          7291 => x"34",
          7292 => x"fc",
          7293 => x"05",
          7294 => x"3f",
          7295 => x"bc",
          7296 => x"31",
          7297 => x"ff",
          7298 => x"fa",
          7299 => x"81",
          7300 => x"76",
          7301 => x"ff",
          7302 => x"17",
          7303 => x"33",
          7304 => x"07",
          7305 => x"10",
          7306 => x"81",
          7307 => x"98",
          7308 => x"2b",
          7309 => x"53",
          7310 => x"45",
          7311 => x"25",
          7312 => x"ff",
          7313 => x"78",
          7314 => x"38",
          7315 => x"8b",
          7316 => x"83",
          7317 => x"5b",
          7318 => x"fc",
          7319 => x"8f",
          7320 => x"f4",
          7321 => x"fc",
          7322 => x"0b",
          7323 => x"23",
          7324 => x"53",
          7325 => x"ff",
          7326 => x"c4",
          7327 => x"b9",
          7328 => x"7e",
          7329 => x"0b",
          7330 => x"84",
          7331 => x"59",
          7332 => x"34",
          7333 => x"1a",
          7334 => x"fc",
          7335 => x"86",
          7336 => x"0b",
          7337 => x"84",
          7338 => x"84",
          7339 => x"ff",
          7340 => x"80",
          7341 => x"ff",
          7342 => x"88",
          7343 => x"57",
          7344 => x"88",
          7345 => x"64",
          7346 => x"84",
          7347 => x"70",
          7348 => x"84",
          7349 => x"05",
          7350 => x"43",
          7351 => x"05",
          7352 => x"83",
          7353 => x"ee",
          7354 => x"24",
          7355 => x"61",
          7356 => x"06",
          7357 => x"27",
          7358 => x"fc",
          7359 => x"80",
          7360 => x"38",
          7361 => x"fb",
          7362 => x"73",
          7363 => x"0c",
          7364 => x"04",
          7365 => x"11",
          7366 => x"33",
          7367 => x"71",
          7368 => x"7a",
          7369 => x"33",
          7370 => x"71",
          7371 => x"83",
          7372 => x"05",
          7373 => x"85",
          7374 => x"88",
          7375 => x"88",
          7376 => x"45",
          7377 => x"58",
          7378 => x"56",
          7379 => x"05",
          7380 => x"85",
          7381 => x"b9",
          7382 => x"17",
          7383 => x"85",
          7384 => x"8b",
          7385 => x"2b",
          7386 => x"86",
          7387 => x"15",
          7388 => x"2b",
          7389 => x"2a",
          7390 => x"48",
          7391 => x"41",
          7392 => x"05",
          7393 => x"87",
          7394 => x"b9",
          7395 => x"70",
          7396 => x"33",
          7397 => x"07",
          7398 => x"06",
          7399 => x"5f",
          7400 => x"7b",
          7401 => x"81",
          7402 => x"b9",
          7403 => x"1f",
          7404 => x"83",
          7405 => x"8b",
          7406 => x"2b",
          7407 => x"73",
          7408 => x"33",
          7409 => x"07",
          7410 => x"5e",
          7411 => x"43",
          7412 => x"76",
          7413 => x"81",
          7414 => x"b9",
          7415 => x"1f",
          7416 => x"12",
          7417 => x"2b",
          7418 => x"07",
          7419 => x"14",
          7420 => x"33",
          7421 => x"07",
          7422 => x"40",
          7423 => x"40",
          7424 => x"78",
          7425 => x"60",
          7426 => x"84",
          7427 => x"70",
          7428 => x"33",
          7429 => x"71",
          7430 => x"66",
          7431 => x"70",
          7432 => x"52",
          7433 => x"05",
          7434 => x"fe",
          7435 => x"84",
          7436 => x"1e",
          7437 => x"83",
          7438 => x"5c",
          7439 => x"39",
          7440 => x"0b",
          7441 => x"0c",
          7442 => x"84",
          7443 => x"82",
          7444 => x"7f",
          7445 => x"f4",
          7446 => x"a4",
          7447 => x"fc",
          7448 => x"76",
          7449 => x"81",
          7450 => x"b9",
          7451 => x"7f",
          7452 => x"81",
          7453 => x"34",
          7454 => x"08",
          7455 => x"15",
          7456 => x"87",
          7457 => x"b9",
          7458 => x"b9",
          7459 => x"05",
          7460 => x"07",
          7461 => x"ff",
          7462 => x"2a",
          7463 => x"5e",
          7464 => x"34",
          7465 => x"34",
          7466 => x"22",
          7467 => x"10",
          7468 => x"08",
          7469 => x"5c",
          7470 => x"1c",
          7471 => x"83",
          7472 => x"51",
          7473 => x"7f",
          7474 => x"39",
          7475 => x"87",
          7476 => x"8b",
          7477 => x"2b",
          7478 => x"84",
          7479 => x"1d",
          7480 => x"2b",
          7481 => x"2a",
          7482 => x"43",
          7483 => x"61",
          7484 => x"63",
          7485 => x"34",
          7486 => x"08",
          7487 => x"11",
          7488 => x"33",
          7489 => x"71",
          7490 => x"74",
          7491 => x"33",
          7492 => x"71",
          7493 => x"70",
          7494 => x"5f",
          7495 => x"56",
          7496 => x"64",
          7497 => x"78",
          7498 => x"34",
          7499 => x"08",
          7500 => x"81",
          7501 => x"88",
          7502 => x"ff",
          7503 => x"88",
          7504 => x"58",
          7505 => x"34",
          7506 => x"34",
          7507 => x"08",
          7508 => x"33",
          7509 => x"71",
          7510 => x"83",
          7511 => x"05",
          7512 => x"12",
          7513 => x"2b",
          7514 => x"2b",
          7515 => x"06",
          7516 => x"88",
          7517 => x"5d",
          7518 => x"5d",
          7519 => x"82",
          7520 => x"83",
          7521 => x"b9",
          7522 => x"1f",
          7523 => x"12",
          7524 => x"2b",
          7525 => x"07",
          7526 => x"33",
          7527 => x"71",
          7528 => x"81",
          7529 => x"70",
          7530 => x"5d",
          7531 => x"5a",
          7532 => x"60",
          7533 => x"81",
          7534 => x"83",
          7535 => x"5b",
          7536 => x"86",
          7537 => x"16",
          7538 => x"2b",
          7539 => x"07",
          7540 => x"18",
          7541 => x"33",
          7542 => x"07",
          7543 => x"5e",
          7544 => x"41",
          7545 => x"1e",
          7546 => x"1e",
          7547 => x"fc",
          7548 => x"84",
          7549 => x"12",
          7550 => x"2b",
          7551 => x"07",
          7552 => x"14",
          7553 => x"33",
          7554 => x"07",
          7555 => x"44",
          7556 => x"5a",
          7557 => x"7c",
          7558 => x"34",
          7559 => x"05",
          7560 => x"fc",
          7561 => x"33",
          7562 => x"71",
          7563 => x"81",
          7564 => x"70",
          7565 => x"5b",
          7566 => x"75",
          7567 => x"16",
          7568 => x"fc",
          7569 => x"70",
          7570 => x"33",
          7571 => x"71",
          7572 => x"74",
          7573 => x"81",
          7574 => x"88",
          7575 => x"83",
          7576 => x"f8",
          7577 => x"63",
          7578 => x"54",
          7579 => x"59",
          7580 => x"7f",
          7581 => x"7b",
          7582 => x"84",
          7583 => x"70",
          7584 => x"81",
          7585 => x"8b",
          7586 => x"2b",
          7587 => x"70",
          7588 => x"33",
          7589 => x"07",
          7590 => x"06",
          7591 => x"5d",
          7592 => x"5b",
          7593 => x"75",
          7594 => x"81",
          7595 => x"b9",
          7596 => x"1f",
          7597 => x"83",
          7598 => x"8b",
          7599 => x"2b",
          7600 => x"86",
          7601 => x"12",
          7602 => x"2b",
          7603 => x"07",
          7604 => x"14",
          7605 => x"33",
          7606 => x"07",
          7607 => x"59",
          7608 => x"5c",
          7609 => x"5d",
          7610 => x"77",
          7611 => x"79",
          7612 => x"84",
          7613 => x"70",
          7614 => x"33",
          7615 => x"71",
          7616 => x"83",
          7617 => x"05",
          7618 => x"87",
          7619 => x"88",
          7620 => x"88",
          7621 => x"5e",
          7622 => x"41",
          7623 => x"16",
          7624 => x"16",
          7625 => x"fc",
          7626 => x"33",
          7627 => x"71",
          7628 => x"81",
          7629 => x"70",
          7630 => x"5c",
          7631 => x"79",
          7632 => x"1a",
          7633 => x"fc",
          7634 => x"82",
          7635 => x"12",
          7636 => x"2b",
          7637 => x"07",
          7638 => x"33",
          7639 => x"71",
          7640 => x"70",
          7641 => x"5c",
          7642 => x"5a",
          7643 => x"79",
          7644 => x"1a",
          7645 => x"fc",
          7646 => x"70",
          7647 => x"33",
          7648 => x"71",
          7649 => x"74",
          7650 => x"33",
          7651 => x"71",
          7652 => x"70",
          7653 => x"5c",
          7654 => x"5a",
          7655 => x"82",
          7656 => x"83",
          7657 => x"b9",
          7658 => x"1f",
          7659 => x"83",
          7660 => x"88",
          7661 => x"57",
          7662 => x"83",
          7663 => x"5a",
          7664 => x"84",
          7665 => x"b5",
          7666 => x"b9",
          7667 => x"84",
          7668 => x"05",
          7669 => x"ff",
          7670 => x"44",
          7671 => x"39",
          7672 => x"87",
          7673 => x"8b",
          7674 => x"2b",
          7675 => x"84",
          7676 => x"1d",
          7677 => x"2b",
          7678 => x"2a",
          7679 => x"43",
          7680 => x"61",
          7681 => x"63",
          7682 => x"34",
          7683 => x"08",
          7684 => x"11",
          7685 => x"33",
          7686 => x"71",
          7687 => x"74",
          7688 => x"33",
          7689 => x"71",
          7690 => x"70",
          7691 => x"41",
          7692 => x"59",
          7693 => x"64",
          7694 => x"7a",
          7695 => x"34",
          7696 => x"08",
          7697 => x"81",
          7698 => x"88",
          7699 => x"ff",
          7700 => x"88",
          7701 => x"42",
          7702 => x"34",
          7703 => x"34",
          7704 => x"08",
          7705 => x"33",
          7706 => x"71",
          7707 => x"83",
          7708 => x"05",
          7709 => x"12",
          7710 => x"2b",
          7711 => x"2b",
          7712 => x"06",
          7713 => x"88",
          7714 => x"5c",
          7715 => x"45",
          7716 => x"82",
          7717 => x"83",
          7718 => x"b9",
          7719 => x"1f",
          7720 => x"12",
          7721 => x"2b",
          7722 => x"07",
          7723 => x"33",
          7724 => x"71",
          7725 => x"81",
          7726 => x"70",
          7727 => x"5f",
          7728 => x"59",
          7729 => x"7d",
          7730 => x"1e",
          7731 => x"ff",
          7732 => x"f3",
          7733 => x"60",
          7734 => x"a1",
          7735 => x"8c",
          7736 => x"ba",
          7737 => x"2e",
          7738 => x"53",
          7739 => x"ba",
          7740 => x"fe",
          7741 => x"73",
          7742 => x"3f",
          7743 => x"7b",
          7744 => x"38",
          7745 => x"f9",
          7746 => x"7a",
          7747 => x"fc",
          7748 => x"76",
          7749 => x"38",
          7750 => x"8a",
          7751 => x"ba",
          7752 => x"3d",
          7753 => x"51",
          7754 => x"84",
          7755 => x"54",
          7756 => x"08",
          7757 => x"38",
          7758 => x"52",
          7759 => x"08",
          7760 => x"bc",
          7761 => x"ba",
          7762 => x"3d",
          7763 => x"ff",
          7764 => x"b9",
          7765 => x"80",
          7766 => x"f8",
          7767 => x"80",
          7768 => x"84",
          7769 => x"fe",
          7770 => x"84",
          7771 => x"55",
          7772 => x"81",
          7773 => x"34",
          7774 => x"08",
          7775 => x"15",
          7776 => x"85",
          7777 => x"b9",
          7778 => x"76",
          7779 => x"81",
          7780 => x"34",
          7781 => x"08",
          7782 => x"22",
          7783 => x"80",
          7784 => x"83",
          7785 => x"70",
          7786 => x"51",
          7787 => x"88",
          7788 => x"89",
          7789 => x"b9",
          7790 => x"10",
          7791 => x"b9",
          7792 => x"f8",
          7793 => x"76",
          7794 => x"81",
          7795 => x"34",
          7796 => x"80",
          7797 => x"38",
          7798 => x"ff",
          7799 => x"8f",
          7800 => x"81",
          7801 => x"26",
          7802 => x"ba",
          7803 => x"52",
          7804 => x"8c",
          7805 => x"0d",
          7806 => x"0d",
          7807 => x"33",
          7808 => x"71",
          7809 => x"38",
          7810 => x"ec",
          7811 => x"8c",
          7812 => x"06",
          7813 => x"38",
          7814 => x"88",
          7815 => x"ba",
          7816 => x"53",
          7817 => x"8c",
          7818 => x"0d",
          7819 => x"0d",
          7820 => x"02",
          7821 => x"05",
          7822 => x"57",
          7823 => x"76",
          7824 => x"38",
          7825 => x"17",
          7826 => x"81",
          7827 => x"55",
          7828 => x"73",
          7829 => x"87",
          7830 => x"0c",
          7831 => x"52",
          7832 => x"8d",
          7833 => x"8c",
          7834 => x"06",
          7835 => x"2e",
          7836 => x"c0",
          7837 => x"54",
          7838 => x"79",
          7839 => x"38",
          7840 => x"80",
          7841 => x"80",
          7842 => x"81",
          7843 => x"74",
          7844 => x"0c",
          7845 => x"04",
          7846 => x"81",
          7847 => x"ff",
          7848 => x"56",
          7849 => x"ff",
          7850 => x"39",
          7851 => x"7c",
          7852 => x"8c",
          7853 => x"33",
          7854 => x"59",
          7855 => x"74",
          7856 => x"84",
          7857 => x"33",
          7858 => x"06",
          7859 => x"73",
          7860 => x"58",
          7861 => x"c0",
          7862 => x"78",
          7863 => x"76",
          7864 => x"3f",
          7865 => x"08",
          7866 => x"55",
          7867 => x"a7",
          7868 => x"98",
          7869 => x"73",
          7870 => x"78",
          7871 => x"74",
          7872 => x"06",
          7873 => x"2e",
          7874 => x"54",
          7875 => x"84",
          7876 => x"8b",
          7877 => x"84",
          7878 => x"19",
          7879 => x"06",
          7880 => x"79",
          7881 => x"ac",
          7882 => x"fc",
          7883 => x"02",
          7884 => x"05",
          7885 => x"05",
          7886 => x"53",
          7887 => x"53",
          7888 => x"87",
          7889 => x"88",
          7890 => x"72",
          7891 => x"83",
          7892 => x"38",
          7893 => x"c0",
          7894 => x"81",
          7895 => x"2e",
          7896 => x"71",
          7897 => x"70",
          7898 => x"38",
          7899 => x"84",
          7900 => x"86",
          7901 => x"88",
          7902 => x"0c",
          7903 => x"8c",
          7904 => x"0d",
          7905 => x"75",
          7906 => x"84",
          7907 => x"86",
          7908 => x"71",
          7909 => x"c0",
          7910 => x"53",
          7911 => x"38",
          7912 => x"81",
          7913 => x"51",
          7914 => x"2e",
          7915 => x"c0",
          7916 => x"55",
          7917 => x"87",
          7918 => x"08",
          7919 => x"38",
          7920 => x"87",
          7921 => x"14",
          7922 => x"82",
          7923 => x"80",
          7924 => x"38",
          7925 => x"06",
          7926 => x"38",
          7927 => x"f6",
          7928 => x"58",
          7929 => x"19",
          7930 => x"56",
          7931 => x"2e",
          7932 => x"a8",
          7933 => x"56",
          7934 => x"81",
          7935 => x"53",
          7936 => x"18",
          7937 => x"a3",
          7938 => x"8c",
          7939 => x"83",
          7940 => x"78",
          7941 => x"0c",
          7942 => x"04",
          7943 => x"18",
          7944 => x"18",
          7945 => x"19",
          7946 => x"fc",
          7947 => x"59",
          7948 => x"08",
          7949 => x"81",
          7950 => x"84",
          7951 => x"83",
          7952 => x"18",
          7953 => x"1a",
          7954 => x"1a",
          7955 => x"8c",
          7956 => x"56",
          7957 => x"27",
          7958 => x"82",
          7959 => x"74",
          7960 => x"81",
          7961 => x"38",
          7962 => x"1b",
          7963 => x"81",
          7964 => x"fc",
          7965 => x"78",
          7966 => x"75",
          7967 => x"81",
          7968 => x"38",
          7969 => x"57",
          7970 => x"09",
          7971 => x"ee",
          7972 => x"5a",
          7973 => x"56",
          7974 => x"70",
          7975 => x"34",
          7976 => x"76",
          7977 => x"d5",
          7978 => x"19",
          7979 => x"0b",
          7980 => x"34",
          7981 => x"34",
          7982 => x"b9",
          7983 => x"e1",
          7984 => x"34",
          7985 => x"bb",
          7986 => x"f2",
          7987 => x"19",
          7988 => x"0b",
          7989 => x"34",
          7990 => x"84",
          7991 => x"80",
          7992 => x"9f",
          7993 => x"18",
          7994 => x"84",
          7995 => x"74",
          7996 => x"7a",
          7997 => x"34",
          7998 => x"56",
          7999 => x"19",
          8000 => x"2a",
          8001 => x"a3",
          8002 => x"18",
          8003 => x"84",
          8004 => x"7a",
          8005 => x"74",
          8006 => x"34",
          8007 => x"56",
          8008 => x"19",
          8009 => x"2a",
          8010 => x"a7",
          8011 => x"18",
          8012 => x"70",
          8013 => x"5b",
          8014 => x"53",
          8015 => x"18",
          8016 => x"e8",
          8017 => x"19",
          8018 => x"80",
          8019 => x"33",
          8020 => x"3f",
          8021 => x"08",
          8022 => x"b7",
          8023 => x"39",
          8024 => x"60",
          8025 => x"59",
          8026 => x"76",
          8027 => x"9c",
          8028 => x"26",
          8029 => x"58",
          8030 => x"8c",
          8031 => x"0d",
          8032 => x"33",
          8033 => x"82",
          8034 => x"38",
          8035 => x"82",
          8036 => x"81",
          8037 => x"06",
          8038 => x"81",
          8039 => x"89",
          8040 => x"08",
          8041 => x"80",
          8042 => x"08",
          8043 => x"38",
          8044 => x"5c",
          8045 => x"09",
          8046 => x"de",
          8047 => x"78",
          8048 => x"52",
          8049 => x"51",
          8050 => x"84",
          8051 => x"80",
          8052 => x"ff",
          8053 => x"78",
          8054 => x"7a",
          8055 => x"79",
          8056 => x"17",
          8057 => x"81",
          8058 => x"2a",
          8059 => x"05",
          8060 => x"59",
          8061 => x"79",
          8062 => x"80",
          8063 => x"33",
          8064 => x"5d",
          8065 => x"09",
          8066 => x"b5",
          8067 => x"78",
          8068 => x"52",
          8069 => x"51",
          8070 => x"84",
          8071 => x"80",
          8072 => x"ff",
          8073 => x"78",
          8074 => x"79",
          8075 => x"7a",
          8076 => x"17",
          8077 => x"70",
          8078 => x"07",
          8079 => x"71",
          8080 => x"5d",
          8081 => x"79",
          8082 => x"76",
          8083 => x"84",
          8084 => x"8f",
          8085 => x"75",
          8086 => x"18",
          8087 => x"b4",
          8088 => x"2e",
          8089 => x"0b",
          8090 => x"71",
          8091 => x"7b",
          8092 => x"81",
          8093 => x"38",
          8094 => x"53",
          8095 => x"81",
          8096 => x"f7",
          8097 => x"ba",
          8098 => x"2e",
          8099 => x"59",
          8100 => x"b4",
          8101 => x"fd",
          8102 => x"10",
          8103 => x"77",
          8104 => x"81",
          8105 => x"33",
          8106 => x"07",
          8107 => x"0c",
          8108 => x"3d",
          8109 => x"83",
          8110 => x"06",
          8111 => x"75",
          8112 => x"18",
          8113 => x"b4",
          8114 => x"2e",
          8115 => x"0b",
          8116 => x"71",
          8117 => x"7c",
          8118 => x"81",
          8119 => x"38",
          8120 => x"53",
          8121 => x"81",
          8122 => x"f6",
          8123 => x"ba",
          8124 => x"2e",
          8125 => x"59",
          8126 => x"b4",
          8127 => x"fc",
          8128 => x"82",
          8129 => x"06",
          8130 => x"05",
          8131 => x"82",
          8132 => x"90",
          8133 => x"2b",
          8134 => x"33",
          8135 => x"88",
          8136 => x"71",
          8137 => x"fe",
          8138 => x"84",
          8139 => x"41",
          8140 => x"5a",
          8141 => x"0d",
          8142 => x"b4",
          8143 => x"b8",
          8144 => x"81",
          8145 => x"5c",
          8146 => x"81",
          8147 => x"8c",
          8148 => x"09",
          8149 => x"be",
          8150 => x"8c",
          8151 => x"34",
          8152 => x"a8",
          8153 => x"84",
          8154 => x"5b",
          8155 => x"18",
          8156 => x"84",
          8157 => x"33",
          8158 => x"2e",
          8159 => x"fd",
          8160 => x"54",
          8161 => x"a0",
          8162 => x"53",
          8163 => x"17",
          8164 => x"98",
          8165 => x"fd",
          8166 => x"54",
          8167 => x"53",
          8168 => x"53",
          8169 => x"52",
          8170 => x"3f",
          8171 => x"08",
          8172 => x"81",
          8173 => x"38",
          8174 => x"08",
          8175 => x"b4",
          8176 => x"18",
          8177 => x"7c",
          8178 => x"27",
          8179 => x"17",
          8180 => x"82",
          8181 => x"38",
          8182 => x"08",
          8183 => x"39",
          8184 => x"17",
          8185 => x"17",
          8186 => x"18",
          8187 => x"f5",
          8188 => x"5a",
          8189 => x"08",
          8190 => x"81",
          8191 => x"38",
          8192 => x"08",
          8193 => x"b4",
          8194 => x"18",
          8195 => x"ba",
          8196 => x"5e",
          8197 => x"08",
          8198 => x"38",
          8199 => x"55",
          8200 => x"09",
          8201 => x"b8",
          8202 => x"b4",
          8203 => x"18",
          8204 => x"7b",
          8205 => x"33",
          8206 => x"3f",
          8207 => x"a0",
          8208 => x"b4",
          8209 => x"b8",
          8210 => x"81",
          8211 => x"5e",
          8212 => x"81",
          8213 => x"8c",
          8214 => x"09",
          8215 => x"cb",
          8216 => x"8c",
          8217 => x"34",
          8218 => x"a8",
          8219 => x"84",
          8220 => x"5b",
          8221 => x"18",
          8222 => x"91",
          8223 => x"33",
          8224 => x"2e",
          8225 => x"fb",
          8226 => x"54",
          8227 => x"a0",
          8228 => x"53",
          8229 => x"17",
          8230 => x"90",
          8231 => x"fa",
          8232 => x"54",
          8233 => x"a0",
          8234 => x"53",
          8235 => x"17",
          8236 => x"f8",
          8237 => x"39",
          8238 => x"f9",
          8239 => x"9f",
          8240 => x"0d",
          8241 => x"5d",
          8242 => x"58",
          8243 => x"9c",
          8244 => x"1a",
          8245 => x"38",
          8246 => x"74",
          8247 => x"38",
          8248 => x"81",
          8249 => x"81",
          8250 => x"38",
          8251 => x"8c",
          8252 => x"0d",
          8253 => x"2a",
          8254 => x"05",
          8255 => x"b4",
          8256 => x"5c",
          8257 => x"86",
          8258 => x"19",
          8259 => x"5d",
          8260 => x"09",
          8261 => x"fa",
          8262 => x"77",
          8263 => x"52",
          8264 => x"51",
          8265 => x"84",
          8266 => x"80",
          8267 => x"ff",
          8268 => x"77",
          8269 => x"79",
          8270 => x"b0",
          8271 => x"83",
          8272 => x"05",
          8273 => x"ff",
          8274 => x"76",
          8275 => x"76",
          8276 => x"79",
          8277 => x"81",
          8278 => x"34",
          8279 => x"8c",
          8280 => x"0d",
          8281 => x"2e",
          8282 => x"fe",
          8283 => x"87",
          8284 => x"08",
          8285 => x"0b",
          8286 => x"58",
          8287 => x"2e",
          8288 => x"83",
          8289 => x"5b",
          8290 => x"2e",
          8291 => x"84",
          8292 => x"54",
          8293 => x"19",
          8294 => x"33",
          8295 => x"3f",
          8296 => x"08",
          8297 => x"38",
          8298 => x"5a",
          8299 => x"0c",
          8300 => x"fe",
          8301 => x"82",
          8302 => x"06",
          8303 => x"11",
          8304 => x"70",
          8305 => x"0a",
          8306 => x"0a",
          8307 => x"57",
          8308 => x"7d",
          8309 => x"2a",
          8310 => x"1d",
          8311 => x"2a",
          8312 => x"1d",
          8313 => x"2a",
          8314 => x"1d",
          8315 => x"83",
          8316 => x"e8",
          8317 => x"2a",
          8318 => x"2a",
          8319 => x"05",
          8320 => x"59",
          8321 => x"78",
          8322 => x"80",
          8323 => x"33",
          8324 => x"5d",
          8325 => x"09",
          8326 => x"d4",
          8327 => x"77",
          8328 => x"52",
          8329 => x"51",
          8330 => x"84",
          8331 => x"80",
          8332 => x"ff",
          8333 => x"77",
          8334 => x"7b",
          8335 => x"ac",
          8336 => x"ff",
          8337 => x"05",
          8338 => x"81",
          8339 => x"57",
          8340 => x"80",
          8341 => x"7a",
          8342 => x"f0",
          8343 => x"8f",
          8344 => x"56",
          8345 => x"34",
          8346 => x"1a",
          8347 => x"2a",
          8348 => x"05",
          8349 => x"b4",
          8350 => x"5f",
          8351 => x"83",
          8352 => x"54",
          8353 => x"19",
          8354 => x"1a",
          8355 => x"f0",
          8356 => x"58",
          8357 => x"08",
          8358 => x"81",
          8359 => x"38",
          8360 => x"08",
          8361 => x"b4",
          8362 => x"a8",
          8363 => x"a0",
          8364 => x"ba",
          8365 => x"5c",
          8366 => x"7a",
          8367 => x"82",
          8368 => x"74",
          8369 => x"e4",
          8370 => x"75",
          8371 => x"81",
          8372 => x"ee",
          8373 => x"ba",
          8374 => x"2e",
          8375 => x"56",
          8376 => x"b4",
          8377 => x"fc",
          8378 => x"83",
          8379 => x"b8",
          8380 => x"2a",
          8381 => x"8f",
          8382 => x"2a",
          8383 => x"f0",
          8384 => x"06",
          8385 => x"74",
          8386 => x"0b",
          8387 => x"fc",
          8388 => x"54",
          8389 => x"19",
          8390 => x"1a",
          8391 => x"ef",
          8392 => x"5a",
          8393 => x"08",
          8394 => x"81",
          8395 => x"38",
          8396 => x"08",
          8397 => x"b4",
          8398 => x"a8",
          8399 => x"a0",
          8400 => x"ba",
          8401 => x"59",
          8402 => x"77",
          8403 => x"38",
          8404 => x"55",
          8405 => x"09",
          8406 => x"bd",
          8407 => x"76",
          8408 => x"52",
          8409 => x"51",
          8410 => x"7b",
          8411 => x"39",
          8412 => x"53",
          8413 => x"53",
          8414 => x"52",
          8415 => x"3f",
          8416 => x"ba",
          8417 => x"2e",
          8418 => x"fd",
          8419 => x"ba",
          8420 => x"1a",
          8421 => x"08",
          8422 => x"08",
          8423 => x"08",
          8424 => x"08",
          8425 => x"5f",
          8426 => x"fc",
          8427 => x"19",
          8428 => x"82",
          8429 => x"06",
          8430 => x"81",
          8431 => x"53",
          8432 => x"19",
          8433 => x"e4",
          8434 => x"fc",
          8435 => x"54",
          8436 => x"19",
          8437 => x"1a",
          8438 => x"ed",
          8439 => x"5a",
          8440 => x"08",
          8441 => x"81",
          8442 => x"38",
          8443 => x"08",
          8444 => x"b4",
          8445 => x"a8",
          8446 => x"a0",
          8447 => x"ba",
          8448 => x"5f",
          8449 => x"7d",
          8450 => x"38",
          8451 => x"55",
          8452 => x"09",
          8453 => x"fa",
          8454 => x"7c",
          8455 => x"52",
          8456 => x"51",
          8457 => x"7b",
          8458 => x"39",
          8459 => x"1c",
          8460 => x"81",
          8461 => x"ec",
          8462 => x"58",
          8463 => x"7b",
          8464 => x"fe",
          8465 => x"7c",
          8466 => x"06",
          8467 => x"76",
          8468 => x"76",
          8469 => x"79",
          8470 => x"f9",
          8471 => x"58",
          8472 => x"7b",
          8473 => x"83",
          8474 => x"05",
          8475 => x"11",
          8476 => x"2b",
          8477 => x"7f",
          8478 => x"07",
          8479 => x"5d",
          8480 => x"34",
          8481 => x"56",
          8482 => x"34",
          8483 => x"5a",
          8484 => x"34",
          8485 => x"5b",
          8486 => x"34",
          8487 => x"f6",
          8488 => x"7e",
          8489 => x"5c",
          8490 => x"8a",
          8491 => x"08",
          8492 => x"2e",
          8493 => x"76",
          8494 => x"27",
          8495 => x"94",
          8496 => x"56",
          8497 => x"2e",
          8498 => x"76",
          8499 => x"93",
          8500 => x"81",
          8501 => x"19",
          8502 => x"89",
          8503 => x"75",
          8504 => x"b2",
          8505 => x"79",
          8506 => x"3f",
          8507 => x"08",
          8508 => x"d0",
          8509 => x"84",
          8510 => x"81",
          8511 => x"84",
          8512 => x"09",
          8513 => x"72",
          8514 => x"70",
          8515 => x"51",
          8516 => x"82",
          8517 => x"77",
          8518 => x"06",
          8519 => x"73",
          8520 => x"ba",
          8521 => x"3d",
          8522 => x"57",
          8523 => x"84",
          8524 => x"58",
          8525 => x"52",
          8526 => x"a4",
          8527 => x"74",
          8528 => x"08",
          8529 => x"84",
          8530 => x"55",
          8531 => x"08",
          8532 => x"38",
          8533 => x"84",
          8534 => x"26",
          8535 => x"57",
          8536 => x"81",
          8537 => x"19",
          8538 => x"83",
          8539 => x"75",
          8540 => x"ef",
          8541 => x"58",
          8542 => x"08",
          8543 => x"a0",
          8544 => x"8c",
          8545 => x"30",
          8546 => x"80",
          8547 => x"07",
          8548 => x"08",
          8549 => x"55",
          8550 => x"85",
          8551 => x"8c",
          8552 => x"9a",
          8553 => x"08",
          8554 => x"27",
          8555 => x"73",
          8556 => x"27",
          8557 => x"73",
          8558 => x"fe",
          8559 => x"80",
          8560 => x"38",
          8561 => x"52",
          8562 => x"f5",
          8563 => x"8c",
          8564 => x"8c",
          8565 => x"84",
          8566 => x"07",
          8567 => x"58",
          8568 => x"c4",
          8569 => x"e3",
          8570 => x"1a",
          8571 => x"08",
          8572 => x"1a",
          8573 => x"74",
          8574 => x"38",
          8575 => x"1a",
          8576 => x"33",
          8577 => x"79",
          8578 => x"75",
          8579 => x"ba",
          8580 => x"3d",
          8581 => x"0b",
          8582 => x"0c",
          8583 => x"04",
          8584 => x"08",
          8585 => x"39",
          8586 => x"ff",
          8587 => x"53",
          8588 => x"51",
          8589 => x"84",
          8590 => x"55",
          8591 => x"84",
          8592 => x"84",
          8593 => x"8c",
          8594 => x"ff",
          8595 => x"2e",
          8596 => x"81",
          8597 => x"39",
          8598 => x"7a",
          8599 => x"59",
          8600 => x"f0",
          8601 => x"80",
          8602 => x"9f",
          8603 => x"80",
          8604 => x"90",
          8605 => x"18",
          8606 => x"80",
          8607 => x"33",
          8608 => x"26",
          8609 => x"73",
          8610 => x"82",
          8611 => x"22",
          8612 => x"79",
          8613 => x"ac",
          8614 => x"19",
          8615 => x"19",
          8616 => x"08",
          8617 => x"72",
          8618 => x"38",
          8619 => x"13",
          8620 => x"73",
          8621 => x"17",
          8622 => x"19",
          8623 => x"75",
          8624 => x"0c",
          8625 => x"04",
          8626 => x"ba",
          8627 => x"3d",
          8628 => x"17",
          8629 => x"80",
          8630 => x"38",
          8631 => x"70",
          8632 => x"59",
          8633 => x"a5",
          8634 => x"08",
          8635 => x"fe",
          8636 => x"80",
          8637 => x"27",
          8638 => x"17",
          8639 => x"29",
          8640 => x"05",
          8641 => x"98",
          8642 => x"91",
          8643 => x"77",
          8644 => x"3f",
          8645 => x"08",
          8646 => x"8c",
          8647 => x"a4",
          8648 => x"84",
          8649 => x"27",
          8650 => x"9c",
          8651 => x"84",
          8652 => x"73",
          8653 => x"38",
          8654 => x"54",
          8655 => x"cd",
          8656 => x"39",
          8657 => x"ba",
          8658 => x"3d",
          8659 => x"3d",
          8660 => x"08",
          8661 => x"a0",
          8662 => x"57",
          8663 => x"7a",
          8664 => x"80",
          8665 => x"0c",
          8666 => x"55",
          8667 => x"80",
          8668 => x"79",
          8669 => x"5b",
          8670 => x"81",
          8671 => x"08",
          8672 => x"a9",
          8673 => x"2a",
          8674 => x"57",
          8675 => x"27",
          8676 => x"77",
          8677 => x"79",
          8678 => x"78",
          8679 => x"9c",
          8680 => x"56",
          8681 => x"8c",
          8682 => x"0d",
          8683 => x"18",
          8684 => x"22",
          8685 => x"89",
          8686 => x"7b",
          8687 => x"52",
          8688 => x"9c",
          8689 => x"8c",
          8690 => x"56",
          8691 => x"ba",
          8692 => x"d0",
          8693 => x"84",
          8694 => x"ff",
          8695 => x"9c",
          8696 => x"ba",
          8697 => x"82",
          8698 => x"80",
          8699 => x"38",
          8700 => x"52",
          8701 => x"a7",
          8702 => x"8c",
          8703 => x"56",
          8704 => x"08",
          8705 => x"9c",
          8706 => x"84",
          8707 => x"81",
          8708 => x"38",
          8709 => x"ba",
          8710 => x"2e",
          8711 => x"84",
          8712 => x"83",
          8713 => x"58",
          8714 => x"38",
          8715 => x"1a",
          8716 => x"59",
          8717 => x"75",
          8718 => x"38",
          8719 => x"76",
          8720 => x"1b",
          8721 => x"5e",
          8722 => x"0c",
          8723 => x"84",
          8724 => x"55",
          8725 => x"81",
          8726 => x"ff",
          8727 => x"f4",
          8728 => x"8a",
          8729 => x"75",
          8730 => x"80",
          8731 => x"75",
          8732 => x"52",
          8733 => x"51",
          8734 => x"84",
          8735 => x"80",
          8736 => x"16",
          8737 => x"7a",
          8738 => x"84",
          8739 => x"8c",
          8740 => x"0d",
          8741 => x"b4",
          8742 => x"b8",
          8743 => x"81",
          8744 => x"56",
          8745 => x"84",
          8746 => x"80",
          8747 => x"ba",
          8748 => x"1a",
          8749 => x"08",
          8750 => x"31",
          8751 => x"1a",
          8752 => x"e8",
          8753 => x"33",
          8754 => x"2e",
          8755 => x"fe",
          8756 => x"54",
          8757 => x"a0",
          8758 => x"53",
          8759 => x"19",
          8760 => x"c8",
          8761 => x"39",
          8762 => x"55",
          8763 => x"ff",
          8764 => x"76",
          8765 => x"06",
          8766 => x"94",
          8767 => x"1d",
          8768 => x"fe",
          8769 => x"80",
          8770 => x"27",
          8771 => x"8a",
          8772 => x"71",
          8773 => x"08",
          8774 => x"0c",
          8775 => x"39",
          8776 => x"ba",
          8777 => x"3d",
          8778 => x"3d",
          8779 => x"41",
          8780 => x"08",
          8781 => x"ff",
          8782 => x"08",
          8783 => x"75",
          8784 => x"d2",
          8785 => x"5f",
          8786 => x"58",
          8787 => x"76",
          8788 => x"38",
          8789 => x"78",
          8790 => x"78",
          8791 => x"06",
          8792 => x"81",
          8793 => x"b8",
          8794 => x"19",
          8795 => x"bd",
          8796 => x"8c",
          8797 => x"85",
          8798 => x"81",
          8799 => x"1a",
          8800 => x"76",
          8801 => x"9c",
          8802 => x"33",
          8803 => x"80",
          8804 => x"38",
          8805 => x"bf",
          8806 => x"ff",
          8807 => x"60",
          8808 => x"76",
          8809 => x"70",
          8810 => x"32",
          8811 => x"80",
          8812 => x"25",
          8813 => x"45",
          8814 => x"93",
          8815 => x"df",
          8816 => x"61",
          8817 => x"bf",
          8818 => x"2e",
          8819 => x"81",
          8820 => x"52",
          8821 => x"f6",
          8822 => x"8c",
          8823 => x"ba",
          8824 => x"b2",
          8825 => x"08",
          8826 => x"dc",
          8827 => x"ba",
          8828 => x"3d",
          8829 => x"54",
          8830 => x"53",
          8831 => x"19",
          8832 => x"a8",
          8833 => x"84",
          8834 => x"78",
          8835 => x"06",
          8836 => x"84",
          8837 => x"83",
          8838 => x"19",
          8839 => x"08",
          8840 => x"8c",
          8841 => x"7a",
          8842 => x"27",
          8843 => x"82",
          8844 => x"60",
          8845 => x"81",
          8846 => x"38",
          8847 => x"19",
          8848 => x"08",
          8849 => x"52",
          8850 => x"51",
          8851 => x"77",
          8852 => x"39",
          8853 => x"09",
          8854 => x"e7",
          8855 => x"2a",
          8856 => x"7a",
          8857 => x"38",
          8858 => x"77",
          8859 => x"70",
          8860 => x"7f",
          8861 => x"59",
          8862 => x"7d",
          8863 => x"81",
          8864 => x"5d",
          8865 => x"81",
          8866 => x"2e",
          8867 => x"fe",
          8868 => x"39",
          8869 => x"0b",
          8870 => x"7a",
          8871 => x"0c",
          8872 => x"04",
          8873 => x"df",
          8874 => x"33",
          8875 => x"2e",
          8876 => x"cb",
          8877 => x"08",
          8878 => x"9a",
          8879 => x"88",
          8880 => x"56",
          8881 => x"b7",
          8882 => x"70",
          8883 => x"8d",
          8884 => x"51",
          8885 => x"58",
          8886 => x"8c",
          8887 => x"05",
          8888 => x"71",
          8889 => x"2b",
          8890 => x"56",
          8891 => x"80",
          8892 => x"81",
          8893 => x"87",
          8894 => x"61",
          8895 => x"42",
          8896 => x"81",
          8897 => x"17",
          8898 => x"27",
          8899 => x"33",
          8900 => x"81",
          8901 => x"77",
          8902 => x"38",
          8903 => x"26",
          8904 => x"79",
          8905 => x"43",
          8906 => x"ff",
          8907 => x"ff",
          8908 => x"fd",
          8909 => x"83",
          8910 => x"ca",
          8911 => x"55",
          8912 => x"7c",
          8913 => x"55",
          8914 => x"81",
          8915 => x"80",
          8916 => x"70",
          8917 => x"33",
          8918 => x"70",
          8919 => x"ff",
          8920 => x"59",
          8921 => x"74",
          8922 => x"81",
          8923 => x"ac",
          8924 => x"84",
          8925 => x"94",
          8926 => x"ef",
          8927 => x"70",
          8928 => x"80",
          8929 => x"f5",
          8930 => x"ba",
          8931 => x"84",
          8932 => x"82",
          8933 => x"ff",
          8934 => x"ff",
          8935 => x"0c",
          8936 => x"98",
          8937 => x"80",
          8938 => x"08",
          8939 => x"cc",
          8940 => x"33",
          8941 => x"74",
          8942 => x"81",
          8943 => x"38",
          8944 => x"53",
          8945 => x"81",
          8946 => x"dc",
          8947 => x"ba",
          8948 => x"2e",
          8949 => x"56",
          8950 => x"b4",
          8951 => x"5a",
          8952 => x"38",
          8953 => x"70",
          8954 => x"76",
          8955 => x"99",
          8956 => x"33",
          8957 => x"81",
          8958 => x"58",
          8959 => x"34",
          8960 => x"2e",
          8961 => x"75",
          8962 => x"06",
          8963 => x"2e",
          8964 => x"74",
          8965 => x"75",
          8966 => x"e5",
          8967 => x"38",
          8968 => x"58",
          8969 => x"81",
          8970 => x"80",
          8971 => x"70",
          8972 => x"33",
          8973 => x"70",
          8974 => x"ff",
          8975 => x"5d",
          8976 => x"74",
          8977 => x"cd",
          8978 => x"33",
          8979 => x"76",
          8980 => x"0b",
          8981 => x"57",
          8982 => x"05",
          8983 => x"70",
          8984 => x"33",
          8985 => x"ff",
          8986 => x"42",
          8987 => x"2e",
          8988 => x"75",
          8989 => x"38",
          8990 => x"ff",
          8991 => x"0c",
          8992 => x"51",
          8993 => x"84",
          8994 => x"5a",
          8995 => x"08",
          8996 => x"8f",
          8997 => x"ba",
          8998 => x"3d",
          8999 => x"54",
          9000 => x"53",
          9001 => x"1b",
          9002 => x"80",
          9003 => x"84",
          9004 => x"78",
          9005 => x"06",
          9006 => x"84",
          9007 => x"83",
          9008 => x"1b",
          9009 => x"08",
          9010 => x"8c",
          9011 => x"78",
          9012 => x"27",
          9013 => x"82",
          9014 => x"79",
          9015 => x"81",
          9016 => x"38",
          9017 => x"1b",
          9018 => x"08",
          9019 => x"52",
          9020 => x"51",
          9021 => x"77",
          9022 => x"39",
          9023 => x"e4",
          9024 => x"33",
          9025 => x"81",
          9026 => x"60",
          9027 => x"76",
          9028 => x"06",
          9029 => x"2e",
          9030 => x"19",
          9031 => x"bf",
          9032 => x"1f",
          9033 => x"05",
          9034 => x"5f",
          9035 => x"af",
          9036 => x"55",
          9037 => x"52",
          9038 => x"92",
          9039 => x"8c",
          9040 => x"ba",
          9041 => x"2e",
          9042 => x"fe",
          9043 => x"80",
          9044 => x"38",
          9045 => x"ff",
          9046 => x"0c",
          9047 => x"8d",
          9048 => x"7e",
          9049 => x"81",
          9050 => x"8c",
          9051 => x"1a",
          9052 => x"33",
          9053 => x"07",
          9054 => x"76",
          9055 => x"78",
          9056 => x"06",
          9057 => x"05",
          9058 => x"77",
          9059 => x"e6",
          9060 => x"79",
          9061 => x"33",
          9062 => x"88",
          9063 => x"42",
          9064 => x"2e",
          9065 => x"79",
          9066 => x"ff",
          9067 => x"51",
          9068 => x"3f",
          9069 => x"08",
          9070 => x"05",
          9071 => x"43",
          9072 => x"56",
          9073 => x"3f",
          9074 => x"8c",
          9075 => x"81",
          9076 => x"38",
          9077 => x"18",
          9078 => x"27",
          9079 => x"78",
          9080 => x"2a",
          9081 => x"59",
          9082 => x"92",
          9083 => x"2e",
          9084 => x"10",
          9085 => x"22",
          9086 => x"fe",
          9087 => x"1d",
          9088 => x"06",
          9089 => x"ae",
          9090 => x"84",
          9091 => x"93",
          9092 => x"76",
          9093 => x"2e",
          9094 => x"81",
          9095 => x"94",
          9096 => x"0d",
          9097 => x"70",
          9098 => x"81",
          9099 => x"5a",
          9100 => x"56",
          9101 => x"38",
          9102 => x"08",
          9103 => x"57",
          9104 => x"2e",
          9105 => x"1d",
          9106 => x"70",
          9107 => x"5d",
          9108 => x"95",
          9109 => x"5b",
          9110 => x"7b",
          9111 => x"75",
          9112 => x"57",
          9113 => x"81",
          9114 => x"ff",
          9115 => x"ef",
          9116 => x"db",
          9117 => x"81",
          9118 => x"76",
          9119 => x"aa",
          9120 => x"0b",
          9121 => x"81",
          9122 => x"40",
          9123 => x"08",
          9124 => x"8b",
          9125 => x"57",
          9126 => x"81",
          9127 => x"76",
          9128 => x"58",
          9129 => x"55",
          9130 => x"85",
          9131 => x"c2",
          9132 => x"22",
          9133 => x"80",
          9134 => x"74",
          9135 => x"56",
          9136 => x"81",
          9137 => x"07",
          9138 => x"70",
          9139 => x"06",
          9140 => x"81",
          9141 => x"56",
          9142 => x"2e",
          9143 => x"84",
          9144 => x"57",
          9145 => x"77",
          9146 => x"38",
          9147 => x"74",
          9148 => x"02",
          9149 => x"cf",
          9150 => x"76",
          9151 => x"06",
          9152 => x"27",
          9153 => x"15",
          9154 => x"34",
          9155 => x"19",
          9156 => x"59",
          9157 => x"e3",
          9158 => x"59",
          9159 => x"34",
          9160 => x"56",
          9161 => x"a0",
          9162 => x"55",
          9163 => x"98",
          9164 => x"56",
          9165 => x"88",
          9166 => x"1a",
          9167 => x"57",
          9168 => x"09",
          9169 => x"38",
          9170 => x"a0",
          9171 => x"26",
          9172 => x"3d",
          9173 => x"05",
          9174 => x"33",
          9175 => x"74",
          9176 => x"76",
          9177 => x"38",
          9178 => x"8f",
          9179 => x"8c",
          9180 => x"81",
          9181 => x"e3",
          9182 => x"91",
          9183 => x"7a",
          9184 => x"82",
          9185 => x"ba",
          9186 => x"84",
          9187 => x"84",
          9188 => x"06",
          9189 => x"02",
          9190 => x"33",
          9191 => x"7d",
          9192 => x"05",
          9193 => x"33",
          9194 => x"81",
          9195 => x"5f",
          9196 => x"80",
          9197 => x"8d",
          9198 => x"51",
          9199 => x"3f",
          9200 => x"08",
          9201 => x"52",
          9202 => x"8c",
          9203 => x"8c",
          9204 => x"ba",
          9205 => x"82",
          9206 => x"8c",
          9207 => x"5e",
          9208 => x"08",
          9209 => x"b4",
          9210 => x"2e",
          9211 => x"83",
          9212 => x"7f",
          9213 => x"81",
          9214 => x"38",
          9215 => x"53",
          9216 => x"81",
          9217 => x"d4",
          9218 => x"ba",
          9219 => x"2e",
          9220 => x"56",
          9221 => x"b4",
          9222 => x"56",
          9223 => x"9c",
          9224 => x"33",
          9225 => x"81",
          9226 => x"c9",
          9227 => x"70",
          9228 => x"07",
          9229 => x"80",
          9230 => x"38",
          9231 => x"78",
          9232 => x"89",
          9233 => x"7d",
          9234 => x"3f",
          9235 => x"08",
          9236 => x"8c",
          9237 => x"ff",
          9238 => x"58",
          9239 => x"81",
          9240 => x"58",
          9241 => x"38",
          9242 => x"7f",
          9243 => x"98",
          9244 => x"b4",
          9245 => x"2e",
          9246 => x"1c",
          9247 => x"40",
          9248 => x"38",
          9249 => x"53",
          9250 => x"81",
          9251 => x"d3",
          9252 => x"ba",
          9253 => x"2e",
          9254 => x"57",
          9255 => x"b4",
          9256 => x"58",
          9257 => x"38",
          9258 => x"1f",
          9259 => x"80",
          9260 => x"05",
          9261 => x"15",
          9262 => x"38",
          9263 => x"1f",
          9264 => x"58",
          9265 => x"81",
          9266 => x"77",
          9267 => x"59",
          9268 => x"55",
          9269 => x"9c",
          9270 => x"1f",
          9271 => x"5e",
          9272 => x"1b",
          9273 => x"83",
          9274 => x"56",
          9275 => x"8c",
          9276 => x"0d",
          9277 => x"30",
          9278 => x"72",
          9279 => x"57",
          9280 => x"38",
          9281 => x"52",
          9282 => x"c2",
          9283 => x"8c",
          9284 => x"ba",
          9285 => x"2e",
          9286 => x"fe",
          9287 => x"54",
          9288 => x"53",
          9289 => x"18",
          9290 => x"80",
          9291 => x"8c",
          9292 => x"09",
          9293 => x"bf",
          9294 => x"8c",
          9295 => x"34",
          9296 => x"a8",
          9297 => x"55",
          9298 => x"08",
          9299 => x"82",
          9300 => x"60",
          9301 => x"ac",
          9302 => x"8c",
          9303 => x"9c",
          9304 => x"2b",
          9305 => x"71",
          9306 => x"7d",
          9307 => x"3f",
          9308 => x"08",
          9309 => x"8c",
          9310 => x"38",
          9311 => x"8c",
          9312 => x"8b",
          9313 => x"2a",
          9314 => x"29",
          9315 => x"81",
          9316 => x"57",
          9317 => x"81",
          9318 => x"19",
          9319 => x"76",
          9320 => x"81",
          9321 => x"1d",
          9322 => x"1e",
          9323 => x"56",
          9324 => x"77",
          9325 => x"83",
          9326 => x"7a",
          9327 => x"81",
          9328 => x"38",
          9329 => x"53",
          9330 => x"81",
          9331 => x"d0",
          9332 => x"ba",
          9333 => x"2e",
          9334 => x"57",
          9335 => x"b4",
          9336 => x"58",
          9337 => x"38",
          9338 => x"9c",
          9339 => x"81",
          9340 => x"5c",
          9341 => x"1c",
          9342 => x"8b",
          9343 => x"8c",
          9344 => x"9a",
          9345 => x"9b",
          9346 => x"8d",
          9347 => x"76",
          9348 => x"59",
          9349 => x"ff",
          9350 => x"78",
          9351 => x"22",
          9352 => x"58",
          9353 => x"8c",
          9354 => x"05",
          9355 => x"70",
          9356 => x"34",
          9357 => x"56",
          9358 => x"76",
          9359 => x"ff",
          9360 => x"18",
          9361 => x"27",
          9362 => x"83",
          9363 => x"81",
          9364 => x"10",
          9365 => x"58",
          9366 => x"2e",
          9367 => x"7c",
          9368 => x"0b",
          9369 => x"80",
          9370 => x"e9",
          9371 => x"ba",
          9372 => x"84",
          9373 => x"fc",
          9374 => x"ff",
          9375 => x"fe",
          9376 => x"eb",
          9377 => x"b4",
          9378 => x"b8",
          9379 => x"81",
          9380 => x"59",
          9381 => x"81",
          9382 => x"8c",
          9383 => x"38",
          9384 => x"08",
          9385 => x"b4",
          9386 => x"1d",
          9387 => x"ba",
          9388 => x"41",
          9389 => x"08",
          9390 => x"38",
          9391 => x"42",
          9392 => x"09",
          9393 => x"bc",
          9394 => x"b4",
          9395 => x"1d",
          9396 => x"78",
          9397 => x"33",
          9398 => x"3f",
          9399 => x"a4",
          9400 => x"1f",
          9401 => x"57",
          9402 => x"81",
          9403 => x"81",
          9404 => x"38",
          9405 => x"81",
          9406 => x"76",
          9407 => x"9f",
          9408 => x"39",
          9409 => x"07",
          9410 => x"39",
          9411 => x"1c",
          9412 => x"52",
          9413 => x"51",
          9414 => x"84",
          9415 => x"76",
          9416 => x"06",
          9417 => x"ba",
          9418 => x"1d",
          9419 => x"08",
          9420 => x"31",
          9421 => x"1d",
          9422 => x"38",
          9423 => x"5f",
          9424 => x"aa",
          9425 => x"8c",
          9426 => x"f8",
          9427 => x"1c",
          9428 => x"80",
          9429 => x"38",
          9430 => x"75",
          9431 => x"e8",
          9432 => x"59",
          9433 => x"2e",
          9434 => x"fa",
          9435 => x"54",
          9436 => x"a0",
          9437 => x"53",
          9438 => x"1c",
          9439 => x"ac",
          9440 => x"39",
          9441 => x"18",
          9442 => x"08",
          9443 => x"52",
          9444 => x"51",
          9445 => x"f8",
          9446 => x"3d",
          9447 => x"71",
          9448 => x"5c",
          9449 => x"1e",
          9450 => x"08",
          9451 => x"b5",
          9452 => x"08",
          9453 => x"d9",
          9454 => x"71",
          9455 => x"08",
          9456 => x"58",
          9457 => x"72",
          9458 => x"38",
          9459 => x"14",
          9460 => x"1b",
          9461 => x"7a",
          9462 => x"80",
          9463 => x"70",
          9464 => x"06",
          9465 => x"8f",
          9466 => x"83",
          9467 => x"1a",
          9468 => x"22",
          9469 => x"5b",
          9470 => x"7a",
          9471 => x"25",
          9472 => x"06",
          9473 => x"7c",
          9474 => x"57",
          9475 => x"18",
          9476 => x"89",
          9477 => x"58",
          9478 => x"16",
          9479 => x"18",
          9480 => x"74",
          9481 => x"38",
          9482 => x"81",
          9483 => x"89",
          9484 => x"70",
          9485 => x"25",
          9486 => x"77",
          9487 => x"38",
          9488 => x"8b",
          9489 => x"70",
          9490 => x"34",
          9491 => x"74",
          9492 => x"05",
          9493 => x"18",
          9494 => x"27",
          9495 => x"7c",
          9496 => x"55",
          9497 => x"16",
          9498 => x"33",
          9499 => x"38",
          9500 => x"38",
          9501 => x"1e",
          9502 => x"7c",
          9503 => x"56",
          9504 => x"17",
          9505 => x"08",
          9506 => x"55",
          9507 => x"38",
          9508 => x"34",
          9509 => x"53",
          9510 => x"88",
          9511 => x"1c",
          9512 => x"83",
          9513 => x"12",
          9514 => x"2b",
          9515 => x"07",
          9516 => x"70",
          9517 => x"2b",
          9518 => x"07",
          9519 => x"97",
          9520 => x"17",
          9521 => x"2b",
          9522 => x"5b",
          9523 => x"5b",
          9524 => x"1e",
          9525 => x"33",
          9526 => x"71",
          9527 => x"5d",
          9528 => x"1e",
          9529 => x"0d",
          9530 => x"55",
          9531 => x"77",
          9532 => x"81",
          9533 => x"58",
          9534 => x"b5",
          9535 => x"2b",
          9536 => x"81",
          9537 => x"84",
          9538 => x"83",
          9539 => x"55",
          9540 => x"27",
          9541 => x"76",
          9542 => x"38",
          9543 => x"54",
          9544 => x"74",
          9545 => x"82",
          9546 => x"80",
          9547 => x"08",
          9548 => x"19",
          9549 => x"22",
          9550 => x"79",
          9551 => x"fd",
          9552 => x"30",
          9553 => x"78",
          9554 => x"72",
          9555 => x"58",
          9556 => x"80",
          9557 => x"7a",
          9558 => x"05",
          9559 => x"8c",
          9560 => x"5b",
          9561 => x"73",
          9562 => x"5a",
          9563 => x"80",
          9564 => x"38",
          9565 => x"7e",
          9566 => x"89",
          9567 => x"bf",
          9568 => x"78",
          9569 => x"38",
          9570 => x"8c",
          9571 => x"5b",
          9572 => x"b4",
          9573 => x"2a",
          9574 => x"06",
          9575 => x"2e",
          9576 => x"14",
          9577 => x"ff",
          9578 => x"73",
          9579 => x"05",
          9580 => x"16",
          9581 => x"19",
          9582 => x"33",
          9583 => x"56",
          9584 => x"b7",
          9585 => x"39",
          9586 => x"53",
          9587 => x"7b",
          9588 => x"25",
          9589 => x"06",
          9590 => x"58",
          9591 => x"ef",
          9592 => x"70",
          9593 => x"57",
          9594 => x"70",
          9595 => x"53",
          9596 => x"83",
          9597 => x"74",
          9598 => x"81",
          9599 => x"80",
          9600 => x"38",
          9601 => x"88",
          9602 => x"33",
          9603 => x"3d",
          9604 => x"9f",
          9605 => x"a7",
          9606 => x"8c",
          9607 => x"80",
          9608 => x"70",
          9609 => x"33",
          9610 => x"81",
          9611 => x"7f",
          9612 => x"2e",
          9613 => x"83",
          9614 => x"27",
          9615 => x"10",
          9616 => x"76",
          9617 => x"57",
          9618 => x"ff",
          9619 => x"32",
          9620 => x"73",
          9621 => x"25",
          9622 => x"5b",
          9623 => x"90",
          9624 => x"dc",
          9625 => x"38",
          9626 => x"26",
          9627 => x"e5",
          9628 => x"e5",
          9629 => x"81",
          9630 => x"54",
          9631 => x"2e",
          9632 => x"73",
          9633 => x"38",
          9634 => x"33",
          9635 => x"06",
          9636 => x"73",
          9637 => x"81",
          9638 => x"7a",
          9639 => x"76",
          9640 => x"80",
          9641 => x"10",
          9642 => x"7d",
          9643 => x"62",
          9644 => x"05",
          9645 => x"54",
          9646 => x"2e",
          9647 => x"80",
          9648 => x"73",
          9649 => x"70",
          9650 => x"25",
          9651 => x"55",
          9652 => x"80",
          9653 => x"81",
          9654 => x"54",
          9655 => x"54",
          9656 => x"2e",
          9657 => x"80",
          9658 => x"30",
          9659 => x"77",
          9660 => x"57",
          9661 => x"72",
          9662 => x"73",
          9663 => x"94",
          9664 => x"55",
          9665 => x"fe",
          9666 => x"39",
          9667 => x"73",
          9668 => x"e7",
          9669 => x"8c",
          9670 => x"ff",
          9671 => x"fe",
          9672 => x"54",
          9673 => x"8c",
          9674 => x"0d",
          9675 => x"a8",
          9676 => x"ff",
          9677 => x"7a",
          9678 => x"e3",
          9679 => x"ff",
          9680 => x"1d",
          9681 => x"7b",
          9682 => x"3f",
          9683 => x"08",
          9684 => x"0c",
          9685 => x"04",
          9686 => x"dc",
          9687 => x"70",
          9688 => x"07",
          9689 => x"56",
          9690 => x"a1",
          9691 => x"42",
          9692 => x"33",
          9693 => x"72",
          9694 => x"38",
          9695 => x"32",
          9696 => x"80",
          9697 => x"40",
          9698 => x"e1",
          9699 => x"0c",
          9700 => x"82",
          9701 => x"81",
          9702 => x"38",
          9703 => x"83",
          9704 => x"17",
          9705 => x"2e",
          9706 => x"17",
          9707 => x"05",
          9708 => x"a0",
          9709 => x"70",
          9710 => x"42",
          9711 => x"59",
          9712 => x"84",
          9713 => x"38",
          9714 => x"76",
          9715 => x"59",
          9716 => x"80",
          9717 => x"80",
          9718 => x"38",
          9719 => x"70",
          9720 => x"06",
          9721 => x"55",
          9722 => x"2e",
          9723 => x"73",
          9724 => x"06",
          9725 => x"2e",
          9726 => x"76",
          9727 => x"38",
          9728 => x"05",
          9729 => x"54",
          9730 => x"9d",
          9731 => x"18",
          9732 => x"ff",
          9733 => x"80",
          9734 => x"fe",
          9735 => x"5e",
          9736 => x"2e",
          9737 => x"eb",
          9738 => x"a0",
          9739 => x"a0",
          9740 => x"05",
          9741 => x"13",
          9742 => x"38",
          9743 => x"5e",
          9744 => x"70",
          9745 => x"59",
          9746 => x"74",
          9747 => x"ed",
          9748 => x"2e",
          9749 => x"74",
          9750 => x"30",
          9751 => x"55",
          9752 => x"77",
          9753 => x"38",
          9754 => x"38",
          9755 => x"7b",
          9756 => x"81",
          9757 => x"32",
          9758 => x"72",
          9759 => x"70",
          9760 => x"51",
          9761 => x"80",
          9762 => x"38",
          9763 => x"86",
          9764 => x"77",
          9765 => x"79",
          9766 => x"75",
          9767 => x"38",
          9768 => x"5b",
          9769 => x"2b",
          9770 => x"77",
          9771 => x"5d",
          9772 => x"22",
          9773 => x"56",
          9774 => x"95",
          9775 => x"33",
          9776 => x"e5",
          9777 => x"38",
          9778 => x"82",
          9779 => x"8c",
          9780 => x"8c",
          9781 => x"38",
          9782 => x"55",
          9783 => x"82",
          9784 => x"81",
          9785 => x"56",
          9786 => x"7d",
          9787 => x"7c",
          9788 => x"38",
          9789 => x"5a",
          9790 => x"81",
          9791 => x"80",
          9792 => x"79",
          9793 => x"79",
          9794 => x"7b",
          9795 => x"3f",
          9796 => x"08",
          9797 => x"56",
          9798 => x"8c",
          9799 => x"81",
          9800 => x"ba",
          9801 => x"2e",
          9802 => x"fb",
          9803 => x"85",
          9804 => x"5a",
          9805 => x"84",
          9806 => x"82",
          9807 => x"59",
          9808 => x"38",
          9809 => x"55",
          9810 => x"8c",
          9811 => x"80",
          9812 => x"39",
          9813 => x"11",
          9814 => x"22",
          9815 => x"56",
          9816 => x"f0",
          9817 => x"2e",
          9818 => x"79",
          9819 => x"fd",
          9820 => x"18",
          9821 => x"ae",
          9822 => x"06",
          9823 => x"77",
          9824 => x"ae",
          9825 => x"06",
          9826 => x"76",
          9827 => x"80",
          9828 => x"0b",
          9829 => x"53",
          9830 => x"73",
          9831 => x"a0",
          9832 => x"70",
          9833 => x"34",
          9834 => x"8a",
          9835 => x"38",
          9836 => x"58",
          9837 => x"34",
          9838 => x"bf",
          9839 => x"8c",
          9840 => x"33",
          9841 => x"ba",
          9842 => x"d6",
          9843 => x"2a",
          9844 => x"77",
          9845 => x"86",
          9846 => x"84",
          9847 => x"56",
          9848 => x"2e",
          9849 => x"90",
          9850 => x"ff",
          9851 => x"80",
          9852 => x"80",
          9853 => x"71",
          9854 => x"62",
          9855 => x"54",
          9856 => x"2e",
          9857 => x"74",
          9858 => x"7b",
          9859 => x"56",
          9860 => x"77",
          9861 => x"ae",
          9862 => x"38",
          9863 => x"76",
          9864 => x"fb",
          9865 => x"83",
          9866 => x"56",
          9867 => x"39",
          9868 => x"81",
          9869 => x"8c",
          9870 => x"77",
          9871 => x"81",
          9872 => x"38",
          9873 => x"5a",
          9874 => x"85",
          9875 => x"34",
          9876 => x"09",
          9877 => x"f6",
          9878 => x"ff",
          9879 => x"1d",
          9880 => x"84",
          9881 => x"93",
          9882 => x"74",
          9883 => x"9d",
          9884 => x"75",
          9885 => x"38",
          9886 => x"78",
          9887 => x"f7",
          9888 => x"07",
          9889 => x"57",
          9890 => x"a4",
          9891 => x"07",
          9892 => x"52",
          9893 => x"85",
          9894 => x"ba",
          9895 => x"ff",
          9896 => x"87",
          9897 => x"5a",
          9898 => x"2e",
          9899 => x"80",
          9900 => x"e6",
          9901 => x"56",
          9902 => x"ff",
          9903 => x"38",
          9904 => x"81",
          9905 => x"e5",
          9906 => x"e5",
          9907 => x"81",
          9908 => x"54",
          9909 => x"2e",
          9910 => x"73",
          9911 => x"38",
          9912 => x"33",
          9913 => x"06",
          9914 => x"73",
          9915 => x"81",
          9916 => x"78",
          9917 => x"ff",
          9918 => x"73",
          9919 => x"38",
          9920 => x"70",
          9921 => x"5f",
          9922 => x"15",
          9923 => x"26",
          9924 => x"81",
          9925 => x"ff",
          9926 => x"70",
          9927 => x"06",
          9928 => x"53",
          9929 => x"05",
          9930 => x"34",
          9931 => x"75",
          9932 => x"fc",
          9933 => x"fa",
          9934 => x"e5",
          9935 => x"81",
          9936 => x"53",
          9937 => x"ff",
          9938 => x"df",
          9939 => x"7d",
          9940 => x"5b",
          9941 => x"79",
          9942 => x"5b",
          9943 => x"cd",
          9944 => x"cc",
          9945 => x"98",
          9946 => x"2b",
          9947 => x"88",
          9948 => x"57",
          9949 => x"7b",
          9950 => x"75",
          9951 => x"54",
          9952 => x"81",
          9953 => x"a0",
          9954 => x"74",
          9955 => x"1b",
          9956 => x"39",
          9957 => x"a0",
          9958 => x"5a",
          9959 => x"2e",
          9960 => x"fa",
          9961 => x"a3",
          9962 => x"2a",
          9963 => x"7b",
          9964 => x"85",
          9965 => x"8c",
          9966 => x"0d",
          9967 => x"0d",
          9968 => x"88",
          9969 => x"05",
          9970 => x"5e",
          9971 => x"ff",
          9972 => x"59",
          9973 => x"80",
          9974 => x"38",
          9975 => x"05",
          9976 => x"9f",
          9977 => x"75",
          9978 => x"d0",
          9979 => x"38",
          9980 => x"85",
          9981 => x"d1",
          9982 => x"80",
          9983 => x"b2",
          9984 => x"10",
          9985 => x"05",
          9986 => x"5a",
          9987 => x"80",
          9988 => x"38",
          9989 => x"7f",
          9990 => x"77",
          9991 => x"7b",
          9992 => x"38",
          9993 => x"51",
          9994 => x"3f",
          9995 => x"08",
          9996 => x"70",
          9997 => x"58",
          9998 => x"86",
          9999 => x"77",
         10000 => x"5d",
         10001 => x"1d",
         10002 => x"34",
         10003 => x"17",
         10004 => x"bb",
         10005 => x"ba",
         10006 => x"ff",
         10007 => x"06",
         10008 => x"58",
         10009 => x"38",
         10010 => x"8d",
         10011 => x"2a",
         10012 => x"8a",
         10013 => x"b1",
         10014 => x"7a",
         10015 => x"ff",
         10016 => x"0c",
         10017 => x"55",
         10018 => x"53",
         10019 => x"53",
         10020 => x"52",
         10021 => x"95",
         10022 => x"8c",
         10023 => x"85",
         10024 => x"81",
         10025 => x"18",
         10026 => x"78",
         10027 => x"b7",
         10028 => x"b6",
         10029 => x"88",
         10030 => x"56",
         10031 => x"82",
         10032 => x"85",
         10033 => x"81",
         10034 => x"84",
         10035 => x"33",
         10036 => x"bf",
         10037 => x"75",
         10038 => x"cd",
         10039 => x"75",
         10040 => x"c5",
         10041 => x"17",
         10042 => x"18",
         10043 => x"2b",
         10044 => x"7c",
         10045 => x"09",
         10046 => x"ad",
         10047 => x"17",
         10048 => x"18",
         10049 => x"2b",
         10050 => x"75",
         10051 => x"dc",
         10052 => x"33",
         10053 => x"71",
         10054 => x"88",
         10055 => x"14",
         10056 => x"07",
         10057 => x"33",
         10058 => x"5a",
         10059 => x"5f",
         10060 => x"18",
         10061 => x"17",
         10062 => x"34",
         10063 => x"33",
         10064 => x"81",
         10065 => x"40",
         10066 => x"7c",
         10067 => x"d9",
         10068 => x"ff",
         10069 => x"29",
         10070 => x"33",
         10071 => x"77",
         10072 => x"77",
         10073 => x"2e",
         10074 => x"ff",
         10075 => x"42",
         10076 => x"38",
         10077 => x"33",
         10078 => x"33",
         10079 => x"07",
         10080 => x"88",
         10081 => x"75",
         10082 => x"5a",
         10083 => x"82",
         10084 => x"cc",
         10085 => x"cb",
         10086 => x"88",
         10087 => x"5c",
         10088 => x"80",
         10089 => x"11",
         10090 => x"33",
         10091 => x"71",
         10092 => x"81",
         10093 => x"72",
         10094 => x"75",
         10095 => x"53",
         10096 => x"42",
         10097 => x"c7",
         10098 => x"c6",
         10099 => x"88",
         10100 => x"58",
         10101 => x"80",
         10102 => x"38",
         10103 => x"84",
         10104 => x"79",
         10105 => x"c1",
         10106 => x"74",
         10107 => x"fd",
         10108 => x"84",
         10109 => x"56",
         10110 => x"08",
         10111 => x"a9",
         10112 => x"8c",
         10113 => x"ff",
         10114 => x"83",
         10115 => x"75",
         10116 => x"26",
         10117 => x"5d",
         10118 => x"26",
         10119 => x"81",
         10120 => x"70",
         10121 => x"7b",
         10122 => x"7b",
         10123 => x"1a",
         10124 => x"b0",
         10125 => x"59",
         10126 => x"8a",
         10127 => x"17",
         10128 => x"58",
         10129 => x"80",
         10130 => x"16",
         10131 => x"78",
         10132 => x"82",
         10133 => x"78",
         10134 => x"81",
         10135 => x"06",
         10136 => x"83",
         10137 => x"2a",
         10138 => x"78",
         10139 => x"26",
         10140 => x"0b",
         10141 => x"ff",
         10142 => x"0c",
         10143 => x"84",
         10144 => x"83",
         10145 => x"38",
         10146 => x"84",
         10147 => x"81",
         10148 => x"84",
         10149 => x"7c",
         10150 => x"84",
         10151 => x"8c",
         10152 => x"0b",
         10153 => x"80",
         10154 => x"ba",
         10155 => x"3d",
         10156 => x"0b",
         10157 => x"0c",
         10158 => x"04",
         10159 => x"11",
         10160 => x"06",
         10161 => x"74",
         10162 => x"38",
         10163 => x"81",
         10164 => x"05",
         10165 => x"7a",
         10166 => x"38",
         10167 => x"83",
         10168 => x"40",
         10169 => x"7f",
         10170 => x"70",
         10171 => x"33",
         10172 => x"05",
         10173 => x"9f",
         10174 => x"56",
         10175 => x"89",
         10176 => x"70",
         10177 => x"57",
         10178 => x"17",
         10179 => x"26",
         10180 => x"17",
         10181 => x"06",
         10182 => x"30",
         10183 => x"59",
         10184 => x"2e",
         10185 => x"85",
         10186 => x"be",
         10187 => x"32",
         10188 => x"72",
         10189 => x"7a",
         10190 => x"55",
         10191 => x"87",
         10192 => x"1c",
         10193 => x"5c",
         10194 => x"ff",
         10195 => x"56",
         10196 => x"78",
         10197 => x"cf",
         10198 => x"2a",
         10199 => x"8a",
         10200 => x"c5",
         10201 => x"fe",
         10202 => x"78",
         10203 => x"75",
         10204 => x"09",
         10205 => x"38",
         10206 => x"81",
         10207 => x"30",
         10208 => x"7b",
         10209 => x"5c",
         10210 => x"38",
         10211 => x"2e",
         10212 => x"93",
         10213 => x"5a",
         10214 => x"fa",
         10215 => x"59",
         10216 => x"2e",
         10217 => x"81",
         10218 => x"80",
         10219 => x"90",
         10220 => x"2b",
         10221 => x"19",
         10222 => x"07",
         10223 => x"fe",
         10224 => x"07",
         10225 => x"40",
         10226 => x"7a",
         10227 => x"5c",
         10228 => x"90",
         10229 => x"78",
         10230 => x"be",
         10231 => x"81",
         10232 => x"30",
         10233 => x"72",
         10234 => x"3d",
         10235 => x"05",
         10236 => x"b6",
         10237 => x"52",
         10238 => x"78",
         10239 => x"56",
         10240 => x"80",
         10241 => x"0b",
         10242 => x"ff",
         10243 => x"0c",
         10244 => x"56",
         10245 => x"a5",
         10246 => x"7a",
         10247 => x"52",
         10248 => x"51",
         10249 => x"3f",
         10250 => x"08",
         10251 => x"38",
         10252 => x"56",
         10253 => x"0c",
         10254 => x"bf",
         10255 => x"33",
         10256 => x"88",
         10257 => x"5e",
         10258 => x"82",
         10259 => x"09",
         10260 => x"38",
         10261 => x"18",
         10262 => x"75",
         10263 => x"82",
         10264 => x"81",
         10265 => x"30",
         10266 => x"7a",
         10267 => x"42",
         10268 => x"75",
         10269 => x"b6",
         10270 => x"77",
         10271 => x"56",
         10272 => x"ba",
         10273 => x"5d",
         10274 => x"2e",
         10275 => x"83",
         10276 => x"81",
         10277 => x"bd",
         10278 => x"2e",
         10279 => x"81",
         10280 => x"5a",
         10281 => x"27",
         10282 => x"f8",
         10283 => x"0b",
         10284 => x"83",
         10285 => x"5d",
         10286 => x"81",
         10287 => x"7e",
         10288 => x"40",
         10289 => x"31",
         10290 => x"52",
         10291 => x"80",
         10292 => x"38",
         10293 => x"e1",
         10294 => x"81",
         10295 => x"e5",
         10296 => x"58",
         10297 => x"05",
         10298 => x"70",
         10299 => x"33",
         10300 => x"ff",
         10301 => x"42",
         10302 => x"2e",
         10303 => x"75",
         10304 => x"38",
         10305 => x"f3",
         10306 => x"7c",
         10307 => x"77",
         10308 => x"0c",
         10309 => x"04",
         10310 => x"80",
         10311 => x"38",
         10312 => x"8a",
         10313 => x"c0",
         10314 => x"ff",
         10315 => x"0b",
         10316 => x"0c",
         10317 => x"04",
         10318 => x"ee",
         10319 => x"bc",
         10320 => x"78",
         10321 => x"5a",
         10322 => x"81",
         10323 => x"71",
         10324 => x"1b",
         10325 => x"5f",
         10326 => x"83",
         10327 => x"80",
         10328 => x"85",
         10329 => x"18",
         10330 => x"5c",
         10331 => x"70",
         10332 => x"33",
         10333 => x"05",
         10334 => x"71",
         10335 => x"5b",
         10336 => x"77",
         10337 => x"91",
         10338 => x"2e",
         10339 => x"3d",
         10340 => x"83",
         10341 => x"39",
         10342 => x"c6",
         10343 => x"17",
         10344 => x"18",
         10345 => x"2b",
         10346 => x"75",
         10347 => x"81",
         10348 => x"38",
         10349 => x"80",
         10350 => x"08",
         10351 => x"38",
         10352 => x"5b",
         10353 => x"09",
         10354 => x"9b",
         10355 => x"77",
         10356 => x"52",
         10357 => x"51",
         10358 => x"3f",
         10359 => x"08",
         10360 => x"38",
         10361 => x"5a",
         10362 => x"0c",
         10363 => x"38",
         10364 => x"34",
         10365 => x"33",
         10366 => x"33",
         10367 => x"07",
         10368 => x"82",
         10369 => x"09",
         10370 => x"fc",
         10371 => x"83",
         10372 => x"12",
         10373 => x"2b",
         10374 => x"07",
         10375 => x"70",
         10376 => x"2b",
         10377 => x"07",
         10378 => x"45",
         10379 => x"77",
         10380 => x"a4",
         10381 => x"81",
         10382 => x"38",
         10383 => x"83",
         10384 => x"12",
         10385 => x"2b",
         10386 => x"07",
         10387 => x"70",
         10388 => x"2b",
         10389 => x"07",
         10390 => x"5b",
         10391 => x"60",
         10392 => x"e4",
         10393 => x"81",
         10394 => x"38",
         10395 => x"83",
         10396 => x"12",
         10397 => x"2b",
         10398 => x"07",
         10399 => x"70",
         10400 => x"2b",
         10401 => x"07",
         10402 => x"5d",
         10403 => x"83",
         10404 => x"12",
         10405 => x"2b",
         10406 => x"07",
         10407 => x"70",
         10408 => x"2b",
         10409 => x"07",
         10410 => x"0c",
         10411 => x"46",
         10412 => x"45",
         10413 => x"7c",
         10414 => x"d1",
         10415 => x"05",
         10416 => x"d1",
         10417 => x"86",
         10418 => x"d1",
         10419 => x"18",
         10420 => x"98",
         10421 => x"cf",
         10422 => x"24",
         10423 => x"7b",
         10424 => x"56",
         10425 => x"75",
         10426 => x"08",
         10427 => x"70",
         10428 => x"33",
         10429 => x"af",
         10430 => x"ba",
         10431 => x"2e",
         10432 => x"81",
         10433 => x"ba",
         10434 => x"18",
         10435 => x"08",
         10436 => x"31",
         10437 => x"18",
         10438 => x"38",
         10439 => x"41",
         10440 => x"81",
         10441 => x"ba",
         10442 => x"fd",
         10443 => x"56",
         10444 => x"f3",
         10445 => x"0b",
         10446 => x"83",
         10447 => x"5a",
         10448 => x"39",
         10449 => x"33",
         10450 => x"33",
         10451 => x"07",
         10452 => x"58",
         10453 => x"38",
         10454 => x"42",
         10455 => x"38",
         10456 => x"83",
         10457 => x"12",
         10458 => x"2b",
         10459 => x"07",
         10460 => x"70",
         10461 => x"2b",
         10462 => x"07",
         10463 => x"5a",
         10464 => x"5a",
         10465 => x"59",
         10466 => x"39",
         10467 => x"80",
         10468 => x"38",
         10469 => x"e3",
         10470 => x"2e",
         10471 => x"93",
         10472 => x"5a",
         10473 => x"f2",
         10474 => x"79",
         10475 => x"fc",
         10476 => x"54",
         10477 => x"a0",
         10478 => x"53",
         10479 => x"17",
         10480 => x"ad",
         10481 => x"85",
         10482 => x"0d",
         10483 => x"05",
         10484 => x"43",
         10485 => x"57",
         10486 => x"5a",
         10487 => x"2e",
         10488 => x"78",
         10489 => x"5a",
         10490 => x"26",
         10491 => x"ba",
         10492 => x"38",
         10493 => x"74",
         10494 => x"d9",
         10495 => x"e8",
         10496 => x"74",
         10497 => x"38",
         10498 => x"84",
         10499 => x"70",
         10500 => x"73",
         10501 => x"38",
         10502 => x"62",
         10503 => x"2e",
         10504 => x"74",
         10505 => x"73",
         10506 => x"54",
         10507 => x"92",
         10508 => x"93",
         10509 => x"84",
         10510 => x"81",
         10511 => x"8c",
         10512 => x"84",
         10513 => x"92",
         10514 => x"8b",
         10515 => x"8c",
         10516 => x"0d",
         10517 => x"d0",
         10518 => x"ff",
         10519 => x"57",
         10520 => x"91",
         10521 => x"77",
         10522 => x"d0",
         10523 => x"77",
         10524 => x"f7",
         10525 => x"08",
         10526 => x"5e",
         10527 => x"08",
         10528 => x"79",
         10529 => x"5b",
         10530 => x"81",
         10531 => x"ff",
         10532 => x"57",
         10533 => x"26",
         10534 => x"15",
         10535 => x"06",
         10536 => x"9f",
         10537 => x"99",
         10538 => x"e0",
         10539 => x"ff",
         10540 => x"74",
         10541 => x"2a",
         10542 => x"76",
         10543 => x"06",
         10544 => x"ff",
         10545 => x"79",
         10546 => x"70",
         10547 => x"2a",
         10548 => x"57",
         10549 => x"2e",
         10550 => x"1b",
         10551 => x"5b",
         10552 => x"ff",
         10553 => x"54",
         10554 => x"7a",
         10555 => x"38",
         10556 => x"0c",
         10557 => x"39",
         10558 => x"6c",
         10559 => x"80",
         10560 => x"56",
         10561 => x"78",
         10562 => x"38",
         10563 => x"70",
         10564 => x"cc",
         10565 => x"3d",
         10566 => x"58",
         10567 => x"84",
         10568 => x"57",
         10569 => x"08",
         10570 => x"38",
         10571 => x"76",
         10572 => x"ba",
         10573 => x"3d",
         10574 => x"40",
         10575 => x"3d",
         10576 => x"e1",
         10577 => x"ba",
         10578 => x"84",
         10579 => x"80",
         10580 => x"38",
         10581 => x"5d",
         10582 => x"81",
         10583 => x"80",
         10584 => x"38",
         10585 => x"83",
         10586 => x"88",
         10587 => x"ff",
         10588 => x"83",
         10589 => x"5b",
         10590 => x"81",
         10591 => x"9b",
         10592 => x"12",
         10593 => x"2b",
         10594 => x"33",
         10595 => x"5e",
         10596 => x"2e",
         10597 => x"80",
         10598 => x"34",
         10599 => x"17",
         10600 => x"90",
         10601 => x"cc",
         10602 => x"34",
         10603 => x"0b",
         10604 => x"7e",
         10605 => x"80",
         10606 => x"34",
         10607 => x"17",
         10608 => x"5d",
         10609 => x"84",
         10610 => x"5b",
         10611 => x"1c",
         10612 => x"9d",
         10613 => x"0b",
         10614 => x"80",
         10615 => x"34",
         10616 => x"0b",
         10617 => x"7b",
         10618 => x"e2",
         10619 => x"11",
         10620 => x"08",
         10621 => x"57",
         10622 => x"89",
         10623 => x"08",
         10624 => x"8a",
         10625 => x"80",
         10626 => x"a3",
         10627 => x"e7",
         10628 => x"98",
         10629 => x"7b",
         10630 => x"b8",
         10631 => x"9c",
         10632 => x"7c",
         10633 => x"76",
         10634 => x"02",
         10635 => x"33",
         10636 => x"81",
         10637 => x"7b",
         10638 => x"77",
         10639 => x"06",
         10640 => x"2e",
         10641 => x"81",
         10642 => x"81",
         10643 => x"83",
         10644 => x"56",
         10645 => x"86",
         10646 => x"c0",
         10647 => x"b4",
         10648 => x"1b",
         10649 => x"1b",
         10650 => x"11",
         10651 => x"33",
         10652 => x"07",
         10653 => x"5e",
         10654 => x"7b",
         10655 => x"f1",
         10656 => x"1a",
         10657 => x"83",
         10658 => x"12",
         10659 => x"2b",
         10660 => x"07",
         10661 => x"70",
         10662 => x"2b",
         10663 => x"07",
         10664 => x"05",
         10665 => x"0c",
         10666 => x"59",
         10667 => x"86",
         10668 => x"1a",
         10669 => x"1a",
         10670 => x"91",
         10671 => x"0b",
         10672 => x"77",
         10673 => x"06",
         10674 => x"2e",
         10675 => x"75",
         10676 => x"f1",
         10677 => x"1a",
         10678 => x"22",
         10679 => x"7c",
         10680 => x"76",
         10681 => x"07",
         10682 => x"5b",
         10683 => x"84",
         10684 => x"70",
         10685 => x"5b",
         10686 => x"84",
         10687 => x"52",
         10688 => x"ac",
         10689 => x"ba",
         10690 => x"84",
         10691 => x"81",
         10692 => x"82",
         10693 => x"8c",
         10694 => x"80",
         10695 => x"7a",
         10696 => x"39",
         10697 => x"05",
         10698 => x"5e",
         10699 => x"77",
         10700 => x"06",
         10701 => x"2e",
         10702 => x"88",
         10703 => x"0c",
         10704 => x"87",
         10705 => x"0c",
         10706 => x"84",
         10707 => x"0c",
         10708 => x"79",
         10709 => x"3f",
         10710 => x"08",
         10711 => x"59",
         10712 => x"c8",
         10713 => x"39",
         10714 => x"31",
         10715 => x"f3",
         10716 => x"33",
         10717 => x"71",
         10718 => x"90",
         10719 => x"07",
         10720 => x"fd",
         10721 => x"55",
         10722 => x"81",
         10723 => x"52",
         10724 => x"ab",
         10725 => x"ba",
         10726 => x"84",
         10727 => x"80",
         10728 => x"38",
         10729 => x"08",
         10730 => x"d9",
         10731 => x"8c",
         10732 => x"83",
         10733 => x"53",
         10734 => x"51",
         10735 => x"3f",
         10736 => x"08",
         10737 => x"9c",
         10738 => x"11",
         10739 => x"58",
         10740 => x"75",
         10741 => x"38",
         10742 => x"18",
         10743 => x"33",
         10744 => x"74",
         10745 => x"7c",
         10746 => x"26",
         10747 => x"80",
         10748 => x"0b",
         10749 => x"80",
         10750 => x"34",
         10751 => x"95",
         10752 => x"17",
         10753 => x"2b",
         10754 => x"07",
         10755 => x"56",
         10756 => x"8e",
         10757 => x"0b",
         10758 => x"a1",
         10759 => x"34",
         10760 => x"91",
         10761 => x"56",
         10762 => x"17",
         10763 => x"57",
         10764 => x"9a",
         10765 => x"0b",
         10766 => x"7d",
         10767 => x"83",
         10768 => x"06",
         10769 => x"ff",
         10770 => x"7f",
         10771 => x"59",
         10772 => x"16",
         10773 => x"ae",
         10774 => x"33",
         10775 => x"2e",
         10776 => x"b5",
         10777 => x"7d",
         10778 => x"52",
         10779 => x"51",
         10780 => x"3f",
         10781 => x"08",
         10782 => x"38",
         10783 => x"5b",
         10784 => x"0c",
         10785 => x"ff",
         10786 => x"0c",
         10787 => x"2e",
         10788 => x"80",
         10789 => x"97",
         10790 => x"b4",
         10791 => x"b8",
         10792 => x"81",
         10793 => x"5a",
         10794 => x"3f",
         10795 => x"08",
         10796 => x"81",
         10797 => x"38",
         10798 => x"08",
         10799 => x"b4",
         10800 => x"17",
         10801 => x"ba",
         10802 => x"55",
         10803 => x"08",
         10804 => x"38",
         10805 => x"55",
         10806 => x"09",
         10807 => x"85",
         10808 => x"b4",
         10809 => x"17",
         10810 => x"79",
         10811 => x"33",
         10812 => x"b8",
         10813 => x"fe",
         10814 => x"94",
         10815 => x"56",
         10816 => x"77",
         10817 => x"76",
         10818 => x"75",
         10819 => x"5a",
         10820 => x"f8",
         10821 => x"fe",
         10822 => x"08",
         10823 => x"59",
         10824 => x"27",
         10825 => x"8a",
         10826 => x"71",
         10827 => x"08",
         10828 => x"74",
         10829 => x"cd",
         10830 => x"2a",
         10831 => x"0c",
         10832 => x"ed",
         10833 => x"1a",
         10834 => x"f7",
         10835 => x"57",
         10836 => x"f7",
         10837 => x"ba",
         10838 => x"80",
         10839 => x"cf",
         10840 => x"57",
         10841 => x"39",
         10842 => x"62",
         10843 => x"40",
         10844 => x"80",
         10845 => x"57",
         10846 => x"9f",
         10847 => x"56",
         10848 => x"97",
         10849 => x"55",
         10850 => x"8f",
         10851 => x"22",
         10852 => x"59",
         10853 => x"2e",
         10854 => x"80",
         10855 => x"76",
         10856 => x"8c",
         10857 => x"33",
         10858 => x"84",
         10859 => x"33",
         10860 => x"87",
         10861 => x"2e",
         10862 => x"94",
         10863 => x"1b",
         10864 => x"56",
         10865 => x"26",
         10866 => x"7b",
         10867 => x"d5",
         10868 => x"75",
         10869 => x"5b",
         10870 => x"38",
         10871 => x"ff",
         10872 => x"2a",
         10873 => x"9b",
         10874 => x"d3",
         10875 => x"08",
         10876 => x"27",
         10877 => x"74",
         10878 => x"f0",
         10879 => x"1b",
         10880 => x"98",
         10881 => x"05",
         10882 => x"fe",
         10883 => x"76",
         10884 => x"e7",
         10885 => x"22",
         10886 => x"b0",
         10887 => x"56",
         10888 => x"2e",
         10889 => x"7a",
         10890 => x"2a",
         10891 => x"80",
         10892 => x"38",
         10893 => x"75",
         10894 => x"38",
         10895 => x"58",
         10896 => x"53",
         10897 => x"19",
         10898 => x"9f",
         10899 => x"ba",
         10900 => x"98",
         10901 => x"11",
         10902 => x"75",
         10903 => x"38",
         10904 => x"77",
         10905 => x"78",
         10906 => x"84",
         10907 => x"29",
         10908 => x"58",
         10909 => x"70",
         10910 => x"33",
         10911 => x"05",
         10912 => x"15",
         10913 => x"38",
         10914 => x"58",
         10915 => x"7e",
         10916 => x"0c",
         10917 => x"1c",
         10918 => x"59",
         10919 => x"5e",
         10920 => x"af",
         10921 => x"75",
         10922 => x"0c",
         10923 => x"04",
         10924 => x"8c",
         10925 => x"0d",
         10926 => x"fe",
         10927 => x"1a",
         10928 => x"83",
         10929 => x"80",
         10930 => x"5b",
         10931 => x"83",
         10932 => x"76",
         10933 => x"08",
         10934 => x"38",
         10935 => x"1a",
         10936 => x"41",
         10937 => x"2e",
         10938 => x"80",
         10939 => x"54",
         10940 => x"19",
         10941 => x"33",
         10942 => x"b1",
         10943 => x"8c",
         10944 => x"85",
         10945 => x"81",
         10946 => x"1a",
         10947 => x"dc",
         10948 => x"1b",
         10949 => x"06",
         10950 => x"5a",
         10951 => x"56",
         10952 => x"2e",
         10953 => x"74",
         10954 => x"56",
         10955 => x"81",
         10956 => x"ff",
         10957 => x"80",
         10958 => x"38",
         10959 => x"05",
         10960 => x"70",
         10961 => x"34",
         10962 => x"75",
         10963 => x"bc",
         10964 => x"b4",
         10965 => x"b8",
         10966 => x"81",
         10967 => x"40",
         10968 => x"3f",
         10969 => x"ba",
         10970 => x"2e",
         10971 => x"ff",
         10972 => x"ba",
         10973 => x"1a",
         10974 => x"08",
         10975 => x"31",
         10976 => x"08",
         10977 => x"a0",
         10978 => x"fe",
         10979 => x"19",
         10980 => x"82",
         10981 => x"06",
         10982 => x"81",
         10983 => x"08",
         10984 => x"05",
         10985 => x"81",
         10986 => x"ff",
         10987 => x"7e",
         10988 => x"39",
         10989 => x"0c",
         10990 => x"56",
         10991 => x"98",
         10992 => x"79",
         10993 => x"98",
         10994 => x"8c",
         10995 => x"a1",
         10996 => x"33",
         10997 => x"83",
         10998 => x"8c",
         10999 => x"55",
         11000 => x"38",
         11001 => x"56",
         11002 => x"39",
         11003 => x"1b",
         11004 => x"84",
         11005 => x"92",
         11006 => x"82",
         11007 => x"34",
         11008 => x"ba",
         11009 => x"3d",
         11010 => x"3d",
         11011 => x"67",
         11012 => x"5c",
         11013 => x"0c",
         11014 => x"80",
         11015 => x"79",
         11016 => x"80",
         11017 => x"75",
         11018 => x"80",
         11019 => x"86",
         11020 => x"1b",
         11021 => x"78",
         11022 => x"fd",
         11023 => x"74",
         11024 => x"76",
         11025 => x"91",
         11026 => x"74",
         11027 => x"90",
         11028 => x"81",
         11029 => x"58",
         11030 => x"76",
         11031 => x"a1",
         11032 => x"08",
         11033 => x"57",
         11034 => x"84",
         11035 => x"5b",
         11036 => x"82",
         11037 => x"83",
         11038 => x"7e",
         11039 => x"60",
         11040 => x"ff",
         11041 => x"2a",
         11042 => x"78",
         11043 => x"84",
         11044 => x"1a",
         11045 => x"80",
         11046 => x"38",
         11047 => x"86",
         11048 => x"ff",
         11049 => x"38",
         11050 => x"0c",
         11051 => x"85",
         11052 => x"1b",
         11053 => x"b4",
         11054 => x"1b",
         11055 => x"d3",
         11056 => x"08",
         11057 => x"17",
         11058 => x"58",
         11059 => x"27",
         11060 => x"8a",
         11061 => x"79",
         11062 => x"08",
         11063 => x"74",
         11064 => x"de",
         11065 => x"7b",
         11066 => x"5c",
         11067 => x"83",
         11068 => x"19",
         11069 => x"27",
         11070 => x"79",
         11071 => x"54",
         11072 => x"52",
         11073 => x"51",
         11074 => x"3f",
         11075 => x"08",
         11076 => x"60",
         11077 => x"7d",
         11078 => x"74",
         11079 => x"38",
         11080 => x"b8",
         11081 => x"29",
         11082 => x"56",
         11083 => x"05",
         11084 => x"70",
         11085 => x"34",
         11086 => x"75",
         11087 => x"59",
         11088 => x"34",
         11089 => x"59",
         11090 => x"7e",
         11091 => x"0c",
         11092 => x"1c",
         11093 => x"71",
         11094 => x"8c",
         11095 => x"5a",
         11096 => x"75",
         11097 => x"38",
         11098 => x"8c",
         11099 => x"fe",
         11100 => x"1a",
         11101 => x"80",
         11102 => x"7a",
         11103 => x"80",
         11104 => x"ba",
         11105 => x"3d",
         11106 => x"84",
         11107 => x"92",
         11108 => x"83",
         11109 => x"74",
         11110 => x"60",
         11111 => x"39",
         11112 => x"08",
         11113 => x"83",
         11114 => x"80",
         11115 => x"5c",
         11116 => x"83",
         11117 => x"77",
         11118 => x"08",
         11119 => x"38",
         11120 => x"17",
         11121 => x"41",
         11122 => x"2e",
         11123 => x"80",
         11124 => x"54",
         11125 => x"16",
         11126 => x"33",
         11127 => x"cd",
         11128 => x"8c",
         11129 => x"85",
         11130 => x"81",
         11131 => x"17",
         11132 => x"bf",
         11133 => x"1b",
         11134 => x"06",
         11135 => x"b8",
         11136 => x"56",
         11137 => x"2e",
         11138 => x"70",
         11139 => x"33",
         11140 => x"05",
         11141 => x"16",
         11142 => x"38",
         11143 => x"0b",
         11144 => x"fe",
         11145 => x"54",
         11146 => x"53",
         11147 => x"53",
         11148 => x"52",
         11149 => x"f4",
         11150 => x"84",
         11151 => x"7f",
         11152 => x"06",
         11153 => x"84",
         11154 => x"83",
         11155 => x"16",
         11156 => x"08",
         11157 => x"8c",
         11158 => x"74",
         11159 => x"27",
         11160 => x"82",
         11161 => x"74",
         11162 => x"81",
         11163 => x"38",
         11164 => x"16",
         11165 => x"08",
         11166 => x"52",
         11167 => x"51",
         11168 => x"3f",
         11169 => x"ca",
         11170 => x"08",
         11171 => x"08",
         11172 => x"38",
         11173 => x"40",
         11174 => x"38",
         11175 => x"12",
         11176 => x"08",
         11177 => x"7c",
         11178 => x"58",
         11179 => x"98",
         11180 => x"79",
         11181 => x"e7",
         11182 => x"8c",
         11183 => x"ba",
         11184 => x"d8",
         11185 => x"33",
         11186 => x"39",
         11187 => x"51",
         11188 => x"3f",
         11189 => x"08",
         11190 => x"8c",
         11191 => x"38",
         11192 => x"54",
         11193 => x"53",
         11194 => x"53",
         11195 => x"52",
         11196 => x"b8",
         11197 => x"8c",
         11198 => x"38",
         11199 => x"08",
         11200 => x"b4",
         11201 => x"17",
         11202 => x"77",
         11203 => x"27",
         11204 => x"82",
         11205 => x"7b",
         11206 => x"81",
         11207 => x"38",
         11208 => x"16",
         11209 => x"08",
         11210 => x"52",
         11211 => x"51",
         11212 => x"3f",
         11213 => x"89",
         11214 => x"33",
         11215 => x"9b",
         11216 => x"8c",
         11217 => x"55",
         11218 => x"38",
         11219 => x"56",
         11220 => x"39",
         11221 => x"16",
         11222 => x"16",
         11223 => x"17",
         11224 => x"ff",
         11225 => x"84",
         11226 => x"80",
         11227 => x"ba",
         11228 => x"17",
         11229 => x"08",
         11230 => x"31",
         11231 => x"17",
         11232 => x"98",
         11233 => x"33",
         11234 => x"2e",
         11235 => x"fe",
         11236 => x"54",
         11237 => x"a0",
         11238 => x"53",
         11239 => x"16",
         11240 => x"96",
         11241 => x"7c",
         11242 => x"94",
         11243 => x"56",
         11244 => x"81",
         11245 => x"34",
         11246 => x"ba",
         11247 => x"3d",
         11248 => x"0b",
         11249 => x"82",
         11250 => x"8c",
         11251 => x"0d",
         11252 => x"0d",
         11253 => x"5a",
         11254 => x"9f",
         11255 => x"56",
         11256 => x"97",
         11257 => x"55",
         11258 => x"8f",
         11259 => x"22",
         11260 => x"58",
         11261 => x"2e",
         11262 => x"80",
         11263 => x"79",
         11264 => x"d8",
         11265 => x"33",
         11266 => x"81",
         11267 => x"7a",
         11268 => x"c8",
         11269 => x"19",
         11270 => x"b4",
         11271 => x"2e",
         11272 => x"17",
         11273 => x"81",
         11274 => x"54",
         11275 => x"17",
         11276 => x"33",
         11277 => x"f5",
         11278 => x"8c",
         11279 => x"85",
         11280 => x"81",
         11281 => x"18",
         11282 => x"90",
         11283 => x"08",
         11284 => x"a0",
         11285 => x"78",
         11286 => x"77",
         11287 => x"08",
         11288 => x"ff",
         11289 => x"56",
         11290 => x"34",
         11291 => x"5a",
         11292 => x"34",
         11293 => x"33",
         11294 => x"56",
         11295 => x"2e",
         11296 => x"8c",
         11297 => x"74",
         11298 => x"88",
         11299 => x"9d",
         11300 => x"90",
         11301 => x"9e",
         11302 => x"98",
         11303 => x"9f",
         11304 => x"7a",
         11305 => x"97",
         11306 => x"0b",
         11307 => x"80",
         11308 => x"18",
         11309 => x"92",
         11310 => x"0b",
         11311 => x"7b",
         11312 => x"83",
         11313 => x"51",
         11314 => x"3f",
         11315 => x"08",
         11316 => x"81",
         11317 => x"56",
         11318 => x"34",
         11319 => x"8c",
         11320 => x"0d",
         11321 => x"b4",
         11322 => x"b8",
         11323 => x"81",
         11324 => x"5b",
         11325 => x"3f",
         11326 => x"ba",
         11327 => x"c9",
         11328 => x"8c",
         11329 => x"34",
         11330 => x"a8",
         11331 => x"84",
         11332 => x"57",
         11333 => x"18",
         11334 => x"8e",
         11335 => x"33",
         11336 => x"2e",
         11337 => x"fe",
         11338 => x"54",
         11339 => x"a0",
         11340 => x"53",
         11341 => x"17",
         11342 => x"92",
         11343 => x"56",
         11344 => x"78",
         11345 => x"74",
         11346 => x"74",
         11347 => x"75",
         11348 => x"8c",
         11349 => x"74",
         11350 => x"88",
         11351 => x"9d",
         11352 => x"90",
         11353 => x"9e",
         11354 => x"98",
         11355 => x"9f",
         11356 => x"7a",
         11357 => x"97",
         11358 => x"0b",
         11359 => x"80",
         11360 => x"18",
         11361 => x"92",
         11362 => x"0b",
         11363 => x"7b",
         11364 => x"83",
         11365 => x"51",
         11366 => x"3f",
         11367 => x"08",
         11368 => x"81",
         11369 => x"56",
         11370 => x"34",
         11371 => x"81",
         11372 => x"ff",
         11373 => x"84",
         11374 => x"81",
         11375 => x"fc",
         11376 => x"78",
         11377 => x"fc",
         11378 => x"3d",
         11379 => x"52",
         11380 => x"3f",
         11381 => x"08",
         11382 => x"8c",
         11383 => x"89",
         11384 => x"2e",
         11385 => x"08",
         11386 => x"2e",
         11387 => x"33",
         11388 => x"2e",
         11389 => x"13",
         11390 => x"22",
         11391 => x"77",
         11392 => x"80",
         11393 => x"75",
         11394 => x"38",
         11395 => x"73",
         11396 => x"0c",
         11397 => x"04",
         11398 => x"51",
         11399 => x"3f",
         11400 => x"08",
         11401 => x"72",
         11402 => x"75",
         11403 => x"d5",
         11404 => x"0d",
         11405 => x"5b",
         11406 => x"80",
         11407 => x"75",
         11408 => x"57",
         11409 => x"26",
         11410 => x"ba",
         11411 => x"70",
         11412 => x"ba",
         11413 => x"84",
         11414 => x"51",
         11415 => x"90",
         11416 => x"d1",
         11417 => x"0b",
         11418 => x"0c",
         11419 => x"04",
         11420 => x"ba",
         11421 => x"3d",
         11422 => x"33",
         11423 => x"81",
         11424 => x"53",
         11425 => x"26",
         11426 => x"19",
         11427 => x"06",
         11428 => x"54",
         11429 => x"80",
         11430 => x"0b",
         11431 => x"5b",
         11432 => x"79",
         11433 => x"70",
         11434 => x"33",
         11435 => x"05",
         11436 => x"9f",
         11437 => x"52",
         11438 => x"89",
         11439 => x"70",
         11440 => x"53",
         11441 => x"13",
         11442 => x"26",
         11443 => x"13",
         11444 => x"06",
         11445 => x"30",
         11446 => x"55",
         11447 => x"2e",
         11448 => x"85",
         11449 => x"be",
         11450 => x"32",
         11451 => x"72",
         11452 => x"76",
         11453 => x"52",
         11454 => x"92",
         11455 => x"84",
         11456 => x"83",
         11457 => x"99",
         11458 => x"fe",
         11459 => x"83",
         11460 => x"77",
         11461 => x"fe",
         11462 => x"3d",
         11463 => x"98",
         11464 => x"52",
         11465 => x"d1",
         11466 => x"ba",
         11467 => x"84",
         11468 => x"80",
         11469 => x"74",
         11470 => x"0c",
         11471 => x"04",
         11472 => x"52",
         11473 => x"05",
         11474 => x"3f",
         11475 => x"08",
         11476 => x"8c",
         11477 => x"38",
         11478 => x"05",
         11479 => x"2b",
         11480 => x"77",
         11481 => x"38",
         11482 => x"33",
         11483 => x"81",
         11484 => x"75",
         11485 => x"38",
         11486 => x"11",
         11487 => x"33",
         11488 => x"07",
         11489 => x"5a",
         11490 => x"79",
         11491 => x"38",
         11492 => x"0c",
         11493 => x"8c",
         11494 => x"0d",
         11495 => x"8c",
         11496 => x"09",
         11497 => x"8f",
         11498 => x"84",
         11499 => x"98",
         11500 => x"95",
         11501 => x"17",
         11502 => x"2b",
         11503 => x"07",
         11504 => x"1b",
         11505 => x"cc",
         11506 => x"98",
         11507 => x"74",
         11508 => x"0c",
         11509 => x"04",
         11510 => x"0d",
         11511 => x"08",
         11512 => x"08",
         11513 => x"7c",
         11514 => x"80",
         11515 => x"b4",
         11516 => x"e5",
         11517 => x"c5",
         11518 => x"8c",
         11519 => x"ba",
         11520 => x"c8",
         11521 => x"d9",
         11522 => x"61",
         11523 => x"80",
         11524 => x"58",
         11525 => x"08",
         11526 => x"80",
         11527 => x"38",
         11528 => x"98",
         11529 => x"a0",
         11530 => x"ff",
         11531 => x"84",
         11532 => x"59",
         11533 => x"08",
         11534 => x"60",
         11535 => x"08",
         11536 => x"16",
         11537 => x"b1",
         11538 => x"8c",
         11539 => x"33",
         11540 => x"83",
         11541 => x"54",
         11542 => x"16",
         11543 => x"33",
         11544 => x"c9",
         11545 => x"8c",
         11546 => x"85",
         11547 => x"81",
         11548 => x"17",
         11549 => x"d4",
         11550 => x"3d",
         11551 => x"33",
         11552 => x"71",
         11553 => x"63",
         11554 => x"40",
         11555 => x"78",
         11556 => x"da",
         11557 => x"db",
         11558 => x"52",
         11559 => x"a3",
         11560 => x"ba",
         11561 => x"84",
         11562 => x"82",
         11563 => x"52",
         11564 => x"a8",
         11565 => x"ba",
         11566 => x"84",
         11567 => x"bb",
         11568 => x"3d",
         11569 => x"33",
         11570 => x"71",
         11571 => x"63",
         11572 => x"58",
         11573 => x"7d",
         11574 => x"fd",
         11575 => x"2e",
         11576 => x"ba",
         11577 => x"7a",
         11578 => x"e2",
         11579 => x"8c",
         11580 => x"ba",
         11581 => x"2e",
         11582 => x"78",
         11583 => x"d8",
         11584 => x"c8",
         11585 => x"3d",
         11586 => x"52",
         11587 => x"bd",
         11588 => x"7f",
         11589 => x"5b",
         11590 => x"2e",
         11591 => x"1f",
         11592 => x"81",
         11593 => x"5f",
         11594 => x"f5",
         11595 => x"56",
         11596 => x"81",
         11597 => x"80",
         11598 => x"7e",
         11599 => x"56",
         11600 => x"e6",
         11601 => x"ff",
         11602 => x"59",
         11603 => x"75",
         11604 => x"76",
         11605 => x"18",
         11606 => x"08",
         11607 => x"af",
         11608 => x"da",
         11609 => x"79",
         11610 => x"77",
         11611 => x"8a",
         11612 => x"84",
         11613 => x"70",
         11614 => x"e5",
         11615 => x"08",
         11616 => x"59",
         11617 => x"7e",
         11618 => x"38",
         11619 => x"17",
         11620 => x"5f",
         11621 => x"38",
         11622 => x"7a",
         11623 => x"38",
         11624 => x"7a",
         11625 => x"76",
         11626 => x"33",
         11627 => x"05",
         11628 => x"17",
         11629 => x"26",
         11630 => x"7c",
         11631 => x"5e",
         11632 => x"2e",
         11633 => x"81",
         11634 => x"59",
         11635 => x"78",
         11636 => x"0c",
         11637 => x"0d",
         11638 => x"33",
         11639 => x"71",
         11640 => x"90",
         11641 => x"07",
         11642 => x"fd",
         11643 => x"16",
         11644 => x"33",
         11645 => x"71",
         11646 => x"79",
         11647 => x"3d",
         11648 => x"80",
         11649 => x"ff",
         11650 => x"84",
         11651 => x"59",
         11652 => x"08",
         11653 => x"96",
         11654 => x"39",
         11655 => x"16",
         11656 => x"16",
         11657 => x"17",
         11658 => x"ff",
         11659 => x"81",
         11660 => x"8c",
         11661 => x"38",
         11662 => x"08",
         11663 => x"b4",
         11664 => x"17",
         11665 => x"ba",
         11666 => x"55",
         11667 => x"08",
         11668 => x"38",
         11669 => x"55",
         11670 => x"09",
         11671 => x"f6",
         11672 => x"b4",
         11673 => x"17",
         11674 => x"7d",
         11675 => x"33",
         11676 => x"b8",
         11677 => x"fb",
         11678 => x"18",
         11679 => x"08",
         11680 => x"af",
         11681 => x"0b",
         11682 => x"33",
         11683 => x"83",
         11684 => x"70",
         11685 => x"43",
         11686 => x"5a",
         11687 => x"09",
         11688 => x"e8",
         11689 => x"39",
         11690 => x"08",
         11691 => x"59",
         11692 => x"7c",
         11693 => x"5e",
         11694 => x"27",
         11695 => x"80",
         11696 => x"18",
         11697 => x"5a",
         11698 => x"70",
         11699 => x"34",
         11700 => x"d4",
         11701 => x"39",
         11702 => x"7c",
         11703 => x"ba",
         11704 => x"e4",
         11705 => x"f7",
         11706 => x"7d",
         11707 => x"56",
         11708 => x"9f",
         11709 => x"54",
         11710 => x"97",
         11711 => x"53",
         11712 => x"8f",
         11713 => x"22",
         11714 => x"59",
         11715 => x"2e",
         11716 => x"80",
         11717 => x"75",
         11718 => x"c2",
         11719 => x"33",
         11720 => x"ba",
         11721 => x"08",
         11722 => x"26",
         11723 => x"94",
         11724 => x"80",
         11725 => x"2e",
         11726 => x"79",
         11727 => x"70",
         11728 => x"5a",
         11729 => x"2e",
         11730 => x"75",
         11731 => x"51",
         11732 => x"3f",
         11733 => x"08",
         11734 => x"54",
         11735 => x"53",
         11736 => x"3f",
         11737 => x"08",
         11738 => x"d5",
         11739 => x"74",
         11740 => x"17",
         11741 => x"31",
         11742 => x"56",
         11743 => x"80",
         11744 => x"38",
         11745 => x"81",
         11746 => x"76",
         11747 => x"08",
         11748 => x"0c",
         11749 => x"70",
         11750 => x"06",
         11751 => x"78",
         11752 => x"fe",
         11753 => x"74",
         11754 => x"f3",
         11755 => x"8c",
         11756 => x"ba",
         11757 => x"2e",
         11758 => x"73",
         11759 => x"38",
         11760 => x"82",
         11761 => x"53",
         11762 => x"08",
         11763 => x"38",
         11764 => x"0c",
         11765 => x"81",
         11766 => x"34",
         11767 => x"84",
         11768 => x"8b",
         11769 => x"90",
         11770 => x"81",
         11771 => x"55",
         11772 => x"bb",
         11773 => x"16",
         11774 => x"80",
         11775 => x"2e",
         11776 => x"fe",
         11777 => x"94",
         11778 => x"15",
         11779 => x"74",
         11780 => x"73",
         11781 => x"90",
         11782 => x"c0",
         11783 => x"90",
         11784 => x"83",
         11785 => x"78",
         11786 => x"38",
         11787 => x"78",
         11788 => x"77",
         11789 => x"80",
         11790 => x"8c",
         11791 => x"0d",
         11792 => x"94",
         11793 => x"15",
         11794 => x"80",
         11795 => x"38",
         11796 => x"0c",
         11797 => x"80",
         11798 => x"a8",
         11799 => x"8c",
         11800 => x"15",
         11801 => x"16",
         11802 => x"ff",
         11803 => x"80",
         11804 => x"79",
         11805 => x"12",
         11806 => x"5a",
         11807 => x"78",
         11808 => x"38",
         11809 => x"74",
         11810 => x"18",
         11811 => x"89",
         11812 => x"5a",
         11813 => x"2e",
         11814 => x"8c",
         11815 => x"fe",
         11816 => x"52",
         11817 => x"89",
         11818 => x"ba",
         11819 => x"fe",
         11820 => x"14",
         11821 => x"82",
         11822 => x"ba",
         11823 => x"06",
         11824 => x"cf",
         11825 => x"08",
         11826 => x"c9",
         11827 => x"74",
         11828 => x"cb",
         11829 => x"8c",
         11830 => x"ba",
         11831 => x"2e",
         11832 => x"ba",
         11833 => x"2e",
         11834 => x"84",
         11835 => x"88",
         11836 => x"98",
         11837 => x"dc",
         11838 => x"91",
         11839 => x"0b",
         11840 => x"0c",
         11841 => x"04",
         11842 => x"7c",
         11843 => x"75",
         11844 => x"38",
         11845 => x"3d",
         11846 => x"8d",
         11847 => x"51",
         11848 => x"84",
         11849 => x"55",
         11850 => x"08",
         11851 => x"38",
         11852 => x"74",
         11853 => x"ba",
         11854 => x"3d",
         11855 => x"76",
         11856 => x"75",
         11857 => x"97",
         11858 => x"8c",
         11859 => x"ba",
         11860 => x"d1",
         11861 => x"33",
         11862 => x"59",
         11863 => x"24",
         11864 => x"16",
         11865 => x"2a",
         11866 => x"54",
         11867 => x"80",
         11868 => x"16",
         11869 => x"33",
         11870 => x"71",
         11871 => x"7d",
         11872 => x"5d",
         11873 => x"78",
         11874 => x"38",
         11875 => x"0c",
         11876 => x"18",
         11877 => x"23",
         11878 => x"51",
         11879 => x"3f",
         11880 => x"08",
         11881 => x"2e",
         11882 => x"80",
         11883 => x"38",
         11884 => x"fe",
         11885 => x"55",
         11886 => x"fe",
         11887 => x"17",
         11888 => x"33",
         11889 => x"71",
         11890 => x"7a",
         11891 => x"0c",
         11892 => x"bc",
         11893 => x"0d",
         11894 => x"54",
         11895 => x"9e",
         11896 => x"53",
         11897 => x"96",
         11898 => x"52",
         11899 => x"8e",
         11900 => x"22",
         11901 => x"57",
         11902 => x"2e",
         11903 => x"52",
         11904 => x"84",
         11905 => x"0c",
         11906 => x"8c",
         11907 => x"0d",
         11908 => x"33",
         11909 => x"c3",
         11910 => x"8c",
         11911 => x"52",
         11912 => x"71",
         11913 => x"54",
         11914 => x"3d",
         11915 => x"58",
         11916 => x"74",
         11917 => x"38",
         11918 => x"73",
         11919 => x"38",
         11920 => x"72",
         11921 => x"38",
         11922 => x"84",
         11923 => x"53",
         11924 => x"81",
         11925 => x"53",
         11926 => x"53",
         11927 => x"38",
         11928 => x"80",
         11929 => x"52",
         11930 => x"9d",
         11931 => x"ba",
         11932 => x"84",
         11933 => x"84",
         11934 => x"84",
         11935 => x"a6",
         11936 => x"74",
         11937 => x"92",
         11938 => x"74",
         11939 => x"be",
         11940 => x"8c",
         11941 => x"70",
         11942 => x"07",
         11943 => x"ba",
         11944 => x"55",
         11945 => x"84",
         11946 => x"8a",
         11947 => x"75",
         11948 => x"52",
         11949 => x"e2",
         11950 => x"74",
         11951 => x"8e",
         11952 => x"8c",
         11953 => x"70",
         11954 => x"07",
         11955 => x"ba",
         11956 => x"55",
         11957 => x"39",
         11958 => x"51",
         11959 => x"3f",
         11960 => x"08",
         11961 => x"0c",
         11962 => x"04",
         11963 => x"51",
         11964 => x"3f",
         11965 => x"08",
         11966 => x"72",
         11967 => x"72",
         11968 => x"56",
         11969 => x"ed",
         11970 => x"57",
         11971 => x"3d",
         11972 => x"3d",
         11973 => x"a5",
         11974 => x"8c",
         11975 => x"ba",
         11976 => x"2e",
         11977 => x"84",
         11978 => x"95",
         11979 => x"65",
         11980 => x"ff",
         11981 => x"84",
         11982 => x"55",
         11983 => x"08",
         11984 => x"80",
         11985 => x"70",
         11986 => x"58",
         11987 => x"97",
         11988 => x"2e",
         11989 => x"52",
         11990 => x"b0",
         11991 => x"84",
         11992 => x"95",
         11993 => x"86",
         11994 => x"8c",
         11995 => x"0d",
         11996 => x"0d",
         11997 => x"5f",
         11998 => x"3d",
         11999 => x"96",
         12000 => x"b9",
         12001 => x"8c",
         12002 => x"ba",
         12003 => x"38",
         12004 => x"74",
         12005 => x"08",
         12006 => x"13",
         12007 => x"59",
         12008 => x"26",
         12009 => x"7f",
         12010 => x"ba",
         12011 => x"3d",
         12012 => x"ba",
         12013 => x"33",
         12014 => x"81",
         12015 => x"38",
         12016 => x"08",
         12017 => x"08",
         12018 => x"77",
         12019 => x"7b",
         12020 => x"5c",
         12021 => x"17",
         12022 => x"82",
         12023 => x"17",
         12024 => x"5d",
         12025 => x"38",
         12026 => x"53",
         12027 => x"81",
         12028 => x"fe",
         12029 => x"84",
         12030 => x"80",
         12031 => x"ff",
         12032 => x"79",
         12033 => x"7f",
         12034 => x"7d",
         12035 => x"76",
         12036 => x"82",
         12037 => x"38",
         12038 => x"05",
         12039 => x"82",
         12040 => x"90",
         12041 => x"2b",
         12042 => x"33",
         12043 => x"88",
         12044 => x"71",
         12045 => x"fe",
         12046 => x"70",
         12047 => x"25",
         12048 => x"84",
         12049 => x"06",
         12050 => x"43",
         12051 => x"54",
         12052 => x"40",
         12053 => x"fe",
         12054 => x"7f",
         12055 => x"18",
         12056 => x"33",
         12057 => x"77",
         12058 => x"79",
         12059 => x"0c",
         12060 => x"04",
         12061 => x"17",
         12062 => x"17",
         12063 => x"18",
         12064 => x"fe",
         12065 => x"81",
         12066 => x"8c",
         12067 => x"38",
         12068 => x"08",
         12069 => x"b4",
         12070 => x"18",
         12071 => x"ba",
         12072 => x"55",
         12073 => x"08",
         12074 => x"38",
         12075 => x"55",
         12076 => x"09",
         12077 => x"b0",
         12078 => x"b4",
         12079 => x"18",
         12080 => x"7c",
         12081 => x"33",
         12082 => x"e0",
         12083 => x"fe",
         12084 => x"77",
         12085 => x"59",
         12086 => x"77",
         12087 => x"80",
         12088 => x"8c",
         12089 => x"80",
         12090 => x"ba",
         12091 => x"2e",
         12092 => x"84",
         12093 => x"30",
         12094 => x"8c",
         12095 => x"25",
         12096 => x"18",
         12097 => x"5c",
         12098 => x"08",
         12099 => x"38",
         12100 => x"7a",
         12101 => x"84",
         12102 => x"07",
         12103 => x"18",
         12104 => x"39",
         12105 => x"05",
         12106 => x"71",
         12107 => x"2b",
         12108 => x"70",
         12109 => x"82",
         12110 => x"06",
         12111 => x"5d",
         12112 => x"5f",
         12113 => x"83",
         12114 => x"39",
         12115 => x"bf",
         12116 => x"58",
         12117 => x"0c",
         12118 => x"0c",
         12119 => x"81",
         12120 => x"84",
         12121 => x"83",
         12122 => x"58",
         12123 => x"f7",
         12124 => x"57",
         12125 => x"80",
         12126 => x"76",
         12127 => x"80",
         12128 => x"74",
         12129 => x"80",
         12130 => x"86",
         12131 => x"18",
         12132 => x"78",
         12133 => x"da",
         12134 => x"73",
         12135 => x"dc",
         12136 => x"33",
         12137 => x"d4",
         12138 => x"33",
         12139 => x"81",
         12140 => x"87",
         12141 => x"2e",
         12142 => x"94",
         12143 => x"73",
         12144 => x"27",
         12145 => x"81",
         12146 => x"17",
         12147 => x"57",
         12148 => x"27",
         12149 => x"16",
         12150 => x"b3",
         12151 => x"80",
         12152 => x"0c",
         12153 => x"8c",
         12154 => x"80",
         12155 => x"78",
         12156 => x"75",
         12157 => x"38",
         12158 => x"34",
         12159 => x"84",
         12160 => x"8b",
         12161 => x"78",
         12162 => x"27",
         12163 => x"73",
         12164 => x"fe",
         12165 => x"84",
         12166 => x"59",
         12167 => x"08",
         12168 => x"e9",
         12169 => x"8c",
         12170 => x"82",
         12171 => x"ba",
         12172 => x"2e",
         12173 => x"80",
         12174 => x"75",
         12175 => x"81",
         12176 => x"8c",
         12177 => x"38",
         12178 => x"fe",
         12179 => x"08",
         12180 => x"74",
         12181 => x"af",
         12182 => x"94",
         12183 => x"16",
         12184 => x"54",
         12185 => x"34",
         12186 => x"79",
         12187 => x"38",
         12188 => x"15",
         12189 => x"f6",
         12190 => x"ba",
         12191 => x"06",
         12192 => x"95",
         12193 => x"08",
         12194 => x"8f",
         12195 => x"90",
         12196 => x"54",
         12197 => x"0b",
         12198 => x"fe",
         12199 => x"17",
         12200 => x"51",
         12201 => x"3f",
         12202 => x"08",
         12203 => x"c2",
         12204 => x"8c",
         12205 => x"81",
         12206 => x"81",
         12207 => x"58",
         12208 => x"08",
         12209 => x"27",
         12210 => x"84",
         12211 => x"98",
         12212 => x"08",
         12213 => x"81",
         12214 => x"8c",
         12215 => x"a1",
         12216 => x"8c",
         12217 => x"08",
         12218 => x"38",
         12219 => x"97",
         12220 => x"74",
         12221 => x"ff",
         12222 => x"84",
         12223 => x"55",
         12224 => x"08",
         12225 => x"73",
         12226 => x"fe",
         12227 => x"84",
         12228 => x"59",
         12229 => x"08",
         12230 => x"cb",
         12231 => x"8c",
         12232 => x"80",
         12233 => x"ba",
         12234 => x"2e",
         12235 => x"80",
         12236 => x"75",
         12237 => x"89",
         12238 => x"8c",
         12239 => x"38",
         12240 => x"fe",
         12241 => x"08",
         12242 => x"74",
         12243 => x"38",
         12244 => x"17",
         12245 => x"33",
         12246 => x"73",
         12247 => x"78",
         12248 => x"26",
         12249 => x"80",
         12250 => x"90",
         12251 => x"fc",
         12252 => x"56",
         12253 => x"82",
         12254 => x"33",
         12255 => x"e4",
         12256 => x"e7",
         12257 => x"90",
         12258 => x"54",
         12259 => x"84",
         12260 => x"90",
         12261 => x"54",
         12262 => x"81",
         12263 => x"33",
         12264 => x"f0",
         12265 => x"8c",
         12266 => x"39",
         12267 => x"bb",
         12268 => x"0d",
         12269 => x"3d",
         12270 => x"52",
         12271 => x"ff",
         12272 => x"84",
         12273 => x"56",
         12274 => x"08",
         12275 => x"38",
         12276 => x"8c",
         12277 => x"0d",
         12278 => x"a8",
         12279 => x"9b",
         12280 => x"59",
         12281 => x"3f",
         12282 => x"08",
         12283 => x"8c",
         12284 => x"02",
         12285 => x"33",
         12286 => x"81",
         12287 => x"86",
         12288 => x"38",
         12289 => x"5b",
         12290 => x"c4",
         12291 => x"ee",
         12292 => x"81",
         12293 => x"87",
         12294 => x"b4",
         12295 => x"3d",
         12296 => x"33",
         12297 => x"71",
         12298 => x"73",
         12299 => x"5c",
         12300 => x"83",
         12301 => x"38",
         12302 => x"81",
         12303 => x"80",
         12304 => x"38",
         12305 => x"18",
         12306 => x"ff",
         12307 => x"5f",
         12308 => x"ba",
         12309 => x"8f",
         12310 => x"55",
         12311 => x"3f",
         12312 => x"08",
         12313 => x"8c",
         12314 => x"38",
         12315 => x"08",
         12316 => x"ff",
         12317 => x"84",
         12318 => x"56",
         12319 => x"08",
         12320 => x"0b",
         12321 => x"0c",
         12322 => x"04",
         12323 => x"94",
         12324 => x"98",
         12325 => x"2b",
         12326 => x"5d",
         12327 => x"98",
         12328 => x"8c",
         12329 => x"88",
         12330 => x"8c",
         12331 => x"38",
         12332 => x"a8",
         12333 => x"5d",
         12334 => x"2e",
         12335 => x"74",
         12336 => x"ff",
         12337 => x"84",
         12338 => x"56",
         12339 => x"08",
         12340 => x"38",
         12341 => x"77",
         12342 => x"56",
         12343 => x"2e",
         12344 => x"80",
         12345 => x"7a",
         12346 => x"55",
         12347 => x"89",
         12348 => x"08",
         12349 => x"fd",
         12350 => x"75",
         12351 => x"7d",
         12352 => x"db",
         12353 => x"8c",
         12354 => x"8c",
         12355 => x"0d",
         12356 => x"5d",
         12357 => x"56",
         12358 => x"17",
         12359 => x"82",
         12360 => x"17",
         12361 => x"55",
         12362 => x"09",
         12363 => x"dd",
         12364 => x"75",
         12365 => x"52",
         12366 => x"51",
         12367 => x"3f",
         12368 => x"08",
         12369 => x"38",
         12370 => x"58",
         12371 => x"0c",
         12372 => x"ab",
         12373 => x"08",
         12374 => x"34",
         12375 => x"18",
         12376 => x"08",
         12377 => x"ec",
         12378 => x"78",
         12379 => x"de",
         12380 => x"8c",
         12381 => x"ba",
         12382 => x"2e",
         12383 => x"75",
         12384 => x"81",
         12385 => x"38",
         12386 => x"c8",
         12387 => x"b4",
         12388 => x"7c",
         12389 => x"33",
         12390 => x"90",
         12391 => x"84",
         12392 => x"7a",
         12393 => x"06",
         12394 => x"84",
         12395 => x"83",
         12396 => x"17",
         12397 => x"08",
         12398 => x"8c",
         12399 => x"74",
         12400 => x"27",
         12401 => x"82",
         12402 => x"74",
         12403 => x"81",
         12404 => x"38",
         12405 => x"17",
         12406 => x"08",
         12407 => x"52",
         12408 => x"51",
         12409 => x"3f",
         12410 => x"c5",
         12411 => x"79",
         12412 => x"e1",
         12413 => x"78",
         12414 => x"e4",
         12415 => x"8c",
         12416 => x"ba",
         12417 => x"2e",
         12418 => x"84",
         12419 => x"81",
         12420 => x"38",
         12421 => x"08",
         12422 => x"cb",
         12423 => x"74",
         12424 => x"fe",
         12425 => x"84",
         12426 => x"b3",
         12427 => x"08",
         12428 => x"19",
         12429 => x"58",
         12430 => x"ff",
         12431 => x"16",
         12432 => x"84",
         12433 => x"07",
         12434 => x"18",
         12435 => x"77",
         12436 => x"a1",
         12437 => x"fd",
         12438 => x"56",
         12439 => x"84",
         12440 => x"56",
         12441 => x"81",
         12442 => x"39",
         12443 => x"82",
         12444 => x"ff",
         12445 => x"a0",
         12446 => x"b2",
         12447 => x"ba",
         12448 => x"84",
         12449 => x"80",
         12450 => x"75",
         12451 => x"0c",
         12452 => x"04",
         12453 => x"52",
         12454 => x"52",
         12455 => x"bf",
         12456 => x"8c",
         12457 => x"ba",
         12458 => x"38",
         12459 => x"ba",
         12460 => x"3d",
         12461 => x"ba",
         12462 => x"2e",
         12463 => x"cb",
         12464 => x"f3",
         12465 => x"85",
         12466 => x"56",
         12467 => x"74",
         12468 => x"7d",
         12469 => x"8f",
         12470 => x"5d",
         12471 => x"3f",
         12472 => x"08",
         12473 => x"84",
         12474 => x"83",
         12475 => x"84",
         12476 => x"81",
         12477 => x"38",
         12478 => x"08",
         12479 => x"cb",
         12480 => x"c9",
         12481 => x"ba",
         12482 => x"12",
         12483 => x"57",
         12484 => x"38",
         12485 => x"18",
         12486 => x"5a",
         12487 => x"75",
         12488 => x"38",
         12489 => x"76",
         12490 => x"19",
         12491 => x"58",
         12492 => x"0c",
         12493 => x"84",
         12494 => x"55",
         12495 => x"81",
         12496 => x"ff",
         12497 => x"f4",
         12498 => x"8a",
         12499 => x"77",
         12500 => x"f9",
         12501 => x"77",
         12502 => x"52",
         12503 => x"51",
         12504 => x"3f",
         12505 => x"08",
         12506 => x"81",
         12507 => x"39",
         12508 => x"84",
         12509 => x"b4",
         12510 => x"b8",
         12511 => x"81",
         12512 => x"58",
         12513 => x"3f",
         12514 => x"ba",
         12515 => x"38",
         12516 => x"08",
         12517 => x"b4",
         12518 => x"18",
         12519 => x"74",
         12520 => x"27",
         12521 => x"82",
         12522 => x"7a",
         12523 => x"81",
         12524 => x"38",
         12525 => x"17",
         12526 => x"08",
         12527 => x"52",
         12528 => x"51",
         12529 => x"3f",
         12530 => x"81",
         12531 => x"08",
         12532 => x"7c",
         12533 => x"38",
         12534 => x"08",
         12535 => x"38",
         12536 => x"51",
         12537 => x"3f",
         12538 => x"08",
         12539 => x"8c",
         12540 => x"fd",
         12541 => x"ba",
         12542 => x"2e",
         12543 => x"84",
         12544 => x"ff",
         12545 => x"38",
         12546 => x"52",
         12547 => x"f9",
         12548 => x"ba",
         12549 => x"f3",
         12550 => x"08",
         12551 => x"19",
         12552 => x"59",
         12553 => x"90",
         12554 => x"94",
         12555 => x"17",
         12556 => x"5c",
         12557 => x"34",
         12558 => x"7a",
         12559 => x"38",
         12560 => x"8c",
         12561 => x"0d",
         12562 => x"22",
         12563 => x"ff",
         12564 => x"81",
         12565 => x"2e",
         12566 => x"fe",
         12567 => x"0b",
         12568 => x"56",
         12569 => x"81",
         12570 => x"ff",
         12571 => x"f4",
         12572 => x"ae",
         12573 => x"34",
         12574 => x"0b",
         12575 => x"34",
         12576 => x"80",
         12577 => x"75",
         12578 => x"34",
         12579 => x"d0",
         12580 => x"cc",
         12581 => x"1a",
         12582 => x"83",
         12583 => x"59",
         12584 => x"d2",
         12585 => x"88",
         12586 => x"80",
         12587 => x"75",
         12588 => x"83",
         12589 => x"38",
         12590 => x"0b",
         12591 => x"b8",
         12592 => x"56",
         12593 => x"05",
         12594 => x"70",
         12595 => x"34",
         12596 => x"75",
         12597 => x"56",
         12598 => x"d9",
         12599 => x"7e",
         12600 => x"ff",
         12601 => x"57",
         12602 => x"17",
         12603 => x"2a",
         12604 => x"f3",
         12605 => x"33",
         12606 => x"2e",
         12607 => x"7d",
         12608 => x"83",
         12609 => x"51",
         12610 => x"3f",
         12611 => x"08",
         12612 => x"8c",
         12613 => x"38",
         12614 => x"ba",
         12615 => x"17",
         12616 => x"8c",
         12617 => x"34",
         12618 => x"17",
         12619 => x"0b",
         12620 => x"7d",
         12621 => x"77",
         12622 => x"77",
         12623 => x"78",
         12624 => x"7c",
         12625 => x"83",
         12626 => x"38",
         12627 => x"0b",
         12628 => x"7d",
         12629 => x"83",
         12630 => x"51",
         12631 => x"3f",
         12632 => x"08",
         12633 => x"ba",
         12634 => x"3d",
         12635 => x"90",
         12636 => x"80",
         12637 => x"74",
         12638 => x"76",
         12639 => x"34",
         12640 => x"7b",
         12641 => x"7a",
         12642 => x"34",
         12643 => x"55",
         12644 => x"17",
         12645 => x"a0",
         12646 => x"1a",
         12647 => x"58",
         12648 => x"39",
         12649 => x"58",
         12650 => x"34",
         12651 => x"5c",
         12652 => x"34",
         12653 => x"0b",
         12654 => x"7d",
         12655 => x"83",
         12656 => x"51",
         12657 => x"3f",
         12658 => x"08",
         12659 => x"39",
         12660 => x"b3",
         12661 => x"08",
         12662 => x"5f",
         12663 => x"9b",
         12664 => x"81",
         12665 => x"70",
         12666 => x"56",
         12667 => x"81",
         12668 => x"ed",
         12669 => x"2e",
         12670 => x"82",
         12671 => x"fe",
         12672 => x"b2",
         12673 => x"ab",
         12674 => x"ba",
         12675 => x"84",
         12676 => x"80",
         12677 => x"75",
         12678 => x"0c",
         12679 => x"04",
         12680 => x"0c",
         12681 => x"52",
         12682 => x"52",
         12683 => x"af",
         12684 => x"8c",
         12685 => x"ba",
         12686 => x"38",
         12687 => x"05",
         12688 => x"06",
         12689 => x"7c",
         12690 => x"0b",
         12691 => x"3d",
         12692 => x"55",
         12693 => x"05",
         12694 => x"70",
         12695 => x"34",
         12696 => x"74",
         12697 => x"3d",
         12698 => x"7a",
         12699 => x"75",
         12700 => x"57",
         12701 => x"81",
         12702 => x"ff",
         12703 => x"ef",
         12704 => x"08",
         12705 => x"ff",
         12706 => x"84",
         12707 => x"56",
         12708 => x"08",
         12709 => x"6a",
         12710 => x"2e",
         12711 => x"88",
         12712 => x"8c",
         12713 => x"0d",
         12714 => x"d0",
         12715 => x"ff",
         12716 => x"58",
         12717 => x"91",
         12718 => x"78",
         12719 => x"d0",
         12720 => x"78",
         12721 => x"fa",
         12722 => x"08",
         12723 => x"70",
         12724 => x"5e",
         12725 => x"7a",
         12726 => x"5c",
         12727 => x"81",
         12728 => x"ff",
         12729 => x"58",
         12730 => x"26",
         12731 => x"16",
         12732 => x"06",
         12733 => x"9f",
         12734 => x"99",
         12735 => x"e0",
         12736 => x"ff",
         12737 => x"75",
         12738 => x"2a",
         12739 => x"77",
         12740 => x"06",
         12741 => x"ff",
         12742 => x"7a",
         12743 => x"70",
         12744 => x"2a",
         12745 => x"58",
         12746 => x"2e",
         12747 => x"1c",
         12748 => x"5c",
         12749 => x"fd",
         12750 => x"08",
         12751 => x"ff",
         12752 => x"83",
         12753 => x"38",
         12754 => x"82",
         12755 => x"fe",
         12756 => x"b2",
         12757 => x"a8",
         12758 => x"ba",
         12759 => x"84",
         12760 => x"fd",
         12761 => x"b8",
         12762 => x"3d",
         12763 => x"81",
         12764 => x"38",
         12765 => x"8d",
         12766 => x"ba",
         12767 => x"84",
         12768 => x"fd",
         12769 => x"58",
         12770 => x"19",
         12771 => x"80",
         12772 => x"56",
         12773 => x"81",
         12774 => x"75",
         12775 => x"57",
         12776 => x"5a",
         12777 => x"02",
         12778 => x"33",
         12779 => x"8b",
         12780 => x"84",
         12781 => x"40",
         12782 => x"38",
         12783 => x"57",
         12784 => x"34",
         12785 => x"0b",
         12786 => x"8b",
         12787 => x"84",
         12788 => x"57",
         12789 => x"2e",
         12790 => x"a7",
         12791 => x"2e",
         12792 => x"7f",
         12793 => x"9a",
         12794 => x"88",
         12795 => x"33",
         12796 => x"57",
         12797 => x"82",
         12798 => x"16",
         12799 => x"fe",
         12800 => x"75",
         12801 => x"c7",
         12802 => x"22",
         12803 => x"b0",
         12804 => x"57",
         12805 => x"2e",
         12806 => x"75",
         12807 => x"b4",
         12808 => x"2e",
         12809 => x"17",
         12810 => x"83",
         12811 => x"54",
         12812 => x"17",
         12813 => x"33",
         12814 => x"f1",
         12815 => x"8c",
         12816 => x"85",
         12817 => x"81",
         12818 => x"18",
         12819 => x"7b",
         12820 => x"56",
         12821 => x"bf",
         12822 => x"33",
         12823 => x"2e",
         12824 => x"bb",
         12825 => x"83",
         12826 => x"5d",
         12827 => x"f2",
         12828 => x"88",
         12829 => x"80",
         12830 => x"76",
         12831 => x"83",
         12832 => x"06",
         12833 => x"90",
         12834 => x"80",
         12835 => x"7d",
         12836 => x"75",
         12837 => x"34",
         12838 => x"0b",
         12839 => x"78",
         12840 => x"08",
         12841 => x"57",
         12842 => x"ff",
         12843 => x"74",
         12844 => x"fe",
         12845 => x"84",
         12846 => x"55",
         12847 => x"08",
         12848 => x"b8",
         12849 => x"19",
         12850 => x"5a",
         12851 => x"77",
         12852 => x"83",
         12853 => x"59",
         12854 => x"2e",
         12855 => x"81",
         12856 => x"54",
         12857 => x"16",
         12858 => x"33",
         12859 => x"bd",
         12860 => x"8c",
         12861 => x"85",
         12862 => x"81",
         12863 => x"17",
         12864 => x"77",
         12865 => x"19",
         12866 => x"7a",
         12867 => x"83",
         12868 => x"19",
         12869 => x"a5",
         12870 => x"78",
         12871 => x"ae",
         12872 => x"8c",
         12873 => x"ba",
         12874 => x"2e",
         12875 => x"82",
         12876 => x"2e",
         12877 => x"74",
         12878 => x"db",
         12879 => x"fe",
         12880 => x"84",
         12881 => x"84",
         12882 => x"b1",
         12883 => x"82",
         12884 => x"8c",
         12885 => x"0d",
         12886 => x"33",
         12887 => x"71",
         12888 => x"90",
         12889 => x"07",
         12890 => x"fd",
         12891 => x"ba",
         12892 => x"2e",
         12893 => x"84",
         12894 => x"80",
         12895 => x"38",
         12896 => x"8c",
         12897 => x"0d",
         12898 => x"b4",
         12899 => x"7b",
         12900 => x"33",
         12901 => x"94",
         12902 => x"84",
         12903 => x"7a",
         12904 => x"06",
         12905 => x"84",
         12906 => x"83",
         12907 => x"16",
         12908 => x"08",
         12909 => x"8c",
         12910 => x"74",
         12911 => x"27",
         12912 => x"82",
         12913 => x"7c",
         12914 => x"81",
         12915 => x"38",
         12916 => x"16",
         12917 => x"08",
         12918 => x"52",
         12919 => x"51",
         12920 => x"3f",
         12921 => x"fa",
         12922 => x"b4",
         12923 => x"b8",
         12924 => x"81",
         12925 => x"5b",
         12926 => x"3f",
         12927 => x"ba",
         12928 => x"c9",
         12929 => x"8c",
         12930 => x"34",
         12931 => x"a8",
         12932 => x"84",
         12933 => x"5d",
         12934 => x"18",
         12935 => x"8e",
         12936 => x"33",
         12937 => x"2e",
         12938 => x"fc",
         12939 => x"54",
         12940 => x"a0",
         12941 => x"53",
         12942 => x"17",
         12943 => x"e0",
         12944 => x"5c",
         12945 => x"ec",
         12946 => x"80",
         12947 => x"02",
         12948 => x"e3",
         12949 => x"57",
         12950 => x"3d",
         12951 => x"97",
         12952 => x"a2",
         12953 => x"ba",
         12954 => x"84",
         12955 => x"80",
         12956 => x"75",
         12957 => x"0c",
         12958 => x"04",
         12959 => x"52",
         12960 => x"05",
         12961 => x"d7",
         12962 => x"8c",
         12963 => x"ba",
         12964 => x"38",
         12965 => x"05",
         12966 => x"06",
         12967 => x"73",
         12968 => x"a7",
         12969 => x"09",
         12970 => x"71",
         12971 => x"06",
         12972 => x"57",
         12973 => x"17",
         12974 => x"81",
         12975 => x"34",
         12976 => x"e2",
         12977 => x"ba",
         12978 => x"ba",
         12979 => x"3d",
         12980 => x"3d",
         12981 => x"82",
         12982 => x"cc",
         12983 => x"3d",
         12984 => x"d9",
         12985 => x"8c",
         12986 => x"ba",
         12987 => x"2e",
         12988 => x"84",
         12989 => x"96",
         12990 => x"78",
         12991 => x"96",
         12992 => x"51",
         12993 => x"3f",
         12994 => x"08",
         12995 => x"8c",
         12996 => x"02",
         12997 => x"33",
         12998 => x"56",
         12999 => x"d2",
         13000 => x"18",
         13001 => x"22",
         13002 => x"07",
         13003 => x"76",
         13004 => x"76",
         13005 => x"74",
         13006 => x"76",
         13007 => x"77",
         13008 => x"76",
         13009 => x"73",
         13010 => x"78",
         13011 => x"83",
         13012 => x"51",
         13013 => x"3f",
         13014 => x"08",
         13015 => x"0c",
         13016 => x"04",
         13017 => x"6b",
         13018 => x"80",
         13019 => x"cc",
         13020 => x"3d",
         13021 => x"c5",
         13022 => x"8c",
         13023 => x"8c",
         13024 => x"84",
         13025 => x"07",
         13026 => x"56",
         13027 => x"2e",
         13028 => x"70",
         13029 => x"56",
         13030 => x"38",
         13031 => x"78",
         13032 => x"56",
         13033 => x"2e",
         13034 => x"81",
         13035 => x"5a",
         13036 => x"2e",
         13037 => x"7c",
         13038 => x"58",
         13039 => x"b4",
         13040 => x"2e",
         13041 => x"83",
         13042 => x"5a",
         13043 => x"2e",
         13044 => x"81",
         13045 => x"54",
         13046 => x"16",
         13047 => x"33",
         13048 => x"c9",
         13049 => x"8c",
         13050 => x"85",
         13051 => x"81",
         13052 => x"17",
         13053 => x"78",
         13054 => x"70",
         13055 => x"80",
         13056 => x"83",
         13057 => x"80",
         13058 => x"84",
         13059 => x"a7",
         13060 => x"b8",
         13061 => x"33",
         13062 => x"71",
         13063 => x"88",
         13064 => x"14",
         13065 => x"07",
         13066 => x"33",
         13067 => x"0c",
         13068 => x"57",
         13069 => x"84",
         13070 => x"9a",
         13071 => x"7c",
         13072 => x"80",
         13073 => x"70",
         13074 => x"f4",
         13075 => x"ba",
         13076 => x"84",
         13077 => x"80",
         13078 => x"38",
         13079 => x"09",
         13080 => x"b8",
         13081 => x"34",
         13082 => x"b0",
         13083 => x"b4",
         13084 => x"b8",
         13085 => x"81",
         13086 => x"5b",
         13087 => x"3f",
         13088 => x"ba",
         13089 => x"2e",
         13090 => x"fe",
         13091 => x"ba",
         13092 => x"17",
         13093 => x"08",
         13094 => x"31",
         13095 => x"08",
         13096 => x"a0",
         13097 => x"fe",
         13098 => x"16",
         13099 => x"82",
         13100 => x"06",
         13101 => x"77",
         13102 => x"08",
         13103 => x"05",
         13104 => x"81",
         13105 => x"fe",
         13106 => x"79",
         13107 => x"76",
         13108 => x"52",
         13109 => x"51",
         13110 => x"3f",
         13111 => x"08",
         13112 => x"8d",
         13113 => x"39",
         13114 => x"51",
         13115 => x"3f",
         13116 => x"08",
         13117 => x"8c",
         13118 => x"38",
         13119 => x"08",
         13120 => x"08",
         13121 => x"59",
         13122 => x"19",
         13123 => x"59",
         13124 => x"75",
         13125 => x"59",
         13126 => x"ec",
         13127 => x"1c",
         13128 => x"76",
         13129 => x"2e",
         13130 => x"ff",
         13131 => x"70",
         13132 => x"58",
         13133 => x"ea",
         13134 => x"39",
         13135 => x"ba",
         13136 => x"0d",
         13137 => x"3d",
         13138 => x"52",
         13139 => x"ff",
         13140 => x"84",
         13141 => x"56",
         13142 => x"08",
         13143 => x"8f",
         13144 => x"7d",
         13145 => x"76",
         13146 => x"58",
         13147 => x"55",
         13148 => x"74",
         13149 => x"70",
         13150 => x"ff",
         13151 => x"58",
         13152 => x"27",
         13153 => x"a2",
         13154 => x"5c",
         13155 => x"ff",
         13156 => x"57",
         13157 => x"f5",
         13158 => x"0c",
         13159 => x"ff",
         13160 => x"38",
         13161 => x"95",
         13162 => x"52",
         13163 => x"08",
         13164 => x"3f",
         13165 => x"08",
         13166 => x"06",
         13167 => x"2e",
         13168 => x"83",
         13169 => x"83",
         13170 => x"70",
         13171 => x"5b",
         13172 => x"80",
         13173 => x"38",
         13174 => x"77",
         13175 => x"81",
         13176 => x"70",
         13177 => x"57",
         13178 => x"80",
         13179 => x"74",
         13180 => x"81",
         13181 => x"75",
         13182 => x"59",
         13183 => x"38",
         13184 => x"27",
         13185 => x"79",
         13186 => x"96",
         13187 => x"77",
         13188 => x"76",
         13189 => x"74",
         13190 => x"05",
         13191 => x"1a",
         13192 => x"70",
         13193 => x"34",
         13194 => x"3d",
         13195 => x"70",
         13196 => x"5b",
         13197 => x"77",
         13198 => x"d1",
         13199 => x"33",
         13200 => x"76",
         13201 => x"bc",
         13202 => x"2e",
         13203 => x"b7",
         13204 => x"16",
         13205 => x"5c",
         13206 => x"09",
         13207 => x"38",
         13208 => x"79",
         13209 => x"45",
         13210 => x"52",
         13211 => x"52",
         13212 => x"e4",
         13213 => x"8c",
         13214 => x"ba",
         13215 => x"2e",
         13216 => x"56",
         13217 => x"8c",
         13218 => x"0d",
         13219 => x"52",
         13220 => x"e7",
         13221 => x"8c",
         13222 => x"ff",
         13223 => x"fd",
         13224 => x"56",
         13225 => x"8c",
         13226 => x"0d",
         13227 => x"9c",
         13228 => x"c3",
         13229 => x"75",
         13230 => x"ee",
         13231 => x"8c",
         13232 => x"ba",
         13233 => x"c1",
         13234 => x"2e",
         13235 => x"8b",
         13236 => x"57",
         13237 => x"81",
         13238 => x"76",
         13239 => x"58",
         13240 => x"55",
         13241 => x"7d",
         13242 => x"83",
         13243 => x"51",
         13244 => x"3f",
         13245 => x"08",
         13246 => x"ff",
         13247 => x"7a",
         13248 => x"38",
         13249 => x"9c",
         13250 => x"8c",
         13251 => x"09",
         13252 => x"ee",
         13253 => x"79",
         13254 => x"e6",
         13255 => x"75",
         13256 => x"58",
         13257 => x"3f",
         13258 => x"08",
         13259 => x"8c",
         13260 => x"09",
         13261 => x"84",
         13262 => x"8c",
         13263 => x"5c",
         13264 => x"08",
         13265 => x"b4",
         13266 => x"2e",
         13267 => x"18",
         13268 => x"79",
         13269 => x"06",
         13270 => x"81",
         13271 => x"b8",
         13272 => x"18",
         13273 => x"d5",
         13274 => x"ba",
         13275 => x"2e",
         13276 => x"57",
         13277 => x"b4",
         13278 => x"57",
         13279 => x"78",
         13280 => x"70",
         13281 => x"57",
         13282 => x"2e",
         13283 => x"74",
         13284 => x"25",
         13285 => x"5c",
         13286 => x"81",
         13287 => x"1a",
         13288 => x"2e",
         13289 => x"52",
         13290 => x"ef",
         13291 => x"ba",
         13292 => x"84",
         13293 => x"80",
         13294 => x"38",
         13295 => x"84",
         13296 => x"38",
         13297 => x"fd",
         13298 => x"6c",
         13299 => x"76",
         13300 => x"58",
         13301 => x"55",
         13302 => x"6b",
         13303 => x"8b",
         13304 => x"6c",
         13305 => x"55",
         13306 => x"05",
         13307 => x"70",
         13308 => x"34",
         13309 => x"74",
         13310 => x"eb",
         13311 => x"81",
         13312 => x"76",
         13313 => x"58",
         13314 => x"55",
         13315 => x"fd",
         13316 => x"5a",
         13317 => x"7d",
         13318 => x"83",
         13319 => x"51",
         13320 => x"3f",
         13321 => x"08",
         13322 => x"39",
         13323 => x"df",
         13324 => x"b4",
         13325 => x"7a",
         13326 => x"33",
         13327 => x"ec",
         13328 => x"8c",
         13329 => x"09",
         13330 => x"c3",
         13331 => x"8c",
         13332 => x"34",
         13333 => x"a8",
         13334 => x"5c",
         13335 => x"08",
         13336 => x"82",
         13337 => x"74",
         13338 => x"38",
         13339 => x"08",
         13340 => x"39",
         13341 => x"52",
         13342 => x"ed",
         13343 => x"ba",
         13344 => x"84",
         13345 => x"80",
         13346 => x"38",
         13347 => x"81",
         13348 => x"78",
         13349 => x"e7",
         13350 => x"39",
         13351 => x"18",
         13352 => x"08",
         13353 => x"52",
         13354 => x"51",
         13355 => x"3f",
         13356 => x"f2",
         13357 => x"62",
         13358 => x"80",
         13359 => x"5e",
         13360 => x"56",
         13361 => x"9f",
         13362 => x"55",
         13363 => x"97",
         13364 => x"54",
         13365 => x"8f",
         13366 => x"22",
         13367 => x"59",
         13368 => x"2e",
         13369 => x"80",
         13370 => x"75",
         13371 => x"91",
         13372 => x"75",
         13373 => x"79",
         13374 => x"a2",
         13375 => x"08",
         13376 => x"90",
         13377 => x"81",
         13378 => x"56",
         13379 => x"2e",
         13380 => x"7e",
         13381 => x"70",
         13382 => x"55",
         13383 => x"5c",
         13384 => x"82",
         13385 => x"7a",
         13386 => x"70",
         13387 => x"2a",
         13388 => x"08",
         13389 => x"08",
         13390 => x"5f",
         13391 => x"78",
         13392 => x"9c",
         13393 => x"26",
         13394 => x"58",
         13395 => x"5b",
         13396 => x"52",
         13397 => x"d8",
         13398 => x"15",
         13399 => x"9c",
         13400 => x"26",
         13401 => x"55",
         13402 => x"08",
         13403 => x"dc",
         13404 => x"8c",
         13405 => x"81",
         13406 => x"ba",
         13407 => x"c5",
         13408 => x"59",
         13409 => x"bb",
         13410 => x"2e",
         13411 => x"c2",
         13412 => x"75",
         13413 => x"ba",
         13414 => x"3d",
         13415 => x"0b",
         13416 => x"0c",
         13417 => x"04",
         13418 => x"51",
         13419 => x"3f",
         13420 => x"08",
         13421 => x"73",
         13422 => x"73",
         13423 => x"56",
         13424 => x"7b",
         13425 => x"8e",
         13426 => x"56",
         13427 => x"2e",
         13428 => x"18",
         13429 => x"2e",
         13430 => x"73",
         13431 => x"7e",
         13432 => x"dd",
         13433 => x"8c",
         13434 => x"ba",
         13435 => x"a3",
         13436 => x"19",
         13437 => x"59",
         13438 => x"38",
         13439 => x"12",
         13440 => x"80",
         13441 => x"38",
         13442 => x"0c",
         13443 => x"0c",
         13444 => x"80",
         13445 => x"7b",
         13446 => x"9c",
         13447 => x"05",
         13448 => x"58",
         13449 => x"26",
         13450 => x"76",
         13451 => x"16",
         13452 => x"33",
         13453 => x"7c",
         13454 => x"75",
         13455 => x"39",
         13456 => x"97",
         13457 => x"80",
         13458 => x"39",
         13459 => x"c5",
         13460 => x"fe",
         13461 => x"1b",
         13462 => x"39",
         13463 => x"08",
         13464 => x"a3",
         13465 => x"3d",
         13466 => x"05",
         13467 => x"33",
         13468 => x"ff",
         13469 => x"08",
         13470 => x"40",
         13471 => x"85",
         13472 => x"70",
         13473 => x"33",
         13474 => x"56",
         13475 => x"2e",
         13476 => x"74",
         13477 => x"ba",
         13478 => x"38",
         13479 => x"33",
         13480 => x"24",
         13481 => x"75",
         13482 => x"d1",
         13483 => x"08",
         13484 => x"80",
         13485 => x"80",
         13486 => x"16",
         13487 => x"11",
         13488 => x"81",
         13489 => x"5b",
         13490 => x"79",
         13491 => x"a9",
         13492 => x"8c",
         13493 => x"06",
         13494 => x"5d",
         13495 => x"7b",
         13496 => x"75",
         13497 => x"06",
         13498 => x"7f",
         13499 => x"9f",
         13500 => x"53",
         13501 => x"51",
         13502 => x"3f",
         13503 => x"08",
         13504 => x"6d",
         13505 => x"2e",
         13506 => x"74",
         13507 => x"26",
         13508 => x"ff",
         13509 => x"55",
         13510 => x"38",
         13511 => x"88",
         13512 => x"7f",
         13513 => x"38",
         13514 => x"0a",
         13515 => x"38",
         13516 => x"06",
         13517 => x"e7",
         13518 => x"2a",
         13519 => x"89",
         13520 => x"2b",
         13521 => x"47",
         13522 => x"2e",
         13523 => x"65",
         13524 => x"25",
         13525 => x"5f",
         13526 => x"83",
         13527 => x"80",
         13528 => x"38",
         13529 => x"53",
         13530 => x"51",
         13531 => x"3f",
         13532 => x"ba",
         13533 => x"95",
         13534 => x"ff",
         13535 => x"83",
         13536 => x"71",
         13537 => x"59",
         13538 => x"77",
         13539 => x"2e",
         13540 => x"82",
         13541 => x"90",
         13542 => x"83",
         13543 => x"44",
         13544 => x"2e",
         13545 => x"83",
         13546 => x"11",
         13547 => x"33",
         13548 => x"71",
         13549 => x"81",
         13550 => x"72",
         13551 => x"75",
         13552 => x"83",
         13553 => x"11",
         13554 => x"33",
         13555 => x"71",
         13556 => x"81",
         13557 => x"72",
         13558 => x"75",
         13559 => x"5c",
         13560 => x"42",
         13561 => x"a3",
         13562 => x"4e",
         13563 => x"4f",
         13564 => x"78",
         13565 => x"80",
         13566 => x"82",
         13567 => x"57",
         13568 => x"26",
         13569 => x"61",
         13570 => x"81",
         13571 => x"63",
         13572 => x"f9",
         13573 => x"06",
         13574 => x"2e",
         13575 => x"81",
         13576 => x"83",
         13577 => x"6e",
         13578 => x"46",
         13579 => x"62",
         13580 => x"c2",
         13581 => x"38",
         13582 => x"57",
         13583 => x"e7",
         13584 => x"58",
         13585 => x"9d",
         13586 => x"26",
         13587 => x"e7",
         13588 => x"10",
         13589 => x"22",
         13590 => x"74",
         13591 => x"38",
         13592 => x"ee",
         13593 => x"78",
         13594 => x"ba",
         13595 => x"8c",
         13596 => x"05",
         13597 => x"8c",
         13598 => x"26",
         13599 => x"0b",
         13600 => x"08",
         13601 => x"8c",
         13602 => x"11",
         13603 => x"05",
         13604 => x"83",
         13605 => x"2a",
         13606 => x"a0",
         13607 => x"7d",
         13608 => x"66",
         13609 => x"70",
         13610 => x"31",
         13611 => x"44",
         13612 => x"89",
         13613 => x"1d",
         13614 => x"29",
         13615 => x"31",
         13616 => x"79",
         13617 => x"38",
         13618 => x"7d",
         13619 => x"70",
         13620 => x"56",
         13621 => x"3f",
         13622 => x"08",
         13623 => x"2e",
         13624 => x"62",
         13625 => x"81",
         13626 => x"38",
         13627 => x"0b",
         13628 => x"08",
         13629 => x"38",
         13630 => x"38",
         13631 => x"74",
         13632 => x"89",
         13633 => x"5b",
         13634 => x"8b",
         13635 => x"ba",
         13636 => x"3d",
         13637 => x"98",
         13638 => x"4e",
         13639 => x"93",
         13640 => x"8c",
         13641 => x"0d",
         13642 => x"0c",
         13643 => x"d0",
         13644 => x"ff",
         13645 => x"57",
         13646 => x"91",
         13647 => x"77",
         13648 => x"d0",
         13649 => x"77",
         13650 => x"b2",
         13651 => x"83",
         13652 => x"5c",
         13653 => x"57",
         13654 => x"81",
         13655 => x"76",
         13656 => x"58",
         13657 => x"12",
         13658 => x"62",
         13659 => x"38",
         13660 => x"81",
         13661 => x"44",
         13662 => x"45",
         13663 => x"89",
         13664 => x"70",
         13665 => x"59",
         13666 => x"70",
         13667 => x"47",
         13668 => x"09",
         13669 => x"38",
         13670 => x"38",
         13671 => x"70",
         13672 => x"07",
         13673 => x"07",
         13674 => x"7a",
         13675 => x"ce",
         13676 => x"84",
         13677 => x"83",
         13678 => x"98",
         13679 => x"f9",
         13680 => x"3d",
         13681 => x"81",
         13682 => x"fe",
         13683 => x"81",
         13684 => x"8c",
         13685 => x"38",
         13686 => x"77",
         13687 => x"8c",
         13688 => x"75",
         13689 => x"5f",
         13690 => x"57",
         13691 => x"fe",
         13692 => x"7f",
         13693 => x"fb",
         13694 => x"fa",
         13695 => x"83",
         13696 => x"38",
         13697 => x"3d",
         13698 => x"95",
         13699 => x"06",
         13700 => x"67",
         13701 => x"f5",
         13702 => x"70",
         13703 => x"43",
         13704 => x"84",
         13705 => x"9f",
         13706 => x"38",
         13707 => x"77",
         13708 => x"80",
         13709 => x"f5",
         13710 => x"76",
         13711 => x"0c",
         13712 => x"84",
         13713 => x"04",
         13714 => x"81",
         13715 => x"38",
         13716 => x"27",
         13717 => x"81",
         13718 => x"57",
         13719 => x"38",
         13720 => x"57",
         13721 => x"70",
         13722 => x"34",
         13723 => x"74",
         13724 => x"61",
         13725 => x"59",
         13726 => x"70",
         13727 => x"33",
         13728 => x"05",
         13729 => x"15",
         13730 => x"38",
         13731 => x"45",
         13732 => x"82",
         13733 => x"34",
         13734 => x"05",
         13735 => x"ff",
         13736 => x"6a",
         13737 => x"34",
         13738 => x"5c",
         13739 => x"05",
         13740 => x"90",
         13741 => x"83",
         13742 => x"5a",
         13743 => x"91",
         13744 => x"9e",
         13745 => x"49",
         13746 => x"05",
         13747 => x"75",
         13748 => x"26",
         13749 => x"75",
         13750 => x"06",
         13751 => x"93",
         13752 => x"88",
         13753 => x"61",
         13754 => x"f8",
         13755 => x"34",
         13756 => x"05",
         13757 => x"99",
         13758 => x"61",
         13759 => x"80",
         13760 => x"34",
         13761 => x"05",
         13762 => x"2a",
         13763 => x"9d",
         13764 => x"90",
         13765 => x"61",
         13766 => x"7e",
         13767 => x"ba",
         13768 => x"ba",
         13769 => x"9f",
         13770 => x"83",
         13771 => x"38",
         13772 => x"05",
         13773 => x"a8",
         13774 => x"61",
         13775 => x"80",
         13776 => x"05",
         13777 => x"ff",
         13778 => x"74",
         13779 => x"34",
         13780 => x"4b",
         13781 => x"05",
         13782 => x"61",
         13783 => x"a9",
         13784 => x"34",
         13785 => x"05",
         13786 => x"59",
         13787 => x"70",
         13788 => x"33",
         13789 => x"05",
         13790 => x"15",
         13791 => x"38",
         13792 => x"05",
         13793 => x"69",
         13794 => x"ff",
         13795 => x"aa",
         13796 => x"54",
         13797 => x"52",
         13798 => x"c6",
         13799 => x"57",
         13800 => x"08",
         13801 => x"60",
         13802 => x"83",
         13803 => x"38",
         13804 => x"55",
         13805 => x"81",
         13806 => x"ff",
         13807 => x"f4",
         13808 => x"41",
         13809 => x"2e",
         13810 => x"87",
         13811 => x"57",
         13812 => x"83",
         13813 => x"76",
         13814 => x"88",
         13815 => x"55",
         13816 => x"81",
         13817 => x"76",
         13818 => x"78",
         13819 => x"05",
         13820 => x"98",
         13821 => x"64",
         13822 => x"65",
         13823 => x"26",
         13824 => x"59",
         13825 => x"53",
         13826 => x"51",
         13827 => x"3f",
         13828 => x"08",
         13829 => x"84",
         13830 => x"55",
         13831 => x"81",
         13832 => x"ff",
         13833 => x"f4",
         13834 => x"77",
         13835 => x"5b",
         13836 => x"7f",
         13837 => x"7f",
         13838 => x"89",
         13839 => x"62",
         13840 => x"38",
         13841 => x"55",
         13842 => x"83",
         13843 => x"74",
         13844 => x"60",
         13845 => x"fe",
         13846 => x"84",
         13847 => x"85",
         13848 => x"1b",
         13849 => x"57",
         13850 => x"38",
         13851 => x"83",
         13852 => x"86",
         13853 => x"ff",
         13854 => x"38",
         13855 => x"82",
         13856 => x"81",
         13857 => x"c1",
         13858 => x"2a",
         13859 => x"7d",
         13860 => x"84",
         13861 => x"59",
         13862 => x"81",
         13863 => x"ff",
         13864 => x"f4",
         13865 => x"69",
         13866 => x"6b",
         13867 => x"be",
         13868 => x"67",
         13869 => x"81",
         13870 => x"67",
         13871 => x"78",
         13872 => x"34",
         13873 => x"05",
         13874 => x"80",
         13875 => x"62",
         13876 => x"f7",
         13877 => x"67",
         13878 => x"84",
         13879 => x"82",
         13880 => x"57",
         13881 => x"05",
         13882 => x"8c",
         13883 => x"05",
         13884 => x"83",
         13885 => x"67",
         13886 => x"05",
         13887 => x"83",
         13888 => x"84",
         13889 => x"61",
         13890 => x"34",
         13891 => x"ca",
         13892 => x"88",
         13893 => x"61",
         13894 => x"34",
         13895 => x"58",
         13896 => x"cc",
         13897 => x"98",
         13898 => x"61",
         13899 => x"34",
         13900 => x"53",
         13901 => x"51",
         13902 => x"3f",
         13903 => x"ba",
         13904 => x"c9",
         13905 => x"80",
         13906 => x"fe",
         13907 => x"81",
         13908 => x"8c",
         13909 => x"38",
         13910 => x"08",
         13911 => x"0c",
         13912 => x"84",
         13913 => x"04",
         13914 => x"e4",
         13915 => x"64",
         13916 => x"f6",
         13917 => x"ae",
         13918 => x"2a",
         13919 => x"83",
         13920 => x"56",
         13921 => x"2e",
         13922 => x"77",
         13923 => x"83",
         13924 => x"77",
         13925 => x"70",
         13926 => x"58",
         13927 => x"86",
         13928 => x"27",
         13929 => x"52",
         13930 => x"f5",
         13931 => x"ba",
         13932 => x"10",
         13933 => x"70",
         13934 => x"5c",
         13935 => x"0b",
         13936 => x"08",
         13937 => x"05",
         13938 => x"ff",
         13939 => x"27",
         13940 => x"8e",
         13941 => x"39",
         13942 => x"08",
         13943 => x"26",
         13944 => x"7a",
         13945 => x"77",
         13946 => x"7a",
         13947 => x"8e",
         13948 => x"39",
         13949 => x"44",
         13950 => x"f8",
         13951 => x"43",
         13952 => x"75",
         13953 => x"34",
         13954 => x"49",
         13955 => x"05",
         13956 => x"2a",
         13957 => x"a2",
         13958 => x"98",
         13959 => x"61",
         13960 => x"f9",
         13961 => x"61",
         13962 => x"34",
         13963 => x"c4",
         13964 => x"61",
         13965 => x"34",
         13966 => x"80",
         13967 => x"7c",
         13968 => x"34",
         13969 => x"5c",
         13970 => x"05",
         13971 => x"2a",
         13972 => x"a6",
         13973 => x"98",
         13974 => x"61",
         13975 => x"82",
         13976 => x"34",
         13977 => x"05",
         13978 => x"ae",
         13979 => x"61",
         13980 => x"81",
         13981 => x"34",
         13982 => x"05",
         13983 => x"b2",
         13984 => x"61",
         13985 => x"ff",
         13986 => x"c0",
         13987 => x"61",
         13988 => x"34",
         13989 => x"c7",
         13990 => x"e8",
         13991 => x"76",
         13992 => x"58",
         13993 => x"81",
         13994 => x"ff",
         13995 => x"80",
         13996 => x"38",
         13997 => x"05",
         13998 => x"70",
         13999 => x"34",
         14000 => x"74",
         14001 => x"b8",
         14002 => x"80",
         14003 => x"79",
         14004 => x"d9",
         14005 => x"84",
         14006 => x"f4",
         14007 => x"90",
         14008 => x"42",
         14009 => x"b2",
         14010 => x"54",
         14011 => x"08",
         14012 => x"79",
         14013 => x"b4",
         14014 => x"39",
         14015 => x"ba",
         14016 => x"3d",
         14017 => x"98",
         14018 => x"61",
         14019 => x"ff",
         14020 => x"05",
         14021 => x"6a",
         14022 => x"4c",
         14023 => x"34",
         14024 => x"05",
         14025 => x"85",
         14026 => x"61",
         14027 => x"ff",
         14028 => x"34",
         14029 => x"05",
         14030 => x"89",
         14031 => x"61",
         14032 => x"8f",
         14033 => x"57",
         14034 => x"76",
         14035 => x"53",
         14036 => x"51",
         14037 => x"3f",
         14038 => x"56",
         14039 => x"70",
         14040 => x"34",
         14041 => x"76",
         14042 => x"5c",
         14043 => x"70",
         14044 => x"34",
         14045 => x"d2",
         14046 => x"05",
         14047 => x"e1",
         14048 => x"05",
         14049 => x"c1",
         14050 => x"f2",
         14051 => x"05",
         14052 => x"61",
         14053 => x"34",
         14054 => x"83",
         14055 => x"80",
         14056 => x"e7",
         14057 => x"ff",
         14058 => x"61",
         14059 => x"34",
         14060 => x"59",
         14061 => x"e9",
         14062 => x"90",
         14063 => x"61",
         14064 => x"34",
         14065 => x"40",
         14066 => x"eb",
         14067 => x"61",
         14068 => x"34",
         14069 => x"ed",
         14070 => x"61",
         14071 => x"34",
         14072 => x"ef",
         14073 => x"d5",
         14074 => x"aa",
         14075 => x"54",
         14076 => x"60",
         14077 => x"fe",
         14078 => x"81",
         14079 => x"53",
         14080 => x"51",
         14081 => x"3f",
         14082 => x"55",
         14083 => x"f4",
         14084 => x"61",
         14085 => x"7b",
         14086 => x"5a",
         14087 => x"78",
         14088 => x"8d",
         14089 => x"3d",
         14090 => x"81",
         14091 => x"79",
         14092 => x"b4",
         14093 => x"2e",
         14094 => x"9e",
         14095 => x"33",
         14096 => x"2e",
         14097 => x"76",
         14098 => x"58",
         14099 => x"57",
         14100 => x"86",
         14101 => x"24",
         14102 => x"76",
         14103 => x"76",
         14104 => x"55",
         14105 => x"8c",
         14106 => x"0d",
         14107 => x"0d",
         14108 => x"05",
         14109 => x"59",
         14110 => x"2e",
         14111 => x"84",
         14112 => x"80",
         14113 => x"38",
         14114 => x"77",
         14115 => x"56",
         14116 => x"34",
         14117 => x"74",
         14118 => x"38",
         14119 => x"0c",
         14120 => x"18",
         14121 => x"0d",
         14122 => x"fc",
         14123 => x"53",
         14124 => x"76",
         14125 => x"9e",
         14126 => x"7a",
         14127 => x"70",
         14128 => x"2a",
         14129 => x"1b",
         14130 => x"88",
         14131 => x"56",
         14132 => x"8d",
         14133 => x"ff",
         14134 => x"a3",
         14135 => x"0d",
         14136 => x"05",
         14137 => x"58",
         14138 => x"77",
         14139 => x"76",
         14140 => x"58",
         14141 => x"55",
         14142 => x"a1",
         14143 => x"0c",
         14144 => x"80",
         14145 => x"56",
         14146 => x"80",
         14147 => x"77",
         14148 => x"56",
         14149 => x"34",
         14150 => x"74",
         14151 => x"38",
         14152 => x"0c",
         14153 => x"18",
         14154 => x"80",
         14155 => x"38",
         14156 => x"ac",
         14157 => x"54",
         14158 => x"76",
         14159 => x"9d",
         14160 => x"ba",
         14161 => x"38",
         14162 => x"ba",
         14163 => x"84",
         14164 => x"9f",
         14165 => x"9f",
         14166 => x"11",
         14167 => x"c0",
         14168 => x"08",
         14169 => x"a2",
         14170 => x"32",
         14171 => x"72",
         14172 => x"70",
         14173 => x"56",
         14174 => x"39",
         14175 => x"51",
         14176 => x"ff",
         14177 => x"84",
         14178 => x"9f",
         14179 => x"fd",
         14180 => x"02",
         14181 => x"05",
         14182 => x"80",
         14183 => x"ff",
         14184 => x"72",
         14185 => x"06",
         14186 => x"ba",
         14187 => x"3d",
         14188 => x"ff",
         14189 => x"54",
         14190 => x"2e",
         14191 => x"e9",
         14192 => x"2e",
         14193 => x"e7",
         14194 => x"72",
         14195 => x"38",
         14196 => x"83",
         14197 => x"53",
         14198 => x"ff",
         14199 => x"71",
         14200 => x"d0",
         14201 => x"51",
         14202 => x"81",
         14203 => x"81",
         14204 => x"ba",
         14205 => x"85",
         14206 => x"fe",
         14207 => x"92",
         14208 => x"84",
         14209 => x"22",
         14210 => x"53",
         14211 => x"26",
         14212 => x"53",
         14213 => x"8c",
         14214 => x"0d",
         14215 => x"b5",
         14216 => x"06",
         14217 => x"81",
         14218 => x"38",
         14219 => x"e5",
         14220 => x"22",
         14221 => x"0c",
         14222 => x"0d",
         14223 => x"0d",
         14224 => x"83",
         14225 => x"80",
         14226 => x"83",
         14227 => x"83",
         14228 => x"56",
         14229 => x"26",
         14230 => x"74",
         14231 => x"56",
         14232 => x"30",
         14233 => x"73",
         14234 => x"54",
         14235 => x"70",
         14236 => x"70",
         14237 => x"22",
         14238 => x"2a",
         14239 => x"ff",
         14240 => x"52",
         14241 => x"24",
         14242 => x"cf",
         14243 => x"15",
         14244 => x"05",
         14245 => x"73",
         14246 => x"25",
         14247 => x"07",
         14248 => x"70",
         14249 => x"38",
         14250 => x"84",
         14251 => x"87",
         14252 => x"83",
         14253 => x"ff",
         14254 => x"88",
         14255 => x"71",
         14256 => x"ca",
         14257 => x"73",
         14258 => x"a0",
         14259 => x"ff",
         14260 => x"51",
         14261 => x"39",
         14262 => x"70",
         14263 => x"06",
         14264 => x"39",
         14265 => x"83",
         14266 => x"57",
         14267 => x"e6",
         14268 => x"ff",
         14269 => x"51",
         14270 => x"16",
         14271 => x"ff",
         14272 => x"d0",
         14273 => x"70",
         14274 => x"06",
         14275 => x"39",
         14276 => x"83",
         14277 => x"57",
         14278 => x"39",
         14279 => x"81",
         14280 => x"31",
         14281 => x"ff",
         14282 => x"55",
         14283 => x"75",
         14284 => x"75",
         14285 => x"52",
         14286 => x"39",
         14287 => x"ff",
         14288 => x"ff",
         14289 => x"00",
         14290 => x"ff",
         14291 => x"19",
         14292 => x"19",
         14293 => x"19",
         14294 => x"19",
         14295 => x"19",
         14296 => x"19",
         14297 => x"19",
         14298 => x"19",
         14299 => x"19",
         14300 => x"19",
         14301 => x"19",
         14302 => x"19",
         14303 => x"19",
         14304 => x"18",
         14305 => x"18",
         14306 => x"18",
         14307 => x"18",
         14308 => x"18",
         14309 => x"18",
         14310 => x"18",
         14311 => x"1e",
         14312 => x"1f",
         14313 => x"1f",
         14314 => x"1f",
         14315 => x"1f",
         14316 => x"1f",
         14317 => x"1f",
         14318 => x"1f",
         14319 => x"1f",
         14320 => x"1f",
         14321 => x"1f",
         14322 => x"1f",
         14323 => x"1f",
         14324 => x"1f",
         14325 => x"1f",
         14326 => x"1f",
         14327 => x"1f",
         14328 => x"1f",
         14329 => x"1f",
         14330 => x"1f",
         14331 => x"1f",
         14332 => x"1f",
         14333 => x"1f",
         14334 => x"1f",
         14335 => x"1f",
         14336 => x"1f",
         14337 => x"1f",
         14338 => x"1f",
         14339 => x"1f",
         14340 => x"1f",
         14341 => x"1f",
         14342 => x"1f",
         14343 => x"1f",
         14344 => x"1f",
         14345 => x"1f",
         14346 => x"1f",
         14347 => x"1f",
         14348 => x"1f",
         14349 => x"1f",
         14350 => x"1f",
         14351 => x"1f",
         14352 => x"1f",
         14353 => x"1f",
         14354 => x"24",
         14355 => x"1f",
         14356 => x"1f",
         14357 => x"1f",
         14358 => x"1f",
         14359 => x"1f",
         14360 => x"1f",
         14361 => x"1f",
         14362 => x"1f",
         14363 => x"1f",
         14364 => x"1f",
         14365 => x"1f",
         14366 => x"1f",
         14367 => x"1f",
         14368 => x"1f",
         14369 => x"1f",
         14370 => x"1f",
         14371 => x"24",
         14372 => x"23",
         14373 => x"1f",
         14374 => x"22",
         14375 => x"24",
         14376 => x"23",
         14377 => x"22",
         14378 => x"21",
         14379 => x"1f",
         14380 => x"1f",
         14381 => x"1f",
         14382 => x"1f",
         14383 => x"1f",
         14384 => x"1f",
         14385 => x"1f",
         14386 => x"1f",
         14387 => x"1f",
         14388 => x"1f",
         14389 => x"1f",
         14390 => x"1f",
         14391 => x"1f",
         14392 => x"1f",
         14393 => x"1f",
         14394 => x"1f",
         14395 => x"1f",
         14396 => x"1f",
         14397 => x"1f",
         14398 => x"1f",
         14399 => x"1f",
         14400 => x"1f",
         14401 => x"1f",
         14402 => x"1f",
         14403 => x"1f",
         14404 => x"1f",
         14405 => x"1f",
         14406 => x"1f",
         14407 => x"1f",
         14408 => x"1f",
         14409 => x"1f",
         14410 => x"1f",
         14411 => x"1f",
         14412 => x"1f",
         14413 => x"1f",
         14414 => x"1f",
         14415 => x"1f",
         14416 => x"1f",
         14417 => x"1f",
         14418 => x"1f",
         14419 => x"1f",
         14420 => x"1f",
         14421 => x"1f",
         14422 => x"1f",
         14423 => x"1f",
         14424 => x"1f",
         14425 => x"1f",
         14426 => x"1f",
         14427 => x"1f",
         14428 => x"1f",
         14429 => x"1f",
         14430 => x"1f",
         14431 => x"21",
         14432 => x"21",
         14433 => x"1f",
         14434 => x"1f",
         14435 => x"1f",
         14436 => x"1f",
         14437 => x"1f",
         14438 => x"1f",
         14439 => x"1f",
         14440 => x"1f",
         14441 => x"21",
         14442 => x"21",
         14443 => x"1f",
         14444 => x"21",
         14445 => x"1f",
         14446 => x"21",
         14447 => x"21",
         14448 => x"21",
         14449 => x"32",
         14450 => x"32",
         14451 => x"32",
         14452 => x"32",
         14453 => x"32",
         14454 => x"32",
         14455 => x"3b",
         14456 => x"3a",
         14457 => x"38",
         14458 => x"36",
         14459 => x"3a",
         14460 => x"34",
         14461 => x"37",
         14462 => x"36",
         14463 => x"39",
         14464 => x"36",
         14465 => x"37",
         14466 => x"39",
         14467 => x"34",
         14468 => x"38",
         14469 => x"38",
         14470 => x"37",
         14471 => x"34",
         14472 => x"34",
         14473 => x"37",
         14474 => x"36",
         14475 => x"36",
         14476 => x"36",
         14477 => x"46",
         14478 => x"46",
         14479 => x"46",
         14480 => x"46",
         14481 => x"46",
         14482 => x"46",
         14483 => x"46",
         14484 => x"47",
         14485 => x"47",
         14486 => x"47",
         14487 => x"47",
         14488 => x"47",
         14489 => x"47",
         14490 => x"47",
         14491 => x"47",
         14492 => x"47",
         14493 => x"47",
         14494 => x"47",
         14495 => x"47",
         14496 => x"47",
         14497 => x"47",
         14498 => x"47",
         14499 => x"47",
         14500 => x"47",
         14501 => x"47",
         14502 => x"47",
         14503 => x"47",
         14504 => x"47",
         14505 => x"47",
         14506 => x"47",
         14507 => x"47",
         14508 => x"47",
         14509 => x"47",
         14510 => x"47",
         14511 => x"47",
         14512 => x"47",
         14513 => x"47",
         14514 => x"48",
         14515 => x"48",
         14516 => x"48",
         14517 => x"48",
         14518 => x"47",
         14519 => x"48",
         14520 => x"48",
         14521 => x"47",
         14522 => x"47",
         14523 => x"47",
         14524 => x"48",
         14525 => x"48",
         14526 => x"47",
         14527 => x"47",
         14528 => x"47",
         14529 => x"47",
         14530 => x"47",
         14531 => x"47",
         14532 => x"47",
         14533 => x"47",
         14534 => x"54",
         14535 => x"55",
         14536 => x"55",
         14537 => x"54",
         14538 => x"54",
         14539 => x"54",
         14540 => x"54",
         14541 => x"55",
         14542 => x"52",
         14543 => x"55",
         14544 => x"57",
         14545 => x"52",
         14546 => x"52",
         14547 => x"52",
         14548 => x"52",
         14549 => x"52",
         14550 => x"52",
         14551 => x"55",
         14552 => x"57",
         14553 => x"56",
         14554 => x"52",
         14555 => x"52",
         14556 => x"52",
         14557 => x"52",
         14558 => x"52",
         14559 => x"52",
         14560 => x"52",
         14561 => x"52",
         14562 => x"52",
         14563 => x"52",
         14564 => x"52",
         14565 => x"52",
         14566 => x"52",
         14567 => x"52",
         14568 => x"52",
         14569 => x"52",
         14570 => x"52",
         14571 => x"52",
         14572 => x"52",
         14573 => x"55",
         14574 => x"52",
         14575 => x"52",
         14576 => x"52",
         14577 => x"54",
         14578 => x"53",
         14579 => x"53",
         14580 => x"52",
         14581 => x"52",
         14582 => x"52",
         14583 => x"52",
         14584 => x"53",
         14585 => x"52",
         14586 => x"53",
         14587 => x"59",
         14588 => x"59",
         14589 => x"59",
         14590 => x"59",
         14591 => x"59",
         14592 => x"59",
         14593 => x"59",
         14594 => x"58",
         14595 => x"59",
         14596 => x"59",
         14597 => x"59",
         14598 => x"59",
         14599 => x"59",
         14600 => x"59",
         14601 => x"59",
         14602 => x"59",
         14603 => x"59",
         14604 => x"59",
         14605 => x"59",
         14606 => x"59",
         14607 => x"59",
         14608 => x"59",
         14609 => x"59",
         14610 => x"59",
         14611 => x"59",
         14612 => x"59",
         14613 => x"59",
         14614 => x"59",
         14615 => x"59",
         14616 => x"59",
         14617 => x"59",
         14618 => x"5a",
         14619 => x"59",
         14620 => x"59",
         14621 => x"59",
         14622 => x"5a",
         14623 => x"5a",
         14624 => x"5a",
         14625 => x"59",
         14626 => x"5a",
         14627 => x"5a",
         14628 => x"5a",
         14629 => x"5a",
         14630 => x"5a",
         14631 => x"59",
         14632 => x"59",
         14633 => x"59",
         14634 => x"59",
         14635 => x"59",
         14636 => x"59",
         14637 => x"63",
         14638 => x"61",
         14639 => x"61",
         14640 => x"61",
         14641 => x"61",
         14642 => x"61",
         14643 => x"61",
         14644 => x"61",
         14645 => x"61",
         14646 => x"61",
         14647 => x"61",
         14648 => x"61",
         14649 => x"61",
         14650 => x"61",
         14651 => x"5e",
         14652 => x"61",
         14653 => x"61",
         14654 => x"61",
         14655 => x"61",
         14656 => x"61",
         14657 => x"61",
         14658 => x"63",
         14659 => x"61",
         14660 => x"61",
         14661 => x"63",
         14662 => x"61",
         14663 => x"63",
         14664 => x"5e",
         14665 => x"63",
         14666 => x"df",
         14667 => x"df",
         14668 => x"df",
         14669 => x"df",
         14670 => x"de",
         14671 => x"de",
         14672 => x"de",
         14673 => x"de",
         14674 => x"de",
         14675 => x"0e",
         14676 => x"0b",
         14677 => x"0b",
         14678 => x"0f",
         14679 => x"0b",
         14680 => x"0b",
         14681 => x"0b",
         14682 => x"0b",
         14683 => x"0b",
         14684 => x"0b",
         14685 => x"0b",
         14686 => x"0d",
         14687 => x"0b",
         14688 => x"0f",
         14689 => x"0f",
         14690 => x"0b",
         14691 => x"0b",
         14692 => x"0b",
         14693 => x"0b",
         14694 => x"0b",
         14695 => x"0b",
         14696 => x"0b",
         14697 => x"0b",
         14698 => x"0b",
         14699 => x"0b",
         14700 => x"0b",
         14701 => x"0b",
         14702 => x"0b",
         14703 => x"0b",
         14704 => x"0b",
         14705 => x"0b",
         14706 => x"0b",
         14707 => x"0b",
         14708 => x"0b",
         14709 => x"0b",
         14710 => x"0b",
         14711 => x"0b",
         14712 => x"0b",
         14713 => x"0b",
         14714 => x"0b",
         14715 => x"0b",
         14716 => x"0b",
         14717 => x"0b",
         14718 => x"0b",
         14719 => x"0b",
         14720 => x"0b",
         14721 => x"0b",
         14722 => x"0b",
         14723 => x"0b",
         14724 => x"0b",
         14725 => x"0b",
         14726 => x"0f",
         14727 => x"0b",
         14728 => x"0b",
         14729 => x"0b",
         14730 => x"0b",
         14731 => x"0e",
         14732 => x"0b",
         14733 => x"0b",
         14734 => x"0b",
         14735 => x"0b",
         14736 => x"0b",
         14737 => x"0b",
         14738 => x"0b",
         14739 => x"0b",
         14740 => x"0b",
         14741 => x"0b",
         14742 => x"0e",
         14743 => x"0e",
         14744 => x"0e",
         14745 => x"0e",
         14746 => x"0e",
         14747 => x"0b",
         14748 => x"0e",
         14749 => x"0b",
         14750 => x"0b",
         14751 => x"0e",
         14752 => x"0b",
         14753 => x"0b",
         14754 => x"0c",
         14755 => x"0e",
         14756 => x"0b",
         14757 => x"0b",
         14758 => x"0f",
         14759 => x"0b",
         14760 => x"0c",
         14761 => x"0b",
         14762 => x"0b",
         14763 => x"0e",
         14764 => x"6e",
         14765 => x"00",
         14766 => x"6f",
         14767 => x"00",
         14768 => x"6e",
         14769 => x"00",
         14770 => x"6f",
         14771 => x"00",
         14772 => x"78",
         14773 => x"00",
         14774 => x"6c",
         14775 => x"00",
         14776 => x"6f",
         14777 => x"00",
         14778 => x"69",
         14779 => x"00",
         14780 => x"75",
         14781 => x"00",
         14782 => x"62",
         14783 => x"68",
         14784 => x"77",
         14785 => x"64",
         14786 => x"65",
         14787 => x"64",
         14788 => x"65",
         14789 => x"6c",
         14790 => x"00",
         14791 => x"70",
         14792 => x"73",
         14793 => x"74",
         14794 => x"73",
         14795 => x"00",
         14796 => x"66",
         14797 => x"00",
         14798 => x"73",
         14799 => x"00",
         14800 => x"73",
         14801 => x"30",
         14802 => x"61",
         14803 => x"00",
         14804 => x"61",
         14805 => x"00",
         14806 => x"6c",
         14807 => x"00",
         14808 => x"00",
         14809 => x"6b",
         14810 => x"6e",
         14811 => x"72",
         14812 => x"00",
         14813 => x"72",
         14814 => x"74",
         14815 => x"20",
         14816 => x"6f",
         14817 => x"63",
         14818 => x"00",
         14819 => x"6f",
         14820 => x"6e",
         14821 => x"70",
         14822 => x"66",
         14823 => x"73",
         14824 => x"00",
         14825 => x"73",
         14826 => x"69",
         14827 => x"6e",
         14828 => x"65",
         14829 => x"79",
         14830 => x"00",
         14831 => x"6c",
         14832 => x"73",
         14833 => x"63",
         14834 => x"2e",
         14835 => x"6d",
         14836 => x"74",
         14837 => x"70",
         14838 => x"74",
         14839 => x"20",
         14840 => x"63",
         14841 => x"65",
         14842 => x"00",
         14843 => x"72",
         14844 => x"20",
         14845 => x"72",
         14846 => x"2e",
         14847 => x"20",
         14848 => x"70",
         14849 => x"62",
         14850 => x"66",
         14851 => x"73",
         14852 => x"65",
         14853 => x"6f",
         14854 => x"20",
         14855 => x"64",
         14856 => x"2e",
         14857 => x"73",
         14858 => x"6f",
         14859 => x"6e",
         14860 => x"65",
         14861 => x"00",
         14862 => x"69",
         14863 => x"6e",
         14864 => x"65",
         14865 => x"73",
         14866 => x"76",
         14867 => x"64",
         14868 => x"00",
         14869 => x"20",
         14870 => x"77",
         14871 => x"65",
         14872 => x"6f",
         14873 => x"74",
         14874 => x"00",
         14875 => x"6c",
         14876 => x"61",
         14877 => x"65",
         14878 => x"76",
         14879 => x"64",
         14880 => x"00",
         14881 => x"6c",
         14882 => x"6c",
         14883 => x"64",
         14884 => x"78",
         14885 => x"73",
         14886 => x"00",
         14887 => x"63",
         14888 => x"20",
         14889 => x"69",
         14890 => x"00",
         14891 => x"76",
         14892 => x"64",
         14893 => x"6c",
         14894 => x"6d",
         14895 => x"00",
         14896 => x"20",
         14897 => x"68",
         14898 => x"75",
         14899 => x"00",
         14900 => x"20",
         14901 => x"65",
         14902 => x"75",
         14903 => x"00",
         14904 => x"73",
         14905 => x"6f",
         14906 => x"65",
         14907 => x"2e",
         14908 => x"74",
         14909 => x"61",
         14910 => x"72",
         14911 => x"2e",
         14912 => x"73",
         14913 => x"72",
         14914 => x"00",
         14915 => x"63",
         14916 => x"73",
         14917 => x"00",
         14918 => x"6c",
         14919 => x"79",
         14920 => x"20",
         14921 => x"61",
         14922 => x"6c",
         14923 => x"79",
         14924 => x"2f",
         14925 => x"2e",
         14926 => x"00",
         14927 => x"61",
         14928 => x"00",
         14929 => x"38",
         14930 => x"00",
         14931 => x"20",
         14932 => x"32",
         14933 => x"00",
         14934 => x"00",
         14935 => x"00",
         14936 => x"00",
         14937 => x"34",
         14938 => x"00",
         14939 => x"20",
         14940 => x"20",
         14941 => x"00",
         14942 => x"53",
         14943 => x"20",
         14944 => x"28",
         14945 => x"2f",
         14946 => x"32",
         14947 => x"00",
         14948 => x"2e",
         14949 => x"00",
         14950 => x"50",
         14951 => x"72",
         14952 => x"25",
         14953 => x"29",
         14954 => x"20",
         14955 => x"2a",
         14956 => x"00",
         14957 => x"55",
         14958 => x"74",
         14959 => x"75",
         14960 => x"48",
         14961 => x"6c",
         14962 => x"00",
         14963 => x"52",
         14964 => x"54",
         14965 => x"6e",
         14966 => x"72",
         14967 => x"00",
         14968 => x"52",
         14969 => x"52",
         14970 => x"6e",
         14971 => x"72",
         14972 => x"00",
         14973 => x"52",
         14974 => x"54",
         14975 => x"6e",
         14976 => x"72",
         14977 => x"00",
         14978 => x"52",
         14979 => x"52",
         14980 => x"6e",
         14981 => x"72",
         14982 => x"00",
         14983 => x"43",
         14984 => x"57",
         14985 => x"6e",
         14986 => x"72",
         14987 => x"00",
         14988 => x"43",
         14989 => x"52",
         14990 => x"6e",
         14991 => x"72",
         14992 => x"00",
         14993 => x"32",
         14994 => x"74",
         14995 => x"75",
         14996 => x"00",
         14997 => x"6d",
         14998 => x"69",
         14999 => x"72",
         15000 => x"74",
         15001 => x"74",
         15002 => x"67",
         15003 => x"20",
         15004 => x"65",
         15005 => x"2e",
         15006 => x"61",
         15007 => x"6e",
         15008 => x"69",
         15009 => x"2e",
         15010 => x"00",
         15011 => x"74",
         15012 => x"65",
         15013 => x"61",
         15014 => x"00",
         15015 => x"53",
         15016 => x"75",
         15017 => x"74",
         15018 => x"69",
         15019 => x"20",
         15020 => x"69",
         15021 => x"69",
         15022 => x"73",
         15023 => x"64",
         15024 => x"72",
         15025 => x"2c",
         15026 => x"65",
         15027 => x"20",
         15028 => x"74",
         15029 => x"6e",
         15030 => x"6c",
         15031 => x"00",
         15032 => x"00",
         15033 => x"3a",
         15034 => x"00",
         15035 => x"73",
         15036 => x"6e",
         15037 => x"61",
         15038 => x"65",
         15039 => x"00",
         15040 => x"00",
         15041 => x"64",
         15042 => x"6d",
         15043 => x"64",
         15044 => x"00",
         15045 => x"55",
         15046 => x"6e",
         15047 => x"3a",
         15048 => x"5c",
         15049 => x"25",
         15050 => x"00",
         15051 => x"6c",
         15052 => x"65",
         15053 => x"74",
         15054 => x"2e",
         15055 => x"00",
         15056 => x"73",
         15057 => x"74",
         15058 => x"20",
         15059 => x"6c",
         15060 => x"74",
         15061 => x"2e",
         15062 => x"00",
         15063 => x"6c",
         15064 => x"67",
         15065 => x"64",
         15066 => x"20",
         15067 => x"6c",
         15068 => x"2e",
         15069 => x"00",
         15070 => x"6c",
         15071 => x"65",
         15072 => x"6e",
         15073 => x"63",
         15074 => x"20",
         15075 => x"29",
         15076 => x"00",
         15077 => x"65",
         15078 => x"69",
         15079 => x"63",
         15080 => x"20",
         15081 => x"30",
         15082 => x"20",
         15083 => x"0a",
         15084 => x"38",
         15085 => x"25",
         15086 => x"58",
         15087 => x"00",
         15088 => x"38",
         15089 => x"25",
         15090 => x"2d",
         15091 => x"6d",
         15092 => x"69",
         15093 => x"2e",
         15094 => x"00",
         15095 => x"38",
         15096 => x"25",
         15097 => x"29",
         15098 => x"30",
         15099 => x"28",
         15100 => x"78",
         15101 => x"00",
         15102 => x"70",
         15103 => x"67",
         15104 => x"00",
         15105 => x"38",
         15106 => x"25",
         15107 => x"2d",
         15108 => x"65",
         15109 => x"6e",
         15110 => x"2e",
         15111 => x"00",
         15112 => x"6d",
         15113 => x"65",
         15114 => x"79",
         15115 => x"6f",
         15116 => x"65",
         15117 => x"00",
         15118 => x"3a",
         15119 => x"5c",
         15120 => x"00",
         15121 => x"6d",
         15122 => x"20",
         15123 => x"61",
         15124 => x"65",
         15125 => x"63",
         15126 => x"6f",
         15127 => x"72",
         15128 => x"73",
         15129 => x"6f",
         15130 => x"6e",
         15131 => x"00",
         15132 => x"3f",
         15133 => x"2f",
         15134 => x"25",
         15135 => x"64",
         15136 => x"3a",
         15137 => x"25",
         15138 => x"0a",
         15139 => x"43",
         15140 => x"6e",
         15141 => x"75",
         15142 => x"69",
         15143 => x"00",
         15144 => x"44",
         15145 => x"63",
         15146 => x"69",
         15147 => x"65",
         15148 => x"74",
         15149 => x"00",
         15150 => x"64",
         15151 => x"73",
         15152 => x"00",
         15153 => x"20",
         15154 => x"55",
         15155 => x"73",
         15156 => x"56",
         15157 => x"6f",
         15158 => x"64",
         15159 => x"73",
         15160 => x"20",
         15161 => x"58",
         15162 => x"00",
         15163 => x"20",
         15164 => x"55",
         15165 => x"6d",
         15166 => x"20",
         15167 => x"72",
         15168 => x"64",
         15169 => x"73",
         15170 => x"20",
         15171 => x"58",
         15172 => x"00",
         15173 => x"20",
         15174 => x"61",
         15175 => x"53",
         15176 => x"74",
         15177 => x"64",
         15178 => x"73",
         15179 => x"20",
         15180 => x"20",
         15181 => x"58",
         15182 => x"00",
         15183 => x"73",
         15184 => x"00",
         15185 => x"20",
         15186 => x"55",
         15187 => x"20",
         15188 => x"20",
         15189 => x"20",
         15190 => x"20",
         15191 => x"20",
         15192 => x"20",
         15193 => x"58",
         15194 => x"00",
         15195 => x"20",
         15196 => x"73",
         15197 => x"20",
         15198 => x"63",
         15199 => x"72",
         15200 => x"20",
         15201 => x"20",
         15202 => x"20",
         15203 => x"25",
         15204 => x"4d",
         15205 => x"00",
         15206 => x"20",
         15207 => x"73",
         15208 => x"6e",
         15209 => x"44",
         15210 => x"20",
         15211 => x"63",
         15212 => x"72",
         15213 => x"20",
         15214 => x"25",
         15215 => x"4d",
         15216 => x"00",
         15217 => x"20",
         15218 => x"52",
         15219 => x"43",
         15220 => x"6b",
         15221 => x"65",
         15222 => x"20",
         15223 => x"20",
         15224 => x"20",
         15225 => x"25",
         15226 => x"4d",
         15227 => x"00",
         15228 => x"20",
         15229 => x"49",
         15230 => x"20",
         15231 => x"32",
         15232 => x"20",
         15233 => x"43",
         15234 => x"00",
         15235 => x"20",
         15236 => x"20",
         15237 => x"00",
         15238 => x"20",
         15239 => x"53",
         15240 => x"4e",
         15241 => x"55",
         15242 => x"00",
         15243 => x"20",
         15244 => x"54",
         15245 => x"54",
         15246 => x"28",
         15247 => x"6e",
         15248 => x"73",
         15249 => x"32",
         15250 => x"0a",
         15251 => x"20",
         15252 => x"4d",
         15253 => x"20",
         15254 => x"28",
         15255 => x"65",
         15256 => x"20",
         15257 => x"32",
         15258 => x"0a",
         15259 => x"20",
         15260 => x"20",
         15261 => x"44",
         15262 => x"28",
         15263 => x"69",
         15264 => x"20",
         15265 => x"32",
         15266 => x"0a",
         15267 => x"20",
         15268 => x"4d",
         15269 => x"20",
         15270 => x"28",
         15271 => x"58",
         15272 => x"38",
         15273 => x"0a",
         15274 => x"20",
         15275 => x"41",
         15276 => x"20",
         15277 => x"28",
         15278 => x"58",
         15279 => x"38",
         15280 => x"0a",
         15281 => x"20",
         15282 => x"53",
         15283 => x"52",
         15284 => x"28",
         15285 => x"58",
         15286 => x"38",
         15287 => x"0a",
         15288 => x"20",
         15289 => x"52",
         15290 => x"20",
         15291 => x"28",
         15292 => x"58",
         15293 => x"38",
         15294 => x"0a",
         15295 => x"20",
         15296 => x"20",
         15297 => x"41",
         15298 => x"28",
         15299 => x"58",
         15300 => x"38",
         15301 => x"0a",
         15302 => x"66",
         15303 => x"20",
         15304 => x"20",
         15305 => x"66",
         15306 => x"00",
         15307 => x"6b",
         15308 => x"6e",
         15309 => x"4f",
         15310 => x"00",
         15311 => x"61",
         15312 => x"00",
         15313 => x"64",
         15314 => x"00",
         15315 => x"65",
         15316 => x"00",
         15317 => x"4f",
         15318 => x"f0",
         15319 => x"00",
         15320 => x"00",
         15321 => x"f0",
         15322 => x"00",
         15323 => x"00",
         15324 => x"f0",
         15325 => x"00",
         15326 => x"00",
         15327 => x"f0",
         15328 => x"00",
         15329 => x"00",
         15330 => x"f0",
         15331 => x"00",
         15332 => x"00",
         15333 => x"f0",
         15334 => x"00",
         15335 => x"00",
         15336 => x"f0",
         15337 => x"00",
         15338 => x"00",
         15339 => x"f0",
         15340 => x"00",
         15341 => x"00",
         15342 => x"f0",
         15343 => x"00",
         15344 => x"00",
         15345 => x"f0",
         15346 => x"00",
         15347 => x"00",
         15348 => x"f0",
         15349 => x"00",
         15350 => x"00",
         15351 => x"f0",
         15352 => x"00",
         15353 => x"00",
         15354 => x"f0",
         15355 => x"00",
         15356 => x"00",
         15357 => x"f0",
         15358 => x"00",
         15359 => x"00",
         15360 => x"f0",
         15361 => x"00",
         15362 => x"00",
         15363 => x"f0",
         15364 => x"00",
         15365 => x"00",
         15366 => x"f0",
         15367 => x"00",
         15368 => x"00",
         15369 => x"f0",
         15370 => x"00",
         15371 => x"00",
         15372 => x"f0",
         15373 => x"00",
         15374 => x"00",
         15375 => x"f0",
         15376 => x"00",
         15377 => x"00",
         15378 => x"f0",
         15379 => x"00",
         15380 => x"00",
         15381 => x"f0",
         15382 => x"00",
         15383 => x"00",
         15384 => x"44",
         15385 => x"43",
         15386 => x"42",
         15387 => x"41",
         15388 => x"36",
         15389 => x"35",
         15390 => x"34",
         15391 => x"46",
         15392 => x"33",
         15393 => x"32",
         15394 => x"31",
         15395 => x"00",
         15396 => x"00",
         15397 => x"00",
         15398 => x"00",
         15399 => x"00",
         15400 => x"00",
         15401 => x"00",
         15402 => x"00",
         15403 => x"00",
         15404 => x"00",
         15405 => x"00",
         15406 => x"6e",
         15407 => x"20",
         15408 => x"6e",
         15409 => x"65",
         15410 => x"20",
         15411 => x"74",
         15412 => x"20",
         15413 => x"65",
         15414 => x"69",
         15415 => x"6c",
         15416 => x"2e",
         15417 => x"73",
         15418 => x"79",
         15419 => x"73",
         15420 => x"00",
         15421 => x"00",
         15422 => x"36",
         15423 => x"20",
         15424 => x"00",
         15425 => x"69",
         15426 => x"20",
         15427 => x"72",
         15428 => x"74",
         15429 => x"65",
         15430 => x"73",
         15431 => x"79",
         15432 => x"6c",
         15433 => x"6f",
         15434 => x"46",
         15435 => x"00",
         15436 => x"73",
         15437 => x"00",
         15438 => x"31",
         15439 => x"00",
         15440 => x"41",
         15441 => x"42",
         15442 => x"43",
         15443 => x"44",
         15444 => x"31",
         15445 => x"00",
         15446 => x"31",
         15447 => x"00",
         15448 => x"31",
         15449 => x"00",
         15450 => x"31",
         15451 => x"00",
         15452 => x"31",
         15453 => x"00",
         15454 => x"31",
         15455 => x"00",
         15456 => x"31",
         15457 => x"00",
         15458 => x"31",
         15459 => x"00",
         15460 => x"31",
         15461 => x"00",
         15462 => x"32",
         15463 => x"00",
         15464 => x"32",
         15465 => x"00",
         15466 => x"33",
         15467 => x"00",
         15468 => x"46",
         15469 => x"35",
         15470 => x"00",
         15471 => x"36",
         15472 => x"00",
         15473 => x"25",
         15474 => x"64",
         15475 => x"2c",
         15476 => x"25",
         15477 => x"64",
         15478 => x"32",
         15479 => x"00",
         15480 => x"25",
         15481 => x"64",
         15482 => x"3a",
         15483 => x"25",
         15484 => x"64",
         15485 => x"3a",
         15486 => x"2c",
         15487 => x"25",
         15488 => x"00",
         15489 => x"32",
         15490 => x"00",
         15491 => x"5b",
         15492 => x"25",
         15493 => x"00",
         15494 => x"70",
         15495 => x"20",
         15496 => x"73",
         15497 => x"00",
         15498 => x"3a",
         15499 => x"78",
         15500 => x"32",
         15501 => x"00",
         15502 => x"3a",
         15503 => x"78",
         15504 => x"32",
         15505 => x"00",
         15506 => x"3a",
         15507 => x"78",
         15508 => x"00",
         15509 => x"64",
         15510 => x"69",
         15511 => x"53",
         15512 => x"6e",
         15513 => x"00",
         15514 => x"64",
         15515 => x"69",
         15516 => x"53",
         15517 => x"65",
         15518 => x"00",
         15519 => x"64",
         15520 => x"69",
         15521 => x"53",
         15522 => x"72",
         15523 => x"00",
         15524 => x"20",
         15525 => x"74",
         15526 => x"66",
         15527 => x"64",
         15528 => x"00",
         15529 => x"00",
         15530 => x"3a",
         15531 => x"7c",
         15532 => x"00",
         15533 => x"3b",
         15534 => x"00",
         15535 => x"54",
         15536 => x"54",
         15537 => x"00",
         15538 => x"90",
         15539 => x"4f",
         15540 => x"30",
         15541 => x"20",
         15542 => x"45",
         15543 => x"20",
         15544 => x"20",
         15545 => x"20",
         15546 => x"20",
         15547 => x"45",
         15548 => x"20",
         15549 => x"33",
         15550 => x"20",
         15551 => x"f2",
         15552 => x"00",
         15553 => x"00",
         15554 => x"00",
         15555 => x"05",
         15556 => x"10",
         15557 => x"18",
         15558 => x"00",
         15559 => x"45",
         15560 => x"8f",
         15561 => x"45",
         15562 => x"8e",
         15563 => x"92",
         15564 => x"55",
         15565 => x"9a",
         15566 => x"9e",
         15567 => x"4f",
         15568 => x"a6",
         15569 => x"aa",
         15570 => x"ae",
         15571 => x"b2",
         15572 => x"b6",
         15573 => x"ba",
         15574 => x"be",
         15575 => x"c2",
         15576 => x"c6",
         15577 => x"ca",
         15578 => x"ce",
         15579 => x"d2",
         15580 => x"d6",
         15581 => x"da",
         15582 => x"de",
         15583 => x"e2",
         15584 => x"e6",
         15585 => x"ea",
         15586 => x"ee",
         15587 => x"f2",
         15588 => x"f6",
         15589 => x"fa",
         15590 => x"fe",
         15591 => x"2c",
         15592 => x"5d",
         15593 => x"2a",
         15594 => x"3f",
         15595 => x"00",
         15596 => x"00",
         15597 => x"00",
         15598 => x"02",
         15599 => x"00",
         15600 => x"00",
         15601 => x"00",
         15602 => x"00",
         15603 => x"00",
         15604 => x"00",
         15605 => x"00",
         15606 => x"00",
         15607 => x"00",
         15608 => x"00",
         15609 => x"00",
         15610 => x"00",
         15611 => x"00",
         15612 => x"00",
         15613 => x"00",
         15614 => x"00",
         15615 => x"00",
         15616 => x"00",
         15617 => x"00",
         15618 => x"00",
         15619 => x"01",
         15620 => x"00",
         15621 => x"00",
         15622 => x"00",
         15623 => x"00",
         15624 => x"23",
         15625 => x"00",
         15626 => x"00",
         15627 => x"00",
         15628 => x"25",
         15629 => x"25",
         15630 => x"25",
         15631 => x"25",
         15632 => x"25",
         15633 => x"25",
         15634 => x"25",
         15635 => x"25",
         15636 => x"25",
         15637 => x"25",
         15638 => x"25",
         15639 => x"25",
         15640 => x"25",
         15641 => x"25",
         15642 => x"25",
         15643 => x"25",
         15644 => x"25",
         15645 => x"25",
         15646 => x"25",
         15647 => x"25",
         15648 => x"25",
         15649 => x"25",
         15650 => x"25",
         15651 => x"25",
         15652 => x"00",
         15653 => x"03",
         15654 => x"03",
         15655 => x"03",
         15656 => x"03",
         15657 => x"03",
         15658 => x"03",
         15659 => x"22",
         15660 => x"00",
         15661 => x"22",
         15662 => x"23",
         15663 => x"22",
         15664 => x"22",
         15665 => x"22",
         15666 => x"00",
         15667 => x"00",
         15668 => x"03",
         15669 => x"03",
         15670 => x"03",
         15671 => x"00",
         15672 => x"01",
         15673 => x"01",
         15674 => x"01",
         15675 => x"01",
         15676 => x"01",
         15677 => x"01",
         15678 => x"02",
         15679 => x"01",
         15680 => x"01",
         15681 => x"01",
         15682 => x"01",
         15683 => x"01",
         15684 => x"01",
         15685 => x"01",
         15686 => x"01",
         15687 => x"01",
         15688 => x"01",
         15689 => x"01",
         15690 => x"01",
         15691 => x"02",
         15692 => x"01",
         15693 => x"02",
         15694 => x"01",
         15695 => x"01",
         15696 => x"01",
         15697 => x"01",
         15698 => x"01",
         15699 => x"01",
         15700 => x"01",
         15701 => x"01",
         15702 => x"01",
         15703 => x"01",
         15704 => x"01",
         15705 => x"01",
         15706 => x"01",
         15707 => x"01",
         15708 => x"01",
         15709 => x"01",
         15710 => x"01",
         15711 => x"01",
         15712 => x"01",
         15713 => x"01",
         15714 => x"01",
         15715 => x"01",
         15716 => x"01",
         15717 => x"01",
         15718 => x"00",
         15719 => x"01",
         15720 => x"01",
         15721 => x"01",
         15722 => x"01",
         15723 => x"01",
         15724 => x"01",
         15725 => x"00",
         15726 => x"02",
         15727 => x"02",
         15728 => x"02",
         15729 => x"02",
         15730 => x"02",
         15731 => x"02",
         15732 => x"01",
         15733 => x"02",
         15734 => x"01",
         15735 => x"01",
         15736 => x"01",
         15737 => x"02",
         15738 => x"02",
         15739 => x"02",
         15740 => x"01",
         15741 => x"02",
         15742 => x"02",
         15743 => x"01",
         15744 => x"2c",
         15745 => x"02",
         15746 => x"01",
         15747 => x"02",
         15748 => x"02",
         15749 => x"01",
         15750 => x"02",
         15751 => x"02",
         15752 => x"02",
         15753 => x"2c",
         15754 => x"02",
         15755 => x"02",
         15756 => x"01",
         15757 => x"02",
         15758 => x"02",
         15759 => x"02",
         15760 => x"01",
         15761 => x"02",
         15762 => x"02",
         15763 => x"02",
         15764 => x"03",
         15765 => x"03",
         15766 => x"03",
         15767 => x"00",
         15768 => x"03",
         15769 => x"03",
         15770 => x"03",
         15771 => x"00",
         15772 => x"03",
         15773 => x"03",
         15774 => x"00",
         15775 => x"03",
         15776 => x"03",
         15777 => x"03",
         15778 => x"03",
         15779 => x"03",
         15780 => x"03",
         15781 => x"03",
         15782 => x"03",
         15783 => x"04",
         15784 => x"04",
         15785 => x"04",
         15786 => x"04",
         15787 => x"04",
         15788 => x"04",
         15789 => x"04",
         15790 => x"01",
         15791 => x"04",
         15792 => x"00",
         15793 => x"00",
         15794 => x"1e",
         15795 => x"1e",
         15796 => x"1f",
         15797 => x"1f",
         15798 => x"1f",
         15799 => x"1f",
         15800 => x"1f",
         15801 => x"1f",
         15802 => x"1f",
         15803 => x"1f",
         15804 => x"1f",
         15805 => x"1f",
         15806 => x"06",
         15807 => x"00",
         15808 => x"1f",
         15809 => x"1f",
         15810 => x"1f",
         15811 => x"1f",
         15812 => x"1f",
         15813 => x"1f",
         15814 => x"1f",
         15815 => x"06",
         15816 => x"06",
         15817 => x"06",
         15818 => x"00",
         15819 => x"1f",
         15820 => x"1f",
         15821 => x"00",
         15822 => x"1f",
         15823 => x"1f",
         15824 => x"1f",
         15825 => x"1f",
         15826 => x"00",
         15827 => x"21",
         15828 => x"21",
         15829 => x"02",
         15830 => x"00",
         15831 => x"24",
         15832 => x"2c",
         15833 => x"2c",
         15834 => x"2c",
         15835 => x"2c",
         15836 => x"2c",
         15837 => x"2d",
         15838 => x"ff",
         15839 => x"00",
         15840 => x"00",
         15841 => x"e6",
         15842 => x"01",
         15843 => x"00",
         15844 => x"00",
         15845 => x"e6",
         15846 => x"01",
         15847 => x"00",
         15848 => x"00",
         15849 => x"e6",
         15850 => x"03",
         15851 => x"00",
         15852 => x"00",
         15853 => x"e6",
         15854 => x"03",
         15855 => x"00",
         15856 => x"00",
         15857 => x"e6",
         15858 => x"03",
         15859 => x"00",
         15860 => x"00",
         15861 => x"e6",
         15862 => x"04",
         15863 => x"00",
         15864 => x"00",
         15865 => x"e6",
         15866 => x"04",
         15867 => x"00",
         15868 => x"00",
         15869 => x"e6",
         15870 => x"04",
         15871 => x"00",
         15872 => x"00",
         15873 => x"e6",
         15874 => x"04",
         15875 => x"00",
         15876 => x"00",
         15877 => x"e6",
         15878 => x"04",
         15879 => x"00",
         15880 => x"00",
         15881 => x"e6",
         15882 => x"04",
         15883 => x"00",
         15884 => x"00",
         15885 => x"e7",
         15886 => x"04",
         15887 => x"00",
         15888 => x"00",
         15889 => x"e7",
         15890 => x"05",
         15891 => x"00",
         15892 => x"00",
         15893 => x"e7",
         15894 => x"05",
         15895 => x"00",
         15896 => x"00",
         15897 => x"e7",
         15898 => x"05",
         15899 => x"00",
         15900 => x"00",
         15901 => x"e7",
         15902 => x"05",
         15903 => x"00",
         15904 => x"00",
         15905 => x"e7",
         15906 => x"07",
         15907 => x"00",
         15908 => x"00",
         15909 => x"e7",
         15910 => x"07",
         15911 => x"00",
         15912 => x"00",
         15913 => x"e7",
         15914 => x"08",
         15915 => x"00",
         15916 => x"00",
         15917 => x"e7",
         15918 => x"08",
         15919 => x"00",
         15920 => x"00",
         15921 => x"e7",
         15922 => x"08",
         15923 => x"00",
         15924 => x"00",
         15925 => x"e7",
         15926 => x"08",
         15927 => x"00",
         15928 => x"00",
         15929 => x"e7",
         15930 => x"08",
         15931 => x"00",
         15932 => x"00",
         15933 => x"e7",
         15934 => x"08",
         15935 => x"00",
         15936 => x"00",
         15937 => x"e7",
         15938 => x"09",
         15939 => x"00",
         15940 => x"00",
         15941 => x"e7",
         15942 => x"09",
         15943 => x"00",
         15944 => x"00",
         15945 => x"e7",
         15946 => x"09",
         15947 => x"00",
         15948 => x"00",
         15949 => x"e7",
         15950 => x"09",
         15951 => x"00",
         15952 => x"00",
         15953 => x"00",
         15954 => x"00",
         15955 => x"7f",
         15956 => x"00",
         15957 => x"7f",
         15958 => x"00",
         15959 => x"7f",
         15960 => x"00",
         15961 => x"00",
         15962 => x"00",
         15963 => x"ff",
         15964 => x"00",
         15965 => x"00",
         15966 => x"78",
         15967 => x"00",
         15968 => x"e1",
         15969 => x"e1",
         15970 => x"e1",
         15971 => x"00",
         15972 => x"01",
         15973 => x"01",
         15974 => x"10",
         15975 => x"00",
         15976 => x"00",
         15977 => x"00",
         15978 => x"00",
         15979 => x"00",
         15980 => x"00",
         15981 => x"00",
         15982 => x"00",
         15983 => x"00",
         15984 => x"00",
         15985 => x"00",
         15986 => x"00",
         15987 => x"00",
         15988 => x"00",
         15989 => x"00",
         15990 => x"00",
         15991 => x"00",
         15992 => x"00",
         15993 => x"00",
         15994 => x"00",
         15995 => x"00",
         15996 => x"00",
         15997 => x"00",
         15998 => x"00",
         15999 => x"00",
         16000 => x"f0",
         16001 => x"00",
         16002 => x"f0",
         16003 => x"00",
         16004 => x"f0",
         16005 => x"00",
         16006 => x"fd",
         16007 => x"5f",
         16008 => x"3a",
         16009 => x"40",
         16010 => x"f0",
         16011 => x"73",
         16012 => x"77",
         16013 => x"6b",
         16014 => x"6f",
         16015 => x"63",
         16016 => x"67",
         16017 => x"33",
         16018 => x"37",
         16019 => x"2d",
         16020 => x"2c",
         16021 => x"f3",
         16022 => x"3f",
         16023 => x"f0",
         16024 => x"f0",
         16025 => x"82",
         16026 => x"f0",
         16027 => x"58",
         16028 => x"3b",
         16029 => x"40",
         16030 => x"f0",
         16031 => x"53",
         16032 => x"57",
         16033 => x"4b",
         16034 => x"4f",
         16035 => x"43",
         16036 => x"47",
         16037 => x"33",
         16038 => x"37",
         16039 => x"2d",
         16040 => x"2c",
         16041 => x"f3",
         16042 => x"3f",
         16043 => x"f0",
         16044 => x"f0",
         16045 => x"82",
         16046 => x"f0",
         16047 => x"58",
         16048 => x"2a",
         16049 => x"60",
         16050 => x"f0",
         16051 => x"53",
         16052 => x"57",
         16053 => x"4b",
         16054 => x"4f",
         16055 => x"43",
         16056 => x"47",
         16057 => x"23",
         16058 => x"27",
         16059 => x"3d",
         16060 => x"3c",
         16061 => x"e0",
         16062 => x"3f",
         16063 => x"f0",
         16064 => x"f0",
         16065 => x"87",
         16066 => x"f0",
         16067 => x"1e",
         16068 => x"f0",
         16069 => x"00",
         16070 => x"f0",
         16071 => x"13",
         16072 => x"17",
         16073 => x"0b",
         16074 => x"0f",
         16075 => x"03",
         16076 => x"07",
         16077 => x"f0",
         16078 => x"f0",
         16079 => x"f0",
         16080 => x"f0",
         16081 => x"f0",
         16082 => x"f0",
         16083 => x"f0",
         16084 => x"f0",
         16085 => x"82",
         16086 => x"f0",
         16087 => x"cf",
         16088 => x"4d",
         16089 => x"d7",
         16090 => x"f0",
         16091 => x"41",
         16092 => x"78",
         16093 => x"6c",
         16094 => x"d5",
         16095 => x"d9",
         16096 => x"4c",
         16097 => x"7e",
         16098 => x"5f",
         16099 => x"d1",
         16100 => x"d0",
         16101 => x"c2",
         16102 => x"bb",
         16103 => x"f0",
         16104 => x"f0",
         16105 => x"82",
         16106 => x"f0",
         16107 => x"00",
         16108 => x"00",
         16109 => x"00",
         16110 => x"00",
         16111 => x"00",
         16112 => x"00",
         16113 => x"00",
         16114 => x"00",
         16115 => x"00",
         16116 => x"00",
         16117 => x"00",
         16118 => x"00",
         16119 => x"00",
         16120 => x"00",
         16121 => x"00",
         16122 => x"00",
         16123 => x"00",
         16124 => x"00",
         16125 => x"00",
         16126 => x"00",
         16127 => x"00",
         16128 => x"00",
         16129 => x"00",
         16130 => x"00",
         16131 => x"00",
         16132 => x"00",
         16133 => x"00",
         16134 => x"00",
         16135 => x"f1",
         16136 => x"00",
         16137 => x"f1",
         16138 => x"00",
         16139 => x"f1",
         16140 => x"00",
         16141 => x"f1",
         16142 => x"00",
         16143 => x"f1",
         16144 => x"00",
         16145 => x"f1",
         16146 => x"00",
         16147 => x"f1",
         16148 => x"00",
         16149 => x"f1",
         16150 => x"00",
         16151 => x"f1",
         16152 => x"00",
         16153 => x"f1",
         16154 => x"00",
         16155 => x"f1",
         16156 => x"00",
         16157 => x"f1",
         16158 => x"00",
         16159 => x"f1",
         16160 => x"00",
         16161 => x"f1",
         16162 => x"00",
         16163 => x"f1",
         16164 => x"00",
         16165 => x"f1",
         16166 => x"00",
         16167 => x"f1",
         16168 => x"00",
         16169 => x"f1",
         16170 => x"00",
         16171 => x"f1",
         16172 => x"00",
         16173 => x"f1",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"00",
         18159 => x"00",
         18160 => x"00",
         18161 => x"00",
         18162 => x"00",
         18163 => x"00",
         18164 => x"00",
         18165 => x"00",
         18166 => x"00",
         18167 => x"00",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"32",
         18176 => x"01",
         18177 => x"00",
         18178 => x"f2",
         18179 => x"f6",
         18180 => x"fa",
         18181 => x"fe",
         18182 => x"c2",
         18183 => x"c6",
         18184 => x"e5",
         18185 => x"ef",
         18186 => x"62",
         18187 => x"66",
         18188 => x"6b",
         18189 => x"2e",
         18190 => x"22",
         18191 => x"26",
         18192 => x"4f",
         18193 => x"57",
         18194 => x"02",
         18195 => x"06",
         18196 => x"0a",
         18197 => x"0e",
         18198 => x"12",
         18199 => x"16",
         18200 => x"1a",
         18201 => x"be",
         18202 => x"82",
         18203 => x"86",
         18204 => x"8a",
         18205 => x"8e",
         18206 => x"92",
         18207 => x"96",
         18208 => x"9a",
         18209 => x"a5",
         18210 => x"00",
         18211 => x"00",
         18212 => x"00",
         18213 => x"00",
         18214 => x"00",
         18215 => x"00",
         18216 => x"00",
         18217 => x"00",
         18218 => x"00",
         18219 => x"00",
         18220 => x"00",
         18221 => x"00",
         18222 => x"00",
         18223 => x"00",
         18224 => x"00",
         18225 => x"00",
         18226 => x"00",
         18227 => x"00",
         18228 => x"00",
         18229 => x"00",
         18230 => x"00",
         18231 => x"00",
         18232 => x"00",
         18233 => x"00",
         18234 => x"00",
         18235 => x"00",
         18236 => x"00",
         18237 => x"00",
         18238 => x"00",
         18239 => x"00",
         18240 => x"00",
         18241 => x"01",
         18242 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"b5",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8e",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8f",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"90",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"91",
           324 => x"0b",
           325 => x"04",
           326 => x"91",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"92",
           336 => x"0b",
           337 => x"04",
           338 => x"92",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"84",
           386 => x"80",
           387 => x"84",
           388 => x"80",
           389 => x"04",
           390 => x"0c",
           391 => x"84",
           392 => x"80",
           393 => x"04",
           394 => x"0c",
           395 => x"84",
           396 => x"80",
           397 => x"04",
           398 => x"0c",
           399 => x"84",
           400 => x"80",
           401 => x"04",
           402 => x"0c",
           403 => x"84",
           404 => x"80",
           405 => x"04",
           406 => x"0c",
           407 => x"84",
           408 => x"80",
           409 => x"04",
           410 => x"0c",
           411 => x"84",
           412 => x"80",
           413 => x"04",
           414 => x"0c",
           415 => x"84",
           416 => x"80",
           417 => x"04",
           418 => x"0c",
           419 => x"84",
           420 => x"80",
           421 => x"04",
           422 => x"0c",
           423 => x"84",
           424 => x"80",
           425 => x"04",
           426 => x"0c",
           427 => x"84",
           428 => x"80",
           429 => x"04",
           430 => x"0c",
           431 => x"84",
           432 => x"80",
           433 => x"04",
           434 => x"0c",
           435 => x"2d",
           436 => x"08",
           437 => x"90",
           438 => x"98",
           439 => x"c0",
           440 => x"98",
           441 => x"80",
           442 => x"ba",
           443 => x"d2",
           444 => x"ba",
           445 => x"c0",
           446 => x"84",
           447 => x"80",
           448 => x"84",
           449 => x"80",
           450 => x"04",
           451 => x"0c",
           452 => x"2d",
           453 => x"08",
           454 => x"90",
           455 => x"98",
           456 => x"c9",
           457 => x"98",
           458 => x"80",
           459 => x"ba",
           460 => x"d2",
           461 => x"ba",
           462 => x"c0",
           463 => x"84",
           464 => x"82",
           465 => x"84",
           466 => x"80",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"90",
           472 => x"98",
           473 => x"ee",
           474 => x"98",
           475 => x"80",
           476 => x"ba",
           477 => x"df",
           478 => x"ba",
           479 => x"c0",
           480 => x"84",
           481 => x"82",
           482 => x"84",
           483 => x"80",
           484 => x"04",
           485 => x"0c",
           486 => x"2d",
           487 => x"08",
           488 => x"90",
           489 => x"98",
           490 => x"a9",
           491 => x"98",
           492 => x"80",
           493 => x"ba",
           494 => x"84",
           495 => x"ba",
           496 => x"c0",
           497 => x"84",
           498 => x"82",
           499 => x"84",
           500 => x"80",
           501 => x"04",
           502 => x"0c",
           503 => x"2d",
           504 => x"08",
           505 => x"90",
           506 => x"98",
           507 => x"86",
           508 => x"98",
           509 => x"80",
           510 => x"ba",
           511 => x"94",
           512 => x"ba",
           513 => x"c0",
           514 => x"84",
           515 => x"83",
           516 => x"84",
           517 => x"80",
           518 => x"04",
           519 => x"0c",
           520 => x"2d",
           521 => x"08",
           522 => x"90",
           523 => x"98",
           524 => x"b0",
           525 => x"98",
           526 => x"80",
           527 => x"ba",
           528 => x"e7",
           529 => x"ba",
           530 => x"c0",
           531 => x"84",
           532 => x"82",
           533 => x"84",
           534 => x"80",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"90",
           540 => x"98",
           541 => x"c0",
           542 => x"98",
           543 => x"80",
           544 => x"ba",
           545 => x"a1",
           546 => x"ba",
           547 => x"c0",
           548 => x"84",
           549 => x"82",
           550 => x"84",
           551 => x"80",
           552 => x"04",
           553 => x"0c",
           554 => x"2d",
           555 => x"08",
           556 => x"90",
           557 => x"98",
           558 => x"dc",
           559 => x"98",
           560 => x"80",
           561 => x"ba",
           562 => x"b8",
           563 => x"ba",
           564 => x"c0",
           565 => x"84",
           566 => x"81",
           567 => x"84",
           568 => x"80",
           569 => x"04",
           570 => x"0c",
           571 => x"2d",
           572 => x"08",
           573 => x"90",
           574 => x"98",
           575 => x"aa",
           576 => x"98",
           577 => x"80",
           578 => x"ba",
           579 => x"d0",
           580 => x"ba",
           581 => x"c0",
           582 => x"84",
           583 => x"80",
           584 => x"84",
           585 => x"80",
           586 => x"04",
           587 => x"0c",
           588 => x"2d",
           589 => x"08",
           590 => x"90",
           591 => x"98",
           592 => x"2d",
           593 => x"08",
           594 => x"90",
           595 => x"98",
           596 => x"ca",
           597 => x"98",
           598 => x"80",
           599 => x"ba",
           600 => x"dd",
           601 => x"ba",
           602 => x"c0",
           603 => x"84",
           604 => x"81",
           605 => x"84",
           606 => x"80",
           607 => x"04",
           608 => x"0c",
           609 => x"2d",
           610 => x"08",
           611 => x"90",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"51",
           621 => x"73",
           622 => x"73",
           623 => x"81",
           624 => x"10",
           625 => x"07",
           626 => x"0c",
           627 => x"72",
           628 => x"81",
           629 => x"09",
           630 => x"71",
           631 => x"0a",
           632 => x"72",
           633 => x"51",
           634 => x"84",
           635 => x"84",
           636 => x"8e",
           637 => x"70",
           638 => x"0c",
           639 => x"93",
           640 => x"81",
           641 => x"c4",
           642 => x"3d",
           643 => x"70",
           644 => x"52",
           645 => x"74",
           646 => x"f0",
           647 => x"c5",
           648 => x"0d",
           649 => x"0d",
           650 => x"85",
           651 => x"32",
           652 => x"73",
           653 => x"58",
           654 => x"52",
           655 => x"09",
           656 => x"d3",
           657 => x"77",
           658 => x"70",
           659 => x"07",
           660 => x"55",
           661 => x"80",
           662 => x"38",
           663 => x"b2",
           664 => x"8e",
           665 => x"ba",
           666 => x"84",
           667 => x"ff",
           668 => x"84",
           669 => x"75",
           670 => x"57",
           671 => x"73",
           672 => x"30",
           673 => x"9f",
           674 => x"54",
           675 => x"24",
           676 => x"75",
           677 => x"71",
           678 => x"0c",
           679 => x"04",
           680 => x"ba",
           681 => x"3d",
           682 => x"3d",
           683 => x"86",
           684 => x"99",
           685 => x"56",
           686 => x"8e",
           687 => x"53",
           688 => x"3d",
           689 => x"9d",
           690 => x"54",
           691 => x"8d",
           692 => x"fd",
           693 => x"3d",
           694 => x"76",
           695 => x"85",
           696 => x"0d",
           697 => x"0d",
           698 => x"42",
           699 => x"70",
           700 => x"85",
           701 => x"81",
           702 => x"81",
           703 => x"5b",
           704 => x"7b",
           705 => x"06",
           706 => x"7b",
           707 => x"7b",
           708 => x"38",
           709 => x"81",
           710 => x"72",
           711 => x"81",
           712 => x"5f",
           713 => x"81",
           714 => x"b0",
           715 => x"70",
           716 => x"54",
           717 => x"38",
           718 => x"a9",
           719 => x"2a",
           720 => x"81",
           721 => x"7e",
           722 => x"38",
           723 => x"07",
           724 => x"57",
           725 => x"38",
           726 => x"54",
           727 => x"8c",
           728 => x"0d",
           729 => x"2a",
           730 => x"10",
           731 => x"05",
           732 => x"70",
           733 => x"70",
           734 => x"29",
           735 => x"70",
           736 => x"5a",
           737 => x"80",
           738 => x"86",
           739 => x"06",
           740 => x"bd",
           741 => x"33",
           742 => x"fe",
           743 => x"b8",
           744 => x"2e",
           745 => x"93",
           746 => x"74",
           747 => x"8a",
           748 => x"5a",
           749 => x"38",
           750 => x"7c",
           751 => x"8b",
           752 => x"33",
           753 => x"cc",
           754 => x"39",
           755 => x"70",
           756 => x"55",
           757 => x"81",
           758 => x"40",
           759 => x"38",
           760 => x"72",
           761 => x"97",
           762 => x"10",
           763 => x"05",
           764 => x"04",
           765 => x"54",
           766 => x"73",
           767 => x"7c",
           768 => x"8a",
           769 => x"7c",
           770 => x"76",
           771 => x"fe",
           772 => x"ff",
           773 => x"39",
           774 => x"60",
           775 => x"08",
           776 => x"cf",
           777 => x"41",
           778 => x"9c",
           779 => x"75",
           780 => x"3f",
           781 => x"08",
           782 => x"84",
           783 => x"18",
           784 => x"53",
           785 => x"88",
           786 => x"8c",
           787 => x"55",
           788 => x"81",
           789 => x"79",
           790 => x"90",
           791 => x"ba",
           792 => x"84",
           793 => x"c5",
           794 => x"ba",
           795 => x"2b",
           796 => x"40",
           797 => x"2e",
           798 => x"84",
           799 => x"fc",
           800 => x"70",
           801 => x"55",
           802 => x"70",
           803 => x"5f",
           804 => x"9e",
           805 => x"80",
           806 => x"80",
           807 => x"79",
           808 => x"38",
           809 => x"80",
           810 => x"80",
           811 => x"90",
           812 => x"83",
           813 => x"06",
           814 => x"80",
           815 => x"75",
           816 => x"81",
           817 => x"54",
           818 => x"86",
           819 => x"83",
           820 => x"70",
           821 => x"86",
           822 => x"5b",
           823 => x"54",
           824 => x"85",
           825 => x"79",
           826 => x"70",
           827 => x"83",
           828 => x"59",
           829 => x"2e",
           830 => x"7a",
           831 => x"06",
           832 => x"eb",
           833 => x"2a",
           834 => x"73",
           835 => x"7a",
           836 => x"06",
           837 => x"97",
           838 => x"06",
           839 => x"8f",
           840 => x"2a",
           841 => x"7e",
           842 => x"38",
           843 => x"80",
           844 => x"80",
           845 => x"90",
           846 => x"54",
           847 => x"9d",
           848 => x"b0",
           849 => x"3f",
           850 => x"80",
           851 => x"80",
           852 => x"90",
           853 => x"54",
           854 => x"e5",
           855 => x"06",
           856 => x"2e",
           857 => x"79",
           858 => x"29",
           859 => x"05",
           860 => x"5b",
           861 => x"75",
           862 => x"7c",
           863 => x"87",
           864 => x"79",
           865 => x"29",
           866 => x"05",
           867 => x"5b",
           868 => x"80",
           869 => x"7a",
           870 => x"81",
           871 => x"7a",
           872 => x"b9",
           873 => x"e3",
           874 => x"38",
           875 => x"2e",
           876 => x"76",
           877 => x"81",
           878 => x"84",
           879 => x"96",
           880 => x"ff",
           881 => x"52",
           882 => x"3f",
           883 => x"9c",
           884 => x"06",
           885 => x"81",
           886 => x"80",
           887 => x"38",
           888 => x"80",
           889 => x"80",
           890 => x"90",
           891 => x"55",
           892 => x"fc",
           893 => x"52",
           894 => x"f4",
           895 => x"7a",
           896 => x"7a",
           897 => x"33",
           898 => x"fa",
           899 => x"c8",
           900 => x"c0",
           901 => x"f8",
           902 => x"61",
           903 => x"08",
           904 => x"cf",
           905 => x"42",
           906 => x"fd",
           907 => x"84",
           908 => x"80",
           909 => x"13",
           910 => x"2b",
           911 => x"84",
           912 => x"fc",
           913 => x"70",
           914 => x"52",
           915 => x"41",
           916 => x"2a",
           917 => x"5c",
           918 => x"c9",
           919 => x"84",
           920 => x"fc",
           921 => x"70",
           922 => x"54",
           923 => x"25",
           924 => x"7c",
           925 => x"85",
           926 => x"39",
           927 => x"83",
           928 => x"5b",
           929 => x"ff",
           930 => x"ca",
           931 => x"75",
           932 => x"57",
           933 => x"d8",
           934 => x"ff",
           935 => x"ff",
           936 => x"54",
           937 => x"ff",
           938 => x"38",
           939 => x"70",
           940 => x"33",
           941 => x"3f",
           942 => x"fc",
           943 => x"fc",
           944 => x"84",
           945 => x"fc",
           946 => x"70",
           947 => x"58",
           948 => x"7b",
           949 => x"81",
           950 => x"57",
           951 => x"38",
           952 => x"7f",
           953 => x"71",
           954 => x"40",
           955 => x"7e",
           956 => x"38",
           957 => x"bf",
           958 => x"ba",
           959 => x"ad",
           960 => x"07",
           961 => x"5b",
           962 => x"38",
           963 => x"7a",
           964 => x"80",
           965 => x"59",
           966 => x"38",
           967 => x"7f",
           968 => x"71",
           969 => x"06",
           970 => x"5f",
           971 => x"38",
           972 => x"f6",
           973 => x"8c",
           974 => x"ff",
           975 => x"31",
           976 => x"5a",
           977 => x"58",
           978 => x"7a",
           979 => x"7c",
           980 => x"76",
           981 => x"f7",
           982 => x"60",
           983 => x"08",
           984 => x"5d",
           985 => x"79",
           986 => x"75",
           987 => x"3f",
           988 => x"08",
           989 => x"06",
           990 => x"90",
           991 => x"c4",
           992 => x"80",
           993 => x"58",
           994 => x"88",
           995 => x"39",
           996 => x"80",
           997 => x"80",
           998 => x"90",
           999 => x"54",
          1000 => x"fa",
          1001 => x"52",
          1002 => x"c4",
          1003 => x"7c",
          1004 => x"83",
          1005 => x"90",
          1006 => x"06",
          1007 => x"7c",
          1008 => x"83",
          1009 => x"88",
          1010 => x"5f",
          1011 => x"fb",
          1012 => x"d8",
          1013 => x"2c",
          1014 => x"90",
          1015 => x"2c",
          1016 => x"06",
          1017 => x"53",
          1018 => x"38",
          1019 => x"7c",
          1020 => x"82",
          1021 => x"81",
          1022 => x"80",
          1023 => x"38",
          1024 => x"7c",
          1025 => x"2a",
          1026 => x"3f",
          1027 => x"5b",
          1028 => x"f7",
          1029 => x"c8",
          1030 => x"31",
          1031 => x"98",
          1032 => x"f9",
          1033 => x"52",
          1034 => x"c4",
          1035 => x"7c",
          1036 => x"82",
          1037 => x"be",
          1038 => x"75",
          1039 => x"3f",
          1040 => x"08",
          1041 => x"06",
          1042 => x"90",
          1043 => x"fd",
          1044 => x"82",
          1045 => x"71",
          1046 => x"06",
          1047 => x"fd",
          1048 => x"3d",
          1049 => x"ec",
          1050 => x"52",
          1051 => x"b5",
          1052 => x"0d",
          1053 => x"0d",
          1054 => x"0b",
          1055 => x"08",
          1056 => x"70",
          1057 => x"32",
          1058 => x"51",
          1059 => x"57",
          1060 => x"77",
          1061 => x"06",
          1062 => x"74",
          1063 => x"56",
          1064 => x"77",
          1065 => x"84",
          1066 => x"52",
          1067 => x"14",
          1068 => x"2d",
          1069 => x"08",
          1070 => x"38",
          1071 => x"70",
          1072 => x"33",
          1073 => x"2e",
          1074 => x"d5",
          1075 => x"d7",
          1076 => x"f0",
          1077 => x"d5",
          1078 => x"8a",
          1079 => x"08",
          1080 => x"84",
          1081 => x"80",
          1082 => x"ff",
          1083 => x"75",
          1084 => x"0c",
          1085 => x"04",
          1086 => x"78",
          1087 => x"80",
          1088 => x"33",
          1089 => x"81",
          1090 => x"06",
          1091 => x"57",
          1092 => x"77",
          1093 => x"06",
          1094 => x"70",
          1095 => x"33",
          1096 => x"2e",
          1097 => x"98",
          1098 => x"75",
          1099 => x"0c",
          1100 => x"04",
          1101 => x"05",
          1102 => x"72",
          1103 => x"38",
          1104 => x"51",
          1105 => x"53",
          1106 => x"ba",
          1107 => x"2e",
          1108 => x"74",
          1109 => x"56",
          1110 => x"72",
          1111 => x"39",
          1112 => x"84",
          1113 => x"52",
          1114 => x"3f",
          1115 => x"04",
          1116 => x"78",
          1117 => x"33",
          1118 => x"81",
          1119 => x"56",
          1120 => x"ff",
          1121 => x"38",
          1122 => x"81",
          1123 => x"80",
          1124 => x"8c",
          1125 => x"72",
          1126 => x"25",
          1127 => x"08",
          1128 => x"34",
          1129 => x"05",
          1130 => x"15",
          1131 => x"13",
          1132 => x"76",
          1133 => x"ba",
          1134 => x"3d",
          1135 => x"52",
          1136 => x"06",
          1137 => x"08",
          1138 => x"ff",
          1139 => x"8c",
          1140 => x"8c",
          1141 => x"05",
          1142 => x"76",
          1143 => x"fb",
          1144 => x"85",
          1145 => x"81",
          1146 => x"81",
          1147 => x"55",
          1148 => x"ff",
          1149 => x"38",
          1150 => x"81",
          1151 => x"b3",
          1152 => x"2a",
          1153 => x"71",
          1154 => x"c3",
          1155 => x"70",
          1156 => x"71",
          1157 => x"f0",
          1158 => x"76",
          1159 => x"08",
          1160 => x"17",
          1161 => x"ff",
          1162 => x"84",
          1163 => x"87",
          1164 => x"74",
          1165 => x"53",
          1166 => x"34",
          1167 => x"81",
          1168 => x"0c",
          1169 => x"84",
          1170 => x"87",
          1171 => x"75",
          1172 => x"08",
          1173 => x"84",
          1174 => x"52",
          1175 => x"08",
          1176 => x"b9",
          1177 => x"33",
          1178 => x"54",
          1179 => x"8c",
          1180 => x"85",
          1181 => x"07",
          1182 => x"17",
          1183 => x"73",
          1184 => x"0c",
          1185 => x"04",
          1186 => x"53",
          1187 => x"34",
          1188 => x"39",
          1189 => x"75",
          1190 => x"54",
          1191 => x"81",
          1192 => x"51",
          1193 => x"ff",
          1194 => x"70",
          1195 => x"33",
          1196 => x"70",
          1197 => x"34",
          1198 => x"73",
          1199 => x"0c",
          1200 => x"04",
          1201 => x"76",
          1202 => x"55",
          1203 => x"70",
          1204 => x"38",
          1205 => x"a1",
          1206 => x"2e",
          1207 => x"70",
          1208 => x"33",
          1209 => x"05",
          1210 => x"11",
          1211 => x"38",
          1212 => x"8c",
          1213 => x"0d",
          1214 => x"55",
          1215 => x"d9",
          1216 => x"75",
          1217 => x"13",
          1218 => x"53",
          1219 => x"34",
          1220 => x"70",
          1221 => x"38",
          1222 => x"13",
          1223 => x"33",
          1224 => x"11",
          1225 => x"38",
          1226 => x"3d",
          1227 => x"53",
          1228 => x"81",
          1229 => x"51",
          1230 => x"ff",
          1231 => x"31",
          1232 => x"0c",
          1233 => x"0d",
          1234 => x"0d",
          1235 => x"54",
          1236 => x"70",
          1237 => x"33",
          1238 => x"70",
          1239 => x"34",
          1240 => x"73",
          1241 => x"0c",
          1242 => x"04",
          1243 => x"75",
          1244 => x"55",
          1245 => x"70",
          1246 => x"38",
          1247 => x"05",
          1248 => x"70",
          1249 => x"34",
          1250 => x"70",
          1251 => x"84",
          1252 => x"85",
          1253 => x"fc",
          1254 => x"78",
          1255 => x"54",
          1256 => x"a1",
          1257 => x"75",
          1258 => x"57",
          1259 => x"71",
          1260 => x"81",
          1261 => x"81",
          1262 => x"80",
          1263 => x"ff",
          1264 => x"e1",
          1265 => x"70",
          1266 => x"0c",
          1267 => x"04",
          1268 => x"f1",
          1269 => x"53",
          1270 => x"80",
          1271 => x"ff",
          1272 => x"81",
          1273 => x"2e",
          1274 => x"72",
          1275 => x"8c",
          1276 => x"0d",
          1277 => x"ba",
          1278 => x"3d",
          1279 => x"3d",
          1280 => x"53",
          1281 => x"80",
          1282 => x"ba",
          1283 => x"ba",
          1284 => x"05",
          1285 => x"b3",
          1286 => x"ba",
          1287 => x"84",
          1288 => x"80",
          1289 => x"84",
          1290 => x"15",
          1291 => x"34",
          1292 => x"52",
          1293 => x"08",
          1294 => x"3f",
          1295 => x"08",
          1296 => x"ba",
          1297 => x"3d",
          1298 => x"3d",
          1299 => x"71",
          1300 => x"53",
          1301 => x"2e",
          1302 => x"70",
          1303 => x"33",
          1304 => x"2e",
          1305 => x"12",
          1306 => x"2e",
          1307 => x"ea",
          1308 => x"70",
          1309 => x"52",
          1310 => x"8c",
          1311 => x"0d",
          1312 => x"0d",
          1313 => x"72",
          1314 => x"54",
          1315 => x"8e",
          1316 => x"70",
          1317 => x"34",
          1318 => x"70",
          1319 => x"84",
          1320 => x"85",
          1321 => x"fa",
          1322 => x"7a",
          1323 => x"52",
          1324 => x"8b",
          1325 => x"80",
          1326 => x"ba",
          1327 => x"e0",
          1328 => x"80",
          1329 => x"73",
          1330 => x"3f",
          1331 => x"8c",
          1332 => x"80",
          1333 => x"26",
          1334 => x"73",
          1335 => x"2e",
          1336 => x"81",
          1337 => x"2a",
          1338 => x"76",
          1339 => x"54",
          1340 => x"56",
          1341 => x"a8",
          1342 => x"74",
          1343 => x"74",
          1344 => x"78",
          1345 => x"11",
          1346 => x"81",
          1347 => x"06",
          1348 => x"ff",
          1349 => x"52",
          1350 => x"55",
          1351 => x"38",
          1352 => x"07",
          1353 => x"ba",
          1354 => x"3d",
          1355 => x"3d",
          1356 => x"fc",
          1357 => x"70",
          1358 => x"07",
          1359 => x"84",
          1360 => x"31",
          1361 => x"70",
          1362 => x"06",
          1363 => x"80",
          1364 => x"88",
          1365 => x"71",
          1366 => x"f0",
          1367 => x"70",
          1368 => x"2b",
          1369 => x"74",
          1370 => x"53",
          1371 => x"73",
          1372 => x"30",
          1373 => x"10",
          1374 => x"77",
          1375 => x"81",
          1376 => x"70",
          1377 => x"30",
          1378 => x"06",
          1379 => x"84",
          1380 => x"51",
          1381 => x"51",
          1382 => x"53",
          1383 => x"51",
          1384 => x"56",
          1385 => x"54",
          1386 => x"0d",
          1387 => x"0d",
          1388 => x"54",
          1389 => x"54",
          1390 => x"84",
          1391 => x"73",
          1392 => x"31",
          1393 => x"0c",
          1394 => x"0d",
          1395 => x"0d",
          1396 => x"54",
          1397 => x"80",
          1398 => x"76",
          1399 => x"3f",
          1400 => x"08",
          1401 => x"52",
          1402 => x"8d",
          1403 => x"fe",
          1404 => x"84",
          1405 => x"31",
          1406 => x"71",
          1407 => x"c5",
          1408 => x"71",
          1409 => x"38",
          1410 => x"71",
          1411 => x"31",
          1412 => x"57",
          1413 => x"80",
          1414 => x"2e",
          1415 => x"10",
          1416 => x"07",
          1417 => x"07",
          1418 => x"ff",
          1419 => x"70",
          1420 => x"72",
          1421 => x"31",
          1422 => x"56",
          1423 => x"58",
          1424 => x"da",
          1425 => x"ba",
          1426 => x"3d",
          1427 => x"3d",
          1428 => x"2c",
          1429 => x"7a",
          1430 => x"32",
          1431 => x"7d",
          1432 => x"32",
          1433 => x"57",
          1434 => x"56",
          1435 => x"55",
          1436 => x"3f",
          1437 => x"08",
          1438 => x"31",
          1439 => x"0c",
          1440 => x"04",
          1441 => x"7b",
          1442 => x"80",
          1443 => x"77",
          1444 => x"56",
          1445 => x"a0",
          1446 => x"06",
          1447 => x"15",
          1448 => x"70",
          1449 => x"73",
          1450 => x"38",
          1451 => x"80",
          1452 => x"b0",
          1453 => x"38",
          1454 => x"80",
          1455 => x"26",
          1456 => x"8a",
          1457 => x"a0",
          1458 => x"c4",
          1459 => x"74",
          1460 => x"e0",
          1461 => x"ff",
          1462 => x"d0",
          1463 => x"ff",
          1464 => x"90",
          1465 => x"38",
          1466 => x"81",
          1467 => x"54",
          1468 => x"81",
          1469 => x"78",
          1470 => x"38",
          1471 => x"13",
          1472 => x"79",
          1473 => x"56",
          1474 => x"a0",
          1475 => x"38",
          1476 => x"84",
          1477 => x"56",
          1478 => x"81",
          1479 => x"ba",
          1480 => x"3d",
          1481 => x"70",
          1482 => x"0c",
          1483 => x"56",
          1484 => x"2e",
          1485 => x"fe",
          1486 => x"15",
          1487 => x"70",
          1488 => x"73",
          1489 => x"a6",
          1490 => x"73",
          1491 => x"a0",
          1492 => x"a0",
          1493 => x"38",
          1494 => x"80",
          1495 => x"89",
          1496 => x"e1",
          1497 => x"ba",
          1498 => x"3d",
          1499 => x"58",
          1500 => x"78",
          1501 => x"55",
          1502 => x"fe",
          1503 => x"0b",
          1504 => x"0c",
          1505 => x"04",
          1506 => x"7b",
          1507 => x"80",
          1508 => x"77",
          1509 => x"56",
          1510 => x"a0",
          1511 => x"06",
          1512 => x"15",
          1513 => x"70",
          1514 => x"73",
          1515 => x"38",
          1516 => x"80",
          1517 => x"b0",
          1518 => x"38",
          1519 => x"80",
          1520 => x"26",
          1521 => x"8a",
          1522 => x"a0",
          1523 => x"c4",
          1524 => x"74",
          1525 => x"e0",
          1526 => x"ff",
          1527 => x"d0",
          1528 => x"ff",
          1529 => x"90",
          1530 => x"38",
          1531 => x"81",
          1532 => x"54",
          1533 => x"81",
          1534 => x"78",
          1535 => x"38",
          1536 => x"13",
          1537 => x"79",
          1538 => x"56",
          1539 => x"a0",
          1540 => x"38",
          1541 => x"84",
          1542 => x"56",
          1543 => x"81",
          1544 => x"ba",
          1545 => x"3d",
          1546 => x"70",
          1547 => x"0c",
          1548 => x"56",
          1549 => x"2e",
          1550 => x"fe",
          1551 => x"15",
          1552 => x"70",
          1553 => x"73",
          1554 => x"a6",
          1555 => x"73",
          1556 => x"a0",
          1557 => x"a0",
          1558 => x"38",
          1559 => x"80",
          1560 => x"89",
          1561 => x"e1",
          1562 => x"ba",
          1563 => x"3d",
          1564 => x"58",
          1565 => x"78",
          1566 => x"55",
          1567 => x"fe",
          1568 => x"0b",
          1569 => x"0c",
          1570 => x"04",
          1571 => x"3f",
          1572 => x"08",
          1573 => x"84",
          1574 => x"04",
          1575 => x"73",
          1576 => x"26",
          1577 => x"10",
          1578 => x"cc",
          1579 => x"08",
          1580 => x"e4",
          1581 => x"3f",
          1582 => x"04",
          1583 => x"51",
          1584 => x"83",
          1585 => x"83",
          1586 => x"ef",
          1587 => x"3d",
          1588 => x"cf",
          1589 => x"9d",
          1590 => x"0d",
          1591 => x"bc",
          1592 => x"3f",
          1593 => x"04",
          1594 => x"51",
          1595 => x"83",
          1596 => x"83",
          1597 => x"ee",
          1598 => x"3d",
          1599 => x"cf",
          1600 => x"f1",
          1601 => x"0d",
          1602 => x"a4",
          1603 => x"3f",
          1604 => x"04",
          1605 => x"51",
          1606 => x"83",
          1607 => x"83",
          1608 => x"ee",
          1609 => x"3d",
          1610 => x"d0",
          1611 => x"c5",
          1612 => x"0d",
          1613 => x"84",
          1614 => x"3f",
          1615 => x"04",
          1616 => x"51",
          1617 => x"83",
          1618 => x"83",
          1619 => x"ee",
          1620 => x"3d",
          1621 => x"d1",
          1622 => x"99",
          1623 => x"0d",
          1624 => x"d0",
          1625 => x"3f",
          1626 => x"04",
          1627 => x"51",
          1628 => x"83",
          1629 => x"83",
          1630 => x"ed",
          1631 => x"3d",
          1632 => x"d2",
          1633 => x"ed",
          1634 => x"0d",
          1635 => x"8c",
          1636 => x"3f",
          1637 => x"04",
          1638 => x"66",
          1639 => x"80",
          1640 => x"5b",
          1641 => x"79",
          1642 => x"07",
          1643 => x"57",
          1644 => x"57",
          1645 => x"26",
          1646 => x"57",
          1647 => x"70",
          1648 => x"51",
          1649 => x"74",
          1650 => x"81",
          1651 => x"8c",
          1652 => x"58",
          1653 => x"3f",
          1654 => x"08",
          1655 => x"8c",
          1656 => x"80",
          1657 => x"51",
          1658 => x"3f",
          1659 => x"78",
          1660 => x"7b",
          1661 => x"2a",
          1662 => x"57",
          1663 => x"80",
          1664 => x"87",
          1665 => x"08",
          1666 => x"e7",
          1667 => x"38",
          1668 => x"87",
          1669 => x"f5",
          1670 => x"ba",
          1671 => x"83",
          1672 => x"78",
          1673 => x"98",
          1674 => x"3f",
          1675 => x"8c",
          1676 => x"0d",
          1677 => x"8c",
          1678 => x"98",
          1679 => x"ba",
          1680 => x"96",
          1681 => x"54",
          1682 => x"75",
          1683 => x"82",
          1684 => x"84",
          1685 => x"57",
          1686 => x"08",
          1687 => x"7a",
          1688 => x"2e",
          1689 => x"74",
          1690 => x"57",
          1691 => x"87",
          1692 => x"51",
          1693 => x"84",
          1694 => x"52",
          1695 => x"a7",
          1696 => x"8c",
          1697 => x"d2",
          1698 => x"52",
          1699 => x"51",
          1700 => x"ff",
          1701 => x"3d",
          1702 => x"84",
          1703 => x"33",
          1704 => x"58",
          1705 => x"52",
          1706 => x"ec",
          1707 => x"8c",
          1708 => x"76",
          1709 => x"38",
          1710 => x"8a",
          1711 => x"ba",
          1712 => x"3d",
          1713 => x"04",
          1714 => x"56",
          1715 => x"54",
          1716 => x"53",
          1717 => x"51",
          1718 => x"ba",
          1719 => x"ba",
          1720 => x"3d",
          1721 => x"3d",
          1722 => x"63",
          1723 => x"80",
          1724 => x"73",
          1725 => x"41",
          1726 => x"5f",
          1727 => x"80",
          1728 => x"38",
          1729 => x"d2",
          1730 => x"fe",
          1731 => x"cc",
          1732 => x"3f",
          1733 => x"79",
          1734 => x"7c",
          1735 => x"ed",
          1736 => x"2e",
          1737 => x"73",
          1738 => x"7a",
          1739 => x"38",
          1740 => x"83",
          1741 => x"dd",
          1742 => x"14",
          1743 => x"08",
          1744 => x"51",
          1745 => x"78",
          1746 => x"38",
          1747 => x"51",
          1748 => x"80",
          1749 => x"27",
          1750 => x"75",
          1751 => x"55",
          1752 => x"72",
          1753 => x"38",
          1754 => x"53",
          1755 => x"83",
          1756 => x"74",
          1757 => x"81",
          1758 => x"57",
          1759 => x"88",
          1760 => x"74",
          1761 => x"38",
          1762 => x"08",
          1763 => x"eb",
          1764 => x"16",
          1765 => x"26",
          1766 => x"d2",
          1767 => x"d5",
          1768 => x"79",
          1769 => x"80",
          1770 => x"3f",
          1771 => x"08",
          1772 => x"98",
          1773 => x"76",
          1774 => x"ee",
          1775 => x"2e",
          1776 => x"7b",
          1777 => x"78",
          1778 => x"38",
          1779 => x"ba",
          1780 => x"3d",
          1781 => x"d2",
          1782 => x"ae",
          1783 => x"84",
          1784 => x"53",
          1785 => x"eb",
          1786 => x"74",
          1787 => x"38",
          1788 => x"83",
          1789 => x"dc",
          1790 => x"14",
          1791 => x"08",
          1792 => x"51",
          1793 => x"73",
          1794 => x"c0",
          1795 => x"53",
          1796 => x"df",
          1797 => x"52",
          1798 => x"51",
          1799 => x"82",
          1800 => x"f0",
          1801 => x"a0",
          1802 => x"3f",
          1803 => x"dd",
          1804 => x"39",
          1805 => x"51",
          1806 => x"84",
          1807 => x"f0",
          1808 => x"a0",
          1809 => x"3f",
          1810 => x"fd",
          1811 => x"18",
          1812 => x"27",
          1813 => x"08",
          1814 => x"c4",
          1815 => x"3f",
          1816 => x"d5",
          1817 => x"54",
          1818 => x"84",
          1819 => x"26",
          1820 => x"d8",
          1821 => x"f0",
          1822 => x"51",
          1823 => x"81",
          1824 => x"91",
          1825 => x"e3",
          1826 => x"8c",
          1827 => x"06",
          1828 => x"72",
          1829 => x"ec",
          1830 => x"72",
          1831 => x"09",
          1832 => x"e0",
          1833 => x"fc",
          1834 => x"51",
          1835 => x"84",
          1836 => x"98",
          1837 => x"2c",
          1838 => x"70",
          1839 => x"32",
          1840 => x"72",
          1841 => x"07",
          1842 => x"58",
          1843 => x"53",
          1844 => x"fd",
          1845 => x"51",
          1846 => x"84",
          1847 => x"98",
          1848 => x"2c",
          1849 => x"70",
          1850 => x"32",
          1851 => x"72",
          1852 => x"07",
          1853 => x"58",
          1854 => x"53",
          1855 => x"ff",
          1856 => x"b9",
          1857 => x"84",
          1858 => x"8f",
          1859 => x"fe",
          1860 => x"c0",
          1861 => x"53",
          1862 => x"81",
          1863 => x"3f",
          1864 => x"51",
          1865 => x"80",
          1866 => x"3f",
          1867 => x"70",
          1868 => x"52",
          1869 => x"38",
          1870 => x"70",
          1871 => x"52",
          1872 => x"38",
          1873 => x"70",
          1874 => x"52",
          1875 => x"38",
          1876 => x"70",
          1877 => x"52",
          1878 => x"38",
          1879 => x"70",
          1880 => x"52",
          1881 => x"38",
          1882 => x"70",
          1883 => x"52",
          1884 => x"38",
          1885 => x"70",
          1886 => x"52",
          1887 => x"72",
          1888 => x"06",
          1889 => x"38",
          1890 => x"84",
          1891 => x"81",
          1892 => x"3f",
          1893 => x"51",
          1894 => x"80",
          1895 => x"3f",
          1896 => x"84",
          1897 => x"81",
          1898 => x"3f",
          1899 => x"51",
          1900 => x"80",
          1901 => x"3f",
          1902 => x"81",
          1903 => x"80",
          1904 => x"cb",
          1905 => x"9b",
          1906 => x"d3",
          1907 => x"de",
          1908 => x"9b",
          1909 => x"87",
          1910 => x"06",
          1911 => x"80",
          1912 => x"38",
          1913 => x"51",
          1914 => x"83",
          1915 => x"9b",
          1916 => x"51",
          1917 => x"72",
          1918 => x"81",
          1919 => x"71",
          1920 => x"f0",
          1921 => x"39",
          1922 => x"8a",
          1923 => x"9c",
          1924 => x"3f",
          1925 => x"fe",
          1926 => x"2a",
          1927 => x"51",
          1928 => x"2e",
          1929 => x"ff",
          1930 => x"51",
          1931 => x"83",
          1932 => x"9a",
          1933 => x"51",
          1934 => x"72",
          1935 => x"81",
          1936 => x"71",
          1937 => x"94",
          1938 => x"39",
          1939 => x"c6",
          1940 => x"c4",
          1941 => x"3f",
          1942 => x"ba",
          1943 => x"2a",
          1944 => x"51",
          1945 => x"2e",
          1946 => x"ff",
          1947 => x"51",
          1948 => x"83",
          1949 => x"9a",
          1950 => x"51",
          1951 => x"72",
          1952 => x"81",
          1953 => x"71",
          1954 => x"b8",
          1955 => x"39",
          1956 => x"80",
          1957 => x"ff",
          1958 => x"98",
          1959 => x"52",
          1960 => x"b6",
          1961 => x"ba",
          1962 => x"ff",
          1963 => x"40",
          1964 => x"2e",
          1965 => x"83",
          1966 => x"e3",
          1967 => x"3d",
          1968 => x"e0",
          1969 => x"3f",
          1970 => x"f8",
          1971 => x"7e",
          1972 => x"3f",
          1973 => x"ef",
          1974 => x"81",
          1975 => x"59",
          1976 => x"82",
          1977 => x"81",
          1978 => x"38",
          1979 => x"06",
          1980 => x"2e",
          1981 => x"67",
          1982 => x"79",
          1983 => x"dc",
          1984 => x"5c",
          1985 => x"09",
          1986 => x"38",
          1987 => x"33",
          1988 => x"a0",
          1989 => x"80",
          1990 => x"26",
          1991 => x"90",
          1992 => x"84",
          1993 => x"52",
          1994 => x"3f",
          1995 => x"08",
          1996 => x"08",
          1997 => x"7b",
          1998 => x"e8",
          1999 => x"ba",
          2000 => x"38",
          2001 => x"5e",
          2002 => x"83",
          2003 => x"1c",
          2004 => x"06",
          2005 => x"7c",
          2006 => x"9a",
          2007 => x"7b",
          2008 => x"dd",
          2009 => x"52",
          2010 => x"92",
          2011 => x"8c",
          2012 => x"ba",
          2013 => x"2e",
          2014 => x"84",
          2015 => x"48",
          2016 => x"80",
          2017 => x"93",
          2018 => x"8c",
          2019 => x"06",
          2020 => x"80",
          2021 => x"38",
          2022 => x"08",
          2023 => x"3f",
          2024 => x"08",
          2025 => x"f3",
          2026 => x"a5",
          2027 => x"7a",
          2028 => x"8f",
          2029 => x"24",
          2030 => x"7a",
          2031 => x"ee",
          2032 => x"80",
          2033 => x"e4",
          2034 => x"d5",
          2035 => x"f2",
          2036 => x"ba",
          2037 => x"56",
          2038 => x"54",
          2039 => x"53",
          2040 => x"52",
          2041 => x"ae",
          2042 => x"8c",
          2043 => x"8c",
          2044 => x"30",
          2045 => x"80",
          2046 => x"5b",
          2047 => x"7a",
          2048 => x"38",
          2049 => x"7a",
          2050 => x"80",
          2051 => x"81",
          2052 => x"ff",
          2053 => x"7a",
          2054 => x"7f",
          2055 => x"81",
          2056 => x"7c",
          2057 => x"61",
          2058 => x"f2",
          2059 => x"81",
          2060 => x"83",
          2061 => x"d3",
          2062 => x"48",
          2063 => x"80",
          2064 => x"e8",
          2065 => x"0b",
          2066 => x"33",
          2067 => x"06",
          2068 => x"fd",
          2069 => x"53",
          2070 => x"52",
          2071 => x"51",
          2072 => x"3f",
          2073 => x"08",
          2074 => x"81",
          2075 => x"83",
          2076 => x"84",
          2077 => x"80",
          2078 => x"51",
          2079 => x"3f",
          2080 => x"08",
          2081 => x"38",
          2082 => x"08",
          2083 => x"3f",
          2084 => x"ef",
          2085 => x"81",
          2086 => x"59",
          2087 => x"09",
          2088 => x"d3",
          2089 => x"84",
          2090 => x"82",
          2091 => x"82",
          2092 => x"83",
          2093 => x"83",
          2094 => x"80",
          2095 => x"51",
          2096 => x"67",
          2097 => x"79",
          2098 => x"90",
          2099 => x"63",
          2100 => x"33",
          2101 => x"89",
          2102 => x"38",
          2103 => x"83",
          2104 => x"5a",
          2105 => x"83",
          2106 => x"df",
          2107 => x"3d",
          2108 => x"83",
          2109 => x"7e",
          2110 => x"3f",
          2111 => x"52",
          2112 => x"51",
          2113 => x"3f",
          2114 => x"08",
          2115 => x"81",
          2116 => x"38",
          2117 => x"3d",
          2118 => x"fb",
          2119 => x"d6",
          2120 => x"d1",
          2121 => x"81",
          2122 => x"fe",
          2123 => x"d6",
          2124 => x"55",
          2125 => x"54",
          2126 => x"d6",
          2127 => x"51",
          2128 => x"fd",
          2129 => x"8c",
          2130 => x"f5",
          2131 => x"3f",
          2132 => x"81",
          2133 => x"bf",
          2134 => x"e5",
          2135 => x"95",
          2136 => x"39",
          2137 => x"51",
          2138 => x"80",
          2139 => x"83",
          2140 => x"de",
          2141 => x"f3",
          2142 => x"39",
          2143 => x"84",
          2144 => x"80",
          2145 => x"80",
          2146 => x"8c",
          2147 => x"fa",
          2148 => x"52",
          2149 => x"51",
          2150 => x"68",
          2151 => x"84",
          2152 => x"80",
          2153 => x"38",
          2154 => x"08",
          2155 => x"f8",
          2156 => x"3f",
          2157 => x"b8",
          2158 => x"11",
          2159 => x"05",
          2160 => x"3f",
          2161 => x"08",
          2162 => x"f5",
          2163 => x"83",
          2164 => x"d0",
          2165 => x"59",
          2166 => x"3d",
          2167 => x"53",
          2168 => x"51",
          2169 => x"84",
          2170 => x"80",
          2171 => x"38",
          2172 => x"f0",
          2173 => x"80",
          2174 => x"88",
          2175 => x"8c",
          2176 => x"38",
          2177 => x"08",
          2178 => x"83",
          2179 => x"cf",
          2180 => x"d5",
          2181 => x"80",
          2182 => x"51",
          2183 => x"7e",
          2184 => x"59",
          2185 => x"f9",
          2186 => x"9f",
          2187 => x"38",
          2188 => x"70",
          2189 => x"39",
          2190 => x"f4",
          2191 => x"80",
          2192 => x"c0",
          2193 => x"8c",
          2194 => x"f8",
          2195 => x"3d",
          2196 => x"53",
          2197 => x"51",
          2198 => x"84",
          2199 => x"86",
          2200 => x"59",
          2201 => x"78",
          2202 => x"c0",
          2203 => x"3f",
          2204 => x"08",
          2205 => x"52",
          2206 => x"a9",
          2207 => x"7e",
          2208 => x"ae",
          2209 => x"38",
          2210 => x"87",
          2211 => x"82",
          2212 => x"59",
          2213 => x"3d",
          2214 => x"53",
          2215 => x"51",
          2216 => x"84",
          2217 => x"80",
          2218 => x"38",
          2219 => x"fc",
          2220 => x"80",
          2221 => x"d0",
          2222 => x"8c",
          2223 => x"f8",
          2224 => x"3d",
          2225 => x"53",
          2226 => x"51",
          2227 => x"84",
          2228 => x"80",
          2229 => x"38",
          2230 => x"51",
          2231 => x"68",
          2232 => x"78",
          2233 => x"8d",
          2234 => x"33",
          2235 => x"5c",
          2236 => x"2e",
          2237 => x"55",
          2238 => x"33",
          2239 => x"83",
          2240 => x"ce",
          2241 => x"66",
          2242 => x"19",
          2243 => x"59",
          2244 => x"3d",
          2245 => x"53",
          2246 => x"51",
          2247 => x"84",
          2248 => x"80",
          2249 => x"38",
          2250 => x"fc",
          2251 => x"80",
          2252 => x"d4",
          2253 => x"8c",
          2254 => x"f7",
          2255 => x"3d",
          2256 => x"53",
          2257 => x"51",
          2258 => x"84",
          2259 => x"80",
          2260 => x"38",
          2261 => x"51",
          2262 => x"68",
          2263 => x"27",
          2264 => x"65",
          2265 => x"81",
          2266 => x"7c",
          2267 => x"05",
          2268 => x"b8",
          2269 => x"11",
          2270 => x"05",
          2271 => x"3f",
          2272 => x"08",
          2273 => x"b9",
          2274 => x"fe",
          2275 => x"ff",
          2276 => x"e7",
          2277 => x"ba",
          2278 => x"38",
          2279 => x"54",
          2280 => x"84",
          2281 => x"3f",
          2282 => x"08",
          2283 => x"52",
          2284 => x"f1",
          2285 => x"7e",
          2286 => x"ae",
          2287 => x"38",
          2288 => x"84",
          2289 => x"81",
          2290 => x"39",
          2291 => x"80",
          2292 => x"79",
          2293 => x"05",
          2294 => x"fe",
          2295 => x"ff",
          2296 => x"e7",
          2297 => x"ba",
          2298 => x"2e",
          2299 => x"68",
          2300 => x"db",
          2301 => x"34",
          2302 => x"49",
          2303 => x"fc",
          2304 => x"80",
          2305 => x"80",
          2306 => x"8c",
          2307 => x"38",
          2308 => x"b8",
          2309 => x"11",
          2310 => x"05",
          2311 => x"3f",
          2312 => x"08",
          2313 => x"99",
          2314 => x"fe",
          2315 => x"ff",
          2316 => x"e6",
          2317 => x"ba",
          2318 => x"2e",
          2319 => x"b8",
          2320 => x"11",
          2321 => x"05",
          2322 => x"3f",
          2323 => x"08",
          2324 => x"ba",
          2325 => x"83",
          2326 => x"cb",
          2327 => x"67",
          2328 => x"7a",
          2329 => x"65",
          2330 => x"70",
          2331 => x"0c",
          2332 => x"f5",
          2333 => x"d9",
          2334 => x"c5",
          2335 => x"ff",
          2336 => x"87",
          2337 => x"ba",
          2338 => x"3d",
          2339 => x"52",
          2340 => x"3f",
          2341 => x"ba",
          2342 => x"78",
          2343 => x"3f",
          2344 => x"08",
          2345 => x"99",
          2346 => x"8c",
          2347 => x"ec",
          2348 => x"39",
          2349 => x"84",
          2350 => x"80",
          2351 => x"c8",
          2352 => x"8c",
          2353 => x"83",
          2354 => x"5a",
          2355 => x"83",
          2356 => x"f2",
          2357 => x"b8",
          2358 => x"11",
          2359 => x"05",
          2360 => x"3f",
          2361 => x"08",
          2362 => x"f3",
          2363 => x"79",
          2364 => x"8a",
          2365 => x"cc",
          2366 => x"3d",
          2367 => x"53",
          2368 => x"51",
          2369 => x"84",
          2370 => x"80",
          2371 => x"80",
          2372 => x"7a",
          2373 => x"38",
          2374 => x"90",
          2375 => x"70",
          2376 => x"2a",
          2377 => x"5f",
          2378 => x"2e",
          2379 => x"a0",
          2380 => x"88",
          2381 => x"a0",
          2382 => x"3f",
          2383 => x"54",
          2384 => x"52",
          2385 => x"9e",
          2386 => x"ac",
          2387 => x"3f",
          2388 => x"64",
          2389 => x"59",
          2390 => x"45",
          2391 => x"f0",
          2392 => x"80",
          2393 => x"9c",
          2394 => x"8c",
          2395 => x"f2",
          2396 => x"64",
          2397 => x"64",
          2398 => x"b8",
          2399 => x"11",
          2400 => x"05",
          2401 => x"3f",
          2402 => x"08",
          2403 => x"b1",
          2404 => x"02",
          2405 => x"22",
          2406 => x"05",
          2407 => x"45",
          2408 => x"f0",
          2409 => x"80",
          2410 => x"d8",
          2411 => x"8c",
          2412 => x"f2",
          2413 => x"5e",
          2414 => x"05",
          2415 => x"82",
          2416 => x"7d",
          2417 => x"fe",
          2418 => x"ff",
          2419 => x"e1",
          2420 => x"ba",
          2421 => x"b9",
          2422 => x"39",
          2423 => x"fc",
          2424 => x"80",
          2425 => x"a0",
          2426 => x"8c",
          2427 => x"81",
          2428 => x"5c",
          2429 => x"05",
          2430 => x"68",
          2431 => x"fb",
          2432 => x"3d",
          2433 => x"53",
          2434 => x"51",
          2435 => x"84",
          2436 => x"80",
          2437 => x"38",
          2438 => x"0c",
          2439 => x"05",
          2440 => x"f7",
          2441 => x"83",
          2442 => x"06",
          2443 => x"7b",
          2444 => x"98",
          2445 => x"83",
          2446 => x"7c",
          2447 => x"3f",
          2448 => x"7b",
          2449 => x"da",
          2450 => x"82",
          2451 => x"c4",
          2452 => x"3f",
          2453 => x"b8",
          2454 => x"11",
          2455 => x"05",
          2456 => x"3f",
          2457 => x"08",
          2458 => x"38",
          2459 => x"80",
          2460 => x"79",
          2461 => x"5b",
          2462 => x"f7",
          2463 => x"f3",
          2464 => x"7b",
          2465 => x"cf",
          2466 => x"d4",
          2467 => x"ea",
          2468 => x"91",
          2469 => x"80",
          2470 => x"83",
          2471 => x"49",
          2472 => x"83",
          2473 => x"d3",
          2474 => x"59",
          2475 => x"83",
          2476 => x"d3",
          2477 => x"59",
          2478 => x"83",
          2479 => x"59",
          2480 => x"a5",
          2481 => x"d8",
          2482 => x"8b",
          2483 => x"f0",
          2484 => x"3f",
          2485 => x"83",
          2486 => x"59",
          2487 => x"9b",
          2488 => x"dc",
          2489 => x"92",
          2490 => x"93",
          2491 => x"80",
          2492 => x"83",
          2493 => x"49",
          2494 => x"83",
          2495 => x"5e",
          2496 => x"9b",
          2497 => x"e4",
          2498 => x"ee",
          2499 => x"8e",
          2500 => x"80",
          2501 => x"83",
          2502 => x"49",
          2503 => x"83",
          2504 => x"5d",
          2505 => x"94",
          2506 => x"ec",
          2507 => x"ca",
          2508 => x"f8",
          2509 => x"05",
          2510 => x"39",
          2511 => x"08",
          2512 => x"fb",
          2513 => x"3d",
          2514 => x"84",
          2515 => x"87",
          2516 => x"70",
          2517 => x"87",
          2518 => x"74",
          2519 => x"3f",
          2520 => x"08",
          2521 => x"08",
          2522 => x"84",
          2523 => x"51",
          2524 => x"74",
          2525 => x"08",
          2526 => x"87",
          2527 => x"70",
          2528 => x"87",
          2529 => x"74",
          2530 => x"3f",
          2531 => x"08",
          2532 => x"08",
          2533 => x"84",
          2534 => x"51",
          2535 => x"74",
          2536 => x"08",
          2537 => x"8c",
          2538 => x"87",
          2539 => x"0c",
          2540 => x"0b",
          2541 => x"94",
          2542 => x"ec",
          2543 => x"eb",
          2544 => x"84",
          2545 => x"34",
          2546 => x"d5",
          2547 => x"3d",
          2548 => x"0c",
          2549 => x"84",
          2550 => x"56",
          2551 => x"89",
          2552 => x"87",
          2553 => x"51",
          2554 => x"83",
          2555 => x"83",
          2556 => x"c4",
          2557 => x"f2",
          2558 => x"52",
          2559 => x"3f",
          2560 => x"54",
          2561 => x"53",
          2562 => x"52",
          2563 => x"51",
          2564 => x"8d",
          2565 => x"f8",
          2566 => x"fb",
          2567 => x"70",
          2568 => x"80",
          2569 => x"74",
          2570 => x"83",
          2571 => x"70",
          2572 => x"52",
          2573 => x"2e",
          2574 => x"91",
          2575 => x"70",
          2576 => x"ff",
          2577 => x"55",
          2578 => x"f1",
          2579 => x"ff",
          2580 => x"a2",
          2581 => x"38",
          2582 => x"81",
          2583 => x"38",
          2584 => x"70",
          2585 => x"53",
          2586 => x"a0",
          2587 => x"81",
          2588 => x"2e",
          2589 => x"80",
          2590 => x"81",
          2591 => x"39",
          2592 => x"ff",
          2593 => x"70",
          2594 => x"81",
          2595 => x"81",
          2596 => x"32",
          2597 => x"80",
          2598 => x"52",
          2599 => x"80",
          2600 => x"80",
          2601 => x"05",
          2602 => x"76",
          2603 => x"70",
          2604 => x"0c",
          2605 => x"04",
          2606 => x"c4",
          2607 => x"2e",
          2608 => x"81",
          2609 => x"72",
          2610 => x"ff",
          2611 => x"54",
          2612 => x"e4",
          2613 => x"e0",
          2614 => x"55",
          2615 => x"53",
          2616 => x"09",
          2617 => x"f8",
          2618 => x"fc",
          2619 => x"53",
          2620 => x"38",
          2621 => x"ba",
          2622 => x"3d",
          2623 => x"3d",
          2624 => x"72",
          2625 => x"3f",
          2626 => x"08",
          2627 => x"38",
          2628 => x"8c",
          2629 => x"0d",
          2630 => x"0d",
          2631 => x"33",
          2632 => x"53",
          2633 => x"8b",
          2634 => x"38",
          2635 => x"ff",
          2636 => x"52",
          2637 => x"81",
          2638 => x"13",
          2639 => x"52",
          2640 => x"80",
          2641 => x"13",
          2642 => x"52",
          2643 => x"80",
          2644 => x"13",
          2645 => x"52",
          2646 => x"80",
          2647 => x"13",
          2648 => x"52",
          2649 => x"26",
          2650 => x"8a",
          2651 => x"87",
          2652 => x"e7",
          2653 => x"38",
          2654 => x"c0",
          2655 => x"72",
          2656 => x"98",
          2657 => x"13",
          2658 => x"98",
          2659 => x"13",
          2660 => x"98",
          2661 => x"13",
          2662 => x"98",
          2663 => x"13",
          2664 => x"98",
          2665 => x"13",
          2666 => x"98",
          2667 => x"87",
          2668 => x"0c",
          2669 => x"98",
          2670 => x"0b",
          2671 => x"9c",
          2672 => x"71",
          2673 => x"0c",
          2674 => x"04",
          2675 => x"7f",
          2676 => x"98",
          2677 => x"7d",
          2678 => x"98",
          2679 => x"7d",
          2680 => x"c0",
          2681 => x"5c",
          2682 => x"34",
          2683 => x"b4",
          2684 => x"83",
          2685 => x"c0",
          2686 => x"5c",
          2687 => x"34",
          2688 => x"ac",
          2689 => x"85",
          2690 => x"c0",
          2691 => x"5c",
          2692 => x"34",
          2693 => x"a4",
          2694 => x"88",
          2695 => x"c0",
          2696 => x"5a",
          2697 => x"23",
          2698 => x"79",
          2699 => x"06",
          2700 => x"ff",
          2701 => x"86",
          2702 => x"85",
          2703 => x"84",
          2704 => x"83",
          2705 => x"82",
          2706 => x"7d",
          2707 => x"06",
          2708 => x"f4",
          2709 => x"b2",
          2710 => x"0d",
          2711 => x"0d",
          2712 => x"33",
          2713 => x"2e",
          2714 => x"51",
          2715 => x"3f",
          2716 => x"08",
          2717 => x"98",
          2718 => x"71",
          2719 => x"81",
          2720 => x"72",
          2721 => x"38",
          2722 => x"8c",
          2723 => x"0d",
          2724 => x"80",
          2725 => x"84",
          2726 => x"98",
          2727 => x"2c",
          2728 => x"ff",
          2729 => x"06",
          2730 => x"51",
          2731 => x"3f",
          2732 => x"08",
          2733 => x"98",
          2734 => x"71",
          2735 => x"38",
          2736 => x"3d",
          2737 => x"54",
          2738 => x"2b",
          2739 => x"80",
          2740 => x"84",
          2741 => x"98",
          2742 => x"2c",
          2743 => x"ff",
          2744 => x"73",
          2745 => x"14",
          2746 => x"73",
          2747 => x"71",
          2748 => x"0c",
          2749 => x"04",
          2750 => x"02",
          2751 => x"83",
          2752 => x"70",
          2753 => x"53",
          2754 => x"80",
          2755 => x"38",
          2756 => x"94",
          2757 => x"2a",
          2758 => x"53",
          2759 => x"80",
          2760 => x"71",
          2761 => x"81",
          2762 => x"70",
          2763 => x"81",
          2764 => x"53",
          2765 => x"8a",
          2766 => x"2a",
          2767 => x"71",
          2768 => x"81",
          2769 => x"87",
          2770 => x"52",
          2771 => x"86",
          2772 => x"94",
          2773 => x"72",
          2774 => x"ba",
          2775 => x"3d",
          2776 => x"91",
          2777 => x"06",
          2778 => x"97",
          2779 => x"32",
          2780 => x"72",
          2781 => x"38",
          2782 => x"81",
          2783 => x"80",
          2784 => x"87",
          2785 => x"08",
          2786 => x"70",
          2787 => x"54",
          2788 => x"38",
          2789 => x"3d",
          2790 => x"05",
          2791 => x"70",
          2792 => x"52",
          2793 => x"f2",
          2794 => x"3d",
          2795 => x"3d",
          2796 => x"80",
          2797 => x"56",
          2798 => x"77",
          2799 => x"38",
          2800 => x"f2",
          2801 => x"81",
          2802 => x"57",
          2803 => x"2e",
          2804 => x"87",
          2805 => x"08",
          2806 => x"70",
          2807 => x"54",
          2808 => x"2e",
          2809 => x"91",
          2810 => x"06",
          2811 => x"e3",
          2812 => x"32",
          2813 => x"72",
          2814 => x"38",
          2815 => x"81",
          2816 => x"cf",
          2817 => x"ff",
          2818 => x"c0",
          2819 => x"70",
          2820 => x"38",
          2821 => x"90",
          2822 => x"0c",
          2823 => x"33",
          2824 => x"ff",
          2825 => x"84",
          2826 => x"88",
          2827 => x"71",
          2828 => x"81",
          2829 => x"70",
          2830 => x"81",
          2831 => x"53",
          2832 => x"c1",
          2833 => x"2a",
          2834 => x"71",
          2835 => x"b5",
          2836 => x"94",
          2837 => x"96",
          2838 => x"06",
          2839 => x"70",
          2840 => x"39",
          2841 => x"87",
          2842 => x"08",
          2843 => x"8a",
          2844 => x"70",
          2845 => x"ab",
          2846 => x"9e",
          2847 => x"f2",
          2848 => x"c0",
          2849 => x"83",
          2850 => x"87",
          2851 => x"08",
          2852 => x"0c",
          2853 => x"98",
          2854 => x"d4",
          2855 => x"9e",
          2856 => x"f2",
          2857 => x"c0",
          2858 => x"83",
          2859 => x"87",
          2860 => x"08",
          2861 => x"0c",
          2862 => x"b0",
          2863 => x"e4",
          2864 => x"9e",
          2865 => x"f2",
          2866 => x"c0",
          2867 => x"83",
          2868 => x"87",
          2869 => x"08",
          2870 => x"0c",
          2871 => x"c0",
          2872 => x"f4",
          2873 => x"9e",
          2874 => x"f2",
          2875 => x"c0",
          2876 => x"52",
          2877 => x"fc",
          2878 => x"9e",
          2879 => x"f3",
          2880 => x"c0",
          2881 => x"83",
          2882 => x"87",
          2883 => x"08",
          2884 => x"0c",
          2885 => x"f3",
          2886 => x"0b",
          2887 => x"90",
          2888 => x"80",
          2889 => x"52",
          2890 => x"fb",
          2891 => x"f3",
          2892 => x"0b",
          2893 => x"90",
          2894 => x"80",
          2895 => x"52",
          2896 => x"2e",
          2897 => x"52",
          2898 => x"8e",
          2899 => x"87",
          2900 => x"08",
          2901 => x"0a",
          2902 => x"52",
          2903 => x"83",
          2904 => x"71",
          2905 => x"34",
          2906 => x"c0",
          2907 => x"70",
          2908 => x"06",
          2909 => x"70",
          2910 => x"38",
          2911 => x"83",
          2912 => x"80",
          2913 => x"9e",
          2914 => x"a0",
          2915 => x"51",
          2916 => x"80",
          2917 => x"81",
          2918 => x"f3",
          2919 => x"0b",
          2920 => x"90",
          2921 => x"80",
          2922 => x"52",
          2923 => x"2e",
          2924 => x"52",
          2925 => x"92",
          2926 => x"87",
          2927 => x"08",
          2928 => x"80",
          2929 => x"52",
          2930 => x"83",
          2931 => x"71",
          2932 => x"34",
          2933 => x"c0",
          2934 => x"70",
          2935 => x"06",
          2936 => x"70",
          2937 => x"38",
          2938 => x"83",
          2939 => x"80",
          2940 => x"9e",
          2941 => x"81",
          2942 => x"51",
          2943 => x"80",
          2944 => x"81",
          2945 => x"f3",
          2946 => x"0b",
          2947 => x"90",
          2948 => x"c0",
          2949 => x"52",
          2950 => x"2e",
          2951 => x"52",
          2952 => x"96",
          2953 => x"87",
          2954 => x"08",
          2955 => x"06",
          2956 => x"70",
          2957 => x"38",
          2958 => x"83",
          2959 => x"87",
          2960 => x"08",
          2961 => x"70",
          2962 => x"51",
          2963 => x"98",
          2964 => x"87",
          2965 => x"08",
          2966 => x"06",
          2967 => x"70",
          2968 => x"38",
          2969 => x"83",
          2970 => x"87",
          2971 => x"08",
          2972 => x"70",
          2973 => x"51",
          2974 => x"9a",
          2975 => x"87",
          2976 => x"08",
          2977 => x"51",
          2978 => x"80",
          2979 => x"81",
          2980 => x"f3",
          2981 => x"c0",
          2982 => x"87",
          2983 => x"83",
          2984 => x"83",
          2985 => x"81",
          2986 => x"39",
          2987 => x"83",
          2988 => x"ff",
          2989 => x"83",
          2990 => x"54",
          2991 => x"38",
          2992 => x"51",
          2993 => x"83",
          2994 => x"55",
          2995 => x"38",
          2996 => x"33",
          2997 => x"d1",
          2998 => x"90",
          2999 => x"85",
          3000 => x"f3",
          3001 => x"74",
          3002 => x"83",
          3003 => x"54",
          3004 => x"38",
          3005 => x"33",
          3006 => x"b3",
          3007 => x"9b",
          3008 => x"84",
          3009 => x"f3",
          3010 => x"74",
          3011 => x"83",
          3012 => x"56",
          3013 => x"38",
          3014 => x"33",
          3015 => x"b1",
          3016 => x"94",
          3017 => x"83",
          3018 => x"f3",
          3019 => x"75",
          3020 => x"83",
          3021 => x"54",
          3022 => x"38",
          3023 => x"51",
          3024 => x"83",
          3025 => x"52",
          3026 => x"51",
          3027 => x"3f",
          3028 => x"08",
          3029 => x"ec",
          3030 => x"ae",
          3031 => x"f8",
          3032 => x"da",
          3033 => x"b5",
          3034 => x"da",
          3035 => x"85",
          3036 => x"fc",
          3037 => x"da",
          3038 => x"b5",
          3039 => x"f3",
          3040 => x"bd",
          3041 => x"75",
          3042 => x"3f",
          3043 => x"08",
          3044 => x"29",
          3045 => x"54",
          3046 => x"8c",
          3047 => x"da",
          3048 => x"b4",
          3049 => x"f3",
          3050 => x"74",
          3051 => x"83",
          3052 => x"55",
          3053 => x"8a",
          3054 => x"3f",
          3055 => x"04",
          3056 => x"08",
          3057 => x"c0",
          3058 => x"c9",
          3059 => x"ba",
          3060 => x"84",
          3061 => x"71",
          3062 => x"84",
          3063 => x"52",
          3064 => x"51",
          3065 => x"3f",
          3066 => x"f4",
          3067 => x"0d",
          3068 => x"84",
          3069 => x"84",
          3070 => x"51",
          3071 => x"84",
          3072 => x"bd",
          3073 => x"76",
          3074 => x"54",
          3075 => x"08",
          3076 => x"c4",
          3077 => x"f2",
          3078 => x"8e",
          3079 => x"80",
          3080 => x"38",
          3081 => x"83",
          3082 => x"c0",
          3083 => x"d9",
          3084 => x"c1",
          3085 => x"f0",
          3086 => x"d9",
          3087 => x"b3",
          3088 => x"f2",
          3089 => x"83",
          3090 => x"ff",
          3091 => x"83",
          3092 => x"52",
          3093 => x"51",
          3094 => x"3f",
          3095 => x"51",
          3096 => x"83",
          3097 => x"52",
          3098 => x"51",
          3099 => x"3f",
          3100 => x"08",
          3101 => x"c0",
          3102 => x"c8",
          3103 => x"ba",
          3104 => x"84",
          3105 => x"71",
          3106 => x"84",
          3107 => x"52",
          3108 => x"51",
          3109 => x"3f",
          3110 => x"33",
          3111 => x"2e",
          3112 => x"fe",
          3113 => x"db",
          3114 => x"bf",
          3115 => x"f3",
          3116 => x"73",
          3117 => x"84",
          3118 => x"39",
          3119 => x"51",
          3120 => x"3f",
          3121 => x"33",
          3122 => x"2e",
          3123 => x"d6",
          3124 => x"8c",
          3125 => x"9d",
          3126 => x"94",
          3127 => x"80",
          3128 => x"38",
          3129 => x"dc",
          3130 => x"bf",
          3131 => x"f3",
          3132 => x"73",
          3133 => x"a9",
          3134 => x"83",
          3135 => x"52",
          3136 => x"51",
          3137 => x"3f",
          3138 => x"33",
          3139 => x"2e",
          3140 => x"d2",
          3141 => x"9c",
          3142 => x"dc",
          3143 => x"b1",
          3144 => x"f3",
          3145 => x"74",
          3146 => x"e3",
          3147 => x"83",
          3148 => x"52",
          3149 => x"51",
          3150 => x"3f",
          3151 => x"33",
          3152 => x"2e",
          3153 => x"cd",
          3154 => x"d8",
          3155 => x"dc",
          3156 => x"52",
          3157 => x"51",
          3158 => x"3f",
          3159 => x"33",
          3160 => x"2e",
          3161 => x"c7",
          3162 => x"d0",
          3163 => x"d4",
          3164 => x"52",
          3165 => x"51",
          3166 => x"3f",
          3167 => x"33",
          3168 => x"2e",
          3169 => x"c1",
          3170 => x"c8",
          3171 => x"cc",
          3172 => x"52",
          3173 => x"51",
          3174 => x"3f",
          3175 => x"33",
          3176 => x"2e",
          3177 => x"c1",
          3178 => x"e0",
          3179 => x"e4",
          3180 => x"52",
          3181 => x"51",
          3182 => x"3f",
          3183 => x"33",
          3184 => x"2e",
          3185 => x"c1",
          3186 => x"e8",
          3187 => x"ec",
          3188 => x"52",
          3189 => x"51",
          3190 => x"3f",
          3191 => x"33",
          3192 => x"2e",
          3193 => x"c1",
          3194 => x"98",
          3195 => x"9a",
          3196 => x"a0",
          3197 => x"fd",
          3198 => x"8e",
          3199 => x"80",
          3200 => x"38",
          3201 => x"3d",
          3202 => x"05",
          3203 => x"85",
          3204 => x"71",
          3205 => x"c3",
          3206 => x"71",
          3207 => x"de",
          3208 => x"af",
          3209 => x"3d",
          3210 => x"de",
          3211 => x"af",
          3212 => x"3d",
          3213 => x"de",
          3214 => x"af",
          3215 => x"3d",
          3216 => x"de",
          3217 => x"af",
          3218 => x"3d",
          3219 => x"de",
          3220 => x"af",
          3221 => x"3d",
          3222 => x"de",
          3223 => x"af",
          3224 => x"3d",
          3225 => x"88",
          3226 => x"80",
          3227 => x"96",
          3228 => x"83",
          3229 => x"87",
          3230 => x"0c",
          3231 => x"0d",
          3232 => x"ad",
          3233 => x"5a",
          3234 => x"58",
          3235 => x"f3",
          3236 => x"82",
          3237 => x"84",
          3238 => x"80",
          3239 => x"3d",
          3240 => x"83",
          3241 => x"54",
          3242 => x"52",
          3243 => x"d2",
          3244 => x"ba",
          3245 => x"2e",
          3246 => x"51",
          3247 => x"84",
          3248 => x"81",
          3249 => x"80",
          3250 => x"8c",
          3251 => x"38",
          3252 => x"08",
          3253 => x"18",
          3254 => x"74",
          3255 => x"70",
          3256 => x"07",
          3257 => x"55",
          3258 => x"2e",
          3259 => x"ff",
          3260 => x"f3",
          3261 => x"11",
          3262 => x"82",
          3263 => x"84",
          3264 => x"8f",
          3265 => x"2e",
          3266 => x"84",
          3267 => x"a9",
          3268 => x"83",
          3269 => x"ff",
          3270 => x"78",
          3271 => x"81",
          3272 => x"76",
          3273 => x"c0",
          3274 => x"51",
          3275 => x"3f",
          3276 => x"56",
          3277 => x"08",
          3278 => x"52",
          3279 => x"51",
          3280 => x"3f",
          3281 => x"ba",
          3282 => x"3d",
          3283 => x"3d",
          3284 => x"08",
          3285 => x"71",
          3286 => x"33",
          3287 => x"57",
          3288 => x"81",
          3289 => x"0b",
          3290 => x"56",
          3291 => x"10",
          3292 => x"05",
          3293 => x"54",
          3294 => x"3f",
          3295 => x"08",
          3296 => x"73",
          3297 => x"8f",
          3298 => x"8c",
          3299 => x"84",
          3300 => x"73",
          3301 => x"88",
          3302 => x"2e",
          3303 => x"16",
          3304 => x"06",
          3305 => x"76",
          3306 => x"80",
          3307 => x"ba",
          3308 => x"3d",
          3309 => x"1a",
          3310 => x"ff",
          3311 => x"ff",
          3312 => x"c7",
          3313 => x"ba",
          3314 => x"2e",
          3315 => x"1b",
          3316 => x"76",
          3317 => x"3f",
          3318 => x"08",
          3319 => x"54",
          3320 => x"c9",
          3321 => x"70",
          3322 => x"57",
          3323 => x"27",
          3324 => x"ff",
          3325 => x"33",
          3326 => x"76",
          3327 => x"e6",
          3328 => x"70",
          3329 => x"55",
          3330 => x"2e",
          3331 => x"fe",
          3332 => x"75",
          3333 => x"80",
          3334 => x"59",
          3335 => x"39",
          3336 => x"8c",
          3337 => x"f3",
          3338 => x"56",
          3339 => x"3f",
          3340 => x"08",
          3341 => x"83",
          3342 => x"53",
          3343 => x"77",
          3344 => x"cc",
          3345 => x"8c",
          3346 => x"ba",
          3347 => x"ff",
          3348 => x"84",
          3349 => x"55",
          3350 => x"ba",
          3351 => x"9d",
          3352 => x"8c",
          3353 => x"70",
          3354 => x"80",
          3355 => x"53",
          3356 => x"16",
          3357 => x"52",
          3358 => x"8e",
          3359 => x"2e",
          3360 => x"ff",
          3361 => x"0b",
          3362 => x"0c",
          3363 => x"04",
          3364 => x"b5",
          3365 => x"3d",
          3366 => x"08",
          3367 => x"80",
          3368 => x"34",
          3369 => x"33",
          3370 => x"08",
          3371 => x"9e",
          3372 => x"f3",
          3373 => x"56",
          3374 => x"82",
          3375 => x"80",
          3376 => x"38",
          3377 => x"06",
          3378 => x"90",
          3379 => x"80",
          3380 => x"38",
          3381 => x"3d",
          3382 => x"51",
          3383 => x"84",
          3384 => x"98",
          3385 => x"2c",
          3386 => x"ff",
          3387 => x"79",
          3388 => x"84",
          3389 => x"70",
          3390 => x"98",
          3391 => x"c4",
          3392 => x"2b",
          3393 => x"71",
          3394 => x"70",
          3395 => x"de",
          3396 => x"08",
          3397 => x"52",
          3398 => x"46",
          3399 => x"5c",
          3400 => x"74",
          3401 => x"cd",
          3402 => x"27",
          3403 => x"75",
          3404 => x"29",
          3405 => x"05",
          3406 => x"57",
          3407 => x"24",
          3408 => x"75",
          3409 => x"82",
          3410 => x"80",
          3411 => x"dc",
          3412 => x"57",
          3413 => x"91",
          3414 => x"d8",
          3415 => x"70",
          3416 => x"78",
          3417 => x"95",
          3418 => x"2e",
          3419 => x"84",
          3420 => x"81",
          3421 => x"2e",
          3422 => x"81",
          3423 => x"2b",
          3424 => x"84",
          3425 => x"70",
          3426 => x"97",
          3427 => x"2c",
          3428 => x"2b",
          3429 => x"11",
          3430 => x"5f",
          3431 => x"57",
          3432 => x"2e",
          3433 => x"76",
          3434 => x"34",
          3435 => x"81",
          3436 => x"ba",
          3437 => x"80",
          3438 => x"80",
          3439 => x"98",
          3440 => x"ff",
          3441 => x"41",
          3442 => x"80",
          3443 => x"10",
          3444 => x"2b",
          3445 => x"0b",
          3446 => x"16",
          3447 => x"77",
          3448 => x"38",
          3449 => x"15",
          3450 => x"33",
          3451 => x"61",
          3452 => x"38",
          3453 => x"ff",
          3454 => x"f2",
          3455 => x"76",
          3456 => x"ab",
          3457 => x"39",
          3458 => x"b2",
          3459 => x"76",
          3460 => x"76",
          3461 => x"34",
          3462 => x"c4",
          3463 => x"34",
          3464 => x"62",
          3465 => x"26",
          3466 => x"74",
          3467 => x"c3",
          3468 => x"76",
          3469 => x"de",
          3470 => x"7f",
          3471 => x"84",
          3472 => x"80",
          3473 => x"c4",
          3474 => x"84",
          3475 => x"56",
          3476 => x"fd",
          3477 => x"d5",
          3478 => x"88",
          3479 => x"90",
          3480 => x"d0",
          3481 => x"57",
          3482 => x"d0",
          3483 => x"39",
          3484 => x"33",
          3485 => x"06",
          3486 => x"33",
          3487 => x"75",
          3488 => x"d6",
          3489 => x"f0",
          3490 => x"15",
          3491 => x"d1",
          3492 => x"16",
          3493 => x"55",
          3494 => x"3f",
          3495 => x"7c",
          3496 => x"da",
          3497 => x"10",
          3498 => x"05",
          3499 => x"59",
          3500 => x"38",
          3501 => x"cc",
          3502 => x"34",
          3503 => x"33",
          3504 => x"33",
          3505 => x"80",
          3506 => x"84",
          3507 => x"52",
          3508 => x"b5",
          3509 => x"d5",
          3510 => x"a0",
          3511 => x"90",
          3512 => x"f0",
          3513 => x"51",
          3514 => x"3f",
          3515 => x"33",
          3516 => x"7a",
          3517 => x"34",
          3518 => x"06",
          3519 => x"38",
          3520 => x"a6",
          3521 => x"84",
          3522 => x"fb",
          3523 => x"8a",
          3524 => x"f0",
          3525 => x"8d",
          3526 => x"10",
          3527 => x"a4",
          3528 => x"08",
          3529 => x"8e",
          3530 => x"08",
          3531 => x"2e",
          3532 => x"75",
          3533 => x"f2",
          3534 => x"8c",
          3535 => x"cc",
          3536 => x"8c",
          3537 => x"06",
          3538 => x"75",
          3539 => x"ff",
          3540 => x"84",
          3541 => x"84",
          3542 => x"56",
          3543 => x"2e",
          3544 => x"84",
          3545 => x"52",
          3546 => x"b4",
          3547 => x"d5",
          3548 => x"a0",
          3549 => x"f8",
          3550 => x"f0",
          3551 => x"51",
          3552 => x"3f",
          3553 => x"33",
          3554 => x"74",
          3555 => x"34",
          3556 => x"06",
          3557 => x"84",
          3558 => x"70",
          3559 => x"84",
          3560 => x"5b",
          3561 => x"79",
          3562 => x"38",
          3563 => x"08",
          3564 => x"57",
          3565 => x"d0",
          3566 => x"70",
          3567 => x"ff",
          3568 => x"84",
          3569 => x"70",
          3570 => x"84",
          3571 => x"5a",
          3572 => x"78",
          3573 => x"38",
          3574 => x"08",
          3575 => x"57",
          3576 => x"d0",
          3577 => x"70",
          3578 => x"ff",
          3579 => x"84",
          3580 => x"70",
          3581 => x"84",
          3582 => x"5a",
          3583 => x"76",
          3584 => x"38",
          3585 => x"84",
          3586 => x"84",
          3587 => x"56",
          3588 => x"2e",
          3589 => x"ff",
          3590 => x"84",
          3591 => x"75",
          3592 => x"98",
          3593 => x"ff",
          3594 => x"5a",
          3595 => x"80",
          3596 => x"d5",
          3597 => x"a0",
          3598 => x"b4",
          3599 => x"d0",
          3600 => x"2b",
          3601 => x"84",
          3602 => x"5a",
          3603 => x"74",
          3604 => x"86",
          3605 => x"f0",
          3606 => x"51",
          3607 => x"3f",
          3608 => x"0a",
          3609 => x"0a",
          3610 => x"2c",
          3611 => x"33",
          3612 => x"74",
          3613 => x"e2",
          3614 => x"f0",
          3615 => x"51",
          3616 => x"3f",
          3617 => x"0a",
          3618 => x"0a",
          3619 => x"2c",
          3620 => x"33",
          3621 => x"7a",
          3622 => x"b9",
          3623 => x"39",
          3624 => x"81",
          3625 => x"34",
          3626 => x"08",
          3627 => x"51",
          3628 => x"3f",
          3629 => x"0a",
          3630 => x"0a",
          3631 => x"2c",
          3632 => x"33",
          3633 => x"75",
          3634 => x"e6",
          3635 => x"58",
          3636 => x"78",
          3637 => x"f0",
          3638 => x"33",
          3639 => x"90",
          3640 => x"80",
          3641 => x"80",
          3642 => x"98",
          3643 => x"cc",
          3644 => x"55",
          3645 => x"ff",
          3646 => x"b6",
          3647 => x"d0",
          3648 => x"80",
          3649 => x"38",
          3650 => x"08",
          3651 => x"ff",
          3652 => x"84",
          3653 => x"ff",
          3654 => x"84",
          3655 => x"76",
          3656 => x"55",
          3657 => x"d1",
          3658 => x"05",
          3659 => x"34",
          3660 => x"08",
          3661 => x"ff",
          3662 => x"84",
          3663 => x"7b",
          3664 => x"3f",
          3665 => x"08",
          3666 => x"58",
          3667 => x"38",
          3668 => x"33",
          3669 => x"2e",
          3670 => x"83",
          3671 => x"70",
          3672 => x"f3",
          3673 => x"08",
          3674 => x"74",
          3675 => x"75",
          3676 => x"fc",
          3677 => x"a4",
          3678 => x"70",
          3679 => x"80",
          3680 => x"84",
          3681 => x"7b",
          3682 => x"fc",
          3683 => x"10",
          3684 => x"05",
          3685 => x"41",
          3686 => x"ad",
          3687 => x"f8",
          3688 => x"80",
          3689 => x"83",
          3690 => x"58",
          3691 => x"8b",
          3692 => x"0b",
          3693 => x"34",
          3694 => x"d1",
          3695 => x"84",
          3696 => x"b4",
          3697 => x"84",
          3698 => x"55",
          3699 => x"b6",
          3700 => x"f0",
          3701 => x"51",
          3702 => x"3f",
          3703 => x"08",
          3704 => x"ff",
          3705 => x"84",
          3706 => x"52",
          3707 => x"ae",
          3708 => x"d1",
          3709 => x"05",
          3710 => x"d1",
          3711 => x"81",
          3712 => x"74",
          3713 => x"d2",
          3714 => x"9f",
          3715 => x"0b",
          3716 => x"34",
          3717 => x"d1",
          3718 => x"be",
          3719 => x"34",
          3720 => x"1d",
          3721 => x"d0",
          3722 => x"80",
          3723 => x"84",
          3724 => x"52",
          3725 => x"ae",
          3726 => x"d5",
          3727 => x"a0",
          3728 => x"ac",
          3729 => x"f0",
          3730 => x"51",
          3731 => x"3f",
          3732 => x"33",
          3733 => x"7c",
          3734 => x"34",
          3735 => x"06",
          3736 => x"38",
          3737 => x"51",
          3738 => x"3f",
          3739 => x"d1",
          3740 => x"0b",
          3741 => x"34",
          3742 => x"8c",
          3743 => x"0d",
          3744 => x"d0",
          3745 => x"ff",
          3746 => x"7a",
          3747 => x"ca",
          3748 => x"cc",
          3749 => x"59",
          3750 => x"cc",
          3751 => x"58",
          3752 => x"d0",
          3753 => x"f0",
          3754 => x"51",
          3755 => x"3f",
          3756 => x"33",
          3757 => x"70",
          3758 => x"d1",
          3759 => x"52",
          3760 => x"76",
          3761 => x"38",
          3762 => x"08",
          3763 => x"ff",
          3764 => x"84",
          3765 => x"70",
          3766 => x"98",
          3767 => x"cc",
          3768 => x"59",
          3769 => x"24",
          3770 => x"84",
          3771 => x"52",
          3772 => x"ac",
          3773 => x"81",
          3774 => x"81",
          3775 => x"70",
          3776 => x"d1",
          3777 => x"51",
          3778 => x"24",
          3779 => x"84",
          3780 => x"52",
          3781 => x"ac",
          3782 => x"81",
          3783 => x"81",
          3784 => x"70",
          3785 => x"d1",
          3786 => x"51",
          3787 => x"25",
          3788 => x"f3",
          3789 => x"16",
          3790 => x"33",
          3791 => x"d5",
          3792 => x"76",
          3793 => x"ac",
          3794 => x"81",
          3795 => x"81",
          3796 => x"70",
          3797 => x"d1",
          3798 => x"57",
          3799 => x"25",
          3800 => x"7b",
          3801 => x"17",
          3802 => x"84",
          3803 => x"52",
          3804 => x"ff",
          3805 => x"75",
          3806 => x"29",
          3807 => x"05",
          3808 => x"84",
          3809 => x"43",
          3810 => x"76",
          3811 => x"38",
          3812 => x"84",
          3813 => x"70",
          3814 => x"58",
          3815 => x"2e",
          3816 => x"84",
          3817 => x"55",
          3818 => x"ae",
          3819 => x"2b",
          3820 => x"57",
          3821 => x"24",
          3822 => x"16",
          3823 => x"81",
          3824 => x"81",
          3825 => x"81",
          3826 => x"70",
          3827 => x"d1",
          3828 => x"57",
          3829 => x"25",
          3830 => x"18",
          3831 => x"d1",
          3832 => x"81",
          3833 => x"05",
          3834 => x"33",
          3835 => x"d1",
          3836 => x"76",
          3837 => x"38",
          3838 => x"75",
          3839 => x"34",
          3840 => x"d1",
          3841 => x"81",
          3842 => x"81",
          3843 => x"70",
          3844 => x"81",
          3845 => x"58",
          3846 => x"76",
          3847 => x"38",
          3848 => x"70",
          3849 => x"81",
          3850 => x"57",
          3851 => x"25",
          3852 => x"84",
          3853 => x"52",
          3854 => x"aa",
          3855 => x"81",
          3856 => x"81",
          3857 => x"70",
          3858 => x"d1",
          3859 => x"57",
          3860 => x"25",
          3861 => x"84",
          3862 => x"52",
          3863 => x"aa",
          3864 => x"81",
          3865 => x"81",
          3866 => x"70",
          3867 => x"d1",
          3868 => x"57",
          3869 => x"24",
          3870 => x"f0",
          3871 => x"f3",
          3872 => x"75",
          3873 => x"9d",
          3874 => x"ff",
          3875 => x"84",
          3876 => x"84",
          3877 => x"84",
          3878 => x"81",
          3879 => x"05",
          3880 => x"7b",
          3881 => x"c4",
          3882 => x"cc",
          3883 => x"d0",
          3884 => x"74",
          3885 => x"c8",
          3886 => x"f0",
          3887 => x"51",
          3888 => x"3f",
          3889 => x"08",
          3890 => x"ff",
          3891 => x"84",
          3892 => x"52",
          3893 => x"a9",
          3894 => x"d1",
          3895 => x"05",
          3896 => x"d1",
          3897 => x"81",
          3898 => x"c7",
          3899 => x"80",
          3900 => x"84",
          3901 => x"83",
          3902 => x"84",
          3903 => x"85",
          3904 => x"83",
          3905 => x"77",
          3906 => x"80",
          3907 => x"d5",
          3908 => x"7b",
          3909 => x"52",
          3910 => x"d4",
          3911 => x"80",
          3912 => x"80",
          3913 => x"98",
          3914 => x"cc",
          3915 => x"57",
          3916 => x"da",
          3917 => x"d0",
          3918 => x"2b",
          3919 => x"79",
          3920 => x"5d",
          3921 => x"75",
          3922 => x"8e",
          3923 => x"39",
          3924 => x"08",
          3925 => x"fc",
          3926 => x"a4",
          3927 => x"76",
          3928 => x"bb",
          3929 => x"84",
          3930 => x"75",
          3931 => x"38",
          3932 => x"f3",
          3933 => x"f3",
          3934 => x"74",
          3935 => x"d4",
          3936 => x"81",
          3937 => x"83",
          3938 => x"51",
          3939 => x"3f",
          3940 => x"f3",
          3941 => x"3d",
          3942 => x"5f",
          3943 => x"74",
          3944 => x"b8",
          3945 => x"0c",
          3946 => x"18",
          3947 => x"80",
          3948 => x"38",
          3949 => x"75",
          3950 => x"ee",
          3951 => x"8c",
          3952 => x"cc",
          3953 => x"8c",
          3954 => x"06",
          3955 => x"75",
          3956 => x"ff",
          3957 => x"93",
          3958 => x"cc",
          3959 => x"d0",
          3960 => x"5d",
          3961 => x"f2",
          3962 => x"d5",
          3963 => x"88",
          3964 => x"fc",
          3965 => x"f0",
          3966 => x"51",
          3967 => x"3f",
          3968 => x"08",
          3969 => x"ff",
          3970 => x"84",
          3971 => x"ff",
          3972 => x"84",
          3973 => x"79",
          3974 => x"55",
          3975 => x"7c",
          3976 => x"84",
          3977 => x"80",
          3978 => x"cc",
          3979 => x"ba",
          3980 => x"3d",
          3981 => x"51",
          3982 => x"3f",
          3983 => x"08",
          3984 => x"34",
          3985 => x"08",
          3986 => x"81",
          3987 => x"52",
          3988 => x"aa",
          3989 => x"1d",
          3990 => x"06",
          3991 => x"33",
          3992 => x"33",
          3993 => x"56",
          3994 => x"f1",
          3995 => x"d5",
          3996 => x"88",
          3997 => x"f8",
          3998 => x"f0",
          3999 => x"51",
          4000 => x"3f",
          4001 => x"08",
          4002 => x"ff",
          4003 => x"84",
          4004 => x"ff",
          4005 => x"84",
          4006 => x"76",
          4007 => x"55",
          4008 => x"51",
          4009 => x"3f",
          4010 => x"08",
          4011 => x"34",
          4012 => x"08",
          4013 => x"81",
          4014 => x"52",
          4015 => x"a9",
          4016 => x"1d",
          4017 => x"06",
          4018 => x"33",
          4019 => x"33",
          4020 => x"58",
          4021 => x"f0",
          4022 => x"d5",
          4023 => x"88",
          4024 => x"8c",
          4025 => x"f0",
          4026 => x"51",
          4027 => x"3f",
          4028 => x"08",
          4029 => x"ff",
          4030 => x"84",
          4031 => x"ff",
          4032 => x"84",
          4033 => x"60",
          4034 => x"55",
          4035 => x"51",
          4036 => x"3f",
          4037 => x"33",
          4038 => x"87",
          4039 => x"f3",
          4040 => x"19",
          4041 => x"5c",
          4042 => x"a0",
          4043 => x"8c",
          4044 => x"83",
          4045 => x"70",
          4046 => x"f3",
          4047 => x"08",
          4048 => x"74",
          4049 => x"d5",
          4050 => x"7b",
          4051 => x"ff",
          4052 => x"83",
          4053 => x"81",
          4054 => x"ff",
          4055 => x"93",
          4056 => x"f2",
          4057 => x"f3",
          4058 => x"b1",
          4059 => x"fe",
          4060 => x"76",
          4061 => x"75",
          4062 => x"8f",
          4063 => x"f8",
          4064 => x"51",
          4065 => x"3f",
          4066 => x"08",
          4067 => x"c2",
          4068 => x"84",
          4069 => x"80",
          4070 => x"cc",
          4071 => x"ba",
          4072 => x"3d",
          4073 => x"53",
          4074 => x"ba",
          4075 => x"81",
          4076 => x"84",
          4077 => x"82",
          4078 => x"ba",
          4079 => x"3d",
          4080 => x"f3",
          4081 => x"80",
          4082 => x"51",
          4083 => x"3f",
          4084 => x"08",
          4085 => x"8c",
          4086 => x"09",
          4087 => x"ee",
          4088 => x"8c",
          4089 => x"a6",
          4090 => x"ba",
          4091 => x"80",
          4092 => x"8c",
          4093 => x"e3",
          4094 => x"8c",
          4095 => x"70",
          4096 => x"80",
          4097 => x"81",
          4098 => x"f3",
          4099 => x"10",
          4100 => x"a4",
          4101 => x"58",
          4102 => x"74",
          4103 => x"76",
          4104 => x"fc",
          4105 => x"a4",
          4106 => x"70",
          4107 => x"80",
          4108 => x"84",
          4109 => x"75",
          4110 => x"fc",
          4111 => x"10",
          4112 => x"05",
          4113 => x"40",
          4114 => x"38",
          4115 => x"81",
          4116 => x"57",
          4117 => x"83",
          4118 => x"75",
          4119 => x"81",
          4120 => x"38",
          4121 => x"38",
          4122 => x"76",
          4123 => x"74",
          4124 => x"f8",
          4125 => x"fc",
          4126 => x"70",
          4127 => x"5b",
          4128 => x"27",
          4129 => x"80",
          4130 => x"fc",
          4131 => x"39",
          4132 => x"d4",
          4133 => x"f3",
          4134 => x"82",
          4135 => x"06",
          4136 => x"05",
          4137 => x"54",
          4138 => x"80",
          4139 => x"84",
          4140 => x"75",
          4141 => x"fc",
          4142 => x"10",
          4143 => x"05",
          4144 => x"40",
          4145 => x"2e",
          4146 => x"ff",
          4147 => x"83",
          4148 => x"fe",
          4149 => x"83",
          4150 => x"f1",
          4151 => x"e1",
          4152 => x"9f",
          4153 => x"e7",
          4154 => x"e4",
          4155 => x"0d",
          4156 => x"05",
          4157 => x"05",
          4158 => x"33",
          4159 => x"83",
          4160 => x"38",
          4161 => x"81",
          4162 => x"73",
          4163 => x"38",
          4164 => x"82",
          4165 => x"a3",
          4166 => x"87",
          4167 => x"70",
          4168 => x"56",
          4169 => x"79",
          4170 => x"38",
          4171 => x"bc",
          4172 => x"f9",
          4173 => x"83",
          4174 => x"83",
          4175 => x"70",
          4176 => x"90",
          4177 => x"88",
          4178 => x"07",
          4179 => x"56",
          4180 => x"77",
          4181 => x"80",
          4182 => x"05",
          4183 => x"73",
          4184 => x"55",
          4185 => x"26",
          4186 => x"78",
          4187 => x"83",
          4188 => x"84",
          4189 => x"79",
          4190 => x"55",
          4191 => x"e0",
          4192 => x"74",
          4193 => x"05",
          4194 => x"13",
          4195 => x"38",
          4196 => x"04",
          4197 => x"80",
          4198 => x"bc",
          4199 => x"10",
          4200 => x"bd",
          4201 => x"29",
          4202 => x"5b",
          4203 => x"59",
          4204 => x"80",
          4205 => x"80",
          4206 => x"ff",
          4207 => x"ff",
          4208 => x"ff",
          4209 => x"ba",
          4210 => x"ff",
          4211 => x"75",
          4212 => x"5d",
          4213 => x"5b",
          4214 => x"26",
          4215 => x"74",
          4216 => x"56",
          4217 => x"06",
          4218 => x"06",
          4219 => x"06",
          4220 => x"ff",
          4221 => x"ff",
          4222 => x"29",
          4223 => x"57",
          4224 => x"74",
          4225 => x"38",
          4226 => x"33",
          4227 => x"05",
          4228 => x"1b",
          4229 => x"83",
          4230 => x"80",
          4231 => x"38",
          4232 => x"53",
          4233 => x"fe",
          4234 => x"73",
          4235 => x"55",
          4236 => x"b8",
          4237 => x"81",
          4238 => x"e8",
          4239 => x"a0",
          4240 => x"a3",
          4241 => x"84",
          4242 => x"70",
          4243 => x"84",
          4244 => x"70",
          4245 => x"83",
          4246 => x"70",
          4247 => x"5b",
          4248 => x"56",
          4249 => x"78",
          4250 => x"38",
          4251 => x"06",
          4252 => x"06",
          4253 => x"18",
          4254 => x"79",
          4255 => x"bb",
          4256 => x"83",
          4257 => x"80",
          4258 => x"bd",
          4259 => x"b8",
          4260 => x"2b",
          4261 => x"07",
          4262 => x"07",
          4263 => x"7f",
          4264 => x"5b",
          4265 => x"fd",
          4266 => x"be",
          4267 => x"e6",
          4268 => x"bc",
          4269 => x"ff",
          4270 => x"10",
          4271 => x"bd",
          4272 => x"29",
          4273 => x"a0",
          4274 => x"57",
          4275 => x"5f",
          4276 => x"80",
          4277 => x"b8",
          4278 => x"81",
          4279 => x"b7",
          4280 => x"81",
          4281 => x"f9",
          4282 => x"83",
          4283 => x"7c",
          4284 => x"05",
          4285 => x"5f",
          4286 => x"5e",
          4287 => x"26",
          4288 => x"7a",
          4289 => x"7d",
          4290 => x"53",
          4291 => x"06",
          4292 => x"06",
          4293 => x"7d",
          4294 => x"06",
          4295 => x"06",
          4296 => x"58",
          4297 => x"5d",
          4298 => x"26",
          4299 => x"75",
          4300 => x"73",
          4301 => x"83",
          4302 => x"79",
          4303 => x"76",
          4304 => x"7b",
          4305 => x"fb",
          4306 => x"78",
          4307 => x"56",
          4308 => x"fb",
          4309 => x"ee",
          4310 => x"80",
          4311 => x"ff",
          4312 => x"86",
          4313 => x"53",
          4314 => x"80",
          4315 => x"ee",
          4316 => x"8a",
          4317 => x"76",
          4318 => x"74",
          4319 => x"80",
          4320 => x"8a",
          4321 => x"75",
          4322 => x"34",
          4323 => x"81",
          4324 => x"fa",
          4325 => x"90",
          4326 => x"08",
          4327 => x"f8",
          4328 => x"81",
          4329 => x"06",
          4330 => x"55",
          4331 => x"73",
          4332 => x"ff",
          4333 => x"07",
          4334 => x"75",
          4335 => x"87",
          4336 => x"77",
          4337 => x"51",
          4338 => x"8c",
          4339 => x"73",
          4340 => x"06",
          4341 => x"72",
          4342 => x"d0",
          4343 => x"80",
          4344 => x"84",
          4345 => x"87",
          4346 => x"84",
          4347 => x"84",
          4348 => x"04",
          4349 => x"02",
          4350 => x"02",
          4351 => x"05",
          4352 => x"ff",
          4353 => x"56",
          4354 => x"79",
          4355 => x"38",
          4356 => x"33",
          4357 => x"33",
          4358 => x"33",
          4359 => x"12",
          4360 => x"80",
          4361 => x"ba",
          4362 => x"57",
          4363 => x"29",
          4364 => x"ff",
          4365 => x"f8",
          4366 => x"57",
          4367 => x"81",
          4368 => x"38",
          4369 => x"22",
          4370 => x"74",
          4371 => x"23",
          4372 => x"33",
          4373 => x"81",
          4374 => x"81",
          4375 => x"5b",
          4376 => x"26",
          4377 => x"ff",
          4378 => x"83",
          4379 => x"83",
          4380 => x"70",
          4381 => x"06",
          4382 => x"33",
          4383 => x"79",
          4384 => x"89",
          4385 => x"80",
          4386 => x"29",
          4387 => x"54",
          4388 => x"26",
          4389 => x"98",
          4390 => x"54",
          4391 => x"13",
          4392 => x"16",
          4393 => x"81",
          4394 => x"75",
          4395 => x"57",
          4396 => x"54",
          4397 => x"73",
          4398 => x"73",
          4399 => x"a1",
          4400 => x"b8",
          4401 => x"de",
          4402 => x"a0",
          4403 => x"14",
          4404 => x"70",
          4405 => x"34",
          4406 => x"9f",
          4407 => x"eb",
          4408 => x"fe",
          4409 => x"56",
          4410 => x"ba",
          4411 => x"78",
          4412 => x"77",
          4413 => x"06",
          4414 => x"73",
          4415 => x"38",
          4416 => x"81",
          4417 => x"80",
          4418 => x"29",
          4419 => x"75",
          4420 => x"a0",
          4421 => x"a3",
          4422 => x"81",
          4423 => x"81",
          4424 => x"71",
          4425 => x"5c",
          4426 => x"79",
          4427 => x"84",
          4428 => x"54",
          4429 => x"33",
          4430 => x"88",
          4431 => x"70",
          4432 => x"34",
          4433 => x"05",
          4434 => x"70",
          4435 => x"34",
          4436 => x"b8",
          4437 => x"b7",
          4438 => x"71",
          4439 => x"5c",
          4440 => x"75",
          4441 => x"80",
          4442 => x"ba",
          4443 => x"3d",
          4444 => x"83",
          4445 => x"83",
          4446 => x"70",
          4447 => x"06",
          4448 => x"33",
          4449 => x"73",
          4450 => x"f9",
          4451 => x"2e",
          4452 => x"78",
          4453 => x"ff",
          4454 => x"bc",
          4455 => x"72",
          4456 => x"81",
          4457 => x"38",
          4458 => x"81",
          4459 => x"80",
          4460 => x"29",
          4461 => x"11",
          4462 => x"54",
          4463 => x"fe",
          4464 => x"f9",
          4465 => x"98",
          4466 => x"76",
          4467 => x"56",
          4468 => x"e0",
          4469 => x"75",
          4470 => x"57",
          4471 => x"53",
          4472 => x"fe",
          4473 => x"0b",
          4474 => x"34",
          4475 => x"81",
          4476 => x"ff",
          4477 => x"d8",
          4478 => x"39",
          4479 => x"b8",
          4480 => x"56",
          4481 => x"83",
          4482 => x"33",
          4483 => x"88",
          4484 => x"34",
          4485 => x"33",
          4486 => x"39",
          4487 => x"76",
          4488 => x"9f",
          4489 => x"51",
          4490 => x"9b",
          4491 => x"10",
          4492 => x"05",
          4493 => x"04",
          4494 => x"33",
          4495 => x"27",
          4496 => x"83",
          4497 => x"80",
          4498 => x"8c",
          4499 => x"0d",
          4500 => x"83",
          4501 => x"83",
          4502 => x"70",
          4503 => x"54",
          4504 => x"2e",
          4505 => x"12",
          4506 => x"f9",
          4507 => x"0b",
          4508 => x"0c",
          4509 => x"04",
          4510 => x"33",
          4511 => x"70",
          4512 => x"2c",
          4513 => x"55",
          4514 => x"83",
          4515 => x"de",
          4516 => x"bc",
          4517 => x"84",
          4518 => x"ff",
          4519 => x"51",
          4520 => x"83",
          4521 => x"72",
          4522 => x"34",
          4523 => x"ba",
          4524 => x"3d",
          4525 => x"f9",
          4526 => x"73",
          4527 => x"70",
          4528 => x"06",
          4529 => x"55",
          4530 => x"bd",
          4531 => x"84",
          4532 => x"86",
          4533 => x"83",
          4534 => x"72",
          4535 => x"80",
          4536 => x"55",
          4537 => x"74",
          4538 => x"70",
          4539 => x"f9",
          4540 => x"0b",
          4541 => x"0c",
          4542 => x"04",
          4543 => x"f9",
          4544 => x"f9",
          4545 => x"b7",
          4546 => x"05",
          4547 => x"75",
          4548 => x"38",
          4549 => x"70",
          4550 => x"34",
          4551 => x"ff",
          4552 => x"8f",
          4553 => x"70",
          4554 => x"38",
          4555 => x"83",
          4556 => x"51",
          4557 => x"83",
          4558 => x"70",
          4559 => x"71",
          4560 => x"f0",
          4561 => x"84",
          4562 => x"52",
          4563 => x"80",
          4564 => x"81",
          4565 => x"80",
          4566 => x"f9",
          4567 => x"0b",
          4568 => x"0c",
          4569 => x"04",
          4570 => x"33",
          4571 => x"90",
          4572 => x"83",
          4573 => x"80",
          4574 => x"8c",
          4575 => x"0d",
          4576 => x"b8",
          4577 => x"07",
          4578 => x"f9",
          4579 => x"39",
          4580 => x"33",
          4581 => x"86",
          4582 => x"83",
          4583 => x"d7",
          4584 => x"0b",
          4585 => x"34",
          4586 => x"ba",
          4587 => x"3d",
          4588 => x"f9",
          4589 => x"fc",
          4590 => x"51",
          4591 => x"b8",
          4592 => x"39",
          4593 => x"33",
          4594 => x"70",
          4595 => x"34",
          4596 => x"83",
          4597 => x"81",
          4598 => x"07",
          4599 => x"f9",
          4600 => x"93",
          4601 => x"b8",
          4602 => x"06",
          4603 => x"70",
          4604 => x"34",
          4605 => x"83",
          4606 => x"81",
          4607 => x"07",
          4608 => x"f9",
          4609 => x"ef",
          4610 => x"b8",
          4611 => x"06",
          4612 => x"f9",
          4613 => x"df",
          4614 => x"b8",
          4615 => x"06",
          4616 => x"51",
          4617 => x"b8",
          4618 => x"39",
          4619 => x"33",
          4620 => x"b0",
          4621 => x"83",
          4622 => x"fe",
          4623 => x"f9",
          4624 => x"ef",
          4625 => x"07",
          4626 => x"f9",
          4627 => x"a7",
          4628 => x"b8",
          4629 => x"06",
          4630 => x"51",
          4631 => x"b8",
          4632 => x"39",
          4633 => x"33",
          4634 => x"a0",
          4635 => x"83",
          4636 => x"fe",
          4637 => x"f9",
          4638 => x"8f",
          4639 => x"83",
          4640 => x"fd",
          4641 => x"f9",
          4642 => x"fa",
          4643 => x"51",
          4644 => x"b8",
          4645 => x"39",
          4646 => x"02",
          4647 => x"02",
          4648 => x"c3",
          4649 => x"f9",
          4650 => x"f9",
          4651 => x"f9",
          4652 => x"b8",
          4653 => x"41",
          4654 => x"59",
          4655 => x"82",
          4656 => x"82",
          4657 => x"78",
          4658 => x"82",
          4659 => x"b8",
          4660 => x"0b",
          4661 => x"34",
          4662 => x"bc",
          4663 => x"f9",
          4664 => x"83",
          4665 => x"8f",
          4666 => x"78",
          4667 => x"81",
          4668 => x"80",
          4669 => x"82",
          4670 => x"84",
          4671 => x"82",
          4672 => x"bc",
          4673 => x"83",
          4674 => x"82",
          4675 => x"ba",
          4676 => x"84",
          4677 => x"57",
          4678 => x"33",
          4679 => x"fe",
          4680 => x"54",
          4681 => x"52",
          4682 => x"51",
          4683 => x"3f",
          4684 => x"82",
          4685 => x"84",
          4686 => x"7a",
          4687 => x"34",
          4688 => x"ba",
          4689 => x"f9",
          4690 => x"3d",
          4691 => x"0b",
          4692 => x"34",
          4693 => x"b8",
          4694 => x"0b",
          4695 => x"34",
          4696 => x"f9",
          4697 => x"0b",
          4698 => x"23",
          4699 => x"33",
          4700 => x"8e",
          4701 => x"b9",
          4702 => x"79",
          4703 => x"7c",
          4704 => x"83",
          4705 => x"ff",
          4706 => x"80",
          4707 => x"8d",
          4708 => x"79",
          4709 => x"38",
          4710 => x"b9",
          4711 => x"22",
          4712 => x"e3",
          4713 => x"80",
          4714 => x"1a",
          4715 => x"06",
          4716 => x"33",
          4717 => x"78",
          4718 => x"38",
          4719 => x"51",
          4720 => x"3f",
          4721 => x"82",
          4722 => x"84",
          4723 => x"7a",
          4724 => x"34",
          4725 => x"ba",
          4726 => x"f9",
          4727 => x"3d",
          4728 => x"0b",
          4729 => x"34",
          4730 => x"b8",
          4731 => x"0b",
          4732 => x"34",
          4733 => x"f9",
          4734 => x"0b",
          4735 => x"23",
          4736 => x"51",
          4737 => x"3f",
          4738 => x"08",
          4739 => x"fc",
          4740 => x"f6",
          4741 => x"83",
          4742 => x"ff",
          4743 => x"78",
          4744 => x"08",
          4745 => x"38",
          4746 => x"19",
          4747 => x"e4",
          4748 => x"ff",
          4749 => x"19",
          4750 => x"06",
          4751 => x"39",
          4752 => x"7a",
          4753 => x"a7",
          4754 => x"b8",
          4755 => x"f9",
          4756 => x"f9",
          4757 => x"71",
          4758 => x"a3",
          4759 => x"83",
          4760 => x"53",
          4761 => x"71",
          4762 => x"70",
          4763 => x"06",
          4764 => x"33",
          4765 => x"55",
          4766 => x"81",
          4767 => x"38",
          4768 => x"81",
          4769 => x"89",
          4770 => x"38",
          4771 => x"83",
          4772 => x"88",
          4773 => x"38",
          4774 => x"33",
          4775 => x"33",
          4776 => x"33",
          4777 => x"05",
          4778 => x"84",
          4779 => x"33",
          4780 => x"80",
          4781 => x"b8",
          4782 => x"f9",
          4783 => x"f9",
          4784 => x"71",
          4785 => x"5a",
          4786 => x"83",
          4787 => x"34",
          4788 => x"33",
          4789 => x"16",
          4790 => x"f9",
          4791 => x"a3",
          4792 => x"34",
          4793 => x"33",
          4794 => x"06",
          4795 => x"22",
          4796 => x"33",
          4797 => x"11",
          4798 => x"55",
          4799 => x"b8",
          4800 => x"de",
          4801 => x"18",
          4802 => x"06",
          4803 => x"78",
          4804 => x"38",
          4805 => x"33",
          4806 => x"ea",
          4807 => x"53",
          4808 => x"bd",
          4809 => x"83",
          4810 => x"80",
          4811 => x"84",
          4812 => x"57",
          4813 => x"80",
          4814 => x"0b",
          4815 => x"0c",
          4816 => x"04",
          4817 => x"97",
          4818 => x"24",
          4819 => x"75",
          4820 => x"81",
          4821 => x"38",
          4822 => x"51",
          4823 => x"80",
          4824 => x"bd",
          4825 => x"39",
          4826 => x"15",
          4827 => x"b8",
          4828 => x"74",
          4829 => x"2e",
          4830 => x"fe",
          4831 => x"53",
          4832 => x"51",
          4833 => x"81",
          4834 => x"ff",
          4835 => x"72",
          4836 => x"91",
          4837 => x"a0",
          4838 => x"3f",
          4839 => x"81",
          4840 => x"54",
          4841 => x"d8",
          4842 => x"39",
          4843 => x"bd",
          4844 => x"39",
          4845 => x"51",
          4846 => x"80",
          4847 => x"8c",
          4848 => x"0d",
          4849 => x"ff",
          4850 => x"06",
          4851 => x"83",
          4852 => x"70",
          4853 => x"55",
          4854 => x"73",
          4855 => x"53",
          4856 => x"bd",
          4857 => x"a0",
          4858 => x"3f",
          4859 => x"33",
          4860 => x"06",
          4861 => x"53",
          4862 => x"38",
          4863 => x"83",
          4864 => x"fe",
          4865 => x"0b",
          4866 => x"34",
          4867 => x"51",
          4868 => x"fe",
          4869 => x"52",
          4870 => x"d8",
          4871 => x"39",
          4872 => x"02",
          4873 => x"33",
          4874 => x"08",
          4875 => x"81",
          4876 => x"38",
          4877 => x"83",
          4878 => x"8a",
          4879 => x"38",
          4880 => x"82",
          4881 => x"88",
          4882 => x"38",
          4883 => x"88",
          4884 => x"b8",
          4885 => x"f9",
          4886 => x"f9",
          4887 => x"72",
          4888 => x"5e",
          4889 => x"88",
          4890 => x"a3",
          4891 => x"34",
          4892 => x"33",
          4893 => x"33",
          4894 => x"22",
          4895 => x"12",
          4896 => x"40",
          4897 => x"be",
          4898 => x"f9",
          4899 => x"71",
          4900 => x"40",
          4901 => x"b8",
          4902 => x"a3",
          4903 => x"34",
          4904 => x"33",
          4905 => x"06",
          4906 => x"22",
          4907 => x"33",
          4908 => x"11",
          4909 => x"58",
          4910 => x"b8",
          4911 => x"de",
          4912 => x"1d",
          4913 => x"06",
          4914 => x"61",
          4915 => x"38",
          4916 => x"33",
          4917 => x"f1",
          4918 => x"56",
          4919 => x"bd",
          4920 => x"84",
          4921 => x"9c",
          4922 => x"78",
          4923 => x"8a",
          4924 => x"25",
          4925 => x"78",
          4926 => x"b3",
          4927 => x"db",
          4928 => x"38",
          4929 => x"b9",
          4930 => x"b8",
          4931 => x"f9",
          4932 => x"f9",
          4933 => x"72",
          4934 => x"40",
          4935 => x"88",
          4936 => x"a3",
          4937 => x"34",
          4938 => x"33",
          4939 => x"33",
          4940 => x"22",
          4941 => x"12",
          4942 => x"56",
          4943 => x"be",
          4944 => x"f9",
          4945 => x"71",
          4946 => x"57",
          4947 => x"33",
          4948 => x"80",
          4949 => x"b8",
          4950 => x"81",
          4951 => x"f9",
          4952 => x"f9",
          4953 => x"72",
          4954 => x"42",
          4955 => x"83",
          4956 => x"60",
          4957 => x"05",
          4958 => x"58",
          4959 => x"06",
          4960 => x"27",
          4961 => x"77",
          4962 => x"34",
          4963 => x"ba",
          4964 => x"3d",
          4965 => x"9b",
          4966 => x"38",
          4967 => x"83",
          4968 => x"8d",
          4969 => x"06",
          4970 => x"80",
          4971 => x"bd",
          4972 => x"84",
          4973 => x"9c",
          4974 => x"78",
          4975 => x"aa",
          4976 => x"56",
          4977 => x"84",
          4978 => x"b9",
          4979 => x"11",
          4980 => x"84",
          4981 => x"78",
          4982 => x"18",
          4983 => x"ff",
          4984 => x"0b",
          4985 => x"1a",
          4986 => x"84",
          4987 => x"9c",
          4988 => x"78",
          4989 => x"e9",
          4990 => x"84",
          4991 => x"84",
          4992 => x"83",
          4993 => x"83",
          4994 => x"72",
          4995 => x"5e",
          4996 => x"b8",
          4997 => x"87",
          4998 => x"1d",
          4999 => x"80",
          5000 => x"bd",
          5001 => x"ba",
          5002 => x"29",
          5003 => x"59",
          5004 => x"f9",
          5005 => x"83",
          5006 => x"76",
          5007 => x"5b",
          5008 => x"b8",
          5009 => x"b0",
          5010 => x"84",
          5011 => x"70",
          5012 => x"83",
          5013 => x"83",
          5014 => x"72",
          5015 => x"44",
          5016 => x"59",
          5017 => x"33",
          5018 => x"de",
          5019 => x"1f",
          5020 => x"39",
          5021 => x"51",
          5022 => x"80",
          5023 => x"bd",
          5024 => x"39",
          5025 => x"33",
          5026 => x"33",
          5027 => x"06",
          5028 => x"33",
          5029 => x"12",
          5030 => x"80",
          5031 => x"ba",
          5032 => x"5d",
          5033 => x"05",
          5034 => x"ff",
          5035 => x"92",
          5036 => x"59",
          5037 => x"81",
          5038 => x"38",
          5039 => x"06",
          5040 => x"57",
          5041 => x"38",
          5042 => x"83",
          5043 => x"fc",
          5044 => x"0b",
          5045 => x"34",
          5046 => x"b9",
          5047 => x"0b",
          5048 => x"34",
          5049 => x"b9",
          5050 => x"0b",
          5051 => x"0c",
          5052 => x"ba",
          5053 => x"3d",
          5054 => x"f9",
          5055 => x"b9",
          5056 => x"f9",
          5057 => x"b9",
          5058 => x"f9",
          5059 => x"b9",
          5060 => x"0b",
          5061 => x"0c",
          5062 => x"ba",
          5063 => x"3d",
          5064 => x"80",
          5065 => x"81",
          5066 => x"38",
          5067 => x"33",
          5068 => x"33",
          5069 => x"06",
          5070 => x"33",
          5071 => x"06",
          5072 => x"11",
          5073 => x"80",
          5074 => x"ba",
          5075 => x"72",
          5076 => x"70",
          5077 => x"06",
          5078 => x"33",
          5079 => x"5c",
          5080 => x"7d",
          5081 => x"fe",
          5082 => x"ff",
          5083 => x"58",
          5084 => x"38",
          5085 => x"83",
          5086 => x"7b",
          5087 => x"7a",
          5088 => x"78",
          5089 => x"72",
          5090 => x"5f",
          5091 => x"b8",
          5092 => x"a3",
          5093 => x"34",
          5094 => x"33",
          5095 => x"33",
          5096 => x"22",
          5097 => x"12",
          5098 => x"40",
          5099 => x"f9",
          5100 => x"83",
          5101 => x"60",
          5102 => x"05",
          5103 => x"f9",
          5104 => x"a3",
          5105 => x"34",
          5106 => x"33",
          5107 => x"06",
          5108 => x"22",
          5109 => x"33",
          5110 => x"11",
          5111 => x"5e",
          5112 => x"b8",
          5113 => x"98",
          5114 => x"81",
          5115 => x"ff",
          5116 => x"7c",
          5117 => x"ea",
          5118 => x"81",
          5119 => x"96",
          5120 => x"19",
          5121 => x"f9",
          5122 => x"f9",
          5123 => x"81",
          5124 => x"ff",
          5125 => x"ac",
          5126 => x"2e",
          5127 => x"78",
          5128 => x"d7",
          5129 => x"2e",
          5130 => x"84",
          5131 => x"5f",
          5132 => x"38",
          5133 => x"56",
          5134 => x"84",
          5135 => x"10",
          5136 => x"98",
          5137 => x"08",
          5138 => x"83",
          5139 => x"80",
          5140 => x"e7",
          5141 => x"0b",
          5142 => x"0c",
          5143 => x"04",
          5144 => x"33",
          5145 => x"33",
          5146 => x"06",
          5147 => x"33",
          5148 => x"06",
          5149 => x"11",
          5150 => x"80",
          5151 => x"ba",
          5152 => x"72",
          5153 => x"70",
          5154 => x"06",
          5155 => x"33",
          5156 => x"5c",
          5157 => x"7f",
          5158 => x"ef",
          5159 => x"7a",
          5160 => x"7a",
          5161 => x"7a",
          5162 => x"72",
          5163 => x"5c",
          5164 => x"b8",
          5165 => x"a3",
          5166 => x"34",
          5167 => x"33",
          5168 => x"33",
          5169 => x"22",
          5170 => x"12",
          5171 => x"56",
          5172 => x"f9",
          5173 => x"83",
          5174 => x"76",
          5175 => x"5a",
          5176 => x"b8",
          5177 => x"b0",
          5178 => x"84",
          5179 => x"70",
          5180 => x"83",
          5181 => x"83",
          5182 => x"72",
          5183 => x"5b",
          5184 => x"59",
          5185 => x"33",
          5186 => x"18",
          5187 => x"05",
          5188 => x"06",
          5189 => x"7a",
          5190 => x"38",
          5191 => x"33",
          5192 => x"fb",
          5193 => x"56",
          5194 => x"bd",
          5195 => x"70",
          5196 => x"5d",
          5197 => x"26",
          5198 => x"83",
          5199 => x"84",
          5200 => x"83",
          5201 => x"72",
          5202 => x"72",
          5203 => x"72",
          5204 => x"72",
          5205 => x"54",
          5206 => x"5b",
          5207 => x"a8",
          5208 => x"a0",
          5209 => x"84",
          5210 => x"83",
          5211 => x"83",
          5212 => x"72",
          5213 => x"5e",
          5214 => x"a0",
          5215 => x"be",
          5216 => x"f9",
          5217 => x"71",
          5218 => x"5e",
          5219 => x"33",
          5220 => x"80",
          5221 => x"b8",
          5222 => x"81",
          5223 => x"f9",
          5224 => x"f9",
          5225 => x"72",
          5226 => x"44",
          5227 => x"83",
          5228 => x"84",
          5229 => x"34",
          5230 => x"70",
          5231 => x"5b",
          5232 => x"27",
          5233 => x"77",
          5234 => x"34",
          5235 => x"82",
          5236 => x"88",
          5237 => x"84",
          5238 => x"9c",
          5239 => x"83",
          5240 => x"33",
          5241 => x"88",
          5242 => x"34",
          5243 => x"33",
          5244 => x"06",
          5245 => x"56",
          5246 => x"81",
          5247 => x"8e",
          5248 => x"84",
          5249 => x"9c",
          5250 => x"83",
          5251 => x"33",
          5252 => x"88",
          5253 => x"34",
          5254 => x"33",
          5255 => x"33",
          5256 => x"33",
          5257 => x"80",
          5258 => x"39",
          5259 => x"42",
          5260 => x"11",
          5261 => x"51",
          5262 => x"3f",
          5263 => x"08",
          5264 => x"f0",
          5265 => x"8d",
          5266 => x"57",
          5267 => x"b9",
          5268 => x"10",
          5269 => x"41",
          5270 => x"05",
          5271 => x"b9",
          5272 => x"fb",
          5273 => x"f9",
          5274 => x"5c",
          5275 => x"1c",
          5276 => x"83",
          5277 => x"84",
          5278 => x"83",
          5279 => x"5b",
          5280 => x"e5",
          5281 => x"80",
          5282 => x"bc",
          5283 => x"bd",
          5284 => x"29",
          5285 => x"5b",
          5286 => x"19",
          5287 => x"a3",
          5288 => x"34",
          5289 => x"33",
          5290 => x"33",
          5291 => x"22",
          5292 => x"12",
          5293 => x"56",
          5294 => x"be",
          5295 => x"f9",
          5296 => x"71",
          5297 => x"5e",
          5298 => x"33",
          5299 => x"b0",
          5300 => x"84",
          5301 => x"70",
          5302 => x"83",
          5303 => x"83",
          5304 => x"72",
          5305 => x"41",
          5306 => x"5a",
          5307 => x"33",
          5308 => x"1e",
          5309 => x"70",
          5310 => x"5c",
          5311 => x"26",
          5312 => x"84",
          5313 => x"58",
          5314 => x"38",
          5315 => x"75",
          5316 => x"34",
          5317 => x"b9",
          5318 => x"b8",
          5319 => x"7f",
          5320 => x"bd",
          5321 => x"84",
          5322 => x"f3",
          5323 => x"52",
          5324 => x"e4",
          5325 => x"84",
          5326 => x"9c",
          5327 => x"84",
          5328 => x"83",
          5329 => x"84",
          5330 => x"83",
          5331 => x"84",
          5332 => x"57",
          5333 => x"ba",
          5334 => x"39",
          5335 => x"33",
          5336 => x"34",
          5337 => x"33",
          5338 => x"34",
          5339 => x"33",
          5340 => x"34",
          5341 => x"84",
          5342 => x"5b",
          5343 => x"ff",
          5344 => x"b9",
          5345 => x"7c",
          5346 => x"81",
          5347 => x"38",
          5348 => x"33",
          5349 => x"83",
          5350 => x"81",
          5351 => x"53",
          5352 => x"52",
          5353 => x"52",
          5354 => x"fe",
          5355 => x"fe",
          5356 => x"84",
          5357 => x"81",
          5358 => x"f8",
          5359 => x"76",
          5360 => x"a0",
          5361 => x"38",
          5362 => x"f7",
          5363 => x"fd",
          5364 => x"c0",
          5365 => x"84",
          5366 => x"5b",
          5367 => x"ff",
          5368 => x"7b",
          5369 => x"38",
          5370 => x"b9",
          5371 => x"11",
          5372 => x"75",
          5373 => x"a5",
          5374 => x"10",
          5375 => x"05",
          5376 => x"04",
          5377 => x"33",
          5378 => x"2e",
          5379 => x"83",
          5380 => x"84",
          5381 => x"71",
          5382 => x"09",
          5383 => x"72",
          5384 => x"59",
          5385 => x"83",
          5386 => x"fd",
          5387 => x"b9",
          5388 => x"75",
          5389 => x"e7",
          5390 => x"e1",
          5391 => x"70",
          5392 => x"84",
          5393 => x"5d",
          5394 => x"7b",
          5395 => x"38",
          5396 => x"bd",
          5397 => x"39",
          5398 => x"f9",
          5399 => x"f9",
          5400 => x"81",
          5401 => x"57",
          5402 => x"fd",
          5403 => x"17",
          5404 => x"f9",
          5405 => x"9c",
          5406 => x"83",
          5407 => x"83",
          5408 => x"84",
          5409 => x"ff",
          5410 => x"76",
          5411 => x"84",
          5412 => x"56",
          5413 => x"bc",
          5414 => x"39",
          5415 => x"33",
          5416 => x"2e",
          5417 => x"83",
          5418 => x"84",
          5419 => x"71",
          5420 => x"09",
          5421 => x"72",
          5422 => x"59",
          5423 => x"83",
          5424 => x"fc",
          5425 => x"b9",
          5426 => x"7a",
          5427 => x"c4",
          5428 => x"e0",
          5429 => x"99",
          5430 => x"06",
          5431 => x"84",
          5432 => x"83",
          5433 => x"83",
          5434 => x"72",
          5435 => x"87",
          5436 => x"11",
          5437 => x"22",
          5438 => x"58",
          5439 => x"05",
          5440 => x"ff",
          5441 => x"90",
          5442 => x"fe",
          5443 => x"5a",
          5444 => x"84",
          5445 => x"92",
          5446 => x"0b",
          5447 => x"34",
          5448 => x"84",
          5449 => x"5a",
          5450 => x"fb",
          5451 => x"b9",
          5452 => x"77",
          5453 => x"81",
          5454 => x"38",
          5455 => x"f8",
          5456 => x"d0",
          5457 => x"8d",
          5458 => x"80",
          5459 => x"38",
          5460 => x"33",
          5461 => x"33",
          5462 => x"84",
          5463 => x"ff",
          5464 => x"56",
          5465 => x"83",
          5466 => x"76",
          5467 => x"34",
          5468 => x"84",
          5469 => x"57",
          5470 => x"8c",
          5471 => x"b9",
          5472 => x"f9",
          5473 => x"61",
          5474 => x"ff",
          5475 => x"59",
          5476 => x"60",
          5477 => x"75",
          5478 => x"f9",
          5479 => x"f4",
          5480 => x"98",
          5481 => x"e2",
          5482 => x"84",
          5483 => x"57",
          5484 => x"27",
          5485 => x"76",
          5486 => x"e0",
          5487 => x"53",
          5488 => x"f8",
          5489 => x"c2",
          5490 => x"70",
          5491 => x"84",
          5492 => x"58",
          5493 => x"39",
          5494 => x"b9",
          5495 => x"57",
          5496 => x"8d",
          5497 => x"e0",
          5498 => x"83",
          5499 => x"75",
          5500 => x"76",
          5501 => x"51",
          5502 => x"fa",
          5503 => x"b9",
          5504 => x"81",
          5505 => x"b7",
          5506 => x"e3",
          5507 => x"70",
          5508 => x"84",
          5509 => x"ff",
          5510 => x"ff",
          5511 => x"ff",
          5512 => x"ff",
          5513 => x"40",
          5514 => x"59",
          5515 => x"7e",
          5516 => x"77",
          5517 => x"f9",
          5518 => x"81",
          5519 => x"18",
          5520 => x"7f",
          5521 => x"77",
          5522 => x"f9",
          5523 => x"b8",
          5524 => x"11",
          5525 => x"60",
          5526 => x"38",
          5527 => x"83",
          5528 => x"f9",
          5529 => x"b9",
          5530 => x"7e",
          5531 => x"ef",
          5532 => x"e1",
          5533 => x"ff",
          5534 => x"7a",
          5535 => x"94",
          5536 => x"bc",
          5537 => x"80",
          5538 => x"ff",
          5539 => x"bd",
          5540 => x"29",
          5541 => x"a0",
          5542 => x"f9",
          5543 => x"40",
          5544 => x"05",
          5545 => x"ff",
          5546 => x"92",
          5547 => x"59",
          5548 => x"60",
          5549 => x"f0",
          5550 => x"ff",
          5551 => x"7c",
          5552 => x"80",
          5553 => x"fe",
          5554 => x"ff",
          5555 => x"76",
          5556 => x"38",
          5557 => x"75",
          5558 => x"23",
          5559 => x"06",
          5560 => x"41",
          5561 => x"24",
          5562 => x"84",
          5563 => x"56",
          5564 => x"8d",
          5565 => x"16",
          5566 => x"f9",
          5567 => x"81",
          5568 => x"f9",
          5569 => x"57",
          5570 => x"76",
          5571 => x"75",
          5572 => x"05",
          5573 => x"06",
          5574 => x"5c",
          5575 => x"58",
          5576 => x"80",
          5577 => x"b0",
          5578 => x"ff",
          5579 => x"ff",
          5580 => x"29",
          5581 => x"42",
          5582 => x"27",
          5583 => x"84",
          5584 => x"57",
          5585 => x"33",
          5586 => x"88",
          5587 => x"70",
          5588 => x"34",
          5589 => x"05",
          5590 => x"70",
          5591 => x"34",
          5592 => x"b8",
          5593 => x"b7",
          5594 => x"71",
          5595 => x"40",
          5596 => x"60",
          5597 => x"38",
          5598 => x"33",
          5599 => x"88",
          5600 => x"70",
          5601 => x"34",
          5602 => x"05",
          5603 => x"70",
          5604 => x"34",
          5605 => x"b8",
          5606 => x"b7",
          5607 => x"71",
          5608 => x"40",
          5609 => x"78",
          5610 => x"38",
          5611 => x"84",
          5612 => x"56",
          5613 => x"87",
          5614 => x"52",
          5615 => x"33",
          5616 => x"3f",
          5617 => x"80",
          5618 => x"80",
          5619 => x"84",
          5620 => x"5d",
          5621 => x"79",
          5622 => x"38",
          5623 => x"22",
          5624 => x"2e",
          5625 => x"8b",
          5626 => x"f9",
          5627 => x"76",
          5628 => x"83",
          5629 => x"79",
          5630 => x"76",
          5631 => x"ed",
          5632 => x"ff",
          5633 => x"60",
          5634 => x"38",
          5635 => x"06",
          5636 => x"26",
          5637 => x"7b",
          5638 => x"7d",
          5639 => x"76",
          5640 => x"7a",
          5641 => x"70",
          5642 => x"05",
          5643 => x"80",
          5644 => x"5d",
          5645 => x"b0",
          5646 => x"83",
          5647 => x"5d",
          5648 => x"38",
          5649 => x"57",
          5650 => x"38",
          5651 => x"33",
          5652 => x"71",
          5653 => x"71",
          5654 => x"71",
          5655 => x"59",
          5656 => x"77",
          5657 => x"38",
          5658 => x"84",
          5659 => x"7d",
          5660 => x"05",
          5661 => x"77",
          5662 => x"84",
          5663 => x"84",
          5664 => x"41",
          5665 => x"ff",
          5666 => x"ff",
          5667 => x"ba",
          5668 => x"29",
          5669 => x"59",
          5670 => x"77",
          5671 => x"76",
          5672 => x"70",
          5673 => x"05",
          5674 => x"76",
          5675 => x"76",
          5676 => x"e0",
          5677 => x"b8",
          5678 => x"de",
          5679 => x"a0",
          5680 => x"19",
          5681 => x"70",
          5682 => x"34",
          5683 => x"76",
          5684 => x"c0",
          5685 => x"e0",
          5686 => x"79",
          5687 => x"05",
          5688 => x"17",
          5689 => x"27",
          5690 => x"a8",
          5691 => x"70",
          5692 => x"5d",
          5693 => x"39",
          5694 => x"33",
          5695 => x"06",
          5696 => x"80",
          5697 => x"84",
          5698 => x"5d",
          5699 => x"f0",
          5700 => x"06",
          5701 => x"f2",
          5702 => x"b8",
          5703 => x"70",
          5704 => x"59",
          5705 => x"39",
          5706 => x"17",
          5707 => x"b8",
          5708 => x"7c",
          5709 => x"bc",
          5710 => x"80",
          5711 => x"ba",
          5712 => x"ff",
          5713 => x"5f",
          5714 => x"39",
          5715 => x"33",
          5716 => x"75",
          5717 => x"34",
          5718 => x"81",
          5719 => x"56",
          5720 => x"83",
          5721 => x"81",
          5722 => x"07",
          5723 => x"f9",
          5724 => x"39",
          5725 => x"33",
          5726 => x"83",
          5727 => x"83",
          5728 => x"d4",
          5729 => x"b8",
          5730 => x"06",
          5731 => x"75",
          5732 => x"34",
          5733 => x"f9",
          5734 => x"9f",
          5735 => x"56",
          5736 => x"b8",
          5737 => x"39",
          5738 => x"83",
          5739 => x"81",
          5740 => x"ff",
          5741 => x"f4",
          5742 => x"f9",
          5743 => x"8f",
          5744 => x"83",
          5745 => x"ff",
          5746 => x"f9",
          5747 => x"9f",
          5748 => x"56",
          5749 => x"b8",
          5750 => x"39",
          5751 => x"33",
          5752 => x"80",
          5753 => x"75",
          5754 => x"34",
          5755 => x"83",
          5756 => x"81",
          5757 => x"c0",
          5758 => x"83",
          5759 => x"fe",
          5760 => x"f9",
          5761 => x"af",
          5762 => x"56",
          5763 => x"b8",
          5764 => x"39",
          5765 => x"33",
          5766 => x"86",
          5767 => x"83",
          5768 => x"fe",
          5769 => x"f9",
          5770 => x"fc",
          5771 => x"56",
          5772 => x"b8",
          5773 => x"39",
          5774 => x"33",
          5775 => x"82",
          5776 => x"83",
          5777 => x"fe",
          5778 => x"f9",
          5779 => x"f8",
          5780 => x"83",
          5781 => x"fd",
          5782 => x"f9",
          5783 => x"f0",
          5784 => x"83",
          5785 => x"fd",
          5786 => x"f9",
          5787 => x"f0",
          5788 => x"83",
          5789 => x"fd",
          5790 => x"f9",
          5791 => x"df",
          5792 => x"07",
          5793 => x"f9",
          5794 => x"cc",
          5795 => x"b8",
          5796 => x"06",
          5797 => x"75",
          5798 => x"34",
          5799 => x"80",
          5800 => x"bd",
          5801 => x"81",
          5802 => x"3f",
          5803 => x"84",
          5804 => x"83",
          5805 => x"84",
          5806 => x"83",
          5807 => x"84",
          5808 => x"59",
          5809 => x"ba",
          5810 => x"84",
          5811 => x"e8",
          5812 => x"0b",
          5813 => x"34",
          5814 => x"ba",
          5815 => x"3d",
          5816 => x"83",
          5817 => x"83",
          5818 => x"70",
          5819 => x"58",
          5820 => x"e7",
          5821 => x"b9",
          5822 => x"3d",
          5823 => x"d8",
          5824 => x"f9",
          5825 => x"ba",
          5826 => x"38",
          5827 => x"08",
          5828 => x"0c",
          5829 => x"b9",
          5830 => x"0b",
          5831 => x"0c",
          5832 => x"04",
          5833 => x"bd",
          5834 => x"39",
          5835 => x"33",
          5836 => x"5c",
          5837 => x"8d",
          5838 => x"83",
          5839 => x"02",
          5840 => x"22",
          5841 => x"1e",
          5842 => x"84",
          5843 => x"ca",
          5844 => x"83",
          5845 => x"80",
          5846 => x"d1",
          5847 => x"f9",
          5848 => x"81",
          5849 => x"ff",
          5850 => x"d8",
          5851 => x"83",
          5852 => x"80",
          5853 => x"d0",
          5854 => x"98",
          5855 => x"fe",
          5856 => x"ef",
          5857 => x"f9",
          5858 => x"05",
          5859 => x"9f",
          5860 => x"58",
          5861 => x"a6",
          5862 => x"81",
          5863 => x"84",
          5864 => x"40",
          5865 => x"ee",
          5866 => x"83",
          5867 => x"ee",
          5868 => x"f9",
          5869 => x"05",
          5870 => x"9f",
          5871 => x"58",
          5872 => x"e2",
          5873 => x"bc",
          5874 => x"84",
          5875 => x"ff",
          5876 => x"56",
          5877 => x"f3",
          5878 => x"57",
          5879 => x"84",
          5880 => x"70",
          5881 => x"58",
          5882 => x"26",
          5883 => x"83",
          5884 => x"84",
          5885 => x"70",
          5886 => x"83",
          5887 => x"71",
          5888 => x"87",
          5889 => x"05",
          5890 => x"22",
          5891 => x"7e",
          5892 => x"83",
          5893 => x"83",
          5894 => x"5d",
          5895 => x"5f",
          5896 => x"2e",
          5897 => x"79",
          5898 => x"06",
          5899 => x"57",
          5900 => x"84",
          5901 => x"b7",
          5902 => x"76",
          5903 => x"98",
          5904 => x"56",
          5905 => x"ba",
          5906 => x"ff",
          5907 => x"57",
          5908 => x"24",
          5909 => x"84",
          5910 => x"56",
          5911 => x"82",
          5912 => x"16",
          5913 => x"f9",
          5914 => x"81",
          5915 => x"f9",
          5916 => x"57",
          5917 => x"76",
          5918 => x"75",
          5919 => x"05",
          5920 => x"06",
          5921 => x"5c",
          5922 => x"58",
          5923 => x"80",
          5924 => x"b0",
          5925 => x"ff",
          5926 => x"ff",
          5927 => x"29",
          5928 => x"42",
          5929 => x"27",
          5930 => x"84",
          5931 => x"57",
          5932 => x"33",
          5933 => x"88",
          5934 => x"70",
          5935 => x"34",
          5936 => x"05",
          5937 => x"70",
          5938 => x"34",
          5939 => x"b8",
          5940 => x"b7",
          5941 => x"71",
          5942 => x"41",
          5943 => x"76",
          5944 => x"38",
          5945 => x"33",
          5946 => x"88",
          5947 => x"70",
          5948 => x"34",
          5949 => x"05",
          5950 => x"70",
          5951 => x"34",
          5952 => x"b8",
          5953 => x"b7",
          5954 => x"71",
          5955 => x"41",
          5956 => x"78",
          5957 => x"38",
          5958 => x"83",
          5959 => x"33",
          5960 => x"88",
          5961 => x"34",
          5962 => x"33",
          5963 => x"33",
          5964 => x"22",
          5965 => x"33",
          5966 => x"5d",
          5967 => x"76",
          5968 => x"84",
          5969 => x"70",
          5970 => x"ff",
          5971 => x"58",
          5972 => x"83",
          5973 => x"79",
          5974 => x"23",
          5975 => x"06",
          5976 => x"5a",
          5977 => x"83",
          5978 => x"76",
          5979 => x"34",
          5980 => x"33",
          5981 => x"06",
          5982 => x"59",
          5983 => x"27",
          5984 => x"80",
          5985 => x"f9",
          5986 => x"88",
          5987 => x"bd",
          5988 => x"84",
          5989 => x"ff",
          5990 => x"56",
          5991 => x"ef",
          5992 => x"57",
          5993 => x"75",
          5994 => x"81",
          5995 => x"38",
          5996 => x"33",
          5997 => x"06",
          5998 => x"33",
          5999 => x"5d",
          6000 => x"2e",
          6001 => x"f4",
          6002 => x"a1",
          6003 => x"56",
          6004 => x"bc",
          6005 => x"39",
          6006 => x"75",
          6007 => x"23",
          6008 => x"7c",
          6009 => x"75",
          6010 => x"34",
          6011 => x"77",
          6012 => x"77",
          6013 => x"8d",
          6014 => x"70",
          6015 => x"34",
          6016 => x"33",
          6017 => x"05",
          6018 => x"7a",
          6019 => x"38",
          6020 => x"81",
          6021 => x"83",
          6022 => x"77",
          6023 => x"59",
          6024 => x"27",
          6025 => x"d3",
          6026 => x"31",
          6027 => x"f9",
          6028 => x"a8",
          6029 => x"83",
          6030 => x"fc",
          6031 => x"83",
          6032 => x"fc",
          6033 => x"0b",
          6034 => x"23",
          6035 => x"80",
          6036 => x"bc",
          6037 => x"39",
          6038 => x"18",
          6039 => x"b8",
          6040 => x"77",
          6041 => x"83",
          6042 => x"e9",
          6043 => x"3d",
          6044 => x"05",
          6045 => x"82",
          6046 => x"72",
          6047 => x"38",
          6048 => x"9c",
          6049 => x"84",
          6050 => x"85",
          6051 => x"76",
          6052 => x"d7",
          6053 => x"0b",
          6054 => x"0c",
          6055 => x"04",
          6056 => x"02",
          6057 => x"5c",
          6058 => x"f8",
          6059 => x"81",
          6060 => x"f7",
          6061 => x"58",
          6062 => x"74",
          6063 => x"d6",
          6064 => x"56",
          6065 => x"90",
          6066 => x"78",
          6067 => x"0c",
          6068 => x"04",
          6069 => x"08",
          6070 => x"73",
          6071 => x"38",
          6072 => x"70",
          6073 => x"70",
          6074 => x"2a",
          6075 => x"58",
          6076 => x"ec",
          6077 => x"80",
          6078 => x"2e",
          6079 => x"83",
          6080 => x"7b",
          6081 => x"30",
          6082 => x"76",
          6083 => x"5d",
          6084 => x"85",
          6085 => x"b8",
          6086 => x"f9",
          6087 => x"f9",
          6088 => x"71",
          6089 => x"a3",
          6090 => x"83",
          6091 => x"5b",
          6092 => x"79",
          6093 => x"83",
          6094 => x"83",
          6095 => x"58",
          6096 => x"74",
          6097 => x"8c",
          6098 => x"54",
          6099 => x"80",
          6100 => x"0b",
          6101 => x"88",
          6102 => x"98",
          6103 => x"75",
          6104 => x"38",
          6105 => x"84",
          6106 => x"83",
          6107 => x"34",
          6108 => x"81",
          6109 => x"55",
          6110 => x"27",
          6111 => x"54",
          6112 => x"14",
          6113 => x"ff",
          6114 => x"b6",
          6115 => x"54",
          6116 => x"2e",
          6117 => x"72",
          6118 => x"86",
          6119 => x"83",
          6120 => x"34",
          6121 => x"06",
          6122 => x"ff",
          6123 => x"38",
          6124 => x"ca",
          6125 => x"f7",
          6126 => x"83",
          6127 => x"34",
          6128 => x"81",
          6129 => x"5e",
          6130 => x"ff",
          6131 => x"f7",
          6132 => x"98",
          6133 => x"25",
          6134 => x"75",
          6135 => x"34",
          6136 => x"06",
          6137 => x"81",
          6138 => x"06",
          6139 => x"72",
          6140 => x"e7",
          6141 => x"83",
          6142 => x"73",
          6143 => x"53",
          6144 => x"85",
          6145 => x"0b",
          6146 => x"34",
          6147 => x"f7",
          6148 => x"f7",
          6149 => x"f7",
          6150 => x"83",
          6151 => x"83",
          6152 => x"5d",
          6153 => x"5c",
          6154 => x"f7",
          6155 => x"55",
          6156 => x"2e",
          6157 => x"f7",
          6158 => x"54",
          6159 => x"82",
          6160 => x"f7",
          6161 => x"53",
          6162 => x"2e",
          6163 => x"f7",
          6164 => x"54",
          6165 => x"38",
          6166 => x"06",
          6167 => x"ff",
          6168 => x"83",
          6169 => x"33",
          6170 => x"2e",
          6171 => x"74",
          6172 => x"53",
          6173 => x"2e",
          6174 => x"83",
          6175 => x"33",
          6176 => x"27",
          6177 => x"83",
          6178 => x"87",
          6179 => x"c0",
          6180 => x"54",
          6181 => x"27",
          6182 => x"81",
          6183 => x"98",
          6184 => x"f7",
          6185 => x"81",
          6186 => x"ff",
          6187 => x"89",
          6188 => x"f6",
          6189 => x"f7",
          6190 => x"83",
          6191 => x"fe",
          6192 => x"72",
          6193 => x"8b",
          6194 => x"10",
          6195 => x"05",
          6196 => x"04",
          6197 => x"08",
          6198 => x"2e",
          6199 => x"f4",
          6200 => x"98",
          6201 => x"5e",
          6202 => x"fc",
          6203 => x"0b",
          6204 => x"33",
          6205 => x"81",
          6206 => x"74",
          6207 => x"f8",
          6208 => x"c0",
          6209 => x"83",
          6210 => x"73",
          6211 => x"58",
          6212 => x"94",
          6213 => x"be",
          6214 => x"84",
          6215 => x"33",
          6216 => x"f0",
          6217 => x"39",
          6218 => x"08",
          6219 => x"2e",
          6220 => x"72",
          6221 => x"f4",
          6222 => x"76",
          6223 => x"54",
          6224 => x"80",
          6225 => x"39",
          6226 => x"57",
          6227 => x"81",
          6228 => x"79",
          6229 => x"81",
          6230 => x"38",
          6231 => x"80",
          6232 => x"81",
          6233 => x"38",
          6234 => x"06",
          6235 => x"27",
          6236 => x"54",
          6237 => x"25",
          6238 => x"80",
          6239 => x"81",
          6240 => x"ff",
          6241 => x"81",
          6242 => x"72",
          6243 => x"2b",
          6244 => x"58",
          6245 => x"24",
          6246 => x"10",
          6247 => x"10",
          6248 => x"83",
          6249 => x"83",
          6250 => x"70",
          6251 => x"54",
          6252 => x"98",
          6253 => x"f7",
          6254 => x"fd",
          6255 => x"59",
          6256 => x"ff",
          6257 => x"81",
          6258 => x"ff",
          6259 => x"59",
          6260 => x"78",
          6261 => x"9f",
          6262 => x"84",
          6263 => x"54",
          6264 => x"2e",
          6265 => x"7b",
          6266 => x"30",
          6267 => x"76",
          6268 => x"56",
          6269 => x"7b",
          6270 => x"81",
          6271 => x"38",
          6272 => x"f9",
          6273 => x"53",
          6274 => x"10",
          6275 => x"05",
          6276 => x"54",
          6277 => x"83",
          6278 => x"13",
          6279 => x"06",
          6280 => x"73",
          6281 => x"84",
          6282 => x"53",
          6283 => x"f9",
          6284 => x"b8",
          6285 => x"74",
          6286 => x"78",
          6287 => x"52",
          6288 => x"d4",
          6289 => x"ba",
          6290 => x"3d",
          6291 => x"76",
          6292 => x"54",
          6293 => x"72",
          6294 => x"92",
          6295 => x"d4",
          6296 => x"05",
          6297 => x"f7",
          6298 => x"fa",
          6299 => x"0b",
          6300 => x"15",
          6301 => x"83",
          6302 => x"34",
          6303 => x"f7",
          6304 => x"fa",
          6305 => x"81",
          6306 => x"72",
          6307 => x"fc",
          6308 => x"f7",
          6309 => x"55",
          6310 => x"fc",
          6311 => x"81",
          6312 => x"73",
          6313 => x"81",
          6314 => x"38",
          6315 => x"08",
          6316 => x"87",
          6317 => x"08",
          6318 => x"73",
          6319 => x"38",
          6320 => x"9c",
          6321 => x"e0",
          6322 => x"ff",
          6323 => x"d7",
          6324 => x"83",
          6325 => x"34",
          6326 => x"72",
          6327 => x"34",
          6328 => x"06",
          6329 => x"9e",
          6330 => x"f7",
          6331 => x"0b",
          6332 => x"33",
          6333 => x"08",
          6334 => x"33",
          6335 => x"e8",
          6336 => x"e7",
          6337 => x"42",
          6338 => x"56",
          6339 => x"79",
          6340 => x"81",
          6341 => x"38",
          6342 => x"81",
          6343 => x"38",
          6344 => x"09",
          6345 => x"c0",
          6346 => x"39",
          6347 => x"81",
          6348 => x"98",
          6349 => x"84",
          6350 => x"57",
          6351 => x"38",
          6352 => x"84",
          6353 => x"ff",
          6354 => x"39",
          6355 => x"b8",
          6356 => x"54",
          6357 => x"81",
          6358 => x"b8",
          6359 => x"59",
          6360 => x"81",
          6361 => x"ec",
          6362 => x"f7",
          6363 => x"0b",
          6364 => x"0c",
          6365 => x"84",
          6366 => x"70",
          6367 => x"ff",
          6368 => x"54",
          6369 => x"83",
          6370 => x"74",
          6371 => x"23",
          6372 => x"06",
          6373 => x"53",
          6374 => x"83",
          6375 => x"73",
          6376 => x"34",
          6377 => x"33",
          6378 => x"06",
          6379 => x"53",
          6380 => x"83",
          6381 => x"72",
          6382 => x"34",
          6383 => x"b7",
          6384 => x"83",
          6385 => x"a5",
          6386 => x"f6",
          6387 => x"54",
          6388 => x"84",
          6389 => x"83",
          6390 => x"fe",
          6391 => x"81",
          6392 => x"90",
          6393 => x"f0",
          6394 => x"bb",
          6395 => x"0d",
          6396 => x"ac",
          6397 => x"0d",
          6398 => x"0d",
          6399 => x"f4",
          6400 => x"58",
          6401 => x"33",
          6402 => x"83",
          6403 => x"52",
          6404 => x"34",
          6405 => x"f4",
          6406 => x"57",
          6407 => x"16",
          6408 => x"86",
          6409 => x"34",
          6410 => x"9c",
          6411 => x"98",
          6412 => x"ce",
          6413 => x"87",
          6414 => x"08",
          6415 => x"98",
          6416 => x"71",
          6417 => x"38",
          6418 => x"87",
          6419 => x"08",
          6420 => x"74",
          6421 => x"72",
          6422 => x"db",
          6423 => x"98",
          6424 => x"ff",
          6425 => x"27",
          6426 => x"72",
          6427 => x"2e",
          6428 => x"87",
          6429 => x"08",
          6430 => x"05",
          6431 => x"98",
          6432 => x"87",
          6433 => x"08",
          6434 => x"2e",
          6435 => x"15",
          6436 => x"98",
          6437 => x"53",
          6438 => x"87",
          6439 => x"ff",
          6440 => x"87",
          6441 => x"08",
          6442 => x"71",
          6443 => x"38",
          6444 => x"ff",
          6445 => x"76",
          6446 => x"38",
          6447 => x"06",
          6448 => x"d8",
          6449 => x"2e",
          6450 => x"84",
          6451 => x"89",
          6452 => x"ff",
          6453 => x"ff",
          6454 => x"76",
          6455 => x"0b",
          6456 => x"52",
          6457 => x"8d",
          6458 => x"ba",
          6459 => x"3d",
          6460 => x"3d",
          6461 => x"84",
          6462 => x"33",
          6463 => x"0b",
          6464 => x"08",
          6465 => x"87",
          6466 => x"06",
          6467 => x"2a",
          6468 => x"56",
          6469 => x"16",
          6470 => x"2a",
          6471 => x"16",
          6472 => x"2a",
          6473 => x"16",
          6474 => x"16",
          6475 => x"98",
          6476 => x"82",
          6477 => x"f4",
          6478 => x"80",
          6479 => x"85",
          6480 => x"98",
          6481 => x"fe",
          6482 => x"34",
          6483 => x"f0",
          6484 => x"87",
          6485 => x"08",
          6486 => x"08",
          6487 => x"90",
          6488 => x"c0",
          6489 => x"53",
          6490 => x"9c",
          6491 => x"73",
          6492 => x"81",
          6493 => x"c0",
          6494 => x"57",
          6495 => x"27",
          6496 => x"81",
          6497 => x"38",
          6498 => x"a4",
          6499 => x"56",
          6500 => x"80",
          6501 => x"56",
          6502 => x"80",
          6503 => x"c0",
          6504 => x"80",
          6505 => x"54",
          6506 => x"9c",
          6507 => x"c0",
          6508 => x"56",
          6509 => x"f6",
          6510 => x"33",
          6511 => x"9c",
          6512 => x"71",
          6513 => x"38",
          6514 => x"2e",
          6515 => x"c0",
          6516 => x"52",
          6517 => x"74",
          6518 => x"38",
          6519 => x"ff",
          6520 => x"38",
          6521 => x"80",
          6522 => x"81",
          6523 => x"72",
          6524 => x"75",
          6525 => x"ff",
          6526 => x"aa",
          6527 => x"15",
          6528 => x"11",
          6529 => x"71",
          6530 => x"38",
          6531 => x"05",
          6532 => x"70",
          6533 => x"34",
          6534 => x"f0",
          6535 => x"ba",
          6536 => x"3d",
          6537 => x"0b",
          6538 => x"52",
          6539 => x"c5",
          6540 => x"ba",
          6541 => x"3d",
          6542 => x"17",
          6543 => x"06",
          6544 => x"ff",
          6545 => x"52",
          6546 => x"f9",
          6547 => x"02",
          6548 => x"05",
          6549 => x"80",
          6550 => x"98",
          6551 => x"2b",
          6552 => x"80",
          6553 => x"98",
          6554 => x"56",
          6555 => x"83",
          6556 => x"90",
          6557 => x"84",
          6558 => x"90",
          6559 => x"85",
          6560 => x"86",
          6561 => x"83",
          6562 => x"80",
          6563 => x"80",
          6564 => x"56",
          6565 => x"27",
          6566 => x"70",
          6567 => x"33",
          6568 => x"05",
          6569 => x"72",
          6570 => x"83",
          6571 => x"55",
          6572 => x"34",
          6573 => x"08",
          6574 => x"76",
          6575 => x"83",
          6576 => x"56",
          6577 => x"81",
          6578 => x"0b",
          6579 => x"e8",
          6580 => x"98",
          6581 => x"f4",
          6582 => x"80",
          6583 => x"54",
          6584 => x"9c",
          6585 => x"c0",
          6586 => x"52",
          6587 => x"f6",
          6588 => x"33",
          6589 => x"9c",
          6590 => x"75",
          6591 => x"38",
          6592 => x"2e",
          6593 => x"c0",
          6594 => x"52",
          6595 => x"74",
          6596 => x"38",
          6597 => x"ff",
          6598 => x"38",
          6599 => x"9c",
          6600 => x"90",
          6601 => x"c0",
          6602 => x"53",
          6603 => x"9c",
          6604 => x"73",
          6605 => x"81",
          6606 => x"c0",
          6607 => x"53",
          6608 => x"27",
          6609 => x"81",
          6610 => x"38",
          6611 => x"a4",
          6612 => x"56",
          6613 => x"a9",
          6614 => x"72",
          6615 => x"38",
          6616 => x"a8",
          6617 => x"ff",
          6618 => x"fe",
          6619 => x"70",
          6620 => x"56",
          6621 => x"38",
          6622 => x"8c",
          6623 => x"0d",
          6624 => x"70",
          6625 => x"58",
          6626 => x"38",
          6627 => x"ff",
          6628 => x"74",
          6629 => x"38",
          6630 => x"e4",
          6631 => x"fe",
          6632 => x"77",
          6633 => x"0c",
          6634 => x"04",
          6635 => x"83",
          6636 => x"51",
          6637 => x"34",
          6638 => x"f4",
          6639 => x"56",
          6640 => x"16",
          6641 => x"86",
          6642 => x"34",
          6643 => x"9c",
          6644 => x"98",
          6645 => x"ce",
          6646 => x"87",
          6647 => x"08",
          6648 => x"98",
          6649 => x"72",
          6650 => x"38",
          6651 => x"87",
          6652 => x"08",
          6653 => x"74",
          6654 => x"71",
          6655 => x"db",
          6656 => x"98",
          6657 => x"ff",
          6658 => x"27",
          6659 => x"71",
          6660 => x"2e",
          6661 => x"87",
          6662 => x"08",
          6663 => x"05",
          6664 => x"98",
          6665 => x"87",
          6666 => x"08",
          6667 => x"2e",
          6668 => x"15",
          6669 => x"98",
          6670 => x"52",
          6671 => x"87",
          6672 => x"ff",
          6673 => x"87",
          6674 => x"08",
          6675 => x"70",
          6676 => x"38",
          6677 => x"ff",
          6678 => x"75",
          6679 => x"38",
          6680 => x"06",
          6681 => x"d8",
          6682 => x"ff",
          6683 => x"ff",
          6684 => x"e7",
          6685 => x"0d",
          6686 => x"51",
          6687 => x"3f",
          6688 => x"04",
          6689 => x"84",
          6690 => x"7a",
          6691 => x"2a",
          6692 => x"ff",
          6693 => x"2b",
          6694 => x"33",
          6695 => x"71",
          6696 => x"83",
          6697 => x"11",
          6698 => x"12",
          6699 => x"2b",
          6700 => x"07",
          6701 => x"53",
          6702 => x"59",
          6703 => x"53",
          6704 => x"81",
          6705 => x"16",
          6706 => x"83",
          6707 => x"8b",
          6708 => x"2b",
          6709 => x"70",
          6710 => x"33",
          6711 => x"71",
          6712 => x"57",
          6713 => x"59",
          6714 => x"71",
          6715 => x"38",
          6716 => x"85",
          6717 => x"8b",
          6718 => x"2b",
          6719 => x"76",
          6720 => x"54",
          6721 => x"86",
          6722 => x"81",
          6723 => x"73",
          6724 => x"84",
          6725 => x"70",
          6726 => x"33",
          6727 => x"71",
          6728 => x"70",
          6729 => x"55",
          6730 => x"77",
          6731 => x"71",
          6732 => x"84",
          6733 => x"16",
          6734 => x"86",
          6735 => x"0b",
          6736 => x"84",
          6737 => x"53",
          6738 => x"34",
          6739 => x"34",
          6740 => x"08",
          6741 => x"81",
          6742 => x"88",
          6743 => x"80",
          6744 => x"88",
          6745 => x"52",
          6746 => x"34",
          6747 => x"34",
          6748 => x"04",
          6749 => x"87",
          6750 => x"8b",
          6751 => x"2b",
          6752 => x"84",
          6753 => x"17",
          6754 => x"2b",
          6755 => x"2a",
          6756 => x"51",
          6757 => x"71",
          6758 => x"72",
          6759 => x"84",
          6760 => x"70",
          6761 => x"33",
          6762 => x"71",
          6763 => x"83",
          6764 => x"5a",
          6765 => x"05",
          6766 => x"87",
          6767 => x"88",
          6768 => x"88",
          6769 => x"59",
          6770 => x"13",
          6771 => x"13",
          6772 => x"fc",
          6773 => x"33",
          6774 => x"71",
          6775 => x"81",
          6776 => x"70",
          6777 => x"5a",
          6778 => x"72",
          6779 => x"13",
          6780 => x"fc",
          6781 => x"70",
          6782 => x"33",
          6783 => x"71",
          6784 => x"74",
          6785 => x"81",
          6786 => x"88",
          6787 => x"83",
          6788 => x"f8",
          6789 => x"7b",
          6790 => x"52",
          6791 => x"5a",
          6792 => x"77",
          6793 => x"73",
          6794 => x"84",
          6795 => x"70",
          6796 => x"81",
          6797 => x"8b",
          6798 => x"2b",
          6799 => x"70",
          6800 => x"33",
          6801 => x"07",
          6802 => x"06",
          6803 => x"5f",
          6804 => x"5a",
          6805 => x"77",
          6806 => x"81",
          6807 => x"b9",
          6808 => x"17",
          6809 => x"83",
          6810 => x"8b",
          6811 => x"2b",
          6812 => x"70",
          6813 => x"33",
          6814 => x"71",
          6815 => x"58",
          6816 => x"5a",
          6817 => x"70",
          6818 => x"e4",
          6819 => x"81",
          6820 => x"88",
          6821 => x"80",
          6822 => x"88",
          6823 => x"54",
          6824 => x"77",
          6825 => x"84",
          6826 => x"70",
          6827 => x"81",
          6828 => x"8b",
          6829 => x"2b",
          6830 => x"82",
          6831 => x"15",
          6832 => x"2b",
          6833 => x"2a",
          6834 => x"52",
          6835 => x"53",
          6836 => x"34",
          6837 => x"34",
          6838 => x"04",
          6839 => x"79",
          6840 => x"08",
          6841 => x"80",
          6842 => x"77",
          6843 => x"38",
          6844 => x"90",
          6845 => x"0d",
          6846 => x"f4",
          6847 => x"fc",
          6848 => x"0b",
          6849 => x"23",
          6850 => x"53",
          6851 => x"ff",
          6852 => x"d2",
          6853 => x"b9",
          6854 => x"76",
          6855 => x"0b",
          6856 => x"84",
          6857 => x"54",
          6858 => x"34",
          6859 => x"15",
          6860 => x"fc",
          6861 => x"86",
          6862 => x"0b",
          6863 => x"84",
          6864 => x"84",
          6865 => x"ff",
          6866 => x"80",
          6867 => x"ff",
          6868 => x"88",
          6869 => x"55",
          6870 => x"17",
          6871 => x"17",
          6872 => x"f8",
          6873 => x"10",
          6874 => x"fc",
          6875 => x"05",
          6876 => x"82",
          6877 => x"0b",
          6878 => x"fe",
          6879 => x"3d",
          6880 => x"80",
          6881 => x"84",
          6882 => x"38",
          6883 => x"2a",
          6884 => x"83",
          6885 => x"51",
          6886 => x"ff",
          6887 => x"b9",
          6888 => x"11",
          6889 => x"33",
          6890 => x"07",
          6891 => x"5a",
          6892 => x"ff",
          6893 => x"80",
          6894 => x"38",
          6895 => x"10",
          6896 => x"81",
          6897 => x"88",
          6898 => x"81",
          6899 => x"79",
          6900 => x"ff",
          6901 => x"7a",
          6902 => x"5c",
          6903 => x"72",
          6904 => x"38",
          6905 => x"85",
          6906 => x"55",
          6907 => x"33",
          6908 => x"71",
          6909 => x"57",
          6910 => x"38",
          6911 => x"ff",
          6912 => x"77",
          6913 => x"80",
          6914 => x"78",
          6915 => x"81",
          6916 => x"88",
          6917 => x"81",
          6918 => x"56",
          6919 => x"59",
          6920 => x"2e",
          6921 => x"59",
          6922 => x"73",
          6923 => x"38",
          6924 => x"80",
          6925 => x"38",
          6926 => x"82",
          6927 => x"16",
          6928 => x"78",
          6929 => x"80",
          6930 => x"88",
          6931 => x"56",
          6932 => x"74",
          6933 => x"15",
          6934 => x"fc",
          6935 => x"88",
          6936 => x"71",
          6937 => x"75",
          6938 => x"84",
          6939 => x"70",
          6940 => x"81",
          6941 => x"88",
          6942 => x"83",
          6943 => x"f8",
          6944 => x"7e",
          6945 => x"06",
          6946 => x"5c",
          6947 => x"59",
          6948 => x"82",
          6949 => x"81",
          6950 => x"72",
          6951 => x"84",
          6952 => x"18",
          6953 => x"34",
          6954 => x"34",
          6955 => x"08",
          6956 => x"11",
          6957 => x"33",
          6958 => x"71",
          6959 => x"74",
          6960 => x"5c",
          6961 => x"84",
          6962 => x"85",
          6963 => x"b9",
          6964 => x"16",
          6965 => x"86",
          6966 => x"12",
          6967 => x"2b",
          6968 => x"2a",
          6969 => x"59",
          6970 => x"34",
          6971 => x"34",
          6972 => x"08",
          6973 => x"11",
          6974 => x"33",
          6975 => x"71",
          6976 => x"74",
          6977 => x"5c",
          6978 => x"86",
          6979 => x"87",
          6980 => x"b9",
          6981 => x"16",
          6982 => x"84",
          6983 => x"12",
          6984 => x"2b",
          6985 => x"2a",
          6986 => x"59",
          6987 => x"34",
          6988 => x"34",
          6989 => x"08",
          6990 => x"51",
          6991 => x"8c",
          6992 => x"0d",
          6993 => x"33",
          6994 => x"71",
          6995 => x"83",
          6996 => x"05",
          6997 => x"85",
          6998 => x"88",
          6999 => x"88",
          7000 => x"59",
          7001 => x"74",
          7002 => x"76",
          7003 => x"84",
          7004 => x"70",
          7005 => x"33",
          7006 => x"71",
          7007 => x"83",
          7008 => x"05",
          7009 => x"87",
          7010 => x"88",
          7011 => x"88",
          7012 => x"5f",
          7013 => x"57",
          7014 => x"1a",
          7015 => x"1a",
          7016 => x"fc",
          7017 => x"33",
          7018 => x"71",
          7019 => x"81",
          7020 => x"70",
          7021 => x"57",
          7022 => x"77",
          7023 => x"18",
          7024 => x"fc",
          7025 => x"05",
          7026 => x"39",
          7027 => x"79",
          7028 => x"08",
          7029 => x"80",
          7030 => x"77",
          7031 => x"38",
          7032 => x"8c",
          7033 => x"0d",
          7034 => x"fb",
          7035 => x"ba",
          7036 => x"ba",
          7037 => x"3d",
          7038 => x"ff",
          7039 => x"b9",
          7040 => x"80",
          7041 => x"f8",
          7042 => x"80",
          7043 => x"84",
          7044 => x"fe",
          7045 => x"84",
          7046 => x"55",
          7047 => x"81",
          7048 => x"34",
          7049 => x"08",
          7050 => x"15",
          7051 => x"85",
          7052 => x"b9",
          7053 => x"76",
          7054 => x"81",
          7055 => x"34",
          7056 => x"08",
          7057 => x"22",
          7058 => x"80",
          7059 => x"83",
          7060 => x"70",
          7061 => x"51",
          7062 => x"88",
          7063 => x"89",
          7064 => x"b9",
          7065 => x"10",
          7066 => x"b9",
          7067 => x"f8",
          7068 => x"76",
          7069 => x"81",
          7070 => x"34",
          7071 => x"80",
          7072 => x"38",
          7073 => x"ed",
          7074 => x"67",
          7075 => x"70",
          7076 => x"08",
          7077 => x"76",
          7078 => x"aa",
          7079 => x"2e",
          7080 => x"7f",
          7081 => x"d7",
          7082 => x"84",
          7083 => x"38",
          7084 => x"83",
          7085 => x"70",
          7086 => x"06",
          7087 => x"83",
          7088 => x"7f",
          7089 => x"2a",
          7090 => x"ff",
          7091 => x"2b",
          7092 => x"33",
          7093 => x"71",
          7094 => x"70",
          7095 => x"83",
          7096 => x"70",
          7097 => x"fc",
          7098 => x"2b",
          7099 => x"33",
          7100 => x"71",
          7101 => x"70",
          7102 => x"90",
          7103 => x"45",
          7104 => x"54",
          7105 => x"48",
          7106 => x"5f",
          7107 => x"24",
          7108 => x"82",
          7109 => x"16",
          7110 => x"2b",
          7111 => x"10",
          7112 => x"33",
          7113 => x"71",
          7114 => x"90",
          7115 => x"5c",
          7116 => x"56",
          7117 => x"85",
          7118 => x"62",
          7119 => x"38",
          7120 => x"77",
          7121 => x"a2",
          7122 => x"2e",
          7123 => x"60",
          7124 => x"62",
          7125 => x"38",
          7126 => x"61",
          7127 => x"f7",
          7128 => x"70",
          7129 => x"33",
          7130 => x"71",
          7131 => x"7a",
          7132 => x"81",
          7133 => x"98",
          7134 => x"2b",
          7135 => x"59",
          7136 => x"5b",
          7137 => x"24",
          7138 => x"76",
          7139 => x"33",
          7140 => x"71",
          7141 => x"83",
          7142 => x"11",
          7143 => x"87",
          7144 => x"8b",
          7145 => x"2b",
          7146 => x"84",
          7147 => x"15",
          7148 => x"2b",
          7149 => x"2a",
          7150 => x"52",
          7151 => x"53",
          7152 => x"77",
          7153 => x"79",
          7154 => x"84",
          7155 => x"70",
          7156 => x"33",
          7157 => x"71",
          7158 => x"83",
          7159 => x"05",
          7160 => x"87",
          7161 => x"88",
          7162 => x"88",
          7163 => x"5e",
          7164 => x"41",
          7165 => x"16",
          7166 => x"16",
          7167 => x"fc",
          7168 => x"33",
          7169 => x"71",
          7170 => x"81",
          7171 => x"70",
          7172 => x"5c",
          7173 => x"79",
          7174 => x"1a",
          7175 => x"fc",
          7176 => x"82",
          7177 => x"12",
          7178 => x"2b",
          7179 => x"07",
          7180 => x"33",
          7181 => x"71",
          7182 => x"70",
          7183 => x"5c",
          7184 => x"5a",
          7185 => x"79",
          7186 => x"1a",
          7187 => x"fc",
          7188 => x"70",
          7189 => x"33",
          7190 => x"71",
          7191 => x"74",
          7192 => x"33",
          7193 => x"71",
          7194 => x"70",
          7195 => x"5c",
          7196 => x"5a",
          7197 => x"82",
          7198 => x"83",
          7199 => x"b9",
          7200 => x"1f",
          7201 => x"83",
          7202 => x"88",
          7203 => x"57",
          7204 => x"83",
          7205 => x"5a",
          7206 => x"84",
          7207 => x"c4",
          7208 => x"b9",
          7209 => x"84",
          7210 => x"05",
          7211 => x"ff",
          7212 => x"44",
          7213 => x"26",
          7214 => x"7e",
          7215 => x"ba",
          7216 => x"3d",
          7217 => x"ff",
          7218 => x"b9",
          7219 => x"80",
          7220 => x"f8",
          7221 => x"80",
          7222 => x"84",
          7223 => x"fe",
          7224 => x"84",
          7225 => x"5e",
          7226 => x"81",
          7227 => x"34",
          7228 => x"08",
          7229 => x"1e",
          7230 => x"85",
          7231 => x"b9",
          7232 => x"60",
          7233 => x"81",
          7234 => x"34",
          7235 => x"08",
          7236 => x"22",
          7237 => x"80",
          7238 => x"83",
          7239 => x"70",
          7240 => x"5a",
          7241 => x"88",
          7242 => x"89",
          7243 => x"b9",
          7244 => x"10",
          7245 => x"b9",
          7246 => x"f8",
          7247 => x"60",
          7248 => x"81",
          7249 => x"34",
          7250 => x"08",
          7251 => x"d3",
          7252 => x"2e",
          7253 => x"7e",
          7254 => x"2e",
          7255 => x"7f",
          7256 => x"3f",
          7257 => x"08",
          7258 => x"0c",
          7259 => x"04",
          7260 => x"b9",
          7261 => x"83",
          7262 => x"5e",
          7263 => x"70",
          7264 => x"33",
          7265 => x"07",
          7266 => x"06",
          7267 => x"48",
          7268 => x"40",
          7269 => x"60",
          7270 => x"61",
          7271 => x"08",
          7272 => x"2a",
          7273 => x"82",
          7274 => x"83",
          7275 => x"b9",
          7276 => x"1f",
          7277 => x"12",
          7278 => x"2b",
          7279 => x"2b",
          7280 => x"06",
          7281 => x"83",
          7282 => x"70",
          7283 => x"5c",
          7284 => x"5b",
          7285 => x"82",
          7286 => x"81",
          7287 => x"60",
          7288 => x"34",
          7289 => x"08",
          7290 => x"7b",
          7291 => x"1c",
          7292 => x"b9",
          7293 => x"84",
          7294 => x"88",
          7295 => x"fd",
          7296 => x"75",
          7297 => x"ff",
          7298 => x"54",
          7299 => x"77",
          7300 => x"06",
          7301 => x"83",
          7302 => x"82",
          7303 => x"18",
          7304 => x"2b",
          7305 => x"10",
          7306 => x"33",
          7307 => x"71",
          7308 => x"90",
          7309 => x"5e",
          7310 => x"58",
          7311 => x"80",
          7312 => x"38",
          7313 => x"61",
          7314 => x"83",
          7315 => x"24",
          7316 => x"77",
          7317 => x"06",
          7318 => x"27",
          7319 => x"fe",
          7320 => x"ff",
          7321 => x"b9",
          7322 => x"80",
          7323 => x"f8",
          7324 => x"80",
          7325 => x"84",
          7326 => x"fe",
          7327 => x"84",
          7328 => x"5a",
          7329 => x"81",
          7330 => x"34",
          7331 => x"08",
          7332 => x"1a",
          7333 => x"85",
          7334 => x"b9",
          7335 => x"7e",
          7336 => x"81",
          7337 => x"34",
          7338 => x"08",
          7339 => x"22",
          7340 => x"80",
          7341 => x"83",
          7342 => x"70",
          7343 => x"56",
          7344 => x"64",
          7345 => x"73",
          7346 => x"34",
          7347 => x"22",
          7348 => x"10",
          7349 => x"08",
          7350 => x"42",
          7351 => x"82",
          7352 => x"61",
          7353 => x"fc",
          7354 => x"7a",
          7355 => x"38",
          7356 => x"ff",
          7357 => x"7b",
          7358 => x"38",
          7359 => x"76",
          7360 => x"bd",
          7361 => x"ea",
          7362 => x"54",
          7363 => x"8c",
          7364 => x"0d",
          7365 => x"82",
          7366 => x"12",
          7367 => x"2b",
          7368 => x"07",
          7369 => x"11",
          7370 => x"33",
          7371 => x"71",
          7372 => x"7e",
          7373 => x"33",
          7374 => x"71",
          7375 => x"70",
          7376 => x"44",
          7377 => x"46",
          7378 => x"45",
          7379 => x"84",
          7380 => x"64",
          7381 => x"84",
          7382 => x"70",
          7383 => x"33",
          7384 => x"71",
          7385 => x"83",
          7386 => x"05",
          7387 => x"87",
          7388 => x"88",
          7389 => x"88",
          7390 => x"42",
          7391 => x"5d",
          7392 => x"86",
          7393 => x"64",
          7394 => x"84",
          7395 => x"16",
          7396 => x"12",
          7397 => x"2b",
          7398 => x"ff",
          7399 => x"2a",
          7400 => x"5d",
          7401 => x"79",
          7402 => x"84",
          7403 => x"70",
          7404 => x"33",
          7405 => x"71",
          7406 => x"83",
          7407 => x"05",
          7408 => x"15",
          7409 => x"2b",
          7410 => x"2a",
          7411 => x"40",
          7412 => x"54",
          7413 => x"75",
          7414 => x"84",
          7415 => x"70",
          7416 => x"81",
          7417 => x"8b",
          7418 => x"2b",
          7419 => x"82",
          7420 => x"15",
          7421 => x"2b",
          7422 => x"2a",
          7423 => x"5b",
          7424 => x"55",
          7425 => x"34",
          7426 => x"34",
          7427 => x"08",
          7428 => x"11",
          7429 => x"33",
          7430 => x"07",
          7431 => x"56",
          7432 => x"42",
          7433 => x"7e",
          7434 => x"51",
          7435 => x"3f",
          7436 => x"08",
          7437 => x"78",
          7438 => x"06",
          7439 => x"99",
          7440 => x"f4",
          7441 => x"fc",
          7442 => x"0b",
          7443 => x"23",
          7444 => x"53",
          7445 => x"ff",
          7446 => x"c0",
          7447 => x"b9",
          7448 => x"7f",
          7449 => x"0b",
          7450 => x"84",
          7451 => x"55",
          7452 => x"34",
          7453 => x"16",
          7454 => x"fc",
          7455 => x"86",
          7456 => x"0b",
          7457 => x"84",
          7458 => x"84",
          7459 => x"ff",
          7460 => x"80",
          7461 => x"ff",
          7462 => x"88",
          7463 => x"44",
          7464 => x"1f",
          7465 => x"1f",
          7466 => x"f8",
          7467 => x"10",
          7468 => x"fc",
          7469 => x"05",
          7470 => x"82",
          7471 => x"0b",
          7472 => x"7e",
          7473 => x"3f",
          7474 => x"c0",
          7475 => x"33",
          7476 => x"71",
          7477 => x"83",
          7478 => x"05",
          7479 => x"85",
          7480 => x"88",
          7481 => x"88",
          7482 => x"5e",
          7483 => x"76",
          7484 => x"34",
          7485 => x"05",
          7486 => x"fc",
          7487 => x"84",
          7488 => x"12",
          7489 => x"2b",
          7490 => x"07",
          7491 => x"14",
          7492 => x"33",
          7493 => x"07",
          7494 => x"41",
          7495 => x"59",
          7496 => x"79",
          7497 => x"34",
          7498 => x"05",
          7499 => x"fc",
          7500 => x"33",
          7501 => x"71",
          7502 => x"81",
          7503 => x"70",
          7504 => x"42",
          7505 => x"78",
          7506 => x"19",
          7507 => x"fc",
          7508 => x"70",
          7509 => x"33",
          7510 => x"71",
          7511 => x"74",
          7512 => x"81",
          7513 => x"88",
          7514 => x"83",
          7515 => x"f8",
          7516 => x"63",
          7517 => x"5d",
          7518 => x"40",
          7519 => x"7f",
          7520 => x"7b",
          7521 => x"84",
          7522 => x"70",
          7523 => x"81",
          7524 => x"8b",
          7525 => x"2b",
          7526 => x"70",
          7527 => x"33",
          7528 => x"07",
          7529 => x"06",
          7530 => x"48",
          7531 => x"46",
          7532 => x"60",
          7533 => x"60",
          7534 => x"61",
          7535 => x"06",
          7536 => x"39",
          7537 => x"87",
          7538 => x"8b",
          7539 => x"2b",
          7540 => x"84",
          7541 => x"19",
          7542 => x"2b",
          7543 => x"2a",
          7544 => x"52",
          7545 => x"84",
          7546 => x"85",
          7547 => x"b9",
          7548 => x"19",
          7549 => x"85",
          7550 => x"8b",
          7551 => x"2b",
          7552 => x"86",
          7553 => x"15",
          7554 => x"2b",
          7555 => x"2a",
          7556 => x"52",
          7557 => x"56",
          7558 => x"05",
          7559 => x"87",
          7560 => x"b9",
          7561 => x"70",
          7562 => x"33",
          7563 => x"07",
          7564 => x"06",
          7565 => x"5b",
          7566 => x"77",
          7567 => x"81",
          7568 => x"b9",
          7569 => x"1f",
          7570 => x"12",
          7571 => x"2b",
          7572 => x"07",
          7573 => x"33",
          7574 => x"71",
          7575 => x"70",
          7576 => x"ff",
          7577 => x"05",
          7578 => x"56",
          7579 => x"58",
          7580 => x"55",
          7581 => x"34",
          7582 => x"34",
          7583 => x"08",
          7584 => x"33",
          7585 => x"71",
          7586 => x"83",
          7587 => x"05",
          7588 => x"12",
          7589 => x"2b",
          7590 => x"ff",
          7591 => x"2a",
          7592 => x"58",
          7593 => x"55",
          7594 => x"76",
          7595 => x"84",
          7596 => x"70",
          7597 => x"33",
          7598 => x"71",
          7599 => x"83",
          7600 => x"11",
          7601 => x"87",
          7602 => x"8b",
          7603 => x"2b",
          7604 => x"84",
          7605 => x"15",
          7606 => x"2b",
          7607 => x"2a",
          7608 => x"52",
          7609 => x"53",
          7610 => x"57",
          7611 => x"34",
          7612 => x"34",
          7613 => x"08",
          7614 => x"11",
          7615 => x"33",
          7616 => x"71",
          7617 => x"74",
          7618 => x"33",
          7619 => x"71",
          7620 => x"70",
          7621 => x"42",
          7622 => x"57",
          7623 => x"86",
          7624 => x"87",
          7625 => x"b9",
          7626 => x"70",
          7627 => x"33",
          7628 => x"07",
          7629 => x"06",
          7630 => x"5a",
          7631 => x"76",
          7632 => x"81",
          7633 => x"b9",
          7634 => x"1f",
          7635 => x"83",
          7636 => x"8b",
          7637 => x"2b",
          7638 => x"73",
          7639 => x"33",
          7640 => x"07",
          7641 => x"41",
          7642 => x"5f",
          7643 => x"79",
          7644 => x"81",
          7645 => x"b9",
          7646 => x"1f",
          7647 => x"12",
          7648 => x"2b",
          7649 => x"07",
          7650 => x"14",
          7651 => x"33",
          7652 => x"07",
          7653 => x"41",
          7654 => x"5f",
          7655 => x"79",
          7656 => x"75",
          7657 => x"84",
          7658 => x"70",
          7659 => x"33",
          7660 => x"71",
          7661 => x"66",
          7662 => x"70",
          7663 => x"52",
          7664 => x"05",
          7665 => x"fe",
          7666 => x"84",
          7667 => x"1e",
          7668 => x"65",
          7669 => x"83",
          7670 => x"5d",
          7671 => x"d5",
          7672 => x"33",
          7673 => x"71",
          7674 => x"83",
          7675 => x"05",
          7676 => x"85",
          7677 => x"88",
          7678 => x"88",
          7679 => x"5d",
          7680 => x"7a",
          7681 => x"34",
          7682 => x"05",
          7683 => x"fc",
          7684 => x"84",
          7685 => x"12",
          7686 => x"2b",
          7687 => x"07",
          7688 => x"14",
          7689 => x"33",
          7690 => x"07",
          7691 => x"5b",
          7692 => x"5c",
          7693 => x"73",
          7694 => x"34",
          7695 => x"05",
          7696 => x"fc",
          7697 => x"33",
          7698 => x"71",
          7699 => x"81",
          7700 => x"70",
          7701 => x"5f",
          7702 => x"75",
          7703 => x"16",
          7704 => x"fc",
          7705 => x"70",
          7706 => x"33",
          7707 => x"71",
          7708 => x"74",
          7709 => x"81",
          7710 => x"88",
          7711 => x"83",
          7712 => x"f8",
          7713 => x"63",
          7714 => x"44",
          7715 => x"5e",
          7716 => x"74",
          7717 => x"7b",
          7718 => x"84",
          7719 => x"70",
          7720 => x"81",
          7721 => x"8b",
          7722 => x"2b",
          7723 => x"70",
          7724 => x"33",
          7725 => x"07",
          7726 => x"06",
          7727 => x"47",
          7728 => x"46",
          7729 => x"7f",
          7730 => x"81",
          7731 => x"83",
          7732 => x"5b",
          7733 => x"7e",
          7734 => x"e5",
          7735 => x"ba",
          7736 => x"84",
          7737 => x"80",
          7738 => x"62",
          7739 => x"84",
          7740 => x"51",
          7741 => x"3f",
          7742 => x"88",
          7743 => x"61",
          7744 => x"b7",
          7745 => x"39",
          7746 => x"7a",
          7747 => x"b9",
          7748 => x"58",
          7749 => x"b7",
          7750 => x"77",
          7751 => x"84",
          7752 => x"89",
          7753 => x"77",
          7754 => x"3f",
          7755 => x"08",
          7756 => x"8c",
          7757 => x"e6",
          7758 => x"80",
          7759 => x"8c",
          7760 => x"b6",
          7761 => x"84",
          7762 => x"89",
          7763 => x"84",
          7764 => x"84",
          7765 => x"a0",
          7766 => x"b9",
          7767 => x"80",
          7768 => x"52",
          7769 => x"51",
          7770 => x"3f",
          7771 => x"08",
          7772 => x"34",
          7773 => x"16",
          7774 => x"fc",
          7775 => x"84",
          7776 => x"0b",
          7777 => x"84",
          7778 => x"56",
          7779 => x"34",
          7780 => x"17",
          7781 => x"fc",
          7782 => x"f8",
          7783 => x"fe",
          7784 => x"70",
          7785 => x"06",
          7786 => x"58",
          7787 => x"74",
          7788 => x"73",
          7789 => x"84",
          7790 => x"70",
          7791 => x"84",
          7792 => x"05",
          7793 => x"55",
          7794 => x"34",
          7795 => x"15",
          7796 => x"77",
          7797 => x"c6",
          7798 => x"39",
          7799 => x"02",
          7800 => x"51",
          7801 => x"72",
          7802 => x"84",
          7803 => x"33",
          7804 => x"ba",
          7805 => x"3d",
          7806 => x"3d",
          7807 => x"05",
          7808 => x"53",
          7809 => x"9d",
          7810 => x"d3",
          7811 => x"ba",
          7812 => x"ff",
          7813 => x"87",
          7814 => x"ba",
          7815 => x"84",
          7816 => x"33",
          7817 => x"ba",
          7818 => x"3d",
          7819 => x"3d",
          7820 => x"60",
          7821 => x"af",
          7822 => x"5c",
          7823 => x"54",
          7824 => x"87",
          7825 => x"88",
          7826 => x"73",
          7827 => x"83",
          7828 => x"38",
          7829 => x"0b",
          7830 => x"8c",
          7831 => x"75",
          7832 => x"d5",
          7833 => x"ba",
          7834 => x"ff",
          7835 => x"80",
          7836 => x"87",
          7837 => x"08",
          7838 => x"38",
          7839 => x"d6",
          7840 => x"80",
          7841 => x"73",
          7842 => x"38",
          7843 => x"55",
          7844 => x"8c",
          7845 => x"0d",
          7846 => x"16",
          7847 => x"81",
          7848 => x"55",
          7849 => x"26",
          7850 => x"d5",
          7851 => x"0d",
          7852 => x"02",
          7853 => x"05",
          7854 => x"57",
          7855 => x"76",
          7856 => x"38",
          7857 => x"17",
          7858 => x"81",
          7859 => x"55",
          7860 => x"73",
          7861 => x"87",
          7862 => x"0c",
          7863 => x"52",
          7864 => x"e7",
          7865 => x"8c",
          7866 => x"06",
          7867 => x"2e",
          7868 => x"c0",
          7869 => x"54",
          7870 => x"79",
          7871 => x"38",
          7872 => x"80",
          7873 => x"80",
          7874 => x"81",
          7875 => x"74",
          7876 => x"0c",
          7877 => x"04",
          7878 => x"81",
          7879 => x"ff",
          7880 => x"56",
          7881 => x"ff",
          7882 => x"39",
          7883 => x"78",
          7884 => x"9b",
          7885 => x"88",
          7886 => x"33",
          7887 => x"81",
          7888 => x"26",
          7889 => x"ba",
          7890 => x"53",
          7891 => x"54",
          7892 => x"9b",
          7893 => x"87",
          7894 => x"0c",
          7895 => x"73",
          7896 => x"72",
          7897 => x"38",
          7898 => x"9a",
          7899 => x"72",
          7900 => x"0c",
          7901 => x"04",
          7902 => x"75",
          7903 => x"ba",
          7904 => x"3d",
          7905 => x"80",
          7906 => x"0b",
          7907 => x"0c",
          7908 => x"04",
          7909 => x"87",
          7910 => x"11",
          7911 => x"cd",
          7912 => x"70",
          7913 => x"06",
          7914 => x"80",
          7915 => x"87",
          7916 => x"08",
          7917 => x"38",
          7918 => x"8c",
          7919 => x"ca",
          7920 => x"0c",
          7921 => x"8c",
          7922 => x"08",
          7923 => x"73",
          7924 => x"9b",
          7925 => x"82",
          7926 => x"ee",
          7927 => x"39",
          7928 => x"7c",
          7929 => x"83",
          7930 => x"5b",
          7931 => x"77",
          7932 => x"06",
          7933 => x"33",
          7934 => x"2e",
          7935 => x"80",
          7936 => x"81",
          7937 => x"fe",
          7938 => x"ba",
          7939 => x"2e",
          7940 => x"59",
          7941 => x"8c",
          7942 => x"0d",
          7943 => x"b4",
          7944 => x"b8",
          7945 => x"81",
          7946 => x"5a",
          7947 => x"81",
          7948 => x"8c",
          7949 => x"09",
          7950 => x"38",
          7951 => x"08",
          7952 => x"b4",
          7953 => x"a8",
          7954 => x"a0",
          7955 => x"ba",
          7956 => x"58",
          7957 => x"76",
          7958 => x"38",
          7959 => x"55",
          7960 => x"09",
          7961 => x"8e",
          7962 => x"75",
          7963 => x"52",
          7964 => x"51",
          7965 => x"76",
          7966 => x"59",
          7967 => x"09",
          7968 => x"fb",
          7969 => x"33",
          7970 => x"2e",
          7971 => x"fe",
          7972 => x"18",
          7973 => x"7a",
          7974 => x"75",
          7975 => x"57",
          7976 => x"57",
          7977 => x"80",
          7978 => x"b6",
          7979 => x"aa",
          7980 => x"19",
          7981 => x"7a",
          7982 => x"0b",
          7983 => x"80",
          7984 => x"19",
          7985 => x"0b",
          7986 => x"80",
          7987 => x"9c",
          7988 => x"f2",
          7989 => x"19",
          7990 => x"0b",
          7991 => x"34",
          7992 => x"84",
          7993 => x"94",
          7994 => x"74",
          7995 => x"34",
          7996 => x"5b",
          7997 => x"19",
          7998 => x"2a",
          7999 => x"a2",
          8000 => x"98",
          8001 => x"84",
          8002 => x"90",
          8003 => x"7a",
          8004 => x"34",
          8005 => x"55",
          8006 => x"19",
          8007 => x"2a",
          8008 => x"a6",
          8009 => x"98",
          8010 => x"84",
          8011 => x"a4",
          8012 => x"05",
          8013 => x"0c",
          8014 => x"7a",
          8015 => x"81",
          8016 => x"fa",
          8017 => x"84",
          8018 => x"53",
          8019 => x"18",
          8020 => x"d8",
          8021 => x"8c",
          8022 => x"fd",
          8023 => x"b2",
          8024 => x"0d",
          8025 => x"08",
          8026 => x"81",
          8027 => x"38",
          8028 => x"76",
          8029 => x"81",
          8030 => x"ba",
          8031 => x"3d",
          8032 => x"77",
          8033 => x"74",
          8034 => x"cc",
          8035 => x"24",
          8036 => x"74",
          8037 => x"81",
          8038 => x"75",
          8039 => x"70",
          8040 => x"19",
          8041 => x"5a",
          8042 => x"17",
          8043 => x"b0",
          8044 => x"33",
          8045 => x"2e",
          8046 => x"83",
          8047 => x"54",
          8048 => x"17",
          8049 => x"33",
          8050 => x"3f",
          8051 => x"08",
          8052 => x"38",
          8053 => x"5b",
          8054 => x"0c",
          8055 => x"38",
          8056 => x"06",
          8057 => x"33",
          8058 => x"89",
          8059 => x"08",
          8060 => x"5d",
          8061 => x"08",
          8062 => x"38",
          8063 => x"18",
          8064 => x"56",
          8065 => x"2e",
          8066 => x"84",
          8067 => x"54",
          8068 => x"17",
          8069 => x"33",
          8070 => x"3f",
          8071 => x"08",
          8072 => x"38",
          8073 => x"5a",
          8074 => x"0c",
          8075 => x"38",
          8076 => x"06",
          8077 => x"33",
          8078 => x"7e",
          8079 => x"06",
          8080 => x"53",
          8081 => x"5d",
          8082 => x"38",
          8083 => x"06",
          8084 => x"0c",
          8085 => x"04",
          8086 => x"a8",
          8087 => x"59",
          8088 => x"79",
          8089 => x"80",
          8090 => x"33",
          8091 => x"5b",
          8092 => x"09",
          8093 => x"c2",
          8094 => x"78",
          8095 => x"52",
          8096 => x"51",
          8097 => x"84",
          8098 => x"80",
          8099 => x"ff",
          8100 => x"78",
          8101 => x"79",
          8102 => x"75",
          8103 => x"06",
          8104 => x"05",
          8105 => x"71",
          8106 => x"2b",
          8107 => x"8c",
          8108 => x"8f",
          8109 => x"74",
          8110 => x"81",
          8111 => x"38",
          8112 => x"a8",
          8113 => x"59",
          8114 => x"79",
          8115 => x"80",
          8116 => x"33",
          8117 => x"5b",
          8118 => x"09",
          8119 => x"81",
          8120 => x"78",
          8121 => x"52",
          8122 => x"51",
          8123 => x"84",
          8124 => x"80",
          8125 => x"ff",
          8126 => x"78",
          8127 => x"79",
          8128 => x"75",
          8129 => x"fc",
          8130 => x"b8",
          8131 => x"33",
          8132 => x"71",
          8133 => x"88",
          8134 => x"14",
          8135 => x"07",
          8136 => x"33",
          8137 => x"ff",
          8138 => x"07",
          8139 => x"0c",
          8140 => x"59",
          8141 => x"3d",
          8142 => x"54",
          8143 => x"53",
          8144 => x"53",
          8145 => x"52",
          8146 => x"3f",
          8147 => x"ba",
          8148 => x"2e",
          8149 => x"fe",
          8150 => x"ba",
          8151 => x"18",
          8152 => x"08",
          8153 => x"31",
          8154 => x"08",
          8155 => x"a0",
          8156 => x"fe",
          8157 => x"17",
          8158 => x"82",
          8159 => x"06",
          8160 => x"81",
          8161 => x"08",
          8162 => x"05",
          8163 => x"81",
          8164 => x"f6",
          8165 => x"5a",
          8166 => x"81",
          8167 => x"08",
          8168 => x"70",
          8169 => x"33",
          8170 => x"81",
          8171 => x"8c",
          8172 => x"09",
          8173 => x"81",
          8174 => x"8c",
          8175 => x"34",
          8176 => x"a8",
          8177 => x"5d",
          8178 => x"08",
          8179 => x"82",
          8180 => x"7d",
          8181 => x"cb",
          8182 => x"8c",
          8183 => x"de",
          8184 => x"b4",
          8185 => x"b8",
          8186 => x"81",
          8187 => x"5c",
          8188 => x"81",
          8189 => x"8c",
          8190 => x"09",
          8191 => x"ff",
          8192 => x"8c",
          8193 => x"34",
          8194 => x"a8",
          8195 => x"84",
          8196 => x"5b",
          8197 => x"18",
          8198 => x"c5",
          8199 => x"33",
          8200 => x"2e",
          8201 => x"fd",
          8202 => x"54",
          8203 => x"a0",
          8204 => x"53",
          8205 => x"17",
          8206 => x"f1",
          8207 => x"fd",
          8208 => x"54",
          8209 => x"53",
          8210 => x"53",
          8211 => x"52",
          8212 => x"3f",
          8213 => x"ba",
          8214 => x"2e",
          8215 => x"fb",
          8216 => x"ba",
          8217 => x"18",
          8218 => x"08",
          8219 => x"31",
          8220 => x"08",
          8221 => x"a0",
          8222 => x"fb",
          8223 => x"17",
          8224 => x"82",
          8225 => x"06",
          8226 => x"81",
          8227 => x"08",
          8228 => x"05",
          8229 => x"81",
          8230 => x"f4",
          8231 => x"5a",
          8232 => x"81",
          8233 => x"08",
          8234 => x"05",
          8235 => x"81",
          8236 => x"f3",
          8237 => x"86",
          8238 => x"7a",
          8239 => x"fa",
          8240 => x"3d",
          8241 => x"64",
          8242 => x"82",
          8243 => x"27",
          8244 => x"9c",
          8245 => x"95",
          8246 => x"55",
          8247 => x"96",
          8248 => x"24",
          8249 => x"74",
          8250 => x"8a",
          8251 => x"ba",
          8252 => x"3d",
          8253 => x"88",
          8254 => x"08",
          8255 => x"0b",
          8256 => x"58",
          8257 => x"2e",
          8258 => x"83",
          8259 => x"5b",
          8260 => x"2e",
          8261 => x"83",
          8262 => x"54",
          8263 => x"19",
          8264 => x"33",
          8265 => x"3f",
          8266 => x"08",
          8267 => x"38",
          8268 => x"5a",
          8269 => x"0c",
          8270 => x"ff",
          8271 => x"10",
          8272 => x"79",
          8273 => x"ff",
          8274 => x"5e",
          8275 => x"34",
          8276 => x"5a",
          8277 => x"34",
          8278 => x"1a",
          8279 => x"ba",
          8280 => x"3d",
          8281 => x"83",
          8282 => x"06",
          8283 => x"75",
          8284 => x"1a",
          8285 => x"80",
          8286 => x"08",
          8287 => x"78",
          8288 => x"38",
          8289 => x"7c",
          8290 => x"7c",
          8291 => x"06",
          8292 => x"81",
          8293 => x"b8",
          8294 => x"19",
          8295 => x"8e",
          8296 => x"8c",
          8297 => x"85",
          8298 => x"81",
          8299 => x"1a",
          8300 => x"79",
          8301 => x"75",
          8302 => x"fc",
          8303 => x"b8",
          8304 => x"33",
          8305 => x"8f",
          8306 => x"f0",
          8307 => x"41",
          8308 => x"7d",
          8309 => x"88",
          8310 => x"b9",
          8311 => x"90",
          8312 => x"ba",
          8313 => x"98",
          8314 => x"bb",
          8315 => x"0b",
          8316 => x"fe",
          8317 => x"81",
          8318 => x"89",
          8319 => x"08",
          8320 => x"08",
          8321 => x"76",
          8322 => x"38",
          8323 => x"1a",
          8324 => x"56",
          8325 => x"2e",
          8326 => x"82",
          8327 => x"54",
          8328 => x"19",
          8329 => x"33",
          8330 => x"3f",
          8331 => x"08",
          8332 => x"38",
          8333 => x"5c",
          8334 => x"0c",
          8335 => x"fd",
          8336 => x"83",
          8337 => x"b8",
          8338 => x"77",
          8339 => x"5f",
          8340 => x"7c",
          8341 => x"38",
          8342 => x"9f",
          8343 => x"33",
          8344 => x"07",
          8345 => x"77",
          8346 => x"83",
          8347 => x"89",
          8348 => x"08",
          8349 => x"0b",
          8350 => x"56",
          8351 => x"2e",
          8352 => x"81",
          8353 => x"b8",
          8354 => x"81",
          8355 => x"57",
          8356 => x"81",
          8357 => x"8c",
          8358 => x"09",
          8359 => x"c7",
          8360 => x"8c",
          8361 => x"34",
          8362 => x"70",
          8363 => x"31",
          8364 => x"84",
          8365 => x"5b",
          8366 => x"74",
          8367 => x"38",
          8368 => x"55",
          8369 => x"82",
          8370 => x"54",
          8371 => x"52",
          8372 => x"51",
          8373 => x"84",
          8374 => x"80",
          8375 => x"ff",
          8376 => x"75",
          8377 => x"77",
          8378 => x"7d",
          8379 => x"19",
          8380 => x"84",
          8381 => x"7c",
          8382 => x"88",
          8383 => x"81",
          8384 => x"8f",
          8385 => x"5c",
          8386 => x"81",
          8387 => x"34",
          8388 => x"81",
          8389 => x"b8",
          8390 => x"81",
          8391 => x"5d",
          8392 => x"81",
          8393 => x"8c",
          8394 => x"09",
          8395 => x"88",
          8396 => x"8c",
          8397 => x"34",
          8398 => x"70",
          8399 => x"31",
          8400 => x"84",
          8401 => x"5d",
          8402 => x"7e",
          8403 => x"ca",
          8404 => x"33",
          8405 => x"2e",
          8406 => x"fb",
          8407 => x"54",
          8408 => x"7c",
          8409 => x"33",
          8410 => x"3f",
          8411 => x"aa",
          8412 => x"76",
          8413 => x"70",
          8414 => x"33",
          8415 => x"ad",
          8416 => x"84",
          8417 => x"7d",
          8418 => x"06",
          8419 => x"84",
          8420 => x"83",
          8421 => x"19",
          8422 => x"1b",
          8423 => x"1b",
          8424 => x"8c",
          8425 => x"56",
          8426 => x"27",
          8427 => x"82",
          8428 => x"74",
          8429 => x"81",
          8430 => x"38",
          8431 => x"1f",
          8432 => x"81",
          8433 => x"ed",
          8434 => x"5c",
          8435 => x"81",
          8436 => x"b8",
          8437 => x"81",
          8438 => x"57",
          8439 => x"81",
          8440 => x"8c",
          8441 => x"09",
          8442 => x"c5",
          8443 => x"8c",
          8444 => x"34",
          8445 => x"70",
          8446 => x"31",
          8447 => x"84",
          8448 => x"5d",
          8449 => x"7e",
          8450 => x"87",
          8451 => x"33",
          8452 => x"2e",
          8453 => x"fa",
          8454 => x"54",
          8455 => x"76",
          8456 => x"33",
          8457 => x"3f",
          8458 => x"e7",
          8459 => x"79",
          8460 => x"52",
          8461 => x"51",
          8462 => x"7e",
          8463 => x"39",
          8464 => x"83",
          8465 => x"05",
          8466 => x"ff",
          8467 => x"58",
          8468 => x"34",
          8469 => x"5a",
          8470 => x"34",
          8471 => x"7e",
          8472 => x"39",
          8473 => x"2b",
          8474 => x"7a",
          8475 => x"83",
          8476 => x"98",
          8477 => x"06",
          8478 => x"06",
          8479 => x"5f",
          8480 => x"7d",
          8481 => x"2a",
          8482 => x"1d",
          8483 => x"2a",
          8484 => x"1d",
          8485 => x"2a",
          8486 => x"1d",
          8487 => x"39",
          8488 => x"7c",
          8489 => x"5b",
          8490 => x"81",
          8491 => x"19",
          8492 => x"80",
          8493 => x"38",
          8494 => x"08",
          8495 => x"38",
          8496 => x"70",
          8497 => x"80",
          8498 => x"38",
          8499 => x"81",
          8500 => x"56",
          8501 => x"9c",
          8502 => x"26",
          8503 => x"56",
          8504 => x"82",
          8505 => x"52",
          8506 => x"f5",
          8507 => x"8c",
          8508 => x"81",
          8509 => x"58",
          8510 => x"08",
          8511 => x"38",
          8512 => x"08",
          8513 => x"70",
          8514 => x"25",
          8515 => x"51",
          8516 => x"73",
          8517 => x"75",
          8518 => x"81",
          8519 => x"38",
          8520 => x"84",
          8521 => x"8c",
          8522 => x"81",
          8523 => x"39",
          8524 => x"08",
          8525 => x"7a",
          8526 => x"f0",
          8527 => x"55",
          8528 => x"8c",
          8529 => x"38",
          8530 => x"08",
          8531 => x"8c",
          8532 => x"ce",
          8533 => x"08",
          8534 => x"08",
          8535 => x"7a",
          8536 => x"39",
          8537 => x"9c",
          8538 => x"26",
          8539 => x"56",
          8540 => x"51",
          8541 => x"80",
          8542 => x"8c",
          8543 => x"81",
          8544 => x"ba",
          8545 => x"70",
          8546 => x"07",
          8547 => x"7b",
          8548 => x"8c",
          8549 => x"51",
          8550 => x"ff",
          8551 => x"ba",
          8552 => x"2e",
          8553 => x"19",
          8554 => x"74",
          8555 => x"38",
          8556 => x"08",
          8557 => x"38",
          8558 => x"57",
          8559 => x"75",
          8560 => x"8e",
          8561 => x"75",
          8562 => x"f5",
          8563 => x"ba",
          8564 => x"ba",
          8565 => x"70",
          8566 => x"08",
          8567 => x"56",
          8568 => x"80",
          8569 => x"80",
          8570 => x"90",
          8571 => x"19",
          8572 => x"94",
          8573 => x"58",
          8574 => x"86",
          8575 => x"94",
          8576 => x"19",
          8577 => x"5a",
          8578 => x"34",
          8579 => x"84",
          8580 => x"8c",
          8581 => x"80",
          8582 => x"8c",
          8583 => x"0d",
          8584 => x"8c",
          8585 => x"da",
          8586 => x"2e",
          8587 => x"75",
          8588 => x"78",
          8589 => x"3f",
          8590 => x"08",
          8591 => x"39",
          8592 => x"08",
          8593 => x"0c",
          8594 => x"04",
          8595 => x"81",
          8596 => x"38",
          8597 => x"b6",
          8598 => x"0d",
          8599 => x"08",
          8600 => x"73",
          8601 => x"26",
          8602 => x"73",
          8603 => x"72",
          8604 => x"73",
          8605 => x"88",
          8606 => x"74",
          8607 => x"76",
          8608 => x"82",
          8609 => x"38",
          8610 => x"53",
          8611 => x"18",
          8612 => x"72",
          8613 => x"38",
          8614 => x"98",
          8615 => x"94",
          8616 => x"18",
          8617 => x"56",
          8618 => x"94",
          8619 => x"2a",
          8620 => x"0c",
          8621 => x"06",
          8622 => x"9c",
          8623 => x"56",
          8624 => x"8c",
          8625 => x"0d",
          8626 => x"84",
          8627 => x"8a",
          8628 => x"ac",
          8629 => x"74",
          8630 => x"ac",
          8631 => x"22",
          8632 => x"57",
          8633 => x"27",
          8634 => x"17",
          8635 => x"15",
          8636 => x"56",
          8637 => x"73",
          8638 => x"8a",
          8639 => x"71",
          8640 => x"08",
          8641 => x"78",
          8642 => x"ff",
          8643 => x"52",
          8644 => x"cd",
          8645 => x"8c",
          8646 => x"ba",
          8647 => x"2e",
          8648 => x"0b",
          8649 => x"08",
          8650 => x"38",
          8651 => x"53",
          8652 => x"08",
          8653 => x"91",
          8654 => x"31",
          8655 => x"27",
          8656 => x"aa",
          8657 => x"84",
          8658 => x"8a",
          8659 => x"f3",
          8660 => x"70",
          8661 => x"08",
          8662 => x"5a",
          8663 => x"0a",
          8664 => x"38",
          8665 => x"18",
          8666 => x"08",
          8667 => x"74",
          8668 => x"38",
          8669 => x"06",
          8670 => x"38",
          8671 => x"18",
          8672 => x"75",
          8673 => x"85",
          8674 => x"22",
          8675 => x"76",
          8676 => x"38",
          8677 => x"0c",
          8678 => x"0c",
          8679 => x"05",
          8680 => x"80",
          8681 => x"ba",
          8682 => x"3d",
          8683 => x"98",
          8684 => x"19",
          8685 => x"7a",
          8686 => x"5c",
          8687 => x"75",
          8688 => x"eb",
          8689 => x"ba",
          8690 => x"82",
          8691 => x"84",
          8692 => x"27",
          8693 => x"56",
          8694 => x"08",
          8695 => x"38",
          8696 => x"84",
          8697 => x"26",
          8698 => x"60",
          8699 => x"98",
          8700 => x"08",
          8701 => x"f9",
          8702 => x"ba",
          8703 => x"87",
          8704 => x"8c",
          8705 => x"ff",
          8706 => x"56",
          8707 => x"08",
          8708 => x"91",
          8709 => x"84",
          8710 => x"ff",
          8711 => x"38",
          8712 => x"08",
          8713 => x"5f",
          8714 => x"ea",
          8715 => x"9c",
          8716 => x"05",
          8717 => x"5c",
          8718 => x"8d",
          8719 => x"22",
          8720 => x"b0",
          8721 => x"5d",
          8722 => x"1a",
          8723 => x"58",
          8724 => x"57",
          8725 => x"70",
          8726 => x"34",
          8727 => x"74",
          8728 => x"56",
          8729 => x"55",
          8730 => x"81",
          8731 => x"54",
          8732 => x"77",
          8733 => x"33",
          8734 => x"3f",
          8735 => x"08",
          8736 => x"81",
          8737 => x"39",
          8738 => x"0c",
          8739 => x"ba",
          8740 => x"3d",
          8741 => x"54",
          8742 => x"53",
          8743 => x"53",
          8744 => x"52",
          8745 => x"3f",
          8746 => x"08",
          8747 => x"84",
          8748 => x"83",
          8749 => x"19",
          8750 => x"08",
          8751 => x"a0",
          8752 => x"fe",
          8753 => x"19",
          8754 => x"82",
          8755 => x"06",
          8756 => x"81",
          8757 => x"08",
          8758 => x"05",
          8759 => x"81",
          8760 => x"e3",
          8761 => x"c5",
          8762 => x"22",
          8763 => x"ff",
          8764 => x"74",
          8765 => x"81",
          8766 => x"7c",
          8767 => x"fe",
          8768 => x"08",
          8769 => x"56",
          8770 => x"7d",
          8771 => x"38",
          8772 => x"76",
          8773 => x"1b",
          8774 => x"19",
          8775 => x"f8",
          8776 => x"84",
          8777 => x"8f",
          8778 => x"ee",
          8779 => x"66",
          8780 => x"7c",
          8781 => x"81",
          8782 => x"1e",
          8783 => x"5e",
          8784 => x"82",
          8785 => x"19",
          8786 => x"80",
          8787 => x"08",
          8788 => x"d1",
          8789 => x"33",
          8790 => x"74",
          8791 => x"81",
          8792 => x"38",
          8793 => x"53",
          8794 => x"81",
          8795 => x"e1",
          8796 => x"ba",
          8797 => x"2e",
          8798 => x"5a",
          8799 => x"b4",
          8800 => x"5b",
          8801 => x"38",
          8802 => x"70",
          8803 => x"76",
          8804 => x"81",
          8805 => x"33",
          8806 => x"81",
          8807 => x"41",
          8808 => x"34",
          8809 => x"32",
          8810 => x"ae",
          8811 => x"72",
          8812 => x"80",
          8813 => x"45",
          8814 => x"74",
          8815 => x"7a",
          8816 => x"56",
          8817 => x"81",
          8818 => x"60",
          8819 => x"38",
          8820 => x"80",
          8821 => x"fa",
          8822 => x"ba",
          8823 => x"84",
          8824 => x"81",
          8825 => x"1c",
          8826 => x"fe",
          8827 => x"84",
          8828 => x"94",
          8829 => x"81",
          8830 => x"08",
          8831 => x"81",
          8832 => x"e1",
          8833 => x"57",
          8834 => x"08",
          8835 => x"81",
          8836 => x"38",
          8837 => x"08",
          8838 => x"b4",
          8839 => x"1a",
          8840 => x"ba",
          8841 => x"5b",
          8842 => x"08",
          8843 => x"38",
          8844 => x"41",
          8845 => x"09",
          8846 => x"a8",
          8847 => x"b4",
          8848 => x"1a",
          8849 => x"7e",
          8850 => x"33",
          8851 => x"3f",
          8852 => x"90",
          8853 => x"2e",
          8854 => x"81",
          8855 => x"86",
          8856 => x"5b",
          8857 => x"93",
          8858 => x"33",
          8859 => x"06",
          8860 => x"08",
          8861 => x"0c",
          8862 => x"76",
          8863 => x"38",
          8864 => x"74",
          8865 => x"39",
          8866 => x"60",
          8867 => x"06",
          8868 => x"c1",
          8869 => x"80",
          8870 => x"0c",
          8871 => x"8c",
          8872 => x"0d",
          8873 => x"fd",
          8874 => x"18",
          8875 => x"77",
          8876 => x"06",
          8877 => x"19",
          8878 => x"33",
          8879 => x"71",
          8880 => x"58",
          8881 => x"ff",
          8882 => x"33",
          8883 => x"06",
          8884 => x"05",
          8885 => x"76",
          8886 => x"e6",
          8887 => x"78",
          8888 => x"33",
          8889 => x"88",
          8890 => x"44",
          8891 => x"2e",
          8892 => x"79",
          8893 => x"ff",
          8894 => x"10",
          8895 => x"5c",
          8896 => x"23",
          8897 => x"81",
          8898 => x"77",
          8899 => x"77",
          8900 => x"2a",
          8901 => x"57",
          8902 => x"90",
          8903 => x"fe",
          8904 => x"38",
          8905 => x"05",
          8906 => x"23",
          8907 => x"81",
          8908 => x"41",
          8909 => x"75",
          8910 => x"2e",
          8911 => x"ff",
          8912 => x"39",
          8913 => x"7c",
          8914 => x"74",
          8915 => x"81",
          8916 => x"78",
          8917 => x"5a",
          8918 => x"05",
          8919 => x"06",
          8920 => x"56",
          8921 => x"38",
          8922 => x"fd",
          8923 => x"0b",
          8924 => x"7a",
          8925 => x"0c",
          8926 => x"04",
          8927 => x"63",
          8928 => x"5c",
          8929 => x"51",
          8930 => x"84",
          8931 => x"5a",
          8932 => x"08",
          8933 => x"81",
          8934 => x"5d",
          8935 => x"1d",
          8936 => x"5e",
          8937 => x"56",
          8938 => x"1b",
          8939 => x"82",
          8940 => x"1b",
          8941 => x"55",
          8942 => x"09",
          8943 => x"df",
          8944 => x"75",
          8945 => x"52",
          8946 => x"51",
          8947 => x"84",
          8948 => x"80",
          8949 => x"ff",
          8950 => x"75",
          8951 => x"76",
          8952 => x"b2",
          8953 => x"08",
          8954 => x"59",
          8955 => x"84",
          8956 => x"19",
          8957 => x"70",
          8958 => x"57",
          8959 => x"1d",
          8960 => x"e5",
          8961 => x"38",
          8962 => x"81",
          8963 => x"8f",
          8964 => x"38",
          8965 => x"38",
          8966 => x"81",
          8967 => x"aa",
          8968 => x"56",
          8969 => x"74",
          8970 => x"81",
          8971 => x"78",
          8972 => x"5a",
          8973 => x"05",
          8974 => x"06",
          8975 => x"56",
          8976 => x"38",
          8977 => x"80",
          8978 => x"1c",
          8979 => x"57",
          8980 => x"8b",
          8981 => x"59",
          8982 => x"81",
          8983 => x"78",
          8984 => x"5a",
          8985 => x"31",
          8986 => x"58",
          8987 => x"80",
          8988 => x"38",
          8989 => x"e1",
          8990 => x"5d",
          8991 => x"1d",
          8992 => x"7b",
          8993 => x"3f",
          8994 => x"08",
          8995 => x"8c",
          8996 => x"fe",
          8997 => x"84",
          8998 => x"93",
          8999 => x"81",
          9000 => x"08",
          9001 => x"81",
          9002 => x"dc",
          9003 => x"57",
          9004 => x"08",
          9005 => x"81",
          9006 => x"38",
          9007 => x"08",
          9008 => x"b4",
          9009 => x"1c",
          9010 => x"ba",
          9011 => x"59",
          9012 => x"08",
          9013 => x"38",
          9014 => x"5a",
          9015 => x"09",
          9016 => x"dd",
          9017 => x"b4",
          9018 => x"1c",
          9019 => x"7d",
          9020 => x"33",
          9021 => x"3f",
          9022 => x"c5",
          9023 => x"fd",
          9024 => x"1c",
          9025 => x"2a",
          9026 => x"55",
          9027 => x"38",
          9028 => x"81",
          9029 => x"80",
          9030 => x"8d",
          9031 => x"81",
          9032 => x"90",
          9033 => x"ac",
          9034 => x"5e",
          9035 => x"2e",
          9036 => x"ff",
          9037 => x"80",
          9038 => x"f4",
          9039 => x"ba",
          9040 => x"84",
          9041 => x"80",
          9042 => x"38",
          9043 => x"75",
          9044 => x"c2",
          9045 => x"5d",
          9046 => x"1d",
          9047 => x"39",
          9048 => x"57",
          9049 => x"09",
          9050 => x"38",
          9051 => x"9b",
          9052 => x"1b",
          9053 => x"2b",
          9054 => x"40",
          9055 => x"38",
          9056 => x"bf",
          9057 => x"f3",
          9058 => x"81",
          9059 => x"83",
          9060 => x"33",
          9061 => x"11",
          9062 => x"71",
          9063 => x"52",
          9064 => x"80",
          9065 => x"38",
          9066 => x"26",
          9067 => x"76",
          9068 => x"8a",
          9069 => x"8c",
          9070 => x"61",
          9071 => x"53",
          9072 => x"5b",
          9073 => x"f6",
          9074 => x"ba",
          9075 => x"09",
          9076 => x"de",
          9077 => x"81",
          9078 => x"78",
          9079 => x"38",
          9080 => x"86",
          9081 => x"56",
          9082 => x"2e",
          9083 => x"80",
          9084 => x"79",
          9085 => x"70",
          9086 => x"7f",
          9087 => x"ff",
          9088 => x"ff",
          9089 => x"fe",
          9090 => x"0b",
          9091 => x"0c",
          9092 => x"04",
          9093 => x"ff",
          9094 => x"38",
          9095 => x"fe",
          9096 => x"3d",
          9097 => x"08",
          9098 => x"33",
          9099 => x"58",
          9100 => x"86",
          9101 => x"b5",
          9102 => x"1d",
          9103 => x"57",
          9104 => x"80",
          9105 => x"81",
          9106 => x"17",
          9107 => x"56",
          9108 => x"38",
          9109 => x"1f",
          9110 => x"60",
          9111 => x"55",
          9112 => x"05",
          9113 => x"70",
          9114 => x"34",
          9115 => x"74",
          9116 => x"80",
          9117 => x"70",
          9118 => x"56",
          9119 => x"82",
          9120 => x"c0",
          9121 => x"34",
          9122 => x"3d",
          9123 => x"1c",
          9124 => x"59",
          9125 => x"5a",
          9126 => x"70",
          9127 => x"33",
          9128 => x"05",
          9129 => x"15",
          9130 => x"38",
          9131 => x"80",
          9132 => x"79",
          9133 => x"74",
          9134 => x"38",
          9135 => x"5a",
          9136 => x"75",
          9137 => x"10",
          9138 => x"2a",
          9139 => x"ff",
          9140 => x"2a",
          9141 => x"58",
          9142 => x"80",
          9143 => x"76",
          9144 => x"32",
          9145 => x"58",
          9146 => x"d7",
          9147 => x"55",
          9148 => x"87",
          9149 => x"80",
          9150 => x"58",
          9151 => x"bf",
          9152 => x"75",
          9153 => x"87",
          9154 => x"76",
          9155 => x"ff",
          9156 => x"2a",
          9157 => x"76",
          9158 => x"1f",
          9159 => x"79",
          9160 => x"58",
          9161 => x"27",
          9162 => x"33",
          9163 => x"2e",
          9164 => x"16",
          9165 => x"27",
          9166 => x"75",
          9167 => x"56",
          9168 => x"2e",
          9169 => x"ea",
          9170 => x"56",
          9171 => x"87",
          9172 => x"98",
          9173 => x"ec",
          9174 => x"71",
          9175 => x"41",
          9176 => x"87",
          9177 => x"f4",
          9178 => x"f8",
          9179 => x"ba",
          9180 => x"38",
          9181 => x"80",
          9182 => x"fe",
          9183 => x"56",
          9184 => x"2e",
          9185 => x"84",
          9186 => x"56",
          9187 => x"08",
          9188 => x"81",
          9189 => x"38",
          9190 => x"05",
          9191 => x"34",
          9192 => x"84",
          9193 => x"05",
          9194 => x"75",
          9195 => x"06",
          9196 => x"7e",
          9197 => x"38",
          9198 => x"1d",
          9199 => x"e7",
          9200 => x"8c",
          9201 => x"80",
          9202 => x"ed",
          9203 => x"ba",
          9204 => x"84",
          9205 => x"81",
          9206 => x"ba",
          9207 => x"19",
          9208 => x"1e",
          9209 => x"57",
          9210 => x"76",
          9211 => x"38",
          9212 => x"40",
          9213 => x"09",
          9214 => x"a3",
          9215 => x"75",
          9216 => x"52",
          9217 => x"51",
          9218 => x"84",
          9219 => x"80",
          9220 => x"ff",
          9221 => x"75",
          9222 => x"76",
          9223 => x"38",
          9224 => x"70",
          9225 => x"74",
          9226 => x"81",
          9227 => x"30",
          9228 => x"78",
          9229 => x"74",
          9230 => x"c9",
          9231 => x"59",
          9232 => x"86",
          9233 => x"52",
          9234 => x"83",
          9235 => x"8c",
          9236 => x"ba",
          9237 => x"2e",
          9238 => x"87",
          9239 => x"2e",
          9240 => x"75",
          9241 => x"83",
          9242 => x"40",
          9243 => x"38",
          9244 => x"57",
          9245 => x"77",
          9246 => x"83",
          9247 => x"57",
          9248 => x"82",
          9249 => x"76",
          9250 => x"52",
          9251 => x"51",
          9252 => x"84",
          9253 => x"80",
          9254 => x"ff",
          9255 => x"76",
          9256 => x"75",
          9257 => x"c3",
          9258 => x"9c",
          9259 => x"55",
          9260 => x"81",
          9261 => x"ff",
          9262 => x"f4",
          9263 => x"9c",
          9264 => x"58",
          9265 => x"70",
          9266 => x"33",
          9267 => x"05",
          9268 => x"15",
          9269 => x"38",
          9270 => x"ab",
          9271 => x"06",
          9272 => x"8c",
          9273 => x"0b",
          9274 => x"77",
          9275 => x"ba",
          9276 => x"3d",
          9277 => x"75",
          9278 => x"25",
          9279 => x"40",
          9280 => x"b9",
          9281 => x"81",
          9282 => x"ec",
          9283 => x"ba",
          9284 => x"84",
          9285 => x"80",
          9286 => x"38",
          9287 => x"81",
          9288 => x"08",
          9289 => x"81",
          9290 => x"d3",
          9291 => x"ba",
          9292 => x"2e",
          9293 => x"83",
          9294 => x"ba",
          9295 => x"19",
          9296 => x"08",
          9297 => x"31",
          9298 => x"19",
          9299 => x"38",
          9300 => x"41",
          9301 => x"84",
          9302 => x"ba",
          9303 => x"fd",
          9304 => x"85",
          9305 => x"08",
          9306 => x"58",
          9307 => x"e9",
          9308 => x"8c",
          9309 => x"ba",
          9310 => x"ef",
          9311 => x"ba",
          9312 => x"58",
          9313 => x"81",
          9314 => x"80",
          9315 => x"70",
          9316 => x"33",
          9317 => x"70",
          9318 => x"ff",
          9319 => x"5d",
          9320 => x"74",
          9321 => x"b8",
          9322 => x"98",
          9323 => x"80",
          9324 => x"08",
          9325 => x"38",
          9326 => x"5b",
          9327 => x"09",
          9328 => x"c9",
          9329 => x"76",
          9330 => x"52",
          9331 => x"51",
          9332 => x"84",
          9333 => x"80",
          9334 => x"ff",
          9335 => x"76",
          9336 => x"75",
          9337 => x"83",
          9338 => x"08",
          9339 => x"61",
          9340 => x"5f",
          9341 => x"8d",
          9342 => x"0b",
          9343 => x"75",
          9344 => x"75",
          9345 => x"75",
          9346 => x"7c",
          9347 => x"05",
          9348 => x"58",
          9349 => x"ff",
          9350 => x"38",
          9351 => x"70",
          9352 => x"5b",
          9353 => x"e6",
          9354 => x"7b",
          9355 => x"75",
          9356 => x"57",
          9357 => x"2a",
          9358 => x"34",
          9359 => x"83",
          9360 => x"81",
          9361 => x"78",
          9362 => x"76",
          9363 => x"2e",
          9364 => x"78",
          9365 => x"22",
          9366 => x"80",
          9367 => x"38",
          9368 => x"81",
          9369 => x"34",
          9370 => x"51",
          9371 => x"84",
          9372 => x"58",
          9373 => x"08",
          9374 => x"7f",
          9375 => x"7f",
          9376 => x"fb",
          9377 => x"54",
          9378 => x"53",
          9379 => x"53",
          9380 => x"52",
          9381 => x"3f",
          9382 => x"ba",
          9383 => x"83",
          9384 => x"8c",
          9385 => x"34",
          9386 => x"a8",
          9387 => x"84",
          9388 => x"57",
          9389 => x"1d",
          9390 => x"c9",
          9391 => x"33",
          9392 => x"2e",
          9393 => x"fb",
          9394 => x"54",
          9395 => x"a0",
          9396 => x"53",
          9397 => x"1c",
          9398 => x"d1",
          9399 => x"fb",
          9400 => x"9c",
          9401 => x"33",
          9402 => x"74",
          9403 => x"09",
          9404 => x"ba",
          9405 => x"39",
          9406 => x"57",
          9407 => x"fa",
          9408 => x"d7",
          9409 => x"c0",
          9410 => x"d4",
          9411 => x"b4",
          9412 => x"61",
          9413 => x"33",
          9414 => x"3f",
          9415 => x"08",
          9416 => x"81",
          9417 => x"84",
          9418 => x"83",
          9419 => x"1c",
          9420 => x"08",
          9421 => x"a0",
          9422 => x"8a",
          9423 => x"33",
          9424 => x"2e",
          9425 => x"ba",
          9426 => x"fc",
          9427 => x"ff",
          9428 => x"7f",
          9429 => x"98",
          9430 => x"39",
          9431 => x"f7",
          9432 => x"70",
          9433 => x"80",
          9434 => x"38",
          9435 => x"81",
          9436 => x"08",
          9437 => x"05",
          9438 => x"81",
          9439 => x"ce",
          9440 => x"c1",
          9441 => x"b4",
          9442 => x"19",
          9443 => x"7c",
          9444 => x"33",
          9445 => x"3f",
          9446 => x"f3",
          9447 => x"61",
          9448 => x"5e",
          9449 => x"96",
          9450 => x"1c",
          9451 => x"82",
          9452 => x"1c",
          9453 => x"80",
          9454 => x"70",
          9455 => x"05",
          9456 => x"57",
          9457 => x"58",
          9458 => x"bc",
          9459 => x"74",
          9460 => x"81",
          9461 => x"56",
          9462 => x"38",
          9463 => x"14",
          9464 => x"ff",
          9465 => x"76",
          9466 => x"82",
          9467 => x"79",
          9468 => x"70",
          9469 => x"55",
          9470 => x"38",
          9471 => x"80",
          9472 => x"7a",
          9473 => x"5e",
          9474 => x"05",
          9475 => x"82",
          9476 => x"70",
          9477 => x"57",
          9478 => x"08",
          9479 => x"81",
          9480 => x"53",
          9481 => x"b2",
          9482 => x"2e",
          9483 => x"75",
          9484 => x"30",
          9485 => x"80",
          9486 => x"54",
          9487 => x"90",
          9488 => x"2e",
          9489 => x"77",
          9490 => x"59",
          9491 => x"58",
          9492 => x"81",
          9493 => x"81",
          9494 => x"76",
          9495 => x"38",
          9496 => x"05",
          9497 => x"81",
          9498 => x"1d",
          9499 => x"a5",
          9500 => x"f3",
          9501 => x"96",
          9502 => x"57",
          9503 => x"05",
          9504 => x"82",
          9505 => x"1c",
          9506 => x"33",
          9507 => x"89",
          9508 => x"1e",
          9509 => x"08",
          9510 => x"33",
          9511 => x"9c",
          9512 => x"11",
          9513 => x"82",
          9514 => x"90",
          9515 => x"2b",
          9516 => x"33",
          9517 => x"88",
          9518 => x"71",
          9519 => x"59",
          9520 => x"96",
          9521 => x"88",
          9522 => x"41",
          9523 => x"56",
          9524 => x"86",
          9525 => x"15",
          9526 => x"33",
          9527 => x"07",
          9528 => x"84",
          9529 => x"3d",
          9530 => x"e5",
          9531 => x"39",
          9532 => x"11",
          9533 => x"31",
          9534 => x"83",
          9535 => x"90",
          9536 => x"51",
          9537 => x"3f",
          9538 => x"08",
          9539 => x"06",
          9540 => x"75",
          9541 => x"81",
          9542 => x"b3",
          9543 => x"2a",
          9544 => x"34",
          9545 => x"34",
          9546 => x"58",
          9547 => x"1f",
          9548 => x"78",
          9549 => x"70",
          9550 => x"54",
          9551 => x"38",
          9552 => x"74",
          9553 => x"70",
          9554 => x"25",
          9555 => x"07",
          9556 => x"75",
          9557 => x"74",
          9558 => x"78",
          9559 => x"0b",
          9560 => x"56",
          9561 => x"72",
          9562 => x"33",
          9563 => x"77",
          9564 => x"88",
          9565 => x"1e",
          9566 => x"54",
          9567 => x"ff",
          9568 => x"54",
          9569 => x"a4",
          9570 => x"08",
          9571 => x"54",
          9572 => x"27",
          9573 => x"84",
          9574 => x"81",
          9575 => x"80",
          9576 => x"a0",
          9577 => x"ff",
          9578 => x"53",
          9579 => x"81",
          9580 => x"81",
          9581 => x"81",
          9582 => x"13",
          9583 => x"59",
          9584 => x"ff",
          9585 => x"b4",
          9586 => x"2a",
          9587 => x"80",
          9588 => x"80",
          9589 => x"73",
          9590 => x"5f",
          9591 => x"39",
          9592 => x"63",
          9593 => x"42",
          9594 => x"65",
          9595 => x"55",
          9596 => x"2e",
          9597 => x"53",
          9598 => x"2e",
          9599 => x"72",
          9600 => x"d9",
          9601 => x"08",
          9602 => x"73",
          9603 => x"94",
          9604 => x"55",
          9605 => x"82",
          9606 => x"42",
          9607 => x"58",
          9608 => x"70",
          9609 => x"52",
          9610 => x"73",
          9611 => x"72",
          9612 => x"ff",
          9613 => x"38",
          9614 => x"74",
          9615 => x"76",
          9616 => x"80",
          9617 => x"17",
          9618 => x"ff",
          9619 => x"af",
          9620 => x"9f",
          9621 => x"80",
          9622 => x"5b",
          9623 => x"82",
          9624 => x"80",
          9625 => x"89",
          9626 => x"ff",
          9627 => x"83",
          9628 => x"83",
          9629 => x"70",
          9630 => x"56",
          9631 => x"80",
          9632 => x"38",
          9633 => x"8f",
          9634 => x"70",
          9635 => x"ff",
          9636 => x"56",
          9637 => x"72",
          9638 => x"5b",
          9639 => x"38",
          9640 => x"26",
          9641 => x"76",
          9642 => x"74",
          9643 => x"17",
          9644 => x"81",
          9645 => x"56",
          9646 => x"80",
          9647 => x"38",
          9648 => x"81",
          9649 => x"32",
          9650 => x"80",
          9651 => x"51",
          9652 => x"72",
          9653 => x"38",
          9654 => x"46",
          9655 => x"33",
          9656 => x"af",
          9657 => x"72",
          9658 => x"70",
          9659 => x"25",
          9660 => x"54",
          9661 => x"38",
          9662 => x"0c",
          9663 => x"3d",
          9664 => x"42",
          9665 => x"26",
          9666 => x"b4",
          9667 => x"52",
          9668 => x"8d",
          9669 => x"ba",
          9670 => x"ff",
          9671 => x"73",
          9672 => x"86",
          9673 => x"ba",
          9674 => x"3d",
          9675 => x"e5",
          9676 => x"81",
          9677 => x"53",
          9678 => x"fe",
          9679 => x"39",
          9680 => x"ab",
          9681 => x"52",
          9682 => x"8d",
          9683 => x"8c",
          9684 => x"8c",
          9685 => x"0d",
          9686 => x"80",
          9687 => x"30",
          9688 => x"73",
          9689 => x"5a",
          9690 => x"2e",
          9691 => x"14",
          9692 => x"70",
          9693 => x"56",
          9694 => x"dd",
          9695 => x"dc",
          9696 => x"70",
          9697 => x"07",
          9698 => x"7d",
          9699 => x"61",
          9700 => x"27",
          9701 => x"76",
          9702 => x"f8",
          9703 => x"2e",
          9704 => x"76",
          9705 => x"80",
          9706 => x"76",
          9707 => x"fe",
          9708 => x"70",
          9709 => x"30",
          9710 => x"52",
          9711 => x"56",
          9712 => x"2e",
          9713 => x"89",
          9714 => x"57",
          9715 => x"76",
          9716 => x"56",
          9717 => x"76",
          9718 => x"c7",
          9719 => x"22",
          9720 => x"ff",
          9721 => x"5d",
          9722 => x"a0",
          9723 => x"38",
          9724 => x"ff",
          9725 => x"ae",
          9726 => x"38",
          9727 => x"aa",
          9728 => x"fe",
          9729 => x"5a",
          9730 => x"2e",
          9731 => x"10",
          9732 => x"54",
          9733 => x"76",
          9734 => x"38",
          9735 => x"22",
          9736 => x"ae",
          9737 => x"06",
          9738 => x"0b",
          9739 => x"53",
          9740 => x"81",
          9741 => x"ff",
          9742 => x"f4",
          9743 => x"5c",
          9744 => x"16",
          9745 => x"19",
          9746 => x"5d",
          9747 => x"80",
          9748 => x"a0",
          9749 => x"38",
          9750 => x"70",
          9751 => x"25",
          9752 => x"75",
          9753 => x"ce",
          9754 => x"bb",
          9755 => x"7c",
          9756 => x"38",
          9757 => x"77",
          9758 => x"70",
          9759 => x"25",
          9760 => x"51",
          9761 => x"72",
          9762 => x"e0",
          9763 => x"2e",
          9764 => x"75",
          9765 => x"38",
          9766 => x"5a",
          9767 => x"9e",
          9768 => x"88",
          9769 => x"82",
          9770 => x"06",
          9771 => x"5f",
          9772 => x"70",
          9773 => x"58",
          9774 => x"ff",
          9775 => x"1c",
          9776 => x"81",
          9777 => x"84",
          9778 => x"2e",
          9779 => x"7d",
          9780 => x"77",
          9781 => x"ed",
          9782 => x"06",
          9783 => x"2e",
          9784 => x"79",
          9785 => x"06",
          9786 => x"38",
          9787 => x"5d",
          9788 => x"85",
          9789 => x"07",
          9790 => x"2a",
          9791 => x"7d",
          9792 => x"38",
          9793 => x"5a",
          9794 => x"34",
          9795 => x"ec",
          9796 => x"8c",
          9797 => x"33",
          9798 => x"ba",
          9799 => x"2e",
          9800 => x"84",
          9801 => x"84",
          9802 => x"06",
          9803 => x"74",
          9804 => x"06",
          9805 => x"2e",
          9806 => x"74",
          9807 => x"06",
          9808 => x"98",
          9809 => x"65",
          9810 => x"42",
          9811 => x"58",
          9812 => x"ce",
          9813 => x"70",
          9814 => x"70",
          9815 => x"56",
          9816 => x"2e",
          9817 => x"80",
          9818 => x"38",
          9819 => x"5a",
          9820 => x"82",
          9821 => x"75",
          9822 => x"81",
          9823 => x"38",
          9824 => x"73",
          9825 => x"81",
          9826 => x"38",
          9827 => x"5b",
          9828 => x"80",
          9829 => x"56",
          9830 => x"76",
          9831 => x"38",
          9832 => x"75",
          9833 => x"57",
          9834 => x"53",
          9835 => x"e9",
          9836 => x"07",
          9837 => x"1d",
          9838 => x"e3",
          9839 => x"ba",
          9840 => x"1d",
          9841 => x"84",
          9842 => x"fe",
          9843 => x"82",
          9844 => x"58",
          9845 => x"38",
          9846 => x"70",
          9847 => x"06",
          9848 => x"80",
          9849 => x"38",
          9850 => x"83",
          9851 => x"05",
          9852 => x"33",
          9853 => x"33",
          9854 => x"07",
          9855 => x"57",
          9856 => x"83",
          9857 => x"38",
          9858 => x"0c",
          9859 => x"55",
          9860 => x"39",
          9861 => x"74",
          9862 => x"f0",
          9863 => x"59",
          9864 => x"38",
          9865 => x"79",
          9866 => x"17",
          9867 => x"81",
          9868 => x"2b",
          9869 => x"70",
          9870 => x"5e",
          9871 => x"09",
          9872 => x"95",
          9873 => x"07",
          9874 => x"39",
          9875 => x"1d",
          9876 => x"2e",
          9877 => x"fc",
          9878 => x"39",
          9879 => x"ab",
          9880 => x"0b",
          9881 => x"0c",
          9882 => x"04",
          9883 => x"26",
          9884 => x"ff",
          9885 => x"c9",
          9886 => x"59",
          9887 => x"81",
          9888 => x"83",
          9889 => x"18",
          9890 => x"fc",
          9891 => x"82",
          9892 => x"b5",
          9893 => x"81",
          9894 => x"84",
          9895 => x"83",
          9896 => x"70",
          9897 => x"06",
          9898 => x"80",
          9899 => x"74",
          9900 => x"83",
          9901 => x"33",
          9902 => x"81",
          9903 => x"b9",
          9904 => x"2e",
          9905 => x"83",
          9906 => x"83",
          9907 => x"70",
          9908 => x"56",
          9909 => x"80",
          9910 => x"38",
          9911 => x"8f",
          9912 => x"70",
          9913 => x"ff",
          9914 => x"59",
          9915 => x"72",
          9916 => x"59",
          9917 => x"38",
          9918 => x"54",
          9919 => x"8a",
          9920 => x"07",
          9921 => x"06",
          9922 => x"9f",
          9923 => x"99",
          9924 => x"7d",
          9925 => x"81",
          9926 => x"17",
          9927 => x"ff",
          9928 => x"5f",
          9929 => x"a0",
          9930 => x"79",
          9931 => x"5b",
          9932 => x"fa",
          9933 => x"53",
          9934 => x"83",
          9935 => x"70",
          9936 => x"5a",
          9937 => x"2e",
          9938 => x"80",
          9939 => x"07",
          9940 => x"05",
          9941 => x"74",
          9942 => x"1b",
          9943 => x"80",
          9944 => x"80",
          9945 => x"71",
          9946 => x"90",
          9947 => x"07",
          9948 => x"5a",
          9949 => x"39",
          9950 => x"05",
          9951 => x"54",
          9952 => x"34",
          9953 => x"11",
          9954 => x"5b",
          9955 => x"81",
          9956 => x"9c",
          9957 => x"07",
          9958 => x"58",
          9959 => x"e5",
          9960 => x"06",
          9961 => x"fd",
          9962 => x"82",
          9963 => x"5c",
          9964 => x"38",
          9965 => x"ba",
          9966 => x"3d",
          9967 => x"3d",
          9968 => x"02",
          9969 => x"e7",
          9970 => x"42",
          9971 => x"0c",
          9972 => x"70",
          9973 => x"79",
          9974 => x"d7",
          9975 => x"81",
          9976 => x"70",
          9977 => x"56",
          9978 => x"85",
          9979 => x"ed",
          9980 => x"2e",
          9981 => x"84",
          9982 => x"56",
          9983 => x"85",
          9984 => x"10",
          9985 => x"d4",
          9986 => x"58",
          9987 => x"76",
          9988 => x"96",
          9989 => x"0c",
          9990 => x"06",
          9991 => x"59",
          9992 => x"9b",
          9993 => x"33",
          9994 => x"b0",
          9995 => x"8c",
          9996 => x"06",
          9997 => x"5e",
          9998 => x"2e",
          9999 => x"80",
         10000 => x"16",
         10001 => x"80",
         10002 => x"18",
         10003 => x"81",
         10004 => x"ff",
         10005 => x"84",
         10006 => x"81",
         10007 => x"81",
         10008 => x"83",
         10009 => x"c2",
         10010 => x"2e",
         10011 => x"82",
         10012 => x"41",
         10013 => x"84",
         10014 => x"5b",
         10015 => x"34",
         10016 => x"18",
         10017 => x"5a",
         10018 => x"7a",
         10019 => x"70",
         10020 => x"33",
         10021 => x"bb",
         10022 => x"ba",
         10023 => x"2e",
         10024 => x"55",
         10025 => x"b4",
         10026 => x"56",
         10027 => x"84",
         10028 => x"84",
         10029 => x"71",
         10030 => x"56",
         10031 => x"74",
         10032 => x"2e",
         10033 => x"75",
         10034 => x"38",
         10035 => x"1d",
         10036 => x"85",
         10037 => x"58",
         10038 => x"83",
         10039 => x"58",
         10040 => x"83",
         10041 => x"c4",
         10042 => x"c3",
         10043 => x"88",
         10044 => x"59",
         10045 => x"2e",
         10046 => x"83",
         10047 => x"cf",
         10048 => x"ce",
         10049 => x"88",
         10050 => x"5a",
         10051 => x"80",
         10052 => x"11",
         10053 => x"33",
         10054 => x"71",
         10055 => x"81",
         10056 => x"72",
         10057 => x"75",
         10058 => x"56",
         10059 => x"5e",
         10060 => x"a0",
         10061 => x"c8",
         10062 => x"18",
         10063 => x"17",
         10064 => x"70",
         10065 => x"5f",
         10066 => x"58",
         10067 => x"82",
         10068 => x"81",
         10069 => x"71",
         10070 => x"19",
         10071 => x"5a",
         10072 => x"23",
         10073 => x"80",
         10074 => x"38",
         10075 => x"06",
         10076 => x"bb",
         10077 => x"17",
         10078 => x"18",
         10079 => x"2b",
         10080 => x"74",
         10081 => x"74",
         10082 => x"5e",
         10083 => x"7c",
         10084 => x"80",
         10085 => x"80",
         10086 => x"71",
         10087 => x"56",
         10088 => x"38",
         10089 => x"83",
         10090 => x"12",
         10091 => x"2b",
         10092 => x"07",
         10093 => x"70",
         10094 => x"2b",
         10095 => x"07",
         10096 => x"58",
         10097 => x"80",
         10098 => x"80",
         10099 => x"71",
         10100 => x"5d",
         10101 => x"7b",
         10102 => x"ce",
         10103 => x"7a",
         10104 => x"5a",
         10105 => x"81",
         10106 => x"52",
         10107 => x"51",
         10108 => x"3f",
         10109 => x"08",
         10110 => x"8c",
         10111 => x"81",
         10112 => x"ba",
         10113 => x"ff",
         10114 => x"26",
         10115 => x"5d",
         10116 => x"f5",
         10117 => x"82",
         10118 => x"f5",
         10119 => x"38",
         10120 => x"16",
         10121 => x"0c",
         10122 => x"0c",
         10123 => x"a8",
         10124 => x"1d",
         10125 => x"57",
         10126 => x"2e",
         10127 => x"88",
         10128 => x"8d",
         10129 => x"2e",
         10130 => x"7d",
         10131 => x"0c",
         10132 => x"7c",
         10133 => x"38",
         10134 => x"70",
         10135 => x"81",
         10136 => x"5a",
         10137 => x"89",
         10138 => x"58",
         10139 => x"08",
         10140 => x"ff",
         10141 => x"0c",
         10142 => x"18",
         10143 => x"0b",
         10144 => x"7c",
         10145 => x"96",
         10146 => x"34",
         10147 => x"22",
         10148 => x"7c",
         10149 => x"23",
         10150 => x"23",
         10151 => x"0b",
         10152 => x"80",
         10153 => x"0c",
         10154 => x"84",
         10155 => x"97",
         10156 => x"8b",
         10157 => x"8c",
         10158 => x"0d",
         10159 => x"d0",
         10160 => x"ff",
         10161 => x"58",
         10162 => x"91",
         10163 => x"78",
         10164 => x"d0",
         10165 => x"78",
         10166 => x"fe",
         10167 => x"08",
         10168 => x"5f",
         10169 => x"08",
         10170 => x"7a",
         10171 => x"5c",
         10172 => x"81",
         10173 => x"ff",
         10174 => x"58",
         10175 => x"26",
         10176 => x"16",
         10177 => x"06",
         10178 => x"9f",
         10179 => x"99",
         10180 => x"e0",
         10181 => x"ff",
         10182 => x"75",
         10183 => x"2a",
         10184 => x"77",
         10185 => x"06",
         10186 => x"ff",
         10187 => x"7a",
         10188 => x"70",
         10189 => x"2a",
         10190 => x"58",
         10191 => x"2e",
         10192 => x"81",
         10193 => x"5e",
         10194 => x"25",
         10195 => x"61",
         10196 => x"39",
         10197 => x"fe",
         10198 => x"82",
         10199 => x"5e",
         10200 => x"fe",
         10201 => x"58",
         10202 => x"7a",
         10203 => x"59",
         10204 => x"2e",
         10205 => x"83",
         10206 => x"75",
         10207 => x"70",
         10208 => x"25",
         10209 => x"5b",
         10210 => x"ad",
         10211 => x"e8",
         10212 => x"38",
         10213 => x"57",
         10214 => x"83",
         10215 => x"70",
         10216 => x"80",
         10217 => x"84",
         10218 => x"84",
         10219 => x"71",
         10220 => x"88",
         10221 => x"ff",
         10222 => x"72",
         10223 => x"83",
         10224 => x"71",
         10225 => x"5b",
         10226 => x"77",
         10227 => x"05",
         10228 => x"19",
         10229 => x"59",
         10230 => x"ff",
         10231 => x"ba",
         10232 => x"70",
         10233 => x"2a",
         10234 => x"9b",
         10235 => x"10",
         10236 => x"84",
         10237 => x"5d",
         10238 => x"42",
         10239 => x"83",
         10240 => x"2e",
         10241 => x"80",
         10242 => x"34",
         10243 => x"18",
         10244 => x"80",
         10245 => x"2e",
         10246 => x"54",
         10247 => x"17",
         10248 => x"33",
         10249 => x"86",
         10250 => x"8c",
         10251 => x"85",
         10252 => x"81",
         10253 => x"18",
         10254 => x"75",
         10255 => x"1f",
         10256 => x"71",
         10257 => x"5d",
         10258 => x"7b",
         10259 => x"2e",
         10260 => x"a8",
         10261 => x"b8",
         10262 => x"58",
         10263 => x"2e",
         10264 => x"75",
         10265 => x"70",
         10266 => x"25",
         10267 => x"42",
         10268 => x"38",
         10269 => x"2e",
         10270 => x"58",
         10271 => x"06",
         10272 => x"84",
         10273 => x"33",
         10274 => x"78",
         10275 => x"06",
         10276 => x"58",
         10277 => x"f8",
         10278 => x"80",
         10279 => x"38",
         10280 => x"1a",
         10281 => x"7a",
         10282 => x"38",
         10283 => x"83",
         10284 => x"18",
         10285 => x"40",
         10286 => x"70",
         10287 => x"33",
         10288 => x"05",
         10289 => x"71",
         10290 => x"5b",
         10291 => x"77",
         10292 => x"c5",
         10293 => x"2e",
         10294 => x"0b",
         10295 => x"83",
         10296 => x"5d",
         10297 => x"81",
         10298 => x"7e",
         10299 => x"40",
         10300 => x"31",
         10301 => x"58",
         10302 => x"80",
         10303 => x"38",
         10304 => x"e1",
         10305 => x"fe",
         10306 => x"58",
         10307 => x"38",
         10308 => x"8c",
         10309 => x"0d",
         10310 => x"75",
         10311 => x"dc",
         10312 => x"81",
         10313 => x"e5",
         10314 => x"58",
         10315 => x"8d",
         10316 => x"8c",
         10317 => x"0d",
         10318 => x"80",
         10319 => x"e5",
         10320 => x"58",
         10321 => x"05",
         10322 => x"70",
         10323 => x"33",
         10324 => x"ff",
         10325 => x"5f",
         10326 => x"2e",
         10327 => x"74",
         10328 => x"38",
         10329 => x"8a",
         10330 => x"c0",
         10331 => x"78",
         10332 => x"5a",
         10333 => x"81",
         10334 => x"71",
         10335 => x"1b",
         10336 => x"40",
         10337 => x"84",
         10338 => x"80",
         10339 => x"93",
         10340 => x"5a",
         10341 => x"83",
         10342 => x"fd",
         10343 => x"e9",
         10344 => x"e8",
         10345 => x"88",
         10346 => x"55",
         10347 => x"09",
         10348 => x"d5",
         10349 => x"58",
         10350 => x"17",
         10351 => x"b1",
         10352 => x"33",
         10353 => x"2e",
         10354 => x"82",
         10355 => x"54",
         10356 => x"17",
         10357 => x"33",
         10358 => x"d2",
         10359 => x"8c",
         10360 => x"85",
         10361 => x"81",
         10362 => x"18",
         10363 => x"99",
         10364 => x"18",
         10365 => x"17",
         10366 => x"18",
         10367 => x"2b",
         10368 => x"75",
         10369 => x"2e",
         10370 => x"f8",
         10371 => x"17",
         10372 => x"82",
         10373 => x"90",
         10374 => x"2b",
         10375 => x"33",
         10376 => x"88",
         10377 => x"71",
         10378 => x"59",
         10379 => x"59",
         10380 => x"85",
         10381 => x"09",
         10382 => x"cd",
         10383 => x"17",
         10384 => x"82",
         10385 => x"90",
         10386 => x"2b",
         10387 => x"33",
         10388 => x"88",
         10389 => x"71",
         10390 => x"40",
         10391 => x"5e",
         10392 => x"85",
         10393 => x"09",
         10394 => x"9d",
         10395 => x"17",
         10396 => x"82",
         10397 => x"90",
         10398 => x"2b",
         10399 => x"33",
         10400 => x"88",
         10401 => x"71",
         10402 => x"0c",
         10403 => x"1c",
         10404 => x"82",
         10405 => x"90",
         10406 => x"2b",
         10407 => x"33",
         10408 => x"88",
         10409 => x"71",
         10410 => x"05",
         10411 => x"49",
         10412 => x"40",
         10413 => x"5a",
         10414 => x"84",
         10415 => x"81",
         10416 => x"84",
         10417 => x"7c",
         10418 => x"84",
         10419 => x"8c",
         10420 => x"0b",
         10421 => x"f7",
         10422 => x"83",
         10423 => x"38",
         10424 => x"0c",
         10425 => x"39",
         10426 => x"17",
         10427 => x"17",
         10428 => x"18",
         10429 => x"ff",
         10430 => x"84",
         10431 => x"7a",
         10432 => x"06",
         10433 => x"84",
         10434 => x"83",
         10435 => x"17",
         10436 => x"08",
         10437 => x"a0",
         10438 => x"8b",
         10439 => x"33",
         10440 => x"2e",
         10441 => x"84",
         10442 => x"5a",
         10443 => x"74",
         10444 => x"2e",
         10445 => x"85",
         10446 => x"18",
         10447 => x"5c",
         10448 => x"ab",
         10449 => x"17",
         10450 => x"18",
         10451 => x"2b",
         10452 => x"8d",
         10453 => x"d2",
         10454 => x"22",
         10455 => x"ca",
         10456 => x"17",
         10457 => x"82",
         10458 => x"90",
         10459 => x"2b",
         10460 => x"33",
         10461 => x"88",
         10462 => x"71",
         10463 => x"0c",
         10464 => x"2b",
         10465 => x"40",
         10466 => x"d8",
         10467 => x"75",
         10468 => x"e8",
         10469 => x"f9",
         10470 => x"80",
         10471 => x"38",
         10472 => x"57",
         10473 => x"f7",
         10474 => x"5a",
         10475 => x"38",
         10476 => x"75",
         10477 => x"08",
         10478 => x"05",
         10479 => x"81",
         10480 => x"ff",
         10481 => x"fc",
         10482 => x"3d",
         10483 => x"d3",
         10484 => x"70",
         10485 => x"41",
         10486 => x"76",
         10487 => x"80",
         10488 => x"38",
         10489 => x"05",
         10490 => x"9f",
         10491 => x"74",
         10492 => x"e2",
         10493 => x"38",
         10494 => x"80",
         10495 => x"d1",
         10496 => x"80",
         10497 => x"c4",
         10498 => x"10",
         10499 => x"05",
         10500 => x"55",
         10501 => x"84",
         10502 => x"34",
         10503 => x"80",
         10504 => x"80",
         10505 => x"54",
         10506 => x"7c",
         10507 => x"2e",
         10508 => x"53",
         10509 => x"53",
         10510 => x"ef",
         10511 => x"ba",
         10512 => x"73",
         10513 => x"0c",
         10514 => x"04",
         10515 => x"ba",
         10516 => x"3d",
         10517 => x"33",
         10518 => x"81",
         10519 => x"56",
         10520 => x"26",
         10521 => x"16",
         10522 => x"06",
         10523 => x"58",
         10524 => x"80",
         10525 => x"7f",
         10526 => x"fc",
         10527 => x"7b",
         10528 => x"5a",
         10529 => x"05",
         10530 => x"70",
         10531 => x"33",
         10532 => x"59",
         10533 => x"99",
         10534 => x"e0",
         10535 => x"ff",
         10536 => x"ff",
         10537 => x"76",
         10538 => x"38",
         10539 => x"81",
         10540 => x"54",
         10541 => x"9f",
         10542 => x"74",
         10543 => x"81",
         10544 => x"76",
         10545 => x"77",
         10546 => x"30",
         10547 => x"9f",
         10548 => x"5c",
         10549 => x"80",
         10550 => x"81",
         10551 => x"5d",
         10552 => x"25",
         10553 => x"7f",
         10554 => x"39",
         10555 => x"f7",
         10556 => x"60",
         10557 => x"8b",
         10558 => x"0d",
         10559 => x"05",
         10560 => x"33",
         10561 => x"56",
         10562 => x"a6",
         10563 => x"06",
         10564 => x"3d",
         10565 => x"9e",
         10566 => x"52",
         10567 => x"3f",
         10568 => x"08",
         10569 => x"8c",
         10570 => x"8f",
         10571 => x"0c",
         10572 => x"84",
         10573 => x"9c",
         10574 => x"7e",
         10575 => x"90",
         10576 => x"5a",
         10577 => x"84",
         10578 => x"57",
         10579 => x"08",
         10580 => x"ba",
         10581 => x"06",
         10582 => x"2e",
         10583 => x"76",
         10584 => x"c1",
         10585 => x"2e",
         10586 => x"77",
         10587 => x"76",
         10588 => x"77",
         10589 => x"06",
         10590 => x"2e",
         10591 => x"66",
         10592 => x"9a",
         10593 => x"88",
         10594 => x"70",
         10595 => x"5e",
         10596 => x"83",
         10597 => x"38",
         10598 => x"17",
         10599 => x"8f",
         10600 => x"0b",
         10601 => x"80",
         10602 => x"17",
         10603 => x"a0",
         10604 => x"34",
         10605 => x"5e",
         10606 => x"17",
         10607 => x"9b",
         10608 => x"33",
         10609 => x"2e",
         10610 => x"66",
         10611 => x"9c",
         10612 => x"0b",
         10613 => x"80",
         10614 => x"34",
         10615 => x"1c",
         10616 => x"81",
         10617 => x"34",
         10618 => x"80",
         10619 => x"b4",
         10620 => x"7c",
         10621 => x"5f",
         10622 => x"27",
         10623 => x"17",
         10624 => x"83",
         10625 => x"57",
         10626 => x"fe",
         10627 => x"80",
         10628 => x"70",
         10629 => x"5b",
         10630 => x"fe",
         10631 => x"78",
         10632 => x"57",
         10633 => x"38",
         10634 => x"38",
         10635 => x"05",
         10636 => x"2a",
         10637 => x"56",
         10638 => x"38",
         10639 => x"81",
         10640 => x"80",
         10641 => x"75",
         10642 => x"79",
         10643 => x"77",
         10644 => x"06",
         10645 => x"2e",
         10646 => x"80",
         10647 => x"7e",
         10648 => x"a0",
         10649 => x"a4",
         10650 => x"9b",
         10651 => x"12",
         10652 => x"2b",
         10653 => x"40",
         10654 => x"5a",
         10655 => x"81",
         10656 => x"88",
         10657 => x"16",
         10658 => x"82",
         10659 => x"90",
         10660 => x"2b",
         10661 => x"33",
         10662 => x"88",
         10663 => x"71",
         10664 => x"8c",
         10665 => x"60",
         10666 => x"41",
         10667 => x"5e",
         10668 => x"84",
         10669 => x"90",
         10670 => x"0b",
         10671 => x"80",
         10672 => x"0c",
         10673 => x"81",
         10674 => x"80",
         10675 => x"38",
         10676 => x"84",
         10677 => x"94",
         10678 => x"1a",
         10679 => x"2b",
         10680 => x"58",
         10681 => x"78",
         10682 => x"56",
         10683 => x"27",
         10684 => x"81",
         10685 => x"5f",
         10686 => x"2e",
         10687 => x"77",
         10688 => x"ff",
         10689 => x"84",
         10690 => x"58",
         10691 => x"08",
         10692 => x"38",
         10693 => x"ba",
         10694 => x"2e",
         10695 => x"75",
         10696 => x"c0",
         10697 => x"c2",
         10698 => x"06",
         10699 => x"38",
         10700 => x"81",
         10701 => x"80",
         10702 => x"38",
         10703 => x"79",
         10704 => x"39",
         10705 => x"79",
         10706 => x"39",
         10707 => x"79",
         10708 => x"39",
         10709 => x"ca",
         10710 => x"8c",
         10711 => x"07",
         10712 => x"fb",
         10713 => x"8b",
         10714 => x"7b",
         10715 => x"fe",
         10716 => x"16",
         10717 => x"33",
         10718 => x"71",
         10719 => x"7d",
         10720 => x"5c",
         10721 => x"7c",
         10722 => x"27",
         10723 => x"74",
         10724 => x"ff",
         10725 => x"84",
         10726 => x"5d",
         10727 => x"08",
         10728 => x"a7",
         10729 => x"8c",
         10730 => x"fc",
         10731 => x"ba",
         10732 => x"2e",
         10733 => x"80",
         10734 => x"76",
         10735 => x"82",
         10736 => x"8c",
         10737 => x"38",
         10738 => x"fe",
         10739 => x"08",
         10740 => x"75",
         10741 => x"af",
         10742 => x"94",
         10743 => x"17",
         10744 => x"55",
         10745 => x"34",
         10746 => x"7d",
         10747 => x"38",
         10748 => x"80",
         10749 => x"34",
         10750 => x"17",
         10751 => x"39",
         10752 => x"94",
         10753 => x"98",
         10754 => x"2b",
         10755 => x"5e",
         10756 => x"0b",
         10757 => x"80",
         10758 => x"34",
         10759 => x"17",
         10760 => x"0b",
         10761 => x"66",
         10762 => x"8b",
         10763 => x"67",
         10764 => x"0b",
         10765 => x"80",
         10766 => x"34",
         10767 => x"7c",
         10768 => x"81",
         10769 => x"38",
         10770 => x"80",
         10771 => x"5e",
         10772 => x"b4",
         10773 => x"2e",
         10774 => x"16",
         10775 => x"7d",
         10776 => x"06",
         10777 => x"54",
         10778 => x"16",
         10779 => x"33",
         10780 => x"ba",
         10781 => x"8c",
         10782 => x"85",
         10783 => x"81",
         10784 => x"17",
         10785 => x"7a",
         10786 => x"18",
         10787 => x"80",
         10788 => x"38",
         10789 => x"f9",
         10790 => x"54",
         10791 => x"53",
         10792 => x"53",
         10793 => x"52",
         10794 => x"81",
         10795 => x"8c",
         10796 => x"09",
         10797 => x"aa",
         10798 => x"8c",
         10799 => x"34",
         10800 => x"a8",
         10801 => x"84",
         10802 => x"5c",
         10803 => x"17",
         10804 => x"92",
         10805 => x"33",
         10806 => x"2e",
         10807 => x"ff",
         10808 => x"54",
         10809 => x"a0",
         10810 => x"53",
         10811 => x"16",
         10812 => x"a3",
         10813 => x"5b",
         10814 => x"74",
         10815 => x"76",
         10816 => x"39",
         10817 => x"0c",
         10818 => x"38",
         10819 => x"06",
         10820 => x"2e",
         10821 => x"7e",
         10822 => x"12",
         10823 => x"5f",
         10824 => x"7d",
         10825 => x"38",
         10826 => x"78",
         10827 => x"1c",
         10828 => x"5c",
         10829 => x"f9",
         10830 => x"89",
         10831 => x"1a",
         10832 => x"f7",
         10833 => x"94",
         10834 => x"56",
         10835 => x"81",
         10836 => x"0c",
         10837 => x"84",
         10838 => x"57",
         10839 => x"f7",
         10840 => x"7f",
         10841 => x"9f",
         10842 => x"0d",
         10843 => x"66",
         10844 => x"5a",
         10845 => x"89",
         10846 => x"2e",
         10847 => x"08",
         10848 => x"2e",
         10849 => x"33",
         10850 => x"2e",
         10851 => x"16",
         10852 => x"22",
         10853 => x"78",
         10854 => x"38",
         10855 => x"41",
         10856 => x"82",
         10857 => x"1a",
         10858 => x"82",
         10859 => x"1a",
         10860 => x"57",
         10861 => x"80",
         10862 => x"38",
         10863 => x"8c",
         10864 => x"31",
         10865 => x"75",
         10866 => x"38",
         10867 => x"81",
         10868 => x"59",
         10869 => x"06",
         10870 => x"e3",
         10871 => x"22",
         10872 => x"89",
         10873 => x"7a",
         10874 => x"83",
         10875 => x"1a",
         10876 => x"75",
         10877 => x"38",
         10878 => x"83",
         10879 => x"98",
         10880 => x"59",
         10881 => x"fe",
         10882 => x"08",
         10883 => x"57",
         10884 => x"83",
         10885 => x"19",
         10886 => x"29",
         10887 => x"05",
         10888 => x"80",
         10889 => x"38",
         10890 => x"89",
         10891 => x"77",
         10892 => x"81",
         10893 => x"55",
         10894 => x"85",
         10895 => x"31",
         10896 => x"76",
         10897 => x"81",
         10898 => x"ff",
         10899 => x"84",
         10900 => x"83",
         10901 => x"83",
         10902 => x"59",
         10903 => x"a9",
         10904 => x"08",
         10905 => x"75",
         10906 => x"38",
         10907 => x"71",
         10908 => x"1b",
         10909 => x"75",
         10910 => x"57",
         10911 => x"81",
         10912 => x"ff",
         10913 => x"ef",
         10914 => x"2b",
         10915 => x"31",
         10916 => x"7f",
         10917 => x"94",
         10918 => x"70",
         10919 => x"0c",
         10920 => x"fe",
         10921 => x"56",
         10922 => x"8c",
         10923 => x"0d",
         10924 => x"ba",
         10925 => x"3d",
         10926 => x"5c",
         10927 => x"9c",
         10928 => x"75",
         10929 => x"84",
         10930 => x"59",
         10931 => x"27",
         10932 => x"58",
         10933 => x"19",
         10934 => x"b6",
         10935 => x"83",
         10936 => x"5d",
         10937 => x"7f",
         10938 => x"06",
         10939 => x"81",
         10940 => x"b8",
         10941 => x"19",
         10942 => x"9e",
         10943 => x"ba",
         10944 => x"2e",
         10945 => x"56",
         10946 => x"b4",
         10947 => x"81",
         10948 => x"94",
         10949 => x"ff",
         10950 => x"7f",
         10951 => x"05",
         10952 => x"80",
         10953 => x"38",
         10954 => x"05",
         10955 => x"70",
         10956 => x"34",
         10957 => x"75",
         10958 => x"d1",
         10959 => x"81",
         10960 => x"77",
         10961 => x"59",
         10962 => x"56",
         10963 => x"fe",
         10964 => x"54",
         10965 => x"53",
         10966 => x"53",
         10967 => x"52",
         10968 => x"c9",
         10969 => x"84",
         10970 => x"7f",
         10971 => x"06",
         10972 => x"84",
         10973 => x"83",
         10974 => x"19",
         10975 => x"08",
         10976 => x"8c",
         10977 => x"74",
         10978 => x"27",
         10979 => x"82",
         10980 => x"74",
         10981 => x"81",
         10982 => x"38",
         10983 => x"19",
         10984 => x"08",
         10985 => x"52",
         10986 => x"51",
         10987 => x"3f",
         10988 => x"bb",
         10989 => x"1b",
         10990 => x"08",
         10991 => x"39",
         10992 => x"52",
         10993 => x"a3",
         10994 => x"ba",
         10995 => x"fc",
         10996 => x"16",
         10997 => x"9c",
         10998 => x"ba",
         10999 => x"06",
         11000 => x"b8",
         11001 => x"08",
         11002 => x"b2",
         11003 => x"91",
         11004 => x"0b",
         11005 => x"0c",
         11006 => x"04",
         11007 => x"1b",
         11008 => x"84",
         11009 => x"92",
         11010 => x"f0",
         11011 => x"65",
         11012 => x"40",
         11013 => x"7e",
         11014 => x"79",
         11015 => x"38",
         11016 => x"75",
         11017 => x"38",
         11018 => x"74",
         11019 => x"38",
         11020 => x"84",
         11021 => x"59",
         11022 => x"85",
         11023 => x"55",
         11024 => x"55",
         11025 => x"38",
         11026 => x"55",
         11027 => x"38",
         11028 => x"70",
         11029 => x"06",
         11030 => x"56",
         11031 => x"82",
         11032 => x"1a",
         11033 => x"5d",
         11034 => x"27",
         11035 => x"09",
         11036 => x"2e",
         11037 => x"76",
         11038 => x"5f",
         11039 => x"38",
         11040 => x"22",
         11041 => x"89",
         11042 => x"56",
         11043 => x"76",
         11044 => x"88",
         11045 => x"74",
         11046 => x"b1",
         11047 => x"2e",
         11048 => x"74",
         11049 => x"8c",
         11050 => x"1b",
         11051 => x"08",
         11052 => x"88",
         11053 => x"56",
         11054 => x"9c",
         11055 => x"81",
         11056 => x"1a",
         11057 => x"9c",
         11058 => x"05",
         11059 => x"77",
         11060 => x"38",
         11061 => x"70",
         11062 => x"18",
         11063 => x"57",
         11064 => x"85",
         11065 => x"15",
         11066 => x"59",
         11067 => x"2e",
         11068 => x"77",
         11069 => x"7f",
         11070 => x"76",
         11071 => x"77",
         11072 => x"7c",
         11073 => x"33",
         11074 => x"a1",
         11075 => x"8c",
         11076 => x"38",
         11077 => x"08",
         11078 => x"57",
         11079 => x"a5",
         11080 => x"0b",
         11081 => x"72",
         11082 => x"58",
         11083 => x"81",
         11084 => x"77",
         11085 => x"59",
         11086 => x"56",
         11087 => x"60",
         11088 => x"1a",
         11089 => x"2b",
         11090 => x"31",
         11091 => x"7f",
         11092 => x"94",
         11093 => x"70",
         11094 => x"0c",
         11095 => x"5a",
         11096 => x"5b",
         11097 => x"83",
         11098 => x"75",
         11099 => x"7a",
         11100 => x"90",
         11101 => x"77",
         11102 => x"5b",
         11103 => x"34",
         11104 => x"84",
         11105 => x"92",
         11106 => x"74",
         11107 => x"0c",
         11108 => x"04",
         11109 => x"55",
         11110 => x"38",
         11111 => x"a2",
         11112 => x"1b",
         11113 => x"76",
         11114 => x"84",
         11115 => x"5a",
         11116 => x"27",
         11117 => x"59",
         11118 => x"16",
         11119 => x"b6",
         11120 => x"83",
         11121 => x"5e",
         11122 => x"7f",
         11123 => x"06",
         11124 => x"81",
         11125 => x"b8",
         11126 => x"16",
         11127 => x"98",
         11128 => x"ba",
         11129 => x"2e",
         11130 => x"57",
         11131 => x"b4",
         11132 => x"83",
         11133 => x"94",
         11134 => x"ff",
         11135 => x"58",
         11136 => x"59",
         11137 => x"80",
         11138 => x"76",
         11139 => x"58",
         11140 => x"81",
         11141 => x"ff",
         11142 => x"ef",
         11143 => x"81",
         11144 => x"34",
         11145 => x"81",
         11146 => x"08",
         11147 => x"70",
         11148 => x"33",
         11149 => x"98",
         11150 => x"5c",
         11151 => x"08",
         11152 => x"81",
         11153 => x"38",
         11154 => x"08",
         11155 => x"b4",
         11156 => x"17",
         11157 => x"ba",
         11158 => x"55",
         11159 => x"08",
         11160 => x"38",
         11161 => x"55",
         11162 => x"09",
         11163 => x"e3",
         11164 => x"b4",
         11165 => x"17",
         11166 => x"7f",
         11167 => x"33",
         11168 => x"a9",
         11169 => x"fe",
         11170 => x"1a",
         11171 => x"1a",
         11172 => x"93",
         11173 => x"33",
         11174 => x"b9",
         11175 => x"b4",
         11176 => x"1b",
         11177 => x"7b",
         11178 => x"0c",
         11179 => x"39",
         11180 => x"52",
         11181 => x"ab",
         11182 => x"ba",
         11183 => x"84",
         11184 => x"fb",
         11185 => x"1a",
         11186 => x"ab",
         11187 => x"79",
         11188 => x"cc",
         11189 => x"8c",
         11190 => x"ba",
         11191 => x"bd",
         11192 => x"81",
         11193 => x"08",
         11194 => x"70",
         11195 => x"33",
         11196 => x"97",
         11197 => x"ba",
         11198 => x"b8",
         11199 => x"8c",
         11200 => x"34",
         11201 => x"a8",
         11202 => x"58",
         11203 => x"08",
         11204 => x"38",
         11205 => x"5c",
         11206 => x"09",
         11207 => x"fc",
         11208 => x"b4",
         11209 => x"17",
         11210 => x"76",
         11211 => x"33",
         11212 => x"f9",
         11213 => x"fb",
         11214 => x"16",
         11215 => x"95",
         11216 => x"ba",
         11217 => x"06",
         11218 => x"f2",
         11219 => x"08",
         11220 => x"ec",
         11221 => x"b4",
         11222 => x"b8",
         11223 => x"81",
         11224 => x"57",
         11225 => x"3f",
         11226 => x"08",
         11227 => x"84",
         11228 => x"83",
         11229 => x"16",
         11230 => x"08",
         11231 => x"a0",
         11232 => x"fe",
         11233 => x"16",
         11234 => x"82",
         11235 => x"06",
         11236 => x"81",
         11237 => x"08",
         11238 => x"05",
         11239 => x"81",
         11240 => x"ff",
         11241 => x"60",
         11242 => x"0c",
         11243 => x"58",
         11244 => x"39",
         11245 => x"1b",
         11246 => x"84",
         11247 => x"92",
         11248 => x"82",
         11249 => x"34",
         11250 => x"ba",
         11251 => x"3d",
         11252 => x"3d",
         11253 => x"89",
         11254 => x"2e",
         11255 => x"08",
         11256 => x"2e",
         11257 => x"33",
         11258 => x"2e",
         11259 => x"16",
         11260 => x"22",
         11261 => x"77",
         11262 => x"38",
         11263 => x"5c",
         11264 => x"81",
         11265 => x"18",
         11266 => x"2a",
         11267 => x"57",
         11268 => x"81",
         11269 => x"a0",
         11270 => x"57",
         11271 => x"79",
         11272 => x"83",
         11273 => x"7a",
         11274 => x"81",
         11275 => x"b8",
         11276 => x"17",
         11277 => x"93",
         11278 => x"ba",
         11279 => x"2e",
         11280 => x"59",
         11281 => x"b4",
         11282 => x"81",
         11283 => x"18",
         11284 => x"33",
         11285 => x"57",
         11286 => x"34",
         11287 => x"19",
         11288 => x"ff",
         11289 => x"5a",
         11290 => x"18",
         11291 => x"2a",
         11292 => x"18",
         11293 => x"76",
         11294 => x"5c",
         11295 => x"83",
         11296 => x"38",
         11297 => x"55",
         11298 => x"74",
         11299 => x"7a",
         11300 => x"74",
         11301 => x"75",
         11302 => x"74",
         11303 => x"78",
         11304 => x"80",
         11305 => x"0b",
         11306 => x"a1",
         11307 => x"34",
         11308 => x"99",
         11309 => x"0b",
         11310 => x"80",
         11311 => x"34",
         11312 => x"0b",
         11313 => x"7b",
         11314 => x"94",
         11315 => x"8c",
         11316 => x"33",
         11317 => x"5b",
         11318 => x"19",
         11319 => x"ba",
         11320 => x"3d",
         11321 => x"54",
         11322 => x"53",
         11323 => x"53",
         11324 => x"52",
         11325 => x"b5",
         11326 => x"84",
         11327 => x"fe",
         11328 => x"ba",
         11329 => x"18",
         11330 => x"08",
         11331 => x"31",
         11332 => x"08",
         11333 => x"a0",
         11334 => x"fe",
         11335 => x"17",
         11336 => x"82",
         11337 => x"06",
         11338 => x"81",
         11339 => x"08",
         11340 => x"05",
         11341 => x"81",
         11342 => x"ff",
         11343 => x"79",
         11344 => x"39",
         11345 => x"55",
         11346 => x"34",
         11347 => x"56",
         11348 => x"34",
         11349 => x"55",
         11350 => x"74",
         11351 => x"7a",
         11352 => x"74",
         11353 => x"75",
         11354 => x"74",
         11355 => x"78",
         11356 => x"80",
         11357 => x"0b",
         11358 => x"a1",
         11359 => x"34",
         11360 => x"99",
         11361 => x"0b",
         11362 => x"80",
         11363 => x"34",
         11364 => x"0b",
         11365 => x"7b",
         11366 => x"c4",
         11367 => x"8c",
         11368 => x"33",
         11369 => x"5b",
         11370 => x"19",
         11371 => x"39",
         11372 => x"51",
         11373 => x"3f",
         11374 => x"08",
         11375 => x"74",
         11376 => x"74",
         11377 => x"5a",
         11378 => x"f9",
         11379 => x"70",
         11380 => x"fe",
         11381 => x"8c",
         11382 => x"ba",
         11383 => x"38",
         11384 => x"80",
         11385 => x"74",
         11386 => x"80",
         11387 => x"72",
         11388 => x"80",
         11389 => x"86",
         11390 => x"16",
         11391 => x"71",
         11392 => x"38",
         11393 => x"58",
         11394 => x"84",
         11395 => x"0c",
         11396 => x"8c",
         11397 => x"0d",
         11398 => x"33",
         11399 => x"bc",
         11400 => x"8c",
         11401 => x"53",
         11402 => x"73",
         11403 => x"56",
         11404 => x"3d",
         11405 => x"70",
         11406 => x"75",
         11407 => x"38",
         11408 => x"05",
         11409 => x"9f",
         11410 => x"71",
         11411 => x"38",
         11412 => x"71",
         11413 => x"38",
         11414 => x"33",
         11415 => x"24",
         11416 => x"84",
         11417 => x"80",
         11418 => x"8c",
         11419 => x"0d",
         11420 => x"84",
         11421 => x"8c",
         11422 => x"78",
         11423 => x"70",
         11424 => x"53",
         11425 => x"89",
         11426 => x"82",
         11427 => x"ff",
         11428 => x"59",
         11429 => x"2e",
         11430 => x"80",
         11431 => x"fc",
         11432 => x"08",
         11433 => x"76",
         11434 => x"58",
         11435 => x"81",
         11436 => x"ff",
         11437 => x"54",
         11438 => x"26",
         11439 => x"12",
         11440 => x"06",
         11441 => x"9f",
         11442 => x"99",
         11443 => x"e0",
         11444 => x"ff",
         11445 => x"71",
         11446 => x"2a",
         11447 => x"73",
         11448 => x"06",
         11449 => x"ff",
         11450 => x"76",
         11451 => x"70",
         11452 => x"2a",
         11453 => x"52",
         11454 => x"2e",
         11455 => x"18",
         11456 => x"58",
         11457 => x"ff",
         11458 => x"51",
         11459 => x"77",
         11460 => x"38",
         11461 => x"51",
         11462 => x"ea",
         11463 => x"53",
         11464 => x"05",
         11465 => x"51",
         11466 => x"84",
         11467 => x"55",
         11468 => x"08",
         11469 => x"38",
         11470 => x"8c",
         11471 => x"0d",
         11472 => x"68",
         11473 => x"d0",
         11474 => x"94",
         11475 => x"8c",
         11476 => x"ba",
         11477 => x"c6",
         11478 => x"d7",
         11479 => x"98",
         11480 => x"80",
         11481 => x"e2",
         11482 => x"05",
         11483 => x"2a",
         11484 => x"59",
         11485 => x"b2",
         11486 => x"9b",
         11487 => x"12",
         11488 => x"2b",
         11489 => x"5e",
         11490 => x"58",
         11491 => x"a4",
         11492 => x"19",
         11493 => x"ba",
         11494 => x"3d",
         11495 => x"ba",
         11496 => x"2e",
         11497 => x"ff",
         11498 => x"0b",
         11499 => x"0c",
         11500 => x"04",
         11501 => x"94",
         11502 => x"98",
         11503 => x"2b",
         11504 => x"98",
         11505 => x"54",
         11506 => x"7e",
         11507 => x"58",
         11508 => x"8c",
         11509 => x"0d",
         11510 => x"3d",
         11511 => x"3d",
         11512 => x"3d",
         11513 => x"80",
         11514 => x"53",
         11515 => x"fd",
         11516 => x"80",
         11517 => x"cf",
         11518 => x"ba",
         11519 => x"84",
         11520 => x"83",
         11521 => x"80",
         11522 => x"7f",
         11523 => x"08",
         11524 => x"0c",
         11525 => x"3d",
         11526 => x"79",
         11527 => x"cc",
         11528 => x"3d",
         11529 => x"5b",
         11530 => x"51",
         11531 => x"3f",
         11532 => x"08",
         11533 => x"8c",
         11534 => x"38",
         11535 => x"3d",
         11536 => x"b4",
         11537 => x"2e",
         11538 => x"ba",
         11539 => x"17",
         11540 => x"7d",
         11541 => x"81",
         11542 => x"b8",
         11543 => x"16",
         11544 => x"8b",
         11545 => x"ba",
         11546 => x"2e",
         11547 => x"57",
         11548 => x"b4",
         11549 => x"82",
         11550 => x"df",
         11551 => x"11",
         11552 => x"33",
         11553 => x"07",
         11554 => x"5d",
         11555 => x"56",
         11556 => x"82",
         11557 => x"80",
         11558 => x"80",
         11559 => x"ff",
         11560 => x"84",
         11561 => x"59",
         11562 => x"08",
         11563 => x"80",
         11564 => x"ff",
         11565 => x"84",
         11566 => x"59",
         11567 => x"08",
         11568 => x"df",
         11569 => x"11",
         11570 => x"33",
         11571 => x"07",
         11572 => x"42",
         11573 => x"56",
         11574 => x"81",
         11575 => x"7a",
         11576 => x"84",
         11577 => x"52",
         11578 => x"a4",
         11579 => x"ba",
         11580 => x"84",
         11581 => x"80",
         11582 => x"38",
         11583 => x"83",
         11584 => x"81",
         11585 => x"e4",
         11586 => x"05",
         11587 => x"ff",
         11588 => x"78",
         11589 => x"33",
         11590 => x"80",
         11591 => x"82",
         11592 => x"17",
         11593 => x"33",
         11594 => x"7c",
         11595 => x"17",
         11596 => x"26",
         11597 => x"76",
         11598 => x"38",
         11599 => x"05",
         11600 => x"80",
         11601 => x"11",
         11602 => x"19",
         11603 => x"58",
         11604 => x"34",
         11605 => x"ff",
         11606 => x"3d",
         11607 => x"58",
         11608 => x"80",
         11609 => x"5a",
         11610 => x"38",
         11611 => x"82",
         11612 => x"0b",
         11613 => x"33",
         11614 => x"83",
         11615 => x"70",
         11616 => x"43",
         11617 => x"5a",
         11618 => x"8d",
         11619 => x"70",
         11620 => x"57",
         11621 => x"f5",
         11622 => x"5b",
         11623 => x"ab",
         11624 => x"76",
         11625 => x"38",
         11626 => x"7e",
         11627 => x"81",
         11628 => x"81",
         11629 => x"77",
         11630 => x"ba",
         11631 => x"05",
         11632 => x"ff",
         11633 => x"06",
         11634 => x"91",
         11635 => x"34",
         11636 => x"8c",
         11637 => x"3d",
         11638 => x"16",
         11639 => x"33",
         11640 => x"71",
         11641 => x"79",
         11642 => x"5e",
         11643 => x"95",
         11644 => x"17",
         11645 => x"2b",
         11646 => x"07",
         11647 => x"dd",
         11648 => x"5d",
         11649 => x"51",
         11650 => x"3f",
         11651 => x"08",
         11652 => x"8c",
         11653 => x"fd",
         11654 => x"b1",
         11655 => x"b4",
         11656 => x"b8",
         11657 => x"81",
         11658 => x"5e",
         11659 => x"3f",
         11660 => x"ba",
         11661 => x"be",
         11662 => x"8c",
         11663 => x"34",
         11664 => x"a8",
         11665 => x"84",
         11666 => x"5a",
         11667 => x"17",
         11668 => x"83",
         11669 => x"33",
         11670 => x"2e",
         11671 => x"fb",
         11672 => x"54",
         11673 => x"a0",
         11674 => x"53",
         11675 => x"16",
         11676 => x"88",
         11677 => x"59",
         11678 => x"ff",
         11679 => x"3d",
         11680 => x"58",
         11681 => x"80",
         11682 => x"e8",
         11683 => x"10",
         11684 => x"05",
         11685 => x"33",
         11686 => x"5e",
         11687 => x"2e",
         11688 => x"fd",
         11689 => x"f1",
         11690 => x"3d",
         11691 => x"19",
         11692 => x"33",
         11693 => x"05",
         11694 => x"60",
         11695 => x"38",
         11696 => x"08",
         11697 => x"59",
         11698 => x"7c",
         11699 => x"5e",
         11700 => x"26",
         11701 => x"f5",
         11702 => x"80",
         11703 => x"84",
         11704 => x"80",
         11705 => x"04",
         11706 => x"7b",
         11707 => x"89",
         11708 => x"2e",
         11709 => x"08",
         11710 => x"2e",
         11711 => x"33",
         11712 => x"2e",
         11713 => x"14",
         11714 => x"22",
         11715 => x"78",
         11716 => x"38",
         11717 => x"5a",
         11718 => x"81",
         11719 => x"15",
         11720 => x"81",
         11721 => x"15",
         11722 => x"76",
         11723 => x"38",
         11724 => x"54",
         11725 => x"78",
         11726 => x"38",
         11727 => x"22",
         11728 => x"52",
         11729 => x"78",
         11730 => x"38",
         11731 => x"17",
         11732 => x"d3",
         11733 => x"8c",
         11734 => x"77",
         11735 => x"55",
         11736 => x"c3",
         11737 => x"8c",
         11738 => x"81",
         11739 => x"30",
         11740 => x"94",
         11741 => x"71",
         11742 => x"08",
         11743 => x"73",
         11744 => x"98",
         11745 => x"27",
         11746 => x"76",
         11747 => x"16",
         11748 => x"17",
         11749 => x"33",
         11750 => x"81",
         11751 => x"57",
         11752 => x"81",
         11753 => x"52",
         11754 => x"99",
         11755 => x"ba",
         11756 => x"84",
         11757 => x"80",
         11758 => x"38",
         11759 => x"98",
         11760 => x"27",
         11761 => x"79",
         11762 => x"14",
         11763 => x"aa",
         11764 => x"16",
         11765 => x"39",
         11766 => x"16",
         11767 => x"72",
         11768 => x"0c",
         11769 => x"04",
         11770 => x"70",
         11771 => x"06",
         11772 => x"fe",
         11773 => x"94",
         11774 => x"57",
         11775 => x"78",
         11776 => x"06",
         11777 => x"77",
         11778 => x"94",
         11779 => x"75",
         11780 => x"38",
         11781 => x"0c",
         11782 => x"80",
         11783 => x"76",
         11784 => x"73",
         11785 => x"59",
         11786 => x"8c",
         11787 => x"08",
         11788 => x"38",
         11789 => x"0c",
         11790 => x"ba",
         11791 => x"3d",
         11792 => x"0b",
         11793 => x"88",
         11794 => x"73",
         11795 => x"fe",
         11796 => x"16",
         11797 => x"2e",
         11798 => x"fe",
         11799 => x"ba",
         11800 => x"94",
         11801 => x"94",
         11802 => x"83",
         11803 => x"75",
         11804 => x"38",
         11805 => x"9c",
         11806 => x"05",
         11807 => x"73",
         11808 => x"f6",
         11809 => x"22",
         11810 => x"b0",
         11811 => x"78",
         11812 => x"5a",
         11813 => x"80",
         11814 => x"38",
         11815 => x"56",
         11816 => x"73",
         11817 => x"ff",
         11818 => x"84",
         11819 => x"54",
         11820 => x"81",
         11821 => x"ff",
         11822 => x"84",
         11823 => x"81",
         11824 => x"fc",
         11825 => x"75",
         11826 => x"fc",
         11827 => x"52",
         11828 => x"97",
         11829 => x"ba",
         11830 => x"84",
         11831 => x"81",
         11832 => x"84",
         11833 => x"ff",
         11834 => x"38",
         11835 => x"08",
         11836 => x"73",
         11837 => x"fe",
         11838 => x"0b",
         11839 => x"82",
         11840 => x"8c",
         11841 => x"0d",
         11842 => x"0d",
         11843 => x"54",
         11844 => x"a2",
         11845 => x"8c",
         11846 => x"52",
         11847 => x"05",
         11848 => x"3f",
         11849 => x"08",
         11850 => x"8c",
         11851 => x"8f",
         11852 => x"0c",
         11853 => x"84",
         11854 => x"8c",
         11855 => x"7a",
         11856 => x"52",
         11857 => x"b9",
         11858 => x"ba",
         11859 => x"84",
         11860 => x"80",
         11861 => x"16",
         11862 => x"2b",
         11863 => x"78",
         11864 => x"86",
         11865 => x"84",
         11866 => x"5b",
         11867 => x"2e",
         11868 => x"9c",
         11869 => x"11",
         11870 => x"33",
         11871 => x"07",
         11872 => x"5d",
         11873 => x"57",
         11874 => x"b3",
         11875 => x"17",
         11876 => x"86",
         11877 => x"17",
         11878 => x"75",
         11879 => x"b9",
         11880 => x"8c",
         11881 => x"84",
         11882 => x"74",
         11883 => x"84",
         11884 => x"0c",
         11885 => x"85",
         11886 => x"0c",
         11887 => x"95",
         11888 => x"18",
         11889 => x"2b",
         11890 => x"07",
         11891 => x"19",
         11892 => x"ff",
         11893 => x"3d",
         11894 => x"89",
         11895 => x"2e",
         11896 => x"08",
         11897 => x"2e",
         11898 => x"33",
         11899 => x"2e",
         11900 => x"13",
         11901 => x"22",
         11902 => x"76",
         11903 => x"80",
         11904 => x"73",
         11905 => x"75",
         11906 => x"ba",
         11907 => x"3d",
         11908 => x"13",
         11909 => x"ff",
         11910 => x"ba",
         11911 => x"06",
         11912 => x"38",
         11913 => x"53",
         11914 => x"f8",
         11915 => x"7c",
         11916 => x"56",
         11917 => x"9f",
         11918 => x"54",
         11919 => x"97",
         11920 => x"53",
         11921 => x"8f",
         11922 => x"22",
         11923 => x"59",
         11924 => x"2e",
         11925 => x"80",
         11926 => x"75",
         11927 => x"c7",
         11928 => x"2e",
         11929 => x"75",
         11930 => x"ff",
         11931 => x"84",
         11932 => x"53",
         11933 => x"08",
         11934 => x"38",
         11935 => x"08",
         11936 => x"52",
         11937 => x"b2",
         11938 => x"52",
         11939 => x"99",
         11940 => x"ba",
         11941 => x"32",
         11942 => x"72",
         11943 => x"84",
         11944 => x"06",
         11945 => x"72",
         11946 => x"0c",
         11947 => x"04",
         11948 => x"75",
         11949 => x"b1",
         11950 => x"52",
         11951 => x"99",
         11952 => x"ba",
         11953 => x"32",
         11954 => x"72",
         11955 => x"84",
         11956 => x"06",
         11957 => x"cf",
         11958 => x"74",
         11959 => x"f9",
         11960 => x"8c",
         11961 => x"8c",
         11962 => x"0d",
         11963 => x"33",
         11964 => x"e8",
         11965 => x"8c",
         11966 => x"53",
         11967 => x"38",
         11968 => x"54",
         11969 => x"39",
         11970 => x"66",
         11971 => x"89",
         11972 => x"97",
         11973 => x"c1",
         11974 => x"ba",
         11975 => x"84",
         11976 => x"80",
         11977 => x"74",
         11978 => x"0c",
         11979 => x"04",
         11980 => x"51",
         11981 => x"3f",
         11982 => x"08",
         11983 => x"8c",
         11984 => x"02",
         11985 => x"33",
         11986 => x"55",
         11987 => x"24",
         11988 => x"80",
         11989 => x"76",
         11990 => x"ff",
         11991 => x"74",
         11992 => x"0c",
         11993 => x"04",
         11994 => x"ba",
         11995 => x"3d",
         11996 => x"3d",
         11997 => x"56",
         11998 => x"95",
         11999 => x"52",
         12000 => x"c0",
         12001 => x"ba",
         12002 => x"84",
         12003 => x"9a",
         12004 => x"0c",
         12005 => x"11",
         12006 => x"94",
         12007 => x"57",
         12008 => x"75",
         12009 => x"75",
         12010 => x"84",
         12011 => x"95",
         12012 => x"84",
         12013 => x"77",
         12014 => x"78",
         12015 => x"93",
         12016 => x"18",
         12017 => x"8c",
         12018 => x"59",
         12019 => x"38",
         12020 => x"71",
         12021 => x"b4",
         12022 => x"2e",
         12023 => x"83",
         12024 => x"5f",
         12025 => x"8d",
         12026 => x"75",
         12027 => x"52",
         12028 => x"51",
         12029 => x"3f",
         12030 => x"08",
         12031 => x"38",
         12032 => x"5e",
         12033 => x"0c",
         12034 => x"57",
         12035 => x"38",
         12036 => x"7d",
         12037 => x"8d",
         12038 => x"b8",
         12039 => x"33",
         12040 => x"71",
         12041 => x"88",
         12042 => x"14",
         12043 => x"07",
         12044 => x"33",
         12045 => x"ff",
         12046 => x"07",
         12047 => x"80",
         12048 => x"60",
         12049 => x"ff",
         12050 => x"05",
         12051 => x"53",
         12052 => x"58",
         12053 => x"78",
         12054 => x"7a",
         12055 => x"94",
         12056 => x"17",
         12057 => x"58",
         12058 => x"34",
         12059 => x"8c",
         12060 => x"0d",
         12061 => x"b4",
         12062 => x"b8",
         12063 => x"81",
         12064 => x"5d",
         12065 => x"3f",
         12066 => x"ba",
         12067 => x"f8",
         12068 => x"8c",
         12069 => x"34",
         12070 => x"a8",
         12071 => x"84",
         12072 => x"5f",
         12073 => x"18",
         12074 => x"bd",
         12075 => x"33",
         12076 => x"2e",
         12077 => x"fe",
         12078 => x"54",
         12079 => x"a0",
         12080 => x"53",
         12081 => x"17",
         12082 => x"fb",
         12083 => x"5e",
         12084 => x"82",
         12085 => x"3d",
         12086 => x"52",
         12087 => x"81",
         12088 => x"ba",
         12089 => x"2e",
         12090 => x"84",
         12091 => x"81",
         12092 => x"38",
         12093 => x"08",
         12094 => x"ba",
         12095 => x"80",
         12096 => x"81",
         12097 => x"58",
         12098 => x"17",
         12099 => x"ca",
         12100 => x"0c",
         12101 => x"0c",
         12102 => x"81",
         12103 => x"84",
         12104 => x"c8",
         12105 => x"b8",
         12106 => x"33",
         12107 => x"88",
         12108 => x"30",
         12109 => x"1f",
         12110 => x"ff",
         12111 => x"5f",
         12112 => x"5f",
         12113 => x"fd",
         12114 => x"8f",
         12115 => x"fd",
         12116 => x"60",
         12117 => x"7f",
         12118 => x"18",
         12119 => x"33",
         12120 => x"77",
         12121 => x"fe",
         12122 => x"60",
         12123 => x"39",
         12124 => x"7b",
         12125 => x"76",
         12126 => x"38",
         12127 => x"74",
         12128 => x"38",
         12129 => x"73",
         12130 => x"38",
         12131 => x"84",
         12132 => x"59",
         12133 => x"81",
         12134 => x"54",
         12135 => x"80",
         12136 => x"17",
         12137 => x"80",
         12138 => x"17",
         12139 => x"2a",
         12140 => x"58",
         12141 => x"80",
         12142 => x"38",
         12143 => x"54",
         12144 => x"08",
         12145 => x"73",
         12146 => x"88",
         12147 => x"08",
         12148 => x"74",
         12149 => x"9c",
         12150 => x"26",
         12151 => x"56",
         12152 => x"18",
         12153 => x"08",
         12154 => x"77",
         12155 => x"59",
         12156 => x"34",
         12157 => x"85",
         12158 => x"18",
         12159 => x"74",
         12160 => x"0c",
         12161 => x"04",
         12162 => x"78",
         12163 => x"38",
         12164 => x"51",
         12165 => x"3f",
         12166 => x"08",
         12167 => x"8c",
         12168 => x"80",
         12169 => x"ba",
         12170 => x"2e",
         12171 => x"84",
         12172 => x"ff",
         12173 => x"38",
         12174 => x"52",
         12175 => x"85",
         12176 => x"ba",
         12177 => x"c8",
         12178 => x"08",
         12179 => x"18",
         12180 => x"58",
         12181 => x"ff",
         12182 => x"15",
         12183 => x"84",
         12184 => x"07",
         12185 => x"17",
         12186 => x"77",
         12187 => x"a0",
         12188 => x"81",
         12189 => x"fe",
         12190 => x"84",
         12191 => x"81",
         12192 => x"fe",
         12193 => x"77",
         12194 => x"fe",
         12195 => x"0b",
         12196 => x"59",
         12197 => x"80",
         12198 => x"0c",
         12199 => x"98",
         12200 => x"76",
         12201 => x"b9",
         12202 => x"8c",
         12203 => x"81",
         12204 => x"ba",
         12205 => x"2e",
         12206 => x"75",
         12207 => x"79",
         12208 => x"8c",
         12209 => x"08",
         12210 => x"38",
         12211 => x"08",
         12212 => x"78",
         12213 => x"54",
         12214 => x"ba",
         12215 => x"81",
         12216 => x"ba",
         12217 => x"17",
         12218 => x"96",
         12219 => x"2e",
         12220 => x"53",
         12221 => x"51",
         12222 => x"3f",
         12223 => x"08",
         12224 => x"8c",
         12225 => x"38",
         12226 => x"51",
         12227 => x"3f",
         12228 => x"08",
         12229 => x"8c",
         12230 => x"80",
         12231 => x"ba",
         12232 => x"2e",
         12233 => x"84",
         12234 => x"ff",
         12235 => x"38",
         12236 => x"52",
         12237 => x"83",
         12238 => x"ba",
         12239 => x"e6",
         12240 => x"08",
         12241 => x"18",
         12242 => x"58",
         12243 => x"90",
         12244 => x"94",
         12245 => x"16",
         12246 => x"54",
         12247 => x"34",
         12248 => x"79",
         12249 => x"38",
         12250 => x"56",
         12251 => x"58",
         12252 => x"81",
         12253 => x"39",
         12254 => x"18",
         12255 => x"fc",
         12256 => x"56",
         12257 => x"0b",
         12258 => x"59",
         12259 => x"39",
         12260 => x"08",
         12261 => x"59",
         12262 => x"39",
         12263 => x"18",
         12264 => x"fd",
         12265 => x"ba",
         12266 => x"c0",
         12267 => x"ff",
         12268 => x"3d",
         12269 => x"a7",
         12270 => x"05",
         12271 => x"51",
         12272 => x"3f",
         12273 => x"08",
         12274 => x"8c",
         12275 => x"8a",
         12276 => x"ba",
         12277 => x"3d",
         12278 => x"4b",
         12279 => x"52",
         12280 => x"52",
         12281 => x"f8",
         12282 => x"8c",
         12283 => x"ba",
         12284 => x"38",
         12285 => x"05",
         12286 => x"2a",
         12287 => x"57",
         12288 => x"cd",
         12289 => x"2b",
         12290 => x"24",
         12291 => x"80",
         12292 => x"70",
         12293 => x"57",
         12294 => x"ff",
         12295 => x"a3",
         12296 => x"11",
         12297 => x"33",
         12298 => x"07",
         12299 => x"5e",
         12300 => x"7c",
         12301 => x"d5",
         12302 => x"2a",
         12303 => x"76",
         12304 => x"ed",
         12305 => x"98",
         12306 => x"2e",
         12307 => x"77",
         12308 => x"84",
         12309 => x"52",
         12310 => x"52",
         12311 => x"f9",
         12312 => x"8c",
         12313 => x"ba",
         12314 => x"e5",
         12315 => x"8c",
         12316 => x"51",
         12317 => x"3f",
         12318 => x"08",
         12319 => x"8c",
         12320 => x"87",
         12321 => x"8c",
         12322 => x"0d",
         12323 => x"33",
         12324 => x"71",
         12325 => x"90",
         12326 => x"07",
         12327 => x"ff",
         12328 => x"ba",
         12329 => x"2e",
         12330 => x"ba",
         12331 => x"a1",
         12332 => x"6f",
         12333 => x"57",
         12334 => x"ff",
         12335 => x"38",
         12336 => x"51",
         12337 => x"3f",
         12338 => x"08",
         12339 => x"8c",
         12340 => x"be",
         12341 => x"70",
         12342 => x"25",
         12343 => x"80",
         12344 => x"74",
         12345 => x"38",
         12346 => x"58",
         12347 => x"27",
         12348 => x"17",
         12349 => x"81",
         12350 => x"56",
         12351 => x"38",
         12352 => x"f5",
         12353 => x"ba",
         12354 => x"ba",
         12355 => x"3d",
         12356 => x"17",
         12357 => x"08",
         12358 => x"b4",
         12359 => x"2e",
         12360 => x"83",
         12361 => x"59",
         12362 => x"2e",
         12363 => x"80",
         12364 => x"54",
         12365 => x"17",
         12366 => x"33",
         12367 => x"ee",
         12368 => x"8c",
         12369 => x"85",
         12370 => x"81",
         12371 => x"18",
         12372 => x"77",
         12373 => x"19",
         12374 => x"78",
         12375 => x"83",
         12376 => x"19",
         12377 => x"fe",
         12378 => x"52",
         12379 => x"8b",
         12380 => x"ba",
         12381 => x"84",
         12382 => x"80",
         12383 => x"38",
         12384 => x"09",
         12385 => x"cd",
         12386 => x"fe",
         12387 => x"54",
         12388 => x"53",
         12389 => x"17",
         12390 => x"f2",
         12391 => x"58",
         12392 => x"08",
         12393 => x"81",
         12394 => x"38",
         12395 => x"08",
         12396 => x"b4",
         12397 => x"18",
         12398 => x"ba",
         12399 => x"55",
         12400 => x"08",
         12401 => x"38",
         12402 => x"55",
         12403 => x"09",
         12404 => x"de",
         12405 => x"b4",
         12406 => x"18",
         12407 => x"7c",
         12408 => x"33",
         12409 => x"c5",
         12410 => x"fe",
         12411 => x"55",
         12412 => x"80",
         12413 => x"52",
         12414 => x"f6",
         12415 => x"ba",
         12416 => x"84",
         12417 => x"80",
         12418 => x"38",
         12419 => x"08",
         12420 => x"e6",
         12421 => x"8c",
         12422 => x"80",
         12423 => x"53",
         12424 => x"51",
         12425 => x"3f",
         12426 => x"08",
         12427 => x"17",
         12428 => x"94",
         12429 => x"5c",
         12430 => x"27",
         12431 => x"81",
         12432 => x"0c",
         12433 => x"81",
         12434 => x"84",
         12435 => x"55",
         12436 => x"ff",
         12437 => x"56",
         12438 => x"79",
         12439 => x"39",
         12440 => x"08",
         12441 => x"39",
         12442 => x"90",
         12443 => x"0d",
         12444 => x"3d",
         12445 => x"52",
         12446 => x"ff",
         12447 => x"84",
         12448 => x"56",
         12449 => x"08",
         12450 => x"38",
         12451 => x"8c",
         12452 => x"0d",
         12453 => x"6f",
         12454 => x"70",
         12455 => x"a6",
         12456 => x"ba",
         12457 => x"84",
         12458 => x"8b",
         12459 => x"84",
         12460 => x"9f",
         12461 => x"84",
         12462 => x"84",
         12463 => x"06",
         12464 => x"80",
         12465 => x"70",
         12466 => x"06",
         12467 => x"56",
         12468 => x"38",
         12469 => x"52",
         12470 => x"52",
         12471 => x"c0",
         12472 => x"8c",
         12473 => x"5c",
         12474 => x"08",
         12475 => x"56",
         12476 => x"08",
         12477 => x"f9",
         12478 => x"8c",
         12479 => x"81",
         12480 => x"81",
         12481 => x"84",
         12482 => x"83",
         12483 => x"5a",
         12484 => x"e2",
         12485 => x"9c",
         12486 => x"05",
         12487 => x"5b",
         12488 => x"8d",
         12489 => x"22",
         12490 => x"b0",
         12491 => x"5c",
         12492 => x"18",
         12493 => x"59",
         12494 => x"57",
         12495 => x"70",
         12496 => x"34",
         12497 => x"74",
         12498 => x"58",
         12499 => x"55",
         12500 => x"81",
         12501 => x"54",
         12502 => x"78",
         12503 => x"33",
         12504 => x"c9",
         12505 => x"8c",
         12506 => x"38",
         12507 => x"dc",
         12508 => x"ff",
         12509 => x"54",
         12510 => x"53",
         12511 => x"53",
         12512 => x"52",
         12513 => x"a5",
         12514 => x"84",
         12515 => x"be",
         12516 => x"8c",
         12517 => x"34",
         12518 => x"a8",
         12519 => x"55",
         12520 => x"08",
         12521 => x"38",
         12522 => x"5b",
         12523 => x"09",
         12524 => x"e1",
         12525 => x"b4",
         12526 => x"18",
         12527 => x"77",
         12528 => x"33",
         12529 => x"e5",
         12530 => x"39",
         12531 => x"7d",
         12532 => x"81",
         12533 => x"b4",
         12534 => x"18",
         12535 => x"ac",
         12536 => x"7c",
         12537 => x"f9",
         12538 => x"8c",
         12539 => x"ba",
         12540 => x"2e",
         12541 => x"84",
         12542 => x"81",
         12543 => x"38",
         12544 => x"08",
         12545 => x"84",
         12546 => x"74",
         12547 => x"fe",
         12548 => x"84",
         12549 => x"fc",
         12550 => x"17",
         12551 => x"94",
         12552 => x"5c",
         12553 => x"27",
         12554 => x"18",
         12555 => x"84",
         12556 => x"07",
         12557 => x"18",
         12558 => x"78",
         12559 => x"a1",
         12560 => x"ba",
         12561 => x"3d",
         12562 => x"17",
         12563 => x"83",
         12564 => x"57",
         12565 => x"78",
         12566 => x"06",
         12567 => x"8b",
         12568 => x"56",
         12569 => x"70",
         12570 => x"34",
         12571 => x"75",
         12572 => x"57",
         12573 => x"18",
         12574 => x"90",
         12575 => x"19",
         12576 => x"75",
         12577 => x"34",
         12578 => x"1a",
         12579 => x"80",
         12580 => x"80",
         12581 => x"d1",
         12582 => x"7c",
         12583 => x"06",
         12584 => x"80",
         12585 => x"77",
         12586 => x"7a",
         12587 => x"34",
         12588 => x"74",
         12589 => x"cc",
         12590 => x"a0",
         12591 => x"1a",
         12592 => x"58",
         12593 => x"81",
         12594 => x"77",
         12595 => x"59",
         12596 => x"56",
         12597 => x"7d",
         12598 => x"80",
         12599 => x"64",
         12600 => x"ff",
         12601 => x"57",
         12602 => x"f2",
         12603 => x"88",
         12604 => x"80",
         12605 => x"75",
         12606 => x"83",
         12607 => x"38",
         12608 => x"0b",
         12609 => x"79",
         12610 => x"96",
         12611 => x"8c",
         12612 => x"ba",
         12613 => x"b6",
         12614 => x"84",
         12615 => x"96",
         12616 => x"ba",
         12617 => x"17",
         12618 => x"98",
         12619 => x"cc",
         12620 => x"34",
         12621 => x"5d",
         12622 => x"34",
         12623 => x"59",
         12624 => x"34",
         12625 => x"79",
         12626 => x"d9",
         12627 => x"90",
         12628 => x"34",
         12629 => x"0b",
         12630 => x"7d",
         12631 => x"80",
         12632 => x"8c",
         12633 => x"84",
         12634 => x"9f",
         12635 => x"76",
         12636 => x"74",
         12637 => x"34",
         12638 => x"57",
         12639 => x"17",
         12640 => x"39",
         12641 => x"5b",
         12642 => x"17",
         12643 => x"2a",
         12644 => x"cd",
         12645 => x"59",
         12646 => x"d8",
         12647 => x"57",
         12648 => x"a1",
         12649 => x"2a",
         12650 => x"18",
         12651 => x"2a",
         12652 => x"18",
         12653 => x"90",
         12654 => x"34",
         12655 => x"0b",
         12656 => x"7d",
         12657 => x"98",
         12658 => x"8c",
         12659 => x"96",
         12660 => x"0d",
         12661 => x"3d",
         12662 => x"5b",
         12663 => x"2e",
         12664 => x"70",
         12665 => x"33",
         12666 => x"56",
         12667 => x"2e",
         12668 => x"74",
         12669 => x"ba",
         12670 => x"38",
         12671 => x"3d",
         12672 => x"52",
         12673 => x"ff",
         12674 => x"84",
         12675 => x"56",
         12676 => x"08",
         12677 => x"38",
         12678 => x"8c",
         12679 => x"0d",
         12680 => x"3d",
         12681 => x"08",
         12682 => x"70",
         12683 => x"9f",
         12684 => x"ba",
         12685 => x"84",
         12686 => x"dc",
         12687 => x"bb",
         12688 => x"a0",
         12689 => x"56",
         12690 => x"a0",
         12691 => x"ae",
         12692 => x"58",
         12693 => x"81",
         12694 => x"77",
         12695 => x"59",
         12696 => x"55",
         12697 => x"99",
         12698 => x"78",
         12699 => x"55",
         12700 => x"05",
         12701 => x"70",
         12702 => x"34",
         12703 => x"74",
         12704 => x"3d",
         12705 => x"51",
         12706 => x"3f",
         12707 => x"08",
         12708 => x"8c",
         12709 => x"38",
         12710 => x"08",
         12711 => x"38",
         12712 => x"ba",
         12713 => x"3d",
         12714 => x"33",
         12715 => x"81",
         12716 => x"57",
         12717 => x"26",
         12718 => x"17",
         12719 => x"06",
         12720 => x"59",
         12721 => x"80",
         12722 => x"7f",
         12723 => x"fc",
         12724 => x"5d",
         12725 => x"5c",
         12726 => x"05",
         12727 => x"70",
         12728 => x"33",
         12729 => x"5a",
         12730 => x"99",
         12731 => x"e0",
         12732 => x"ff",
         12733 => x"ff",
         12734 => x"77",
         12735 => x"38",
         12736 => x"81",
         12737 => x"55",
         12738 => x"9f",
         12739 => x"75",
         12740 => x"81",
         12741 => x"77",
         12742 => x"78",
         12743 => x"30",
         12744 => x"9f",
         12745 => x"5d",
         12746 => x"80",
         12747 => x"81",
         12748 => x"5e",
         12749 => x"24",
         12750 => x"7c",
         12751 => x"5b",
         12752 => x"7b",
         12753 => x"b4",
         12754 => x"0c",
         12755 => x"3d",
         12756 => x"52",
         12757 => x"ff",
         12758 => x"84",
         12759 => x"56",
         12760 => x"08",
         12761 => x"fd",
         12762 => x"aa",
         12763 => x"09",
         12764 => x"ac",
         12765 => x"ff",
         12766 => x"84",
         12767 => x"56",
         12768 => x"08",
         12769 => x"6f",
         12770 => x"8d",
         12771 => x"05",
         12772 => x"58",
         12773 => x"70",
         12774 => x"33",
         12775 => x"05",
         12776 => x"1a",
         12777 => x"38",
         12778 => x"05",
         12779 => x"34",
         12780 => x"70",
         12781 => x"06",
         12782 => x"89",
         12783 => x"07",
         12784 => x"19",
         12785 => x"81",
         12786 => x"34",
         12787 => x"70",
         12788 => x"06",
         12789 => x"80",
         12790 => x"38",
         12791 => x"6b",
         12792 => x"38",
         12793 => x"33",
         12794 => x"71",
         12795 => x"72",
         12796 => x"5c",
         12797 => x"2e",
         12798 => x"fe",
         12799 => x"08",
         12800 => x"56",
         12801 => x"82",
         12802 => x"17",
         12803 => x"29",
         12804 => x"05",
         12805 => x"80",
         12806 => x"38",
         12807 => x"58",
         12808 => x"76",
         12809 => x"83",
         12810 => x"7e",
         12811 => x"81",
         12812 => x"b8",
         12813 => x"17",
         12814 => x"e3",
         12815 => x"ba",
         12816 => x"2e",
         12817 => x"58",
         12818 => x"b4",
         12819 => x"57",
         12820 => x"18",
         12821 => x"fb",
         12822 => x"15",
         12823 => x"ae",
         12824 => x"06",
         12825 => x"70",
         12826 => x"06",
         12827 => x"80",
         12828 => x"7b",
         12829 => x"77",
         12830 => x"34",
         12831 => x"7a",
         12832 => x"81",
         12833 => x"75",
         12834 => x"7d",
         12835 => x"34",
         12836 => x"56",
         12837 => x"18",
         12838 => x"81",
         12839 => x"34",
         12840 => x"3d",
         12841 => x"08",
         12842 => x"74",
         12843 => x"38",
         12844 => x"51",
         12845 => x"3f",
         12846 => x"08",
         12847 => x"8c",
         12848 => x"38",
         12849 => x"98",
         12850 => x"80",
         12851 => x"08",
         12852 => x"38",
         12853 => x"7a",
         12854 => x"7a",
         12855 => x"06",
         12856 => x"81",
         12857 => x"b8",
         12858 => x"16",
         12859 => x"e2",
         12860 => x"ba",
         12861 => x"2e",
         12862 => x"57",
         12863 => x"b4",
         12864 => x"55",
         12865 => x"9c",
         12866 => x"e5",
         12867 => x"0b",
         12868 => x"90",
         12869 => x"27",
         12870 => x"52",
         12871 => x"fc",
         12872 => x"ba",
         12873 => x"84",
         12874 => x"80",
         12875 => x"38",
         12876 => x"84",
         12877 => x"38",
         12878 => x"f9",
         12879 => x"51",
         12880 => x"3f",
         12881 => x"08",
         12882 => x"0c",
         12883 => x"04",
         12884 => x"ba",
         12885 => x"3d",
         12886 => x"18",
         12887 => x"33",
         12888 => x"71",
         12889 => x"78",
         12890 => x"5c",
         12891 => x"84",
         12892 => x"84",
         12893 => x"38",
         12894 => x"08",
         12895 => x"a0",
         12896 => x"ba",
         12897 => x"3d",
         12898 => x"54",
         12899 => x"53",
         12900 => x"16",
         12901 => x"e2",
         12902 => x"58",
         12903 => x"08",
         12904 => x"81",
         12905 => x"38",
         12906 => x"08",
         12907 => x"b4",
         12908 => x"17",
         12909 => x"ba",
         12910 => x"55",
         12911 => x"08",
         12912 => x"38",
         12913 => x"5d",
         12914 => x"09",
         12915 => x"93",
         12916 => x"b4",
         12917 => x"17",
         12918 => x"7b",
         12919 => x"33",
         12920 => x"c9",
         12921 => x"fd",
         12922 => x"54",
         12923 => x"53",
         12924 => x"53",
         12925 => x"52",
         12926 => x"b1",
         12927 => x"84",
         12928 => x"fc",
         12929 => x"ba",
         12930 => x"18",
         12931 => x"08",
         12932 => x"31",
         12933 => x"08",
         12934 => x"a0",
         12935 => x"fc",
         12936 => x"17",
         12937 => x"82",
         12938 => x"06",
         12939 => x"81",
         12940 => x"08",
         12941 => x"05",
         12942 => x"81",
         12943 => x"fe",
         12944 => x"79",
         12945 => x"39",
         12946 => x"02",
         12947 => x"33",
         12948 => x"80",
         12949 => x"56",
         12950 => x"96",
         12951 => x"52",
         12952 => x"ff",
         12953 => x"84",
         12954 => x"56",
         12955 => x"08",
         12956 => x"38",
         12957 => x"8c",
         12958 => x"0d",
         12959 => x"66",
         12960 => x"d0",
         12961 => x"96",
         12962 => x"ba",
         12963 => x"84",
         12964 => x"e0",
         12965 => x"cf",
         12966 => x"a0",
         12967 => x"56",
         12968 => x"74",
         12969 => x"71",
         12970 => x"33",
         12971 => x"74",
         12972 => x"56",
         12973 => x"8b",
         12974 => x"55",
         12975 => x"16",
         12976 => x"fe",
         12977 => x"84",
         12978 => x"84",
         12979 => x"96",
         12980 => x"ec",
         12981 => x"57",
         12982 => x"3d",
         12983 => x"97",
         12984 => x"a1",
         12985 => x"ba",
         12986 => x"84",
         12987 => x"80",
         12988 => x"74",
         12989 => x"0c",
         12990 => x"04",
         12991 => x"52",
         12992 => x"05",
         12993 => x"d8",
         12994 => x"8c",
         12995 => x"ba",
         12996 => x"38",
         12997 => x"05",
         12998 => x"06",
         12999 => x"75",
         13000 => x"84",
         13001 => x"19",
         13002 => x"2b",
         13003 => x"56",
         13004 => x"34",
         13005 => x"55",
         13006 => x"34",
         13007 => x"58",
         13008 => x"34",
         13009 => x"54",
         13010 => x"34",
         13011 => x"0b",
         13012 => x"78",
         13013 => x"88",
         13014 => x"8c",
         13015 => x"8c",
         13016 => x"0d",
         13017 => x"0d",
         13018 => x"5b",
         13019 => x"3d",
         13020 => x"9b",
         13021 => x"a0",
         13022 => x"ba",
         13023 => x"ba",
         13024 => x"70",
         13025 => x"08",
         13026 => x"51",
         13027 => x"80",
         13028 => x"81",
         13029 => x"5a",
         13030 => x"a4",
         13031 => x"70",
         13032 => x"25",
         13033 => x"80",
         13034 => x"38",
         13035 => x"06",
         13036 => x"80",
         13037 => x"38",
         13038 => x"08",
         13039 => x"5a",
         13040 => x"77",
         13041 => x"38",
         13042 => x"7a",
         13043 => x"7a",
         13044 => x"06",
         13045 => x"81",
         13046 => x"b8",
         13047 => x"16",
         13048 => x"dc",
         13049 => x"ba",
         13050 => x"2e",
         13051 => x"57",
         13052 => x"b4",
         13053 => x"57",
         13054 => x"7c",
         13055 => x"58",
         13056 => x"74",
         13057 => x"38",
         13058 => x"74",
         13059 => x"38",
         13060 => x"18",
         13061 => x"11",
         13062 => x"33",
         13063 => x"71",
         13064 => x"81",
         13065 => x"72",
         13066 => x"75",
         13067 => x"62",
         13068 => x"5e",
         13069 => x"76",
         13070 => x"0c",
         13071 => x"04",
         13072 => x"40",
         13073 => x"3d",
         13074 => x"fe",
         13075 => x"84",
         13076 => x"57",
         13077 => x"08",
         13078 => x"8d",
         13079 => x"2e",
         13080 => x"fe",
         13081 => x"7b",
         13082 => x"fe",
         13083 => x"54",
         13084 => x"53",
         13085 => x"53",
         13086 => x"52",
         13087 => x"ad",
         13088 => x"84",
         13089 => x"7a",
         13090 => x"06",
         13091 => x"84",
         13092 => x"83",
         13093 => x"16",
         13094 => x"08",
         13095 => x"8c",
         13096 => x"74",
         13097 => x"27",
         13098 => x"82",
         13099 => x"74",
         13100 => x"81",
         13101 => x"38",
         13102 => x"16",
         13103 => x"08",
         13104 => x"52",
         13105 => x"51",
         13106 => x"3f",
         13107 => x"54",
         13108 => x"16",
         13109 => x"33",
         13110 => x"d2",
         13111 => x"8c",
         13112 => x"fe",
         13113 => x"86",
         13114 => x"74",
         13115 => x"bb",
         13116 => x"8c",
         13117 => x"ba",
         13118 => x"e1",
         13119 => x"8c",
         13120 => x"8c",
         13121 => x"59",
         13122 => x"81",
         13123 => x"57",
         13124 => x"33",
         13125 => x"19",
         13126 => x"27",
         13127 => x"70",
         13128 => x"80",
         13129 => x"80",
         13130 => x"38",
         13131 => x"11",
         13132 => x"57",
         13133 => x"2e",
         13134 => x"e1",
         13135 => x"fd",
         13136 => x"3d",
         13137 => x"a1",
         13138 => x"05",
         13139 => x"51",
         13140 => x"3f",
         13141 => x"08",
         13142 => x"8c",
         13143 => x"38",
         13144 => x"8b",
         13145 => x"a0",
         13146 => x"05",
         13147 => x"15",
         13148 => x"38",
         13149 => x"08",
         13150 => x"81",
         13151 => x"58",
         13152 => x"78",
         13153 => x"38",
         13154 => x"3d",
         13155 => x"81",
         13156 => x"18",
         13157 => x"81",
         13158 => x"7c",
         13159 => x"ff",
         13160 => x"ff",
         13161 => x"a1",
         13162 => x"b5",
         13163 => x"8c",
         13164 => x"dc",
         13165 => x"8c",
         13166 => x"ff",
         13167 => x"80",
         13168 => x"38",
         13169 => x"0b",
         13170 => x"33",
         13171 => x"06",
         13172 => x"78",
         13173 => x"d6",
         13174 => x"78",
         13175 => x"38",
         13176 => x"33",
         13177 => x"06",
         13178 => x"74",
         13179 => x"38",
         13180 => x"09",
         13181 => x"38",
         13182 => x"06",
         13183 => x"a3",
         13184 => x"77",
         13185 => x"38",
         13186 => x"81",
         13187 => x"ff",
         13188 => x"38",
         13189 => x"55",
         13190 => x"81",
         13191 => x"81",
         13192 => x"7b",
         13193 => x"5d",
         13194 => x"a3",
         13195 => x"33",
         13196 => x"06",
         13197 => x"5a",
         13198 => x"fe",
         13199 => x"3d",
         13200 => x"56",
         13201 => x"2e",
         13202 => x"80",
         13203 => x"02",
         13204 => x"79",
         13205 => x"5c",
         13206 => x"2e",
         13207 => x"87",
         13208 => x"5a",
         13209 => x"7d",
         13210 => x"80",
         13211 => x"70",
         13212 => x"ef",
         13213 => x"ba",
         13214 => x"84",
         13215 => x"80",
         13216 => x"74",
         13217 => x"ba",
         13218 => x"3d",
         13219 => x"b5",
         13220 => x"9e",
         13221 => x"ba",
         13222 => x"ff",
         13223 => x"74",
         13224 => x"86",
         13225 => x"ba",
         13226 => x"3d",
         13227 => x"e7",
         13228 => x"fe",
         13229 => x"52",
         13230 => x"f4",
         13231 => x"ba",
         13232 => x"84",
         13233 => x"80",
         13234 => x"80",
         13235 => x"38",
         13236 => x"59",
         13237 => x"70",
         13238 => x"33",
         13239 => x"05",
         13240 => x"15",
         13241 => x"38",
         13242 => x"0b",
         13243 => x"7d",
         13244 => x"ec",
         13245 => x"8c",
         13246 => x"56",
         13247 => x"8a",
         13248 => x"8a",
         13249 => x"ff",
         13250 => x"ba",
         13251 => x"2e",
         13252 => x"fe",
         13253 => x"55",
         13254 => x"fe",
         13255 => x"08",
         13256 => x"52",
         13257 => x"b1",
         13258 => x"8c",
         13259 => x"ba",
         13260 => x"2e",
         13261 => x"81",
         13262 => x"ba",
         13263 => x"19",
         13264 => x"16",
         13265 => x"59",
         13266 => x"77",
         13267 => x"83",
         13268 => x"74",
         13269 => x"81",
         13270 => x"38",
         13271 => x"53",
         13272 => x"81",
         13273 => x"fe",
         13274 => x"84",
         13275 => x"80",
         13276 => x"ff",
         13277 => x"76",
         13278 => x"78",
         13279 => x"38",
         13280 => x"08",
         13281 => x"5a",
         13282 => x"e5",
         13283 => x"38",
         13284 => x"80",
         13285 => x"56",
         13286 => x"2e",
         13287 => x"81",
         13288 => x"81",
         13289 => x"81",
         13290 => x"fe",
         13291 => x"84",
         13292 => x"57",
         13293 => x"08",
         13294 => x"86",
         13295 => x"76",
         13296 => x"bf",
         13297 => x"76",
         13298 => x"a0",
         13299 => x"80",
         13300 => x"05",
         13301 => x"15",
         13302 => x"38",
         13303 => x"0b",
         13304 => x"8b",
         13305 => x"57",
         13306 => x"81",
         13307 => x"76",
         13308 => x"58",
         13309 => x"55",
         13310 => x"fd",
         13311 => x"70",
         13312 => x"33",
         13313 => x"05",
         13314 => x"15",
         13315 => x"38",
         13316 => x"6b",
         13317 => x"34",
         13318 => x"0b",
         13319 => x"7d",
         13320 => x"bc",
         13321 => x"8c",
         13322 => x"ce",
         13323 => x"fe",
         13324 => x"54",
         13325 => x"53",
         13326 => x"18",
         13327 => x"d4",
         13328 => x"ba",
         13329 => x"2e",
         13330 => x"80",
         13331 => x"ba",
         13332 => x"19",
         13333 => x"08",
         13334 => x"31",
         13335 => x"19",
         13336 => x"38",
         13337 => x"55",
         13338 => x"b1",
         13339 => x"8c",
         13340 => x"e8",
         13341 => x"81",
         13342 => x"fe",
         13343 => x"84",
         13344 => x"57",
         13345 => x"08",
         13346 => x"b6",
         13347 => x"39",
         13348 => x"59",
         13349 => x"fd",
         13350 => x"a1",
         13351 => x"b4",
         13352 => x"19",
         13353 => x"7a",
         13354 => x"33",
         13355 => x"fd",
         13356 => x"39",
         13357 => x"60",
         13358 => x"05",
         13359 => x"33",
         13360 => x"89",
         13361 => x"2e",
         13362 => x"08",
         13363 => x"2e",
         13364 => x"33",
         13365 => x"2e",
         13366 => x"15",
         13367 => x"22",
         13368 => x"78",
         13369 => x"38",
         13370 => x"5f",
         13371 => x"38",
         13372 => x"56",
         13373 => x"38",
         13374 => x"81",
         13375 => x"17",
         13376 => x"38",
         13377 => x"70",
         13378 => x"06",
         13379 => x"80",
         13380 => x"38",
         13381 => x"22",
         13382 => x"70",
         13383 => x"57",
         13384 => x"87",
         13385 => x"15",
         13386 => x"30",
         13387 => x"9f",
         13388 => x"8c",
         13389 => x"1c",
         13390 => x"53",
         13391 => x"81",
         13392 => x"38",
         13393 => x"78",
         13394 => x"82",
         13395 => x"56",
         13396 => x"74",
         13397 => x"fe",
         13398 => x"81",
         13399 => x"55",
         13400 => x"75",
         13401 => x"82",
         13402 => x"8c",
         13403 => x"81",
         13404 => x"ba",
         13405 => x"2e",
         13406 => x"84",
         13407 => x"81",
         13408 => x"19",
         13409 => x"2e",
         13410 => x"78",
         13411 => x"06",
         13412 => x"56",
         13413 => x"84",
         13414 => x"90",
         13415 => x"87",
         13416 => x"8c",
         13417 => x"0d",
         13418 => x"33",
         13419 => x"ac",
         13420 => x"8c",
         13421 => x"54",
         13422 => x"38",
         13423 => x"55",
         13424 => x"39",
         13425 => x"81",
         13426 => x"7d",
         13427 => x"80",
         13428 => x"81",
         13429 => x"81",
         13430 => x"38",
         13431 => x"52",
         13432 => x"dd",
         13433 => x"ba",
         13434 => x"84",
         13435 => x"ff",
         13436 => x"81",
         13437 => x"57",
         13438 => x"d7",
         13439 => x"90",
         13440 => x"7b",
         13441 => x"8c",
         13442 => x"18",
         13443 => x"18",
         13444 => x"33",
         13445 => x"5c",
         13446 => x"34",
         13447 => x"fe",
         13448 => x"08",
         13449 => x"7a",
         13450 => x"38",
         13451 => x"94",
         13452 => x"15",
         13453 => x"5d",
         13454 => x"34",
         13455 => x"d6",
         13456 => x"ff",
         13457 => x"5b",
         13458 => x"be",
         13459 => x"fe",
         13460 => x"54",
         13461 => x"ff",
         13462 => x"a1",
         13463 => x"98",
         13464 => x"0d",
         13465 => x"a5",
         13466 => x"88",
         13467 => x"05",
         13468 => x"5f",
         13469 => x"3d",
         13470 => x"5b",
         13471 => x"2e",
         13472 => x"79",
         13473 => x"5b",
         13474 => x"26",
         13475 => x"ba",
         13476 => x"38",
         13477 => x"75",
         13478 => x"92",
         13479 => x"e8",
         13480 => x"76",
         13481 => x"38",
         13482 => x"84",
         13483 => x"70",
         13484 => x"74",
         13485 => x"38",
         13486 => x"75",
         13487 => x"80",
         13488 => x"ba",
         13489 => x"40",
         13490 => x"52",
         13491 => x"ce",
         13492 => x"ba",
         13493 => x"ff",
         13494 => x"06",
         13495 => x"57",
         13496 => x"38",
         13497 => x"81",
         13498 => x"57",
         13499 => x"38",
         13500 => x"05",
         13501 => x"79",
         13502 => x"b0",
         13503 => x"8c",
         13504 => x"38",
         13505 => x"80",
         13506 => x"38",
         13507 => x"80",
         13508 => x"38",
         13509 => x"06",
         13510 => x"ff",
         13511 => x"2e",
         13512 => x"80",
         13513 => x"f8",
         13514 => x"80",
         13515 => x"f0",
         13516 => x"7f",
         13517 => x"83",
         13518 => x"89",
         13519 => x"08",
         13520 => x"89",
         13521 => x"4c",
         13522 => x"80",
         13523 => x"38",
         13524 => x"80",
         13525 => x"56",
         13526 => x"74",
         13527 => x"7d",
         13528 => x"df",
         13529 => x"74",
         13530 => x"79",
         13531 => x"be",
         13532 => x"84",
         13533 => x"83",
         13534 => x"83",
         13535 => x"61",
         13536 => x"33",
         13537 => x"07",
         13538 => x"57",
         13539 => x"d5",
         13540 => x"06",
         13541 => x"7d",
         13542 => x"05",
         13543 => x"33",
         13544 => x"80",
         13545 => x"38",
         13546 => x"83",
         13547 => x"12",
         13548 => x"2b",
         13549 => x"07",
         13550 => x"70",
         13551 => x"2b",
         13552 => x"07",
         13553 => x"83",
         13554 => x"12",
         13555 => x"2b",
         13556 => x"07",
         13557 => x"70",
         13558 => x"2b",
         13559 => x"07",
         13560 => x"0c",
         13561 => x"0c",
         13562 => x"44",
         13563 => x"59",
         13564 => x"4b",
         13565 => x"57",
         13566 => x"27",
         13567 => x"93",
         13568 => x"80",
         13569 => x"38",
         13570 => x"70",
         13571 => x"49",
         13572 => x"83",
         13573 => x"87",
         13574 => x"82",
         13575 => x"61",
         13576 => x"66",
         13577 => x"83",
         13578 => x"4a",
         13579 => x"58",
         13580 => x"8a",
         13581 => x"ae",
         13582 => x"2a",
         13583 => x"83",
         13584 => x"56",
         13585 => x"2e",
         13586 => x"77",
         13587 => x"83",
         13588 => x"77",
         13589 => x"70",
         13590 => x"58",
         13591 => x"86",
         13592 => x"27",
         13593 => x"52",
         13594 => x"80",
         13595 => x"ba",
         13596 => x"84",
         13597 => x"ba",
         13598 => x"f5",
         13599 => x"81",
         13600 => x"8c",
         13601 => x"ba",
         13602 => x"71",
         13603 => x"83",
         13604 => x"43",
         13605 => x"89",
         13606 => x"5c",
         13607 => x"1f",
         13608 => x"05",
         13609 => x"05",
         13610 => x"72",
         13611 => x"57",
         13612 => x"2e",
         13613 => x"74",
         13614 => x"90",
         13615 => x"60",
         13616 => x"74",
         13617 => x"f2",
         13618 => x"31",
         13619 => x"53",
         13620 => x"52",
         13621 => x"cf",
         13622 => x"8c",
         13623 => x"83",
         13624 => x"38",
         13625 => x"09",
         13626 => x"dd",
         13627 => x"f5",
         13628 => x"8c",
         13629 => x"ac",
         13630 => x"f9",
         13631 => x"55",
         13632 => x"26",
         13633 => x"74",
         13634 => x"39",
         13635 => x"84",
         13636 => x"9f",
         13637 => x"ba",
         13638 => x"81",
         13639 => x"39",
         13640 => x"ba",
         13641 => x"3d",
         13642 => x"98",
         13643 => x"33",
         13644 => x"81",
         13645 => x"57",
         13646 => x"26",
         13647 => x"1d",
         13648 => x"06",
         13649 => x"58",
         13650 => x"81",
         13651 => x"0b",
         13652 => x"5f",
         13653 => x"7d",
         13654 => x"70",
         13655 => x"33",
         13656 => x"05",
         13657 => x"9f",
         13658 => x"57",
         13659 => x"89",
         13660 => x"70",
         13661 => x"58",
         13662 => x"18",
         13663 => x"26",
         13664 => x"18",
         13665 => x"06",
         13666 => x"30",
         13667 => x"5a",
         13668 => x"2e",
         13669 => x"85",
         13670 => x"be",
         13671 => x"32",
         13672 => x"72",
         13673 => x"7b",
         13674 => x"4a",
         13675 => x"80",
         13676 => x"1c",
         13677 => x"5c",
         13678 => x"ff",
         13679 => x"56",
         13680 => x"9f",
         13681 => x"53",
         13682 => x"51",
         13683 => x"3f",
         13684 => x"ba",
         13685 => x"b6",
         13686 => x"2a",
         13687 => x"ba",
         13688 => x"56",
         13689 => x"bf",
         13690 => x"8e",
         13691 => x"26",
         13692 => x"74",
         13693 => x"fb",
         13694 => x"56",
         13695 => x"7b",
         13696 => x"ba",
         13697 => x"a3",
         13698 => x"f9",
         13699 => x"81",
         13700 => x"57",
         13701 => x"fd",
         13702 => x"6e",
         13703 => x"46",
         13704 => x"39",
         13705 => x"08",
         13706 => x"9d",
         13707 => x"38",
         13708 => x"81",
         13709 => x"fb",
         13710 => x"57",
         13711 => x"8c",
         13712 => x"0d",
         13713 => x"0c",
         13714 => x"62",
         13715 => x"99",
         13716 => x"60",
         13717 => x"74",
         13718 => x"8e",
         13719 => x"ae",
         13720 => x"61",
         13721 => x"76",
         13722 => x"58",
         13723 => x"55",
         13724 => x"8b",
         13725 => x"c8",
         13726 => x"76",
         13727 => x"58",
         13728 => x"81",
         13729 => x"ff",
         13730 => x"ef",
         13731 => x"05",
         13732 => x"34",
         13733 => x"05",
         13734 => x"8d",
         13735 => x"83",
         13736 => x"4b",
         13737 => x"05",
         13738 => x"2a",
         13739 => x"8f",
         13740 => x"61",
         13741 => x"62",
         13742 => x"30",
         13743 => x"61",
         13744 => x"78",
         13745 => x"06",
         13746 => x"92",
         13747 => x"56",
         13748 => x"ff",
         13749 => x"38",
         13750 => x"ff",
         13751 => x"61",
         13752 => x"74",
         13753 => x"6b",
         13754 => x"34",
         13755 => x"05",
         13756 => x"98",
         13757 => x"61",
         13758 => x"ff",
         13759 => x"34",
         13760 => x"05",
         13761 => x"9c",
         13762 => x"88",
         13763 => x"61",
         13764 => x"7e",
         13765 => x"6b",
         13766 => x"34",
         13767 => x"84",
         13768 => x"84",
         13769 => x"61",
         13770 => x"62",
         13771 => x"f7",
         13772 => x"a7",
         13773 => x"61",
         13774 => x"a1",
         13775 => x"34",
         13776 => x"aa",
         13777 => x"83",
         13778 => x"55",
         13779 => x"05",
         13780 => x"2a",
         13781 => x"97",
         13782 => x"80",
         13783 => x"34",
         13784 => x"05",
         13785 => x"ab",
         13786 => x"d4",
         13787 => x"76",
         13788 => x"58",
         13789 => x"81",
         13790 => x"ff",
         13791 => x"ef",
         13792 => x"fe",
         13793 => x"d5",
         13794 => x"83",
         13795 => x"ff",
         13796 => x"81",
         13797 => x"60",
         13798 => x"fe",
         13799 => x"81",
         13800 => x"8c",
         13801 => x"38",
         13802 => x"62",
         13803 => x"9c",
         13804 => x"57",
         13805 => x"70",
         13806 => x"34",
         13807 => x"74",
         13808 => x"75",
         13809 => x"83",
         13810 => x"38",
         13811 => x"f8",
         13812 => x"2e",
         13813 => x"57",
         13814 => x"76",
         13815 => x"45",
         13816 => x"70",
         13817 => x"34",
         13818 => x"59",
         13819 => x"81",
         13820 => x"76",
         13821 => x"75",
         13822 => x"57",
         13823 => x"66",
         13824 => x"76",
         13825 => x"7a",
         13826 => x"79",
         13827 => x"9d",
         13828 => x"8c",
         13829 => x"38",
         13830 => x"57",
         13831 => x"70",
         13832 => x"34",
         13833 => x"74",
         13834 => x"1b",
         13835 => x"58",
         13836 => x"38",
         13837 => x"40",
         13838 => x"ff",
         13839 => x"56",
         13840 => x"83",
         13841 => x"65",
         13842 => x"26",
         13843 => x"55",
         13844 => x"53",
         13845 => x"51",
         13846 => x"3f",
         13847 => x"08",
         13848 => x"74",
         13849 => x"31",
         13850 => x"db",
         13851 => x"62",
         13852 => x"38",
         13853 => x"83",
         13854 => x"8a",
         13855 => x"62",
         13856 => x"38",
         13857 => x"84",
         13858 => x"83",
         13859 => x"5e",
         13860 => x"38",
         13861 => x"56",
         13862 => x"70",
         13863 => x"34",
         13864 => x"78",
         13865 => x"d5",
         13866 => x"aa",
         13867 => x"83",
         13868 => x"78",
         13869 => x"67",
         13870 => x"81",
         13871 => x"34",
         13872 => x"05",
         13873 => x"84",
         13874 => x"43",
         13875 => x"52",
         13876 => x"fc",
         13877 => x"fe",
         13878 => x"34",
         13879 => x"08",
         13880 => x"07",
         13881 => x"86",
         13882 => x"ba",
         13883 => x"87",
         13884 => x"61",
         13885 => x"34",
         13886 => x"c7",
         13887 => x"61",
         13888 => x"34",
         13889 => x"08",
         13890 => x"05",
         13891 => x"83",
         13892 => x"62",
         13893 => x"64",
         13894 => x"05",
         13895 => x"2a",
         13896 => x"83",
         13897 => x"62",
         13898 => x"7e",
         13899 => x"05",
         13900 => x"78",
         13901 => x"79",
         13902 => x"f1",
         13903 => x"84",
         13904 => x"f7",
         13905 => x"53",
         13906 => x"51",
         13907 => x"3f",
         13908 => x"ba",
         13909 => x"b6",
         13910 => x"8c",
         13911 => x"8c",
         13912 => x"0d",
         13913 => x"0c",
         13914 => x"f9",
         13915 => x"1c",
         13916 => x"5c",
         13917 => x"7a",
         13918 => x"91",
         13919 => x"0b",
         13920 => x"22",
         13921 => x"80",
         13922 => x"74",
         13923 => x"38",
         13924 => x"56",
         13925 => x"17",
         13926 => x"57",
         13927 => x"2e",
         13928 => x"75",
         13929 => x"77",
         13930 => x"fc",
         13931 => x"84",
         13932 => x"10",
         13933 => x"05",
         13934 => x"5e",
         13935 => x"80",
         13936 => x"8c",
         13937 => x"8a",
         13938 => x"fd",
         13939 => x"77",
         13940 => x"38",
         13941 => x"e4",
         13942 => x"8c",
         13943 => x"f5",
         13944 => x"38",
         13945 => x"38",
         13946 => x"5b",
         13947 => x"38",
         13948 => x"c8",
         13949 => x"06",
         13950 => x"2e",
         13951 => x"83",
         13952 => x"39",
         13953 => x"05",
         13954 => x"2a",
         13955 => x"a1",
         13956 => x"90",
         13957 => x"61",
         13958 => x"75",
         13959 => x"76",
         13960 => x"34",
         13961 => x"80",
         13962 => x"05",
         13963 => x"80",
         13964 => x"a1",
         13965 => x"05",
         13966 => x"61",
         13967 => x"34",
         13968 => x"05",
         13969 => x"2a",
         13970 => x"a5",
         13971 => x"90",
         13972 => x"61",
         13973 => x"7c",
         13974 => x"75",
         13975 => x"34",
         13976 => x"05",
         13977 => x"ad",
         13978 => x"61",
         13979 => x"80",
         13980 => x"34",
         13981 => x"05",
         13982 => x"b1",
         13983 => x"61",
         13984 => x"80",
         13985 => x"34",
         13986 => x"80",
         13987 => x"a9",
         13988 => x"05",
         13989 => x"80",
         13990 => x"e5",
         13991 => x"55",
         13992 => x"05",
         13993 => x"70",
         13994 => x"34",
         13995 => x"74",
         13996 => x"cd",
         13997 => x"81",
         13998 => x"76",
         13999 => x"58",
         14000 => x"55",
         14001 => x"f9",
         14002 => x"54",
         14003 => x"52",
         14004 => x"be",
         14005 => x"57",
         14006 => x"08",
         14007 => x"7d",
         14008 => x"05",
         14009 => x"83",
         14010 => x"76",
         14011 => x"8c",
         14012 => x"52",
         14013 => x"bf",
         14014 => x"c3",
         14015 => x"84",
         14016 => x"9f",
         14017 => x"ba",
         14018 => x"f8",
         14019 => x"4a",
         14020 => x"81",
         14021 => x"ff",
         14022 => x"05",
         14023 => x"6a",
         14024 => x"84",
         14025 => x"61",
         14026 => x"ff",
         14027 => x"34",
         14028 => x"05",
         14029 => x"88",
         14030 => x"61",
         14031 => x"ff",
         14032 => x"34",
         14033 => x"7c",
         14034 => x"39",
         14035 => x"1f",
         14036 => x"79",
         14037 => x"d5",
         14038 => x"61",
         14039 => x"75",
         14040 => x"57",
         14041 => x"57",
         14042 => x"60",
         14043 => x"7c",
         14044 => x"5e",
         14045 => x"80",
         14046 => x"81",
         14047 => x"80",
         14048 => x"81",
         14049 => x"80",
         14050 => x"80",
         14051 => x"e4",
         14052 => x"f2",
         14053 => x"05",
         14054 => x"61",
         14055 => x"34",
         14056 => x"83",
         14057 => x"7f",
         14058 => x"7a",
         14059 => x"05",
         14060 => x"2a",
         14061 => x"83",
         14062 => x"7a",
         14063 => x"75",
         14064 => x"05",
         14065 => x"2a",
         14066 => x"83",
         14067 => x"82",
         14068 => x"05",
         14069 => x"83",
         14070 => x"76",
         14071 => x"05",
         14072 => x"83",
         14073 => x"80",
         14074 => x"ff",
         14075 => x"81",
         14076 => x"53",
         14077 => x"51",
         14078 => x"3f",
         14079 => x"1f",
         14080 => x"79",
         14081 => x"a5",
         14082 => x"57",
         14083 => x"39",
         14084 => x"7e",
         14085 => x"80",
         14086 => x"05",
         14087 => x"76",
         14088 => x"38",
         14089 => x"8e",
         14090 => x"54",
         14091 => x"52",
         14092 => x"9a",
         14093 => x"81",
         14094 => x"06",
         14095 => x"3d",
         14096 => x"8d",
         14097 => x"74",
         14098 => x"05",
         14099 => x"17",
         14100 => x"2e",
         14101 => x"77",
         14102 => x"80",
         14103 => x"55",
         14104 => x"76",
         14105 => x"ba",
         14106 => x"3d",
         14107 => x"3d",
         14108 => x"84",
         14109 => x"33",
         14110 => x"8a",
         14111 => x"38",
         14112 => x"56",
         14113 => x"9e",
         14114 => x"08",
         14115 => x"05",
         14116 => x"75",
         14117 => x"55",
         14118 => x"8e",
         14119 => x"18",
         14120 => x"88",
         14121 => x"3d",
         14122 => x"3d",
         14123 => x"74",
         14124 => x"52",
         14125 => x"ff",
         14126 => x"74",
         14127 => x"30",
         14128 => x"9f",
         14129 => x"84",
         14130 => x"1c",
         14131 => x"5a",
         14132 => x"39",
         14133 => x"51",
         14134 => x"ff",
         14135 => x"3d",
         14136 => x"ff",
         14137 => x"3d",
         14138 => x"cc",
         14139 => x"80",
         14140 => x"05",
         14141 => x"15",
         14142 => x"38",
         14143 => x"77",
         14144 => x"2e",
         14145 => x"7c",
         14146 => x"24",
         14147 => x"7d",
         14148 => x"05",
         14149 => x"75",
         14150 => x"55",
         14151 => x"b8",
         14152 => x"18",
         14153 => x"88",
         14154 => x"55",
         14155 => x"9e",
         14156 => x"ff",
         14157 => x"75",
         14158 => x"52",
         14159 => x"ff",
         14160 => x"84",
         14161 => x"86",
         14162 => x"2e",
         14163 => x"0b",
         14164 => x"0c",
         14165 => x"04",
         14166 => x"b0",
         14167 => x"54",
         14168 => x"76",
         14169 => x"9d",
         14170 => x"7b",
         14171 => x"70",
         14172 => x"2a",
         14173 => x"5a",
         14174 => x"a5",
         14175 => x"76",
         14176 => x"3f",
         14177 => x"7d",
         14178 => x"0c",
         14179 => x"04",
         14180 => x"75",
         14181 => x"9a",
         14182 => x"53",
         14183 => x"80",
         14184 => x"38",
         14185 => x"ff",
         14186 => x"84",
         14187 => x"85",
         14188 => x"83",
         14189 => x"27",
         14190 => x"b5",
         14191 => x"06",
         14192 => x"80",
         14193 => x"83",
         14194 => x"51",
         14195 => x"9c",
         14196 => x"70",
         14197 => x"06",
         14198 => x"80",
         14199 => x"38",
         14200 => x"e7",
         14201 => x"22",
         14202 => x"39",
         14203 => x"70",
         14204 => x"84",
         14205 => x"53",
         14206 => x"04",
         14207 => x"02",
         14208 => x"02",
         14209 => x"05",
         14210 => x"80",
         14211 => x"ff",
         14212 => x"70",
         14213 => x"ba",
         14214 => x"3d",
         14215 => x"83",
         14216 => x"81",
         14217 => x"70",
         14218 => x"e9",
         14219 => x"83",
         14220 => x"70",
         14221 => x"8c",
         14222 => x"3d",
         14223 => x"3d",
         14224 => x"70",
         14225 => x"26",
         14226 => x"70",
         14227 => x"06",
         14228 => x"56",
         14229 => x"ff",
         14230 => x"38",
         14231 => x"05",
         14232 => x"71",
         14233 => x"25",
         14234 => x"07",
         14235 => x"53",
         14236 => x"71",
         14237 => x"53",
         14238 => x"88",
         14239 => x"81",
         14240 => x"14",
         14241 => x"76",
         14242 => x"71",
         14243 => x"10",
         14244 => x"82",
         14245 => x"54",
         14246 => x"80",
         14247 => x"26",
         14248 => x"52",
         14249 => x"cb",
         14250 => x"70",
         14251 => x"0c",
         14252 => x"04",
         14253 => x"55",
         14254 => x"71",
         14255 => x"38",
         14256 => x"83",
         14257 => x"54",
         14258 => x"c7",
         14259 => x"83",
         14260 => x"57",
         14261 => x"d3",
         14262 => x"16",
         14263 => x"ff",
         14264 => x"f1",
         14265 => x"70",
         14266 => x"06",
         14267 => x"39",
         14268 => x"83",
         14269 => x"57",
         14270 => x"d0",
         14271 => x"ff",
         14272 => x"51",
         14273 => x"16",
         14274 => x"ff",
         14275 => x"c5",
         14276 => x"70",
         14277 => x"06",
         14278 => x"b9",
         14279 => x"31",
         14280 => x"71",
         14281 => x"ff",
         14282 => x"52",
         14283 => x"39",
         14284 => x"10",
         14285 => x"22",
         14286 => x"ef",
         14287 => x"ff",
         14288 => x"00",
         14289 => x"ff",
         14290 => x"ff",
         14291 => x"00",
         14292 => x"00",
         14293 => x"00",
         14294 => x"00",
         14295 => x"00",
         14296 => x"00",
         14297 => x"00",
         14298 => x"00",
         14299 => x"00",
         14300 => x"00",
         14301 => x"00",
         14302 => x"00",
         14303 => x"00",
         14304 => x"00",
         14305 => x"00",
         14306 => x"00",
         14307 => x"00",
         14308 => x"00",
         14309 => x"00",
         14310 => x"00",
         14311 => x"00",
         14312 => x"00",
         14313 => x"00",
         14314 => x"00",
         14315 => x"00",
         14316 => x"00",
         14317 => x"00",
         14318 => x"00",
         14319 => x"00",
         14320 => x"00",
         14321 => x"00",
         14322 => x"00",
         14323 => x"00",
         14324 => x"00",
         14325 => x"00",
         14326 => x"00",
         14327 => x"00",
         14328 => x"00",
         14329 => x"00",
         14330 => x"00",
         14331 => x"00",
         14332 => x"00",
         14333 => x"00",
         14334 => x"00",
         14335 => x"00",
         14336 => x"00",
         14337 => x"00",
         14338 => x"00",
         14339 => x"00",
         14340 => x"00",
         14341 => x"00",
         14342 => x"00",
         14343 => x"00",
         14344 => x"00",
         14345 => x"00",
         14346 => x"00",
         14347 => x"00",
         14348 => x"00",
         14349 => x"00",
         14350 => x"00",
         14351 => x"00",
         14352 => x"00",
         14353 => x"00",
         14354 => x"00",
         14355 => x"00",
         14356 => x"00",
         14357 => x"00",
         14358 => x"00",
         14359 => x"00",
         14360 => x"00",
         14361 => x"00",
         14362 => x"00",
         14363 => x"00",
         14364 => x"00",
         14365 => x"00",
         14366 => x"00",
         14367 => x"00",
         14368 => x"00",
         14369 => x"00",
         14370 => x"00",
         14371 => x"00",
         14372 => x"00",
         14373 => x"00",
         14374 => x"00",
         14375 => x"00",
         14376 => x"00",
         14377 => x"00",
         14378 => x"00",
         14379 => x"00",
         14380 => x"00",
         14381 => x"00",
         14382 => x"00",
         14383 => x"00",
         14384 => x"00",
         14385 => x"00",
         14386 => x"00",
         14387 => x"00",
         14388 => x"00",
         14389 => x"00",
         14390 => x"00",
         14391 => x"00",
         14392 => x"00",
         14393 => x"00",
         14394 => x"00",
         14395 => x"00",
         14396 => x"00",
         14397 => x"00",
         14398 => x"00",
         14399 => x"00",
         14400 => x"00",
         14401 => x"00",
         14402 => x"00",
         14403 => x"00",
         14404 => x"00",
         14405 => x"00",
         14406 => x"00",
         14407 => x"00",
         14408 => x"00",
         14409 => x"00",
         14410 => x"00",
         14411 => x"00",
         14412 => x"00",
         14413 => x"00",
         14414 => x"00",
         14415 => x"00",
         14416 => x"00",
         14417 => x"00",
         14418 => x"00",
         14419 => x"00",
         14420 => x"00",
         14421 => x"00",
         14422 => x"00",
         14423 => x"00",
         14424 => x"00",
         14425 => x"00",
         14426 => x"00",
         14427 => x"00",
         14428 => x"00",
         14429 => x"00",
         14430 => x"00",
         14431 => x"00",
         14432 => x"00",
         14433 => x"00",
         14434 => x"00",
         14435 => x"00",
         14436 => x"00",
         14437 => x"00",
         14438 => x"00",
         14439 => x"00",
         14440 => x"00",
         14441 => x"00",
         14442 => x"00",
         14443 => x"00",
         14444 => x"00",
         14445 => x"00",
         14446 => x"00",
         14447 => x"00",
         14448 => x"00",
         14449 => x"00",
         14450 => x"00",
         14451 => x"00",
         14452 => x"00",
         14453 => x"00",
         14454 => x"00",
         14455 => x"00",
         14456 => x"00",
         14457 => x"00",
         14458 => x"00",
         14459 => x"00",
         14460 => x"00",
         14461 => x"00",
         14462 => x"00",
         14463 => x"00",
         14464 => x"00",
         14465 => x"00",
         14466 => x"00",
         14467 => x"00",
         14468 => x"00",
         14469 => x"00",
         14470 => x"00",
         14471 => x"00",
         14472 => x"00",
         14473 => x"00",
         14474 => x"00",
         14475 => x"00",
         14476 => x"00",
         14477 => x"00",
         14478 => x"00",
         14479 => x"00",
         14480 => x"00",
         14481 => x"00",
         14482 => x"00",
         14483 => x"00",
         14484 => x"00",
         14485 => x"00",
         14486 => x"00",
         14487 => x"00",
         14488 => x"00",
         14489 => x"00",
         14490 => x"00",
         14491 => x"00",
         14492 => x"00",
         14493 => x"00",
         14494 => x"00",
         14495 => x"00",
         14496 => x"00",
         14497 => x"00",
         14498 => x"00",
         14499 => x"00",
         14500 => x"00",
         14501 => x"00",
         14502 => x"00",
         14503 => x"00",
         14504 => x"00",
         14505 => x"00",
         14506 => x"00",
         14507 => x"00",
         14508 => x"00",
         14509 => x"00",
         14510 => x"00",
         14511 => x"00",
         14512 => x"00",
         14513 => x"00",
         14514 => x"00",
         14515 => x"00",
         14516 => x"00",
         14517 => x"00",
         14518 => x"00",
         14519 => x"00",
         14520 => x"00",
         14521 => x"00",
         14522 => x"00",
         14523 => x"00",
         14524 => x"00",
         14525 => x"00",
         14526 => x"00",
         14527 => x"00",
         14528 => x"00",
         14529 => x"00",
         14530 => x"00",
         14531 => x"00",
         14532 => x"00",
         14533 => x"00",
         14534 => x"00",
         14535 => x"00",
         14536 => x"00",
         14537 => x"00",
         14538 => x"00",
         14539 => x"00",
         14540 => x"00",
         14541 => x"00",
         14542 => x"00",
         14543 => x"00",
         14544 => x"00",
         14545 => x"00",
         14546 => x"00",
         14547 => x"00",
         14548 => x"00",
         14549 => x"00",
         14550 => x"00",
         14551 => x"00",
         14552 => x"00",
         14553 => x"00",
         14554 => x"00",
         14555 => x"00",
         14556 => x"00",
         14557 => x"00",
         14558 => x"00",
         14559 => x"00",
         14560 => x"00",
         14561 => x"00",
         14562 => x"00",
         14563 => x"00",
         14564 => x"00",
         14565 => x"00",
         14566 => x"00",
         14567 => x"00",
         14568 => x"00",
         14569 => x"00",
         14570 => x"00",
         14571 => x"00",
         14572 => x"00",
         14573 => x"00",
         14574 => x"00",
         14575 => x"00",
         14576 => x"00",
         14577 => x"00",
         14578 => x"00",
         14579 => x"00",
         14580 => x"00",
         14581 => x"00",
         14582 => x"00",
         14583 => x"00",
         14584 => x"00",
         14585 => x"00",
         14586 => x"00",
         14587 => x"00",
         14588 => x"00",
         14589 => x"00",
         14590 => x"00",
         14591 => x"00",
         14592 => x"00",
         14593 => x"00",
         14594 => x"00",
         14595 => x"00",
         14596 => x"00",
         14597 => x"00",
         14598 => x"00",
         14599 => x"00",
         14600 => x"00",
         14601 => x"00",
         14602 => x"00",
         14603 => x"00",
         14604 => x"00",
         14605 => x"00",
         14606 => x"00",
         14607 => x"00",
         14608 => x"00",
         14609 => x"00",
         14610 => x"00",
         14611 => x"00",
         14612 => x"00",
         14613 => x"00",
         14614 => x"00",
         14615 => x"00",
         14616 => x"00",
         14617 => x"00",
         14618 => x"00",
         14619 => x"00",
         14620 => x"00",
         14621 => x"00",
         14622 => x"00",
         14623 => x"00",
         14624 => x"00",
         14625 => x"00",
         14626 => x"00",
         14627 => x"00",
         14628 => x"00",
         14629 => x"00",
         14630 => x"00",
         14631 => x"00",
         14632 => x"00",
         14633 => x"00",
         14634 => x"00",
         14635 => x"00",
         14636 => x"00",
         14637 => x"00",
         14638 => x"00",
         14639 => x"00",
         14640 => x"00",
         14641 => x"00",
         14642 => x"00",
         14643 => x"00",
         14644 => x"00",
         14645 => x"00",
         14646 => x"00",
         14647 => x"00",
         14648 => x"00",
         14649 => x"00",
         14650 => x"00",
         14651 => x"00",
         14652 => x"00",
         14653 => x"00",
         14654 => x"00",
         14655 => x"00",
         14656 => x"00",
         14657 => x"00",
         14658 => x"00",
         14659 => x"00",
         14660 => x"00",
         14661 => x"00",
         14662 => x"00",
         14663 => x"00",
         14664 => x"00",
         14665 => x"00",
         14666 => x"00",
         14667 => x"00",
         14668 => x"00",
         14669 => x"00",
         14670 => x"00",
         14671 => x"00",
         14672 => x"00",
         14673 => x"00",
         14674 => x"00",
         14675 => x"00",
         14676 => x"00",
         14677 => x"00",
         14678 => x"00",
         14679 => x"00",
         14680 => x"00",
         14681 => x"00",
         14682 => x"00",
         14683 => x"00",
         14684 => x"00",
         14685 => x"00",
         14686 => x"00",
         14687 => x"00",
         14688 => x"00",
         14689 => x"00",
         14690 => x"00",
         14691 => x"00",
         14692 => x"00",
         14693 => x"00",
         14694 => x"00",
         14695 => x"00",
         14696 => x"00",
         14697 => x"00",
         14698 => x"00",
         14699 => x"00",
         14700 => x"00",
         14701 => x"00",
         14702 => x"00",
         14703 => x"00",
         14704 => x"00",
         14705 => x"00",
         14706 => x"00",
         14707 => x"00",
         14708 => x"00",
         14709 => x"00",
         14710 => x"00",
         14711 => x"00",
         14712 => x"00",
         14713 => x"00",
         14714 => x"00",
         14715 => x"00",
         14716 => x"00",
         14717 => x"00",
         14718 => x"00",
         14719 => x"00",
         14720 => x"00",
         14721 => x"00",
         14722 => x"00",
         14723 => x"00",
         14724 => x"00",
         14725 => x"00",
         14726 => x"00",
         14727 => x"00",
         14728 => x"00",
         14729 => x"00",
         14730 => x"00",
         14731 => x"00",
         14732 => x"00",
         14733 => x"00",
         14734 => x"00",
         14735 => x"00",
         14736 => x"00",
         14737 => x"00",
         14738 => x"00",
         14739 => x"00",
         14740 => x"00",
         14741 => x"00",
         14742 => x"00",
         14743 => x"00",
         14744 => x"00",
         14745 => x"00",
         14746 => x"00",
         14747 => x"00",
         14748 => x"00",
         14749 => x"00",
         14750 => x"00",
         14751 => x"00",
         14752 => x"00",
         14753 => x"00",
         14754 => x"00",
         14755 => x"00",
         14756 => x"00",
         14757 => x"00",
         14758 => x"00",
         14759 => x"00",
         14760 => x"00",
         14761 => x"00",
         14762 => x"00",
         14763 => x"00",
         14764 => x"69",
         14765 => x"00",
         14766 => x"69",
         14767 => x"6c",
         14768 => x"69",
         14769 => x"00",
         14770 => x"6c",
         14771 => x"00",
         14772 => x"65",
         14773 => x"00",
         14774 => x"63",
         14775 => x"72",
         14776 => x"63",
         14777 => x"00",
         14778 => x"64",
         14779 => x"00",
         14780 => x"64",
         14781 => x"00",
         14782 => x"65",
         14783 => x"65",
         14784 => x"65",
         14785 => x"69",
         14786 => x"69",
         14787 => x"66",
         14788 => x"66",
         14789 => x"61",
         14790 => x"00",
         14791 => x"6d",
         14792 => x"65",
         14793 => x"72",
         14794 => x"65",
         14795 => x"00",
         14796 => x"6e",
         14797 => x"00",
         14798 => x"65",
         14799 => x"00",
         14800 => x"6c",
         14801 => x"38",
         14802 => x"62",
         14803 => x"63",
         14804 => x"62",
         14805 => x"63",
         14806 => x"69",
         14807 => x"00",
         14808 => x"64",
         14809 => x"6e",
         14810 => x"77",
         14811 => x"72",
         14812 => x"2e",
         14813 => x"61",
         14814 => x"65",
         14815 => x"73",
         14816 => x"63",
         14817 => x"65",
         14818 => x"00",
         14819 => x"6f",
         14820 => x"61",
         14821 => x"6f",
         14822 => x"20",
         14823 => x"65",
         14824 => x"00",
         14825 => x"6e",
         14826 => x"66",
         14827 => x"65",
         14828 => x"6d",
         14829 => x"72",
         14830 => x"00",
         14831 => x"69",
         14832 => x"69",
         14833 => x"6f",
         14834 => x"64",
         14835 => x"69",
         14836 => x"75",
         14837 => x"6f",
         14838 => x"61",
         14839 => x"6e",
         14840 => x"6e",
         14841 => x"6c",
         14842 => x"00",
         14843 => x"6f",
         14844 => x"74",
         14845 => x"6f",
         14846 => x"64",
         14847 => x"6f",
         14848 => x"6d",
         14849 => x"69",
         14850 => x"20",
         14851 => x"65",
         14852 => x"74",
         14853 => x"66",
         14854 => x"64",
         14855 => x"20",
         14856 => x"6b",
         14857 => x"69",
         14858 => x"6e",
         14859 => x"65",
         14860 => x"6c",
         14861 => x"00",
         14862 => x"72",
         14863 => x"20",
         14864 => x"62",
         14865 => x"69",
         14866 => x"6e",
         14867 => x"69",
         14868 => x"00",
         14869 => x"44",
         14870 => x"20",
         14871 => x"74",
         14872 => x"72",
         14873 => x"63",
         14874 => x"2e",
         14875 => x"69",
         14876 => x"68",
         14877 => x"6c",
         14878 => x"6e",
         14879 => x"69",
         14880 => x"00",
         14881 => x"69",
         14882 => x"61",
         14883 => x"61",
         14884 => x"65",
         14885 => x"74",
         14886 => x"00",
         14887 => x"63",
         14888 => x"73",
         14889 => x"6e",
         14890 => x"2e",
         14891 => x"6e",
         14892 => x"69",
         14893 => x"69",
         14894 => x"61",
         14895 => x"00",
         14896 => x"6f",
         14897 => x"74",
         14898 => x"6f",
         14899 => x"2e",
         14900 => x"6f",
         14901 => x"6c",
         14902 => x"6f",
         14903 => x"2e",
         14904 => x"69",
         14905 => x"6e",
         14906 => x"72",
         14907 => x"79",
         14908 => x"6e",
         14909 => x"6e",
         14910 => x"65",
         14911 => x"72",
         14912 => x"69",
         14913 => x"45",
         14914 => x"72",
         14915 => x"75",
         14916 => x"73",
         14917 => x"00",
         14918 => x"25",
         14919 => x"62",
         14920 => x"73",
         14921 => x"20",
         14922 => x"25",
         14923 => x"62",
         14924 => x"73",
         14925 => x"63",
         14926 => x"00",
         14927 => x"65",
         14928 => x"00",
         14929 => x"30",
         14930 => x"00",
         14931 => x"20",
         14932 => x"30",
         14933 => x"00",
         14934 => x"7c",
         14935 => x"00",
         14936 => x"20",
         14937 => x"30",
         14938 => x"00",
         14939 => x"20",
         14940 => x"20",
         14941 => x"00",
         14942 => x"4f",
         14943 => x"2a",
         14944 => x"20",
         14945 => x"31",
         14946 => x"2f",
         14947 => x"30",
         14948 => x"31",
         14949 => x"00",
         14950 => x"5a",
         14951 => x"20",
         14952 => x"20",
         14953 => x"78",
         14954 => x"73",
         14955 => x"20",
         14956 => x"0a",
         14957 => x"50",
         14958 => x"6e",
         14959 => x"72",
         14960 => x"20",
         14961 => x"64",
         14962 => x"00",
         14963 => x"41",
         14964 => x"20",
         14965 => x"69",
         14966 => x"72",
         14967 => x"74",
         14968 => x"41",
         14969 => x"20",
         14970 => x"69",
         14971 => x"72",
         14972 => x"74",
         14973 => x"41",
         14974 => x"20",
         14975 => x"69",
         14976 => x"72",
         14977 => x"74",
         14978 => x"41",
         14979 => x"20",
         14980 => x"69",
         14981 => x"72",
         14982 => x"74",
         14983 => x"4f",
         14984 => x"20",
         14985 => x"69",
         14986 => x"72",
         14987 => x"74",
         14988 => x"4f",
         14989 => x"20",
         14990 => x"69",
         14991 => x"72",
         14992 => x"74",
         14993 => x"53",
         14994 => x"6e",
         14995 => x"72",
         14996 => x"00",
         14997 => x"69",
         14998 => x"20",
         14999 => x"65",
         15000 => x"70",
         15001 => x"65",
         15002 => x"6e",
         15003 => x"70",
         15004 => x"6d",
         15005 => x"2e",
         15006 => x"6e",
         15007 => x"69",
         15008 => x"74",
         15009 => x"72",
         15010 => x"00",
         15011 => x"75",
         15012 => x"78",
         15013 => x"62",
         15014 => x"00",
         15015 => x"4f",
         15016 => x"70",
         15017 => x"73",
         15018 => x"61",
         15019 => x"64",
         15020 => x"20",
         15021 => x"74",
         15022 => x"69",
         15023 => x"73",
         15024 => x"61",
         15025 => x"30",
         15026 => x"6c",
         15027 => x"65",
         15028 => x"69",
         15029 => x"61",
         15030 => x"6c",
         15031 => x"00",
         15032 => x"20",
         15033 => x"64",
         15034 => x"73",
         15035 => x"69",
         15036 => x"69",
         15037 => x"69",
         15038 => x"73",
         15039 => x"00",
         15040 => x"3a",
         15041 => x"61",
         15042 => x"6f",
         15043 => x"6e",
         15044 => x"00",
         15045 => x"50",
         15046 => x"69",
         15047 => x"64",
         15048 => x"73",
         15049 => x"2e",
         15050 => x"00",
         15051 => x"6f",
         15052 => x"72",
         15053 => x"6f",
         15054 => x"67",
         15055 => x"00",
         15056 => x"65",
         15057 => x"72",
         15058 => x"67",
         15059 => x"70",
         15060 => x"61",
         15061 => x"6e",
         15062 => x"00",
         15063 => x"61",
         15064 => x"6e",
         15065 => x"6f",
         15066 => x"40",
         15067 => x"38",
         15068 => x"2e",
         15069 => x"00",
         15070 => x"61",
         15071 => x"72",
         15072 => x"72",
         15073 => x"20",
         15074 => x"65",
         15075 => x"64",
         15076 => x"00",
         15077 => x"78",
         15078 => x"74",
         15079 => x"20",
         15080 => x"65",
         15081 => x"25",
         15082 => x"78",
         15083 => x"2e",
         15084 => x"30",
         15085 => x"20",
         15086 => x"6c",
         15087 => x"00",
         15088 => x"30",
         15089 => x"20",
         15090 => x"58",
         15091 => x"6f",
         15092 => x"72",
         15093 => x"2e",
         15094 => x"00",
         15095 => x"30",
         15096 => x"28",
         15097 => x"78",
         15098 => x"25",
         15099 => x"78",
         15100 => x"38",
         15101 => x"00",
         15102 => x"6f",
         15103 => x"6e",
         15104 => x"2e",
         15105 => x"30",
         15106 => x"20",
         15107 => x"58",
         15108 => x"6c",
         15109 => x"69",
         15110 => x"2e",
         15111 => x"00",
         15112 => x"75",
         15113 => x"4d",
         15114 => x"72",
         15115 => x"43",
         15116 => x"6c",
         15117 => x"2e",
         15118 => x"64",
         15119 => x"73",
         15120 => x"00",
         15121 => x"65",
         15122 => x"79",
         15123 => x"68",
         15124 => x"74",
         15125 => x"20",
         15126 => x"6e",
         15127 => x"70",
         15128 => x"65",
         15129 => x"63",
         15130 => x"61",
         15131 => x"00",
         15132 => x"3f",
         15133 => x"64",
         15134 => x"2f",
         15135 => x"25",
         15136 => x"64",
         15137 => x"2e",
         15138 => x"64",
         15139 => x"6f",
         15140 => x"6f",
         15141 => x"67",
         15142 => x"74",
         15143 => x"00",
         15144 => x"0a",
         15145 => x"69",
         15146 => x"20",
         15147 => x"6c",
         15148 => x"6e",
         15149 => x"3a",
         15150 => x"64",
         15151 => x"73",
         15152 => x"3a",
         15153 => x"20",
         15154 => x"50",
         15155 => x"65",
         15156 => x"20",
         15157 => x"74",
         15158 => x"41",
         15159 => x"65",
         15160 => x"3d",
         15161 => x"38",
         15162 => x"00",
         15163 => x"20",
         15164 => x"50",
         15165 => x"65",
         15166 => x"79",
         15167 => x"61",
         15168 => x"41",
         15169 => x"65",
         15170 => x"3d",
         15171 => x"38",
         15172 => x"00",
         15173 => x"20",
         15174 => x"74",
         15175 => x"20",
         15176 => x"72",
         15177 => x"64",
         15178 => x"73",
         15179 => x"20",
         15180 => x"3d",
         15181 => x"38",
         15182 => x"00",
         15183 => x"69",
         15184 => x"00",
         15185 => x"20",
         15186 => x"50",
         15187 => x"64",
         15188 => x"20",
         15189 => x"20",
         15190 => x"20",
         15191 => x"20",
         15192 => x"3d",
         15193 => x"34",
         15194 => x"00",
         15195 => x"20",
         15196 => x"79",
         15197 => x"6d",
         15198 => x"6f",
         15199 => x"46",
         15200 => x"20",
         15201 => x"20",
         15202 => x"3d",
         15203 => x"2e",
         15204 => x"64",
         15205 => x"0a",
         15206 => x"20",
         15207 => x"69",
         15208 => x"6f",
         15209 => x"53",
         15210 => x"4d",
         15211 => x"6f",
         15212 => x"46",
         15213 => x"3d",
         15214 => x"2e",
         15215 => x"64",
         15216 => x"0a",
         15217 => x"20",
         15218 => x"44",
         15219 => x"20",
         15220 => x"63",
         15221 => x"72",
         15222 => x"20",
         15223 => x"20",
         15224 => x"3d",
         15225 => x"2e",
         15226 => x"64",
         15227 => x"0a",
         15228 => x"20",
         15229 => x"50",
         15230 => x"20",
         15231 => x"53",
         15232 => x"20",
         15233 => x"4f",
         15234 => x"00",
         15235 => x"20",
         15236 => x"42",
         15237 => x"43",
         15238 => x"20",
         15239 => x"49",
         15240 => x"4f",
         15241 => x"42",
         15242 => x"00",
         15243 => x"20",
         15244 => x"4e",
         15245 => x"43",
         15246 => x"20",
         15247 => x"61",
         15248 => x"6c",
         15249 => x"30",
         15250 => x"2e",
         15251 => x"20",
         15252 => x"49",
         15253 => x"31",
         15254 => x"20",
         15255 => x"6d",
         15256 => x"20",
         15257 => x"30",
         15258 => x"2e",
         15259 => x"20",
         15260 => x"44",
         15261 => x"52",
         15262 => x"20",
         15263 => x"76",
         15264 => x"73",
         15265 => x"30",
         15266 => x"2e",
         15267 => x"20",
         15268 => x"41",
         15269 => x"20",
         15270 => x"20",
         15271 => x"38",
         15272 => x"30",
         15273 => x"2e",
         15274 => x"20",
         15275 => x"52",
         15276 => x"20",
         15277 => x"20",
         15278 => x"38",
         15279 => x"30",
         15280 => x"2e",
         15281 => x"20",
         15282 => x"4e",
         15283 => x"42",
         15284 => x"20",
         15285 => x"38",
         15286 => x"30",
         15287 => x"2e",
         15288 => x"20",
         15289 => x"44",
         15290 => x"20",
         15291 => x"20",
         15292 => x"38",
         15293 => x"30",
         15294 => x"2e",
         15295 => x"20",
         15296 => x"42",
         15297 => x"52",
         15298 => x"20",
         15299 => x"38",
         15300 => x"30",
         15301 => x"2e",
         15302 => x"28",
         15303 => x"6d",
         15304 => x"43",
         15305 => x"6e",
         15306 => x"29",
         15307 => x"6e",
         15308 => x"77",
         15309 => x"56",
         15310 => x"00",
         15311 => x"6d",
         15312 => x"00",
         15313 => x"65",
         15314 => x"6d",
         15315 => x"6c",
         15316 => x"00",
         15317 => x"56",
         15318 => x"00",
         15319 => x"00",
         15320 => x"00",
         15321 => x"00",
         15322 => x"00",
         15323 => x"00",
         15324 => x"00",
         15325 => x"00",
         15326 => x"00",
         15327 => x"00",
         15328 => x"00",
         15329 => x"00",
         15330 => x"00",
         15331 => x"00",
         15332 => x"00",
         15333 => x"00",
         15334 => x"00",
         15335 => x"00",
         15336 => x"00",
         15337 => x"00",
         15338 => x"00",
         15339 => x"00",
         15340 => x"00",
         15341 => x"00",
         15342 => x"00",
         15343 => x"00",
         15344 => x"00",
         15345 => x"00",
         15346 => x"00",
         15347 => x"00",
         15348 => x"00",
         15349 => x"00",
         15350 => x"00",
         15351 => x"00",
         15352 => x"00",
         15353 => x"00",
         15354 => x"00",
         15355 => x"00",
         15356 => x"00",
         15357 => x"00",
         15358 => x"00",
         15359 => x"00",
         15360 => x"00",
         15361 => x"00",
         15362 => x"00",
         15363 => x"00",
         15364 => x"00",
         15365 => x"00",
         15366 => x"00",
         15367 => x"00",
         15368 => x"00",
         15369 => x"00",
         15370 => x"00",
         15371 => x"00",
         15372 => x"00",
         15373 => x"00",
         15374 => x"00",
         15375 => x"00",
         15376 => x"00",
         15377 => x"00",
         15378 => x"00",
         15379 => x"00",
         15380 => x"00",
         15381 => x"00",
         15382 => x"00",
         15383 => x"00",
         15384 => x"5b",
         15385 => x"5b",
         15386 => x"5b",
         15387 => x"5b",
         15388 => x"5b",
         15389 => x"5b",
         15390 => x"5b",
         15391 => x"30",
         15392 => x"5b",
         15393 => x"5b",
         15394 => x"5b",
         15395 => x"00",
         15396 => x"00",
         15397 => x"00",
         15398 => x"00",
         15399 => x"00",
         15400 => x"00",
         15401 => x"00",
         15402 => x"00",
         15403 => x"00",
         15404 => x"00",
         15405 => x"00",
         15406 => x"61",
         15407 => x"74",
         15408 => x"65",
         15409 => x"72",
         15410 => x"65",
         15411 => x"73",
         15412 => x"79",
         15413 => x"6c",
         15414 => x"64",
         15415 => x"62",
         15416 => x"67",
         15417 => x"69",
         15418 => x"72",
         15419 => x"69",
         15420 => x"00",
         15421 => x"00",
         15422 => x"30",
         15423 => x"20",
         15424 => x"0a",
         15425 => x"61",
         15426 => x"64",
         15427 => x"20",
         15428 => x"65",
         15429 => x"68",
         15430 => x"69",
         15431 => x"72",
         15432 => x"69",
         15433 => x"74",
         15434 => x"4f",
         15435 => x"00",
         15436 => x"25",
         15437 => x"00",
         15438 => x"5b",
         15439 => x"00",
         15440 => x"5b",
         15441 => x"5b",
         15442 => x"5b",
         15443 => x"5b",
         15444 => x"5b",
         15445 => x"00",
         15446 => x"5b",
         15447 => x"00",
         15448 => x"5b",
         15449 => x"00",
         15450 => x"5b",
         15451 => x"00",
         15452 => x"5b",
         15453 => x"00",
         15454 => x"5b",
         15455 => x"00",
         15456 => x"5b",
         15457 => x"00",
         15458 => x"5b",
         15459 => x"00",
         15460 => x"5b",
         15461 => x"00",
         15462 => x"5b",
         15463 => x"00",
         15464 => x"5b",
         15465 => x"00",
         15466 => x"5b",
         15467 => x"00",
         15468 => x"5b",
         15469 => x"5b",
         15470 => x"00",
         15471 => x"5b",
         15472 => x"00",
         15473 => x"3a",
         15474 => x"25",
         15475 => x"64",
         15476 => x"2c",
         15477 => x"25",
         15478 => x"30",
         15479 => x"00",
         15480 => x"3a",
         15481 => x"25",
         15482 => x"64",
         15483 => x"3a",
         15484 => x"25",
         15485 => x"64",
         15486 => x"64",
         15487 => x"3a",
         15488 => x"00",
         15489 => x"30",
         15490 => x"00",
         15491 => x"63",
         15492 => x"3b",
         15493 => x"00",
         15494 => x"65",
         15495 => x"74",
         15496 => x"72",
         15497 => x"3a",
         15498 => x"70",
         15499 => x"32",
         15500 => x"30",
         15501 => x"00",
         15502 => x"77",
         15503 => x"32",
         15504 => x"30",
         15505 => x"00",
         15506 => x"64",
         15507 => x"32",
         15508 => x"00",
         15509 => x"61",
         15510 => x"78",
         15511 => x"20",
         15512 => x"49",
         15513 => x"00",
         15514 => x"61",
         15515 => x"78",
         15516 => x"20",
         15517 => x"52",
         15518 => x"00",
         15519 => x"61",
         15520 => x"78",
         15521 => x"20",
         15522 => x"57",
         15523 => x"65",
         15524 => x"6f",
         15525 => x"73",
         15526 => x"65",
         15527 => x"65",
         15528 => x"00",
         15529 => x"44",
         15530 => x"2a",
         15531 => x"3f",
         15532 => x"00",
         15533 => x"2c",
         15534 => x"5d",
         15535 => x"41",
         15536 => x"41",
         15537 => x"00",
         15538 => x"fe",
         15539 => x"44",
         15540 => x"2e",
         15541 => x"4f",
         15542 => x"4d",
         15543 => x"20",
         15544 => x"54",
         15545 => x"20",
         15546 => x"4f",
         15547 => x"4d",
         15548 => x"20",
         15549 => x"54",
         15550 => x"20",
         15551 => x"00",
         15552 => x"00",
         15553 => x"00",
         15554 => x"00",
         15555 => x"03",
         15556 => x"0e",
         15557 => x"16",
         15558 => x"00",
         15559 => x"9a",
         15560 => x"41",
         15561 => x"45",
         15562 => x"49",
         15563 => x"92",
         15564 => x"4f",
         15565 => x"99",
         15566 => x"9d",
         15567 => x"49",
         15568 => x"a5",
         15569 => x"a9",
         15570 => x"ad",
         15571 => x"b1",
         15572 => x"b5",
         15573 => x"b9",
         15574 => x"bd",
         15575 => x"c1",
         15576 => x"c5",
         15577 => x"c9",
         15578 => x"cd",
         15579 => x"d1",
         15580 => x"d5",
         15581 => x"d9",
         15582 => x"dd",
         15583 => x"e1",
         15584 => x"e5",
         15585 => x"e9",
         15586 => x"ed",
         15587 => x"f1",
         15588 => x"f5",
         15589 => x"f9",
         15590 => x"fd",
         15591 => x"2e",
         15592 => x"5b",
         15593 => x"22",
         15594 => x"3e",
         15595 => x"00",
         15596 => x"01",
         15597 => x"10",
         15598 => x"00",
         15599 => x"00",
         15600 => x"01",
         15601 => x"04",
         15602 => x"10",
         15603 => x"00",
         15604 => x"c7",
         15605 => x"e9",
         15606 => x"e4",
         15607 => x"e5",
         15608 => x"ea",
         15609 => x"e8",
         15610 => x"ee",
         15611 => x"c4",
         15612 => x"c9",
         15613 => x"c6",
         15614 => x"f6",
         15615 => x"fb",
         15616 => x"ff",
         15617 => x"dc",
         15618 => x"a3",
         15619 => x"a7",
         15620 => x"e1",
         15621 => x"f3",
         15622 => x"f1",
         15623 => x"aa",
         15624 => x"bf",
         15625 => x"ac",
         15626 => x"bc",
         15627 => x"ab",
         15628 => x"91",
         15629 => x"93",
         15630 => x"24",
         15631 => x"62",
         15632 => x"55",
         15633 => x"51",
         15634 => x"5d",
         15635 => x"5b",
         15636 => x"14",
         15637 => x"2c",
         15638 => x"00",
         15639 => x"5e",
         15640 => x"5a",
         15641 => x"69",
         15642 => x"60",
         15643 => x"6c",
         15644 => x"68",
         15645 => x"65",
         15646 => x"58",
         15647 => x"53",
         15648 => x"6a",
         15649 => x"0c",
         15650 => x"84",
         15651 => x"90",
         15652 => x"b1",
         15653 => x"93",
         15654 => x"a3",
         15655 => x"b5",
         15656 => x"a6",
         15657 => x"a9",
         15658 => x"1e",
         15659 => x"b5",
         15660 => x"61",
         15661 => x"65",
         15662 => x"20",
         15663 => x"f7",
         15664 => x"b0",
         15665 => x"b7",
         15666 => x"7f",
         15667 => x"a0",
         15668 => x"61",
         15669 => x"e0",
         15670 => x"f8",
         15671 => x"ff",
         15672 => x"78",
         15673 => x"30",
         15674 => x"06",
         15675 => x"10",
         15676 => x"2e",
         15677 => x"06",
         15678 => x"4d",
         15679 => x"81",
         15680 => x"82",
         15681 => x"84",
         15682 => x"87",
         15683 => x"89",
         15684 => x"8b",
         15685 => x"8d",
         15686 => x"8f",
         15687 => x"91",
         15688 => x"93",
         15689 => x"f6",
         15690 => x"97",
         15691 => x"98",
         15692 => x"9b",
         15693 => x"9d",
         15694 => x"9f",
         15695 => x"a0",
         15696 => x"a2",
         15697 => x"a4",
         15698 => x"a7",
         15699 => x"a9",
         15700 => x"ab",
         15701 => x"ac",
         15702 => x"af",
         15703 => x"b1",
         15704 => x"b3",
         15705 => x"b5",
         15706 => x"b7",
         15707 => x"b8",
         15708 => x"bb",
         15709 => x"bc",
         15710 => x"f7",
         15711 => x"c1",
         15712 => x"c3",
         15713 => x"c5",
         15714 => x"c7",
         15715 => x"c7",
         15716 => x"cb",
         15717 => x"cd",
         15718 => x"dd",
         15719 => x"8e",
         15720 => x"12",
         15721 => x"03",
         15722 => x"f4",
         15723 => x"f8",
         15724 => x"22",
         15725 => x"3a",
         15726 => x"65",
         15727 => x"3b",
         15728 => x"66",
         15729 => x"40",
         15730 => x"41",
         15731 => x"0a",
         15732 => x"40",
         15733 => x"86",
         15734 => x"89",
         15735 => x"58",
         15736 => x"5a",
         15737 => x"5c",
         15738 => x"5e",
         15739 => x"93",
         15740 => x"62",
         15741 => x"64",
         15742 => x"66",
         15743 => x"97",
         15744 => x"6a",
         15745 => x"6c",
         15746 => x"6e",
         15747 => x"70",
         15748 => x"9d",
         15749 => x"74",
         15750 => x"76",
         15751 => x"78",
         15752 => x"7a",
         15753 => x"7c",
         15754 => x"7e",
         15755 => x"a6",
         15756 => x"82",
         15757 => x"84",
         15758 => x"86",
         15759 => x"ae",
         15760 => x"b1",
         15761 => x"45",
         15762 => x"8e",
         15763 => x"90",
         15764 => x"b7",
         15765 => x"03",
         15766 => x"fe",
         15767 => x"ac",
         15768 => x"86",
         15769 => x"89",
         15770 => x"b1",
         15771 => x"c2",
         15772 => x"a3",
         15773 => x"c4",
         15774 => x"cc",
         15775 => x"8c",
         15776 => x"8f",
         15777 => x"18",
         15778 => x"0a",
         15779 => x"f3",
         15780 => x"f5",
         15781 => x"f7",
         15782 => x"f9",
         15783 => x"fa",
         15784 => x"20",
         15785 => x"10",
         15786 => x"22",
         15787 => x"36",
         15788 => x"0e",
         15789 => x"01",
         15790 => x"d0",
         15791 => x"61",
         15792 => x"00",
         15793 => x"7d",
         15794 => x"63",
         15795 => x"96",
         15796 => x"5a",
         15797 => x"08",
         15798 => x"06",
         15799 => x"08",
         15800 => x"08",
         15801 => x"06",
         15802 => x"07",
         15803 => x"52",
         15804 => x"54",
         15805 => x"56",
         15806 => x"60",
         15807 => x"70",
         15808 => x"ba",
         15809 => x"c8",
         15810 => x"ca",
         15811 => x"da",
         15812 => x"f8",
         15813 => x"ea",
         15814 => x"fa",
         15815 => x"80",
         15816 => x"90",
         15817 => x"a0",
         15818 => x"b0",
         15819 => x"b8",
         15820 => x"b2",
         15821 => x"cc",
         15822 => x"c3",
         15823 => x"02",
         15824 => x"02",
         15825 => x"01",
         15826 => x"f3",
         15827 => x"fc",
         15828 => x"01",
         15829 => x"70",
         15830 => x"84",
         15831 => x"83",
         15832 => x"1a",
         15833 => x"2f",
         15834 => x"02",
         15835 => x"06",
         15836 => x"02",
         15837 => x"64",
         15838 => x"26",
         15839 => x"1a",
         15840 => x"00",
         15841 => x"00",
         15842 => x"02",
         15843 => x"00",
         15844 => x"00",
         15845 => x"00",
         15846 => x"04",
         15847 => x"00",
         15848 => x"00",
         15849 => x"00",
         15850 => x"14",
         15851 => x"00",
         15852 => x"00",
         15853 => x"00",
         15854 => x"2b",
         15855 => x"00",
         15856 => x"00",
         15857 => x"00",
         15858 => x"30",
         15859 => x"00",
         15860 => x"00",
         15861 => x"00",
         15862 => x"3c",
         15863 => x"00",
         15864 => x"00",
         15865 => x"00",
         15866 => x"3d",
         15867 => x"00",
         15868 => x"00",
         15869 => x"00",
         15870 => x"3f",
         15871 => x"00",
         15872 => x"00",
         15873 => x"00",
         15874 => x"40",
         15875 => x"00",
         15876 => x"00",
         15877 => x"00",
         15878 => x"41",
         15879 => x"00",
         15880 => x"00",
         15881 => x"00",
         15882 => x"42",
         15883 => x"00",
         15884 => x"00",
         15885 => x"00",
         15886 => x"43",
         15887 => x"00",
         15888 => x"00",
         15889 => x"00",
         15890 => x"50",
         15891 => x"00",
         15892 => x"00",
         15893 => x"00",
         15894 => x"51",
         15895 => x"00",
         15896 => x"00",
         15897 => x"00",
         15898 => x"54",
         15899 => x"00",
         15900 => x"00",
         15901 => x"00",
         15902 => x"55",
         15903 => x"00",
         15904 => x"00",
         15905 => x"00",
         15906 => x"79",
         15907 => x"00",
         15908 => x"00",
         15909 => x"00",
         15910 => x"78",
         15911 => x"00",
         15912 => x"00",
         15913 => x"00",
         15914 => x"82",
         15915 => x"00",
         15916 => x"00",
         15917 => x"00",
         15918 => x"83",
         15919 => x"00",
         15920 => x"00",
         15921 => x"00",
         15922 => x"85",
         15923 => x"00",
         15924 => x"00",
         15925 => x"00",
         15926 => x"87",
         15927 => x"00",
         15928 => x"00",
         15929 => x"00",
         15930 => x"88",
         15931 => x"00",
         15932 => x"00",
         15933 => x"00",
         15934 => x"89",
         15935 => x"00",
         15936 => x"00",
         15937 => x"00",
         15938 => x"8c",
         15939 => x"00",
         15940 => x"00",
         15941 => x"00",
         15942 => x"8d",
         15943 => x"00",
         15944 => x"00",
         15945 => x"00",
         15946 => x"8e",
         15947 => x"00",
         15948 => x"00",
         15949 => x"00",
         15950 => x"8f",
         15951 => x"00",
         15952 => x"00",
         15953 => x"00",
         15954 => x"00",
         15955 => x"00",
         15956 => x"00",
         15957 => x"00",
         15958 => x"01",
         15959 => x"00",
         15960 => x"01",
         15961 => x"81",
         15962 => x"00",
         15963 => x"7f",
         15964 => x"00",
         15965 => x"00",
         15966 => x"00",
         15967 => x"00",
         15968 => x"f5",
         15969 => x"f5",
         15970 => x"f5",
         15971 => x"00",
         15972 => x"01",
         15973 => x"01",
         15974 => x"01",
         15975 => x"00",
         15976 => x"00",
         15977 => x"00",
         15978 => x"00",
         15979 => x"00",
         15980 => x"00",
         15981 => x"00",
         15982 => x"00",
         15983 => x"00",
         15984 => x"00",
         15985 => x"00",
         15986 => x"00",
         15987 => x"00",
         15988 => x"00",
         15989 => x"00",
         15990 => x"00",
         15991 => x"00",
         15992 => x"00",
         15993 => x"00",
         15994 => x"00",
         15995 => x"00",
         15996 => x"00",
         15997 => x"00",
         15998 => x"00",
         15999 => x"00",
         16000 => x"00",
         16001 => x"00",
         16002 => x"00",
         16003 => x"00",
         16004 => x"00",
         16005 => x"00",
         16006 => x"01",
         16007 => x"fc",
         16008 => x"3b",
         16009 => x"7a",
         16010 => x"f0",
         16011 => x"72",
         16012 => x"76",
         16013 => x"6a",
         16014 => x"6e",
         16015 => x"62",
         16016 => x"66",
         16017 => x"32",
         16018 => x"36",
         16019 => x"f3",
         16020 => x"39",
         16021 => x"7f",
         16022 => x"f2",
         16023 => x"f0",
         16024 => x"f0",
         16025 => x"81",
         16026 => x"f0",
         16027 => x"fc",
         16028 => x"3a",
         16029 => x"5a",
         16030 => x"f0",
         16031 => x"52",
         16032 => x"56",
         16033 => x"4a",
         16034 => x"4e",
         16035 => x"42",
         16036 => x"46",
         16037 => x"32",
         16038 => x"36",
         16039 => x"f3",
         16040 => x"39",
         16041 => x"7f",
         16042 => x"f2",
         16043 => x"f0",
         16044 => x"f0",
         16045 => x"81",
         16046 => x"f0",
         16047 => x"fc",
         16048 => x"2b",
         16049 => x"5a",
         16050 => x"f0",
         16051 => x"52",
         16052 => x"56",
         16053 => x"4a",
         16054 => x"4e",
         16055 => x"42",
         16056 => x"46",
         16057 => x"22",
         16058 => x"26",
         16059 => x"7e",
         16060 => x"29",
         16061 => x"e2",
         16062 => x"f8",
         16063 => x"f0",
         16064 => x"f0",
         16065 => x"86",
         16066 => x"f0",
         16067 => x"fe",
         16068 => x"f0",
         16069 => x"1a",
         16070 => x"f0",
         16071 => x"12",
         16072 => x"16",
         16073 => x"0a",
         16074 => x"0e",
         16075 => x"02",
         16076 => x"06",
         16077 => x"f0",
         16078 => x"f0",
         16079 => x"1e",
         16080 => x"1f",
         16081 => x"f0",
         16082 => x"f0",
         16083 => x"f0",
         16084 => x"f0",
         16085 => x"81",
         16086 => x"f0",
         16087 => x"f0",
         16088 => x"b5",
         16089 => x"77",
         16090 => x"f0",
         16091 => x"70",
         16092 => x"a6",
         16093 => x"5d",
         16094 => x"33",
         16095 => x"6e",
         16096 => x"43",
         16097 => x"36",
         16098 => x"1e",
         16099 => x"9f",
         16100 => x"a3",
         16101 => x"c5",
         16102 => x"c4",
         16103 => x"f0",
         16104 => x"f0",
         16105 => x"81",
         16106 => x"f0",
         16107 => x"00",
         16108 => x"00",
         16109 => x"00",
         16110 => x"00",
         16111 => x"00",
         16112 => x"00",
         16113 => x"00",
         16114 => x"00",
         16115 => x"00",
         16116 => x"00",
         16117 => x"00",
         16118 => x"00",
         16119 => x"00",
         16120 => x"00",
         16121 => x"00",
         16122 => x"00",
         16123 => x"00",
         16124 => x"00",
         16125 => x"00",
         16126 => x"00",
         16127 => x"00",
         16128 => x"00",
         16129 => x"00",
         16130 => x"00",
         16131 => x"00",
         16132 => x"01",
         16133 => x"00",
         16134 => x"00",
         16135 => x"00",
         16136 => x"00",
         16137 => x"00",
         16138 => x"00",
         16139 => x"00",
         16140 => x"00",
         16141 => x"00",
         16142 => x"00",
         16143 => x"00",
         16144 => x"00",
         16145 => x"00",
         16146 => x"00",
         16147 => x"00",
         16148 => x"00",
         16149 => x"00",
         16150 => x"00",
         16151 => x"00",
         16152 => x"00",
         16153 => x"00",
         16154 => x"00",
         16155 => x"00",
         16156 => x"00",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"00",
         16166 => x"00",
         16167 => x"00",
         16168 => x"00",
         16169 => x"00",
         16170 => x"00",
         16171 => x"00",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"00",
         18159 => x"00",
         18160 => x"00",
         18161 => x"00",
         18162 => x"00",
         18163 => x"00",
         18164 => x"00",
         18165 => x"00",
         18166 => x"00",
         18167 => x"00",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"00",
         18176 => x"00",
         18177 => x"00",
         18178 => x"e0",
         18179 => x"cf",
         18180 => x"f9",
         18181 => x"fd",
         18182 => x"c1",
         18183 => x"c5",
         18184 => x"e4",
         18185 => x"ee",
         18186 => x"61",
         18187 => x"65",
         18188 => x"69",
         18189 => x"2a",
         18190 => x"21",
         18191 => x"25",
         18192 => x"29",
         18193 => x"2b",
         18194 => x"01",
         18195 => x"05",
         18196 => x"09",
         18197 => x"0d",
         18198 => x"11",
         18199 => x"15",
         18200 => x"19",
         18201 => x"54",
         18202 => x"81",
         18203 => x"85",
         18204 => x"89",
         18205 => x"8d",
         18206 => x"91",
         18207 => x"95",
         18208 => x"99",
         18209 => x"40",
         18210 => x"00",
         18211 => x"00",
         18212 => x"00",
         18213 => x"00",
         18214 => x"00",
         18215 => x"00",
         18216 => x"00",
         18217 => x"00",
         18218 => x"00",
         18219 => x"00",
         18220 => x"00",
         18221 => x"00",
         18222 => x"00",
         18223 => x"00",
         18224 => x"00",
         18225 => x"00",
         18226 => x"00",
         18227 => x"00",
         18228 => x"00",
         18229 => x"00",
         18230 => x"00",
         18231 => x"00",
         18232 => x"00",
         18233 => x"00",
         18234 => x"00",
         18235 => x"00",
         18236 => x"00",
         18237 => x"00",
         18238 => x"00",
         18239 => x"00",
         18240 => x"02",
         18241 => x"04",
         18242 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"cd",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"bc",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"cc",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"ab",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"96",
           269 => x"0b",
           270 => x"0b",
           271 => x"b6",
           272 => x"0b",
           273 => x"0b",
           274 => x"d6",
           275 => x"0b",
           276 => x"0b",
           277 => x"f6",
           278 => x"0b",
           279 => x"0b",
           280 => x"96",
           281 => x"0b",
           282 => x"0b",
           283 => x"b6",
           284 => x"0b",
           285 => x"0b",
           286 => x"d7",
           287 => x"0b",
           288 => x"0b",
           289 => x"f9",
           290 => x"0b",
           291 => x"0b",
           292 => x"9b",
           293 => x"0b",
           294 => x"0b",
           295 => x"bd",
           296 => x"0b",
           297 => x"0b",
           298 => x"df",
           299 => x"0b",
           300 => x"0b",
           301 => x"81",
           302 => x"0b",
           303 => x"0b",
           304 => x"a3",
           305 => x"0b",
           306 => x"0b",
           307 => x"c5",
           308 => x"0b",
           309 => x"0b",
           310 => x"e7",
           311 => x"0b",
           312 => x"0b",
           313 => x"89",
           314 => x"0b",
           315 => x"0b",
           316 => x"ab",
           317 => x"0b",
           318 => x"0b",
           319 => x"cd",
           320 => x"0b",
           321 => x"0b",
           322 => x"ef",
           323 => x"0b",
           324 => x"0b",
           325 => x"91",
           326 => x"0b",
           327 => x"0b",
           328 => x"b3",
           329 => x"0b",
           330 => x"0b",
           331 => x"d5",
           332 => x"0b",
           333 => x"0b",
           334 => x"f7",
           335 => x"0b",
           336 => x"0b",
           337 => x"99",
           338 => x"0b",
           339 => x"0b",
           340 => x"bb",
           341 => x"0b",
           342 => x"0b",
           343 => x"dc",
           344 => x"0b",
           345 => x"0b",
           346 => x"fe",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"90",
           390 => x"98",
           391 => x"2d",
           392 => x"08",
           393 => x"90",
           394 => x"98",
           395 => x"2d",
           396 => x"08",
           397 => x"90",
           398 => x"98",
           399 => x"2d",
           400 => x"08",
           401 => x"90",
           402 => x"98",
           403 => x"2d",
           404 => x"08",
           405 => x"90",
           406 => x"98",
           407 => x"2d",
           408 => x"08",
           409 => x"90",
           410 => x"98",
           411 => x"2d",
           412 => x"08",
           413 => x"90",
           414 => x"98",
           415 => x"2d",
           416 => x"08",
           417 => x"90",
           418 => x"98",
           419 => x"2d",
           420 => x"08",
           421 => x"90",
           422 => x"98",
           423 => x"2d",
           424 => x"08",
           425 => x"90",
           426 => x"98",
           427 => x"2d",
           428 => x"08",
           429 => x"90",
           430 => x"98",
           431 => x"2d",
           432 => x"08",
           433 => x"90",
           434 => x"98",
           435 => x"db",
           436 => x"98",
           437 => x"80",
           438 => x"ba",
           439 => x"d5",
           440 => x"ba",
           441 => x"c0",
           442 => x"84",
           443 => x"80",
           444 => x"84",
           445 => x"80",
           446 => x"04",
           447 => x"0c",
           448 => x"2d",
           449 => x"08",
           450 => x"90",
           451 => x"98",
           452 => x"f7",
           453 => x"98",
           454 => x"80",
           455 => x"ba",
           456 => x"e3",
           457 => x"ba",
           458 => x"c0",
           459 => x"84",
           460 => x"82",
           461 => x"84",
           462 => x"80",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"90",
           468 => x"98",
           469 => x"e6",
           470 => x"98",
           471 => x"80",
           472 => x"ba",
           473 => x"fa",
           474 => x"ba",
           475 => x"c0",
           476 => x"84",
           477 => x"82",
           478 => x"84",
           479 => x"80",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"90",
           485 => x"98",
           486 => x"d4",
           487 => x"98",
           488 => x"80",
           489 => x"ba",
           490 => x"f4",
           491 => x"ba",
           492 => x"c0",
           493 => x"84",
           494 => x"83",
           495 => x"84",
           496 => x"80",
           497 => x"04",
           498 => x"0c",
           499 => x"2d",
           500 => x"08",
           501 => x"90",
           502 => x"98",
           503 => x"cf",
           504 => x"98",
           505 => x"80",
           506 => x"ba",
           507 => x"f6",
           508 => x"ba",
           509 => x"c0",
           510 => x"84",
           511 => x"83",
           512 => x"84",
           513 => x"80",
           514 => x"04",
           515 => x"0c",
           516 => x"2d",
           517 => x"08",
           518 => x"90",
           519 => x"98",
           520 => x"99",
           521 => x"98",
           522 => x"80",
           523 => x"ba",
           524 => x"e4",
           525 => x"ba",
           526 => x"c0",
           527 => x"84",
           528 => x"82",
           529 => x"84",
           530 => x"80",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"90",
           536 => x"98",
           537 => x"e3",
           538 => x"98",
           539 => x"80",
           540 => x"ba",
           541 => x"9a",
           542 => x"ba",
           543 => x"c0",
           544 => x"84",
           545 => x"83",
           546 => x"84",
           547 => x"80",
           548 => x"04",
           549 => x"0c",
           550 => x"2d",
           551 => x"08",
           552 => x"90",
           553 => x"98",
           554 => x"db",
           555 => x"98",
           556 => x"80",
           557 => x"ba",
           558 => x"b9",
           559 => x"ba",
           560 => x"c0",
           561 => x"84",
           562 => x"83",
           563 => x"84",
           564 => x"80",
           565 => x"04",
           566 => x"0c",
           567 => x"2d",
           568 => x"08",
           569 => x"90",
           570 => x"98",
           571 => x"ab",
           572 => x"98",
           573 => x"80",
           574 => x"ba",
           575 => x"f6",
           576 => x"ba",
           577 => x"c0",
           578 => x"84",
           579 => x"80",
           580 => x"84",
           581 => x"80",
           582 => x"04",
           583 => x"0c",
           584 => x"2d",
           585 => x"08",
           586 => x"90",
           587 => x"98",
           588 => x"94",
           589 => x"98",
           590 => x"80",
           591 => x"ba",
           592 => x"9a",
           593 => x"98",
           594 => x"80",
           595 => x"ba",
           596 => x"db",
           597 => x"ba",
           598 => x"c0",
           599 => x"84",
           600 => x"81",
           601 => x"84",
           602 => x"80",
           603 => x"04",
           604 => x"0c",
           605 => x"2d",
           606 => x"08",
           607 => x"90",
           608 => x"98",
           609 => x"da",
           610 => x"98",
           611 => x"80",
           612 => x"04",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"53",
           621 => x"00",
           622 => x"06",
           623 => x"09",
           624 => x"05",
           625 => x"2b",
           626 => x"06",
           627 => x"04",
           628 => x"72",
           629 => x"05",
           630 => x"05",
           631 => x"72",
           632 => x"53",
           633 => x"51",
           634 => x"04",
           635 => x"70",
           636 => x"27",
           637 => x"71",
           638 => x"53",
           639 => x"0b",
           640 => x"8c",
           641 => x"ce",
           642 => x"fc",
           643 => x"3d",
           644 => x"05",
           645 => x"53",
           646 => x"d5",
           647 => x"81",
           648 => x"3d",
           649 => x"3d",
           650 => x"7c",
           651 => x"81",
           652 => x"80",
           653 => x"56",
           654 => x"80",
           655 => x"2e",
           656 => x"80",
           657 => x"14",
           658 => x"32",
           659 => x"72",
           660 => x"51",
           661 => x"54",
           662 => x"b7",
           663 => x"2e",
           664 => x"51",
           665 => x"84",
           666 => x"53",
           667 => x"08",
           668 => x"38",
           669 => x"08",
           670 => x"05",
           671 => x"14",
           672 => x"70",
           673 => x"07",
           674 => x"54",
           675 => x"80",
           676 => x"80",
           677 => x"52",
           678 => x"8c",
           679 => x"0d",
           680 => x"84",
           681 => x"88",
           682 => x"f5",
           683 => x"54",
           684 => x"05",
           685 => x"73",
           686 => x"58",
           687 => x"05",
           688 => x"8d",
           689 => x"51",
           690 => x"19",
           691 => x"34",
           692 => x"04",
           693 => x"86",
           694 => x"53",
           695 => x"51",
           696 => x"3d",
           697 => x"3d",
           698 => x"65",
           699 => x"80",
           700 => x"0c",
           701 => x"70",
           702 => x"32",
           703 => x"55",
           704 => x"72",
           705 => x"81",
           706 => x"38",
           707 => x"76",
           708 => x"c5",
           709 => x"7b",
           710 => x"5c",
           711 => x"81",
           712 => x"17",
           713 => x"26",
           714 => x"76",
           715 => x"30",
           716 => x"51",
           717 => x"ae",
           718 => x"2e",
           719 => x"83",
           720 => x"32",
           721 => x"54",
           722 => x"9e",
           723 => x"80",
           724 => x"33",
           725 => x"bd",
           726 => x"08",
           727 => x"ba",
           728 => x"3d",
           729 => x"83",
           730 => x"10",
           731 => x"10",
           732 => x"2b",
           733 => x"19",
           734 => x"0a",
           735 => x"05",
           736 => x"52",
           737 => x"5f",
           738 => x"81",
           739 => x"81",
           740 => x"ff",
           741 => x"7c",
           742 => x"76",
           743 => x"ff",
           744 => x"a5",
           745 => x"06",
           746 => x"73",
           747 => x"5b",
           748 => x"58",
           749 => x"dd",
           750 => x"39",
           751 => x"51",
           752 => x"7b",
           753 => x"fe",
           754 => x"8d",
           755 => x"2a",
           756 => x"54",
           757 => x"38",
           758 => x"06",
           759 => x"95",
           760 => x"53",
           761 => x"26",
           762 => x"10",
           763 => x"cc",
           764 => x"08",
           765 => x"18",
           766 => x"d8",
           767 => x"38",
           768 => x"51",
           769 => x"80",
           770 => x"5b",
           771 => x"38",
           772 => x"80",
           773 => x"f6",
           774 => x"7f",
           775 => x"71",
           776 => x"ff",
           777 => x"58",
           778 => x"ba",
           779 => x"52",
           780 => x"9a",
           781 => x"8c",
           782 => x"06",
           783 => x"08",
           784 => x"56",
           785 => x"26",
           786 => x"ba",
           787 => x"05",
           788 => x"70",
           789 => x"34",
           790 => x"51",
           791 => x"84",
           792 => x"56",
           793 => x"08",
           794 => x"84",
           795 => x"98",
           796 => x"06",
           797 => x"80",
           798 => x"77",
           799 => x"29",
           800 => x"05",
           801 => x"59",
           802 => x"2a",
           803 => x"55",
           804 => x"2e",
           805 => x"84",
           806 => x"f8",
           807 => x"53",
           808 => x"8b",
           809 => x"80",
           810 => x"80",
           811 => x"72",
           812 => x"7a",
           813 => x"81",
           814 => x"72",
           815 => x"38",
           816 => x"70",
           817 => x"54",
           818 => x"24",
           819 => x"7a",
           820 => x"06",
           821 => x"71",
           822 => x"56",
           823 => x"06",
           824 => x"2e",
           825 => x"77",
           826 => x"2b",
           827 => x"7c",
           828 => x"56",
           829 => x"80",
           830 => x"38",
           831 => x"81",
           832 => x"85",
           833 => x"84",
           834 => x"54",
           835 => x"38",
           836 => x"81",
           837 => x"86",
           838 => x"81",
           839 => x"85",
           840 => x"88",
           841 => x"5f",
           842 => x"b2",
           843 => x"84",
           844 => x"fc",
           845 => x"70",
           846 => x"40",
           847 => x"25",
           848 => x"52",
           849 => x"a9",
           850 => x"84",
           851 => x"fc",
           852 => x"70",
           853 => x"40",
           854 => x"24",
           855 => x"81",
           856 => x"80",
           857 => x"78",
           858 => x"0a",
           859 => x"0a",
           860 => x"2c",
           861 => x"80",
           862 => x"38",
           863 => x"51",
           864 => x"78",
           865 => x"0a",
           866 => x"0a",
           867 => x"2c",
           868 => x"74",
           869 => x"38",
           870 => x"70",
           871 => x"55",
           872 => x"81",
           873 => x"80",
           874 => x"d8",
           875 => x"f3",
           876 => x"38",
           877 => x"2e",
           878 => x"7d",
           879 => x"2e",
           880 => x"52",
           881 => x"33",
           882 => x"a5",
           883 => x"ba",
           884 => x"81",
           885 => x"74",
           886 => x"7a",
           887 => x"a7",
           888 => x"84",
           889 => x"fc",
           890 => x"70",
           891 => x"40",
           892 => x"25",
           893 => x"7c",
           894 => x"86",
           895 => x"39",
           896 => x"5b",
           897 => x"7c",
           898 => x"76",
           899 => x"fa",
           900 => x"80",
           901 => x"80",
           902 => x"60",
           903 => x"71",
           904 => x"ff",
           905 => x"59",
           906 => x"fb",
           907 => x"60",
           908 => x"fe",
           909 => x"83",
           910 => x"98",
           911 => x"7c",
           912 => x"29",
           913 => x"05",
           914 => x"5e",
           915 => x"57",
           916 => x"87",
           917 => x"06",
           918 => x"fe",
           919 => x"78",
           920 => x"29",
           921 => x"05",
           922 => x"5a",
           923 => x"7f",
           924 => x"38",
           925 => x"51",
           926 => x"e2",
           927 => x"70",
           928 => x"06",
           929 => x"83",
           930 => x"fe",
           931 => x"52",
           932 => x"05",
           933 => x"85",
           934 => x"39",
           935 => x"83",
           936 => x"5b",
           937 => x"ff",
           938 => x"ab",
           939 => x"75",
           940 => x"57",
           941 => x"b9",
           942 => x"75",
           943 => x"81",
           944 => x"78",
           945 => x"29",
           946 => x"05",
           947 => x"5a",
           948 => x"e3",
           949 => x"70",
           950 => x"56",
           951 => x"c6",
           952 => x"39",
           953 => x"05",
           954 => x"53",
           955 => x"80",
           956 => x"df",
           957 => x"ff",
           958 => x"84",
           959 => x"fa",
           960 => x"84",
           961 => x"58",
           962 => x"89",
           963 => x"39",
           964 => x"5b",
           965 => x"58",
           966 => x"f9",
           967 => x"39",
           968 => x"05",
           969 => x"81",
           970 => x"41",
           971 => x"8a",
           972 => x"87",
           973 => x"ba",
           974 => x"ff",
           975 => x"71",
           976 => x"54",
           977 => x"2c",
           978 => x"39",
           979 => x"07",
           980 => x"5b",
           981 => x"38",
           982 => x"7f",
           983 => x"71",
           984 => x"06",
           985 => x"54",
           986 => x"38",
           987 => x"bb",
           988 => x"8c",
           989 => x"ff",
           990 => x"31",
           991 => x"5a",
           992 => x"81",
           993 => x"33",
           994 => x"f7",
           995 => x"c9",
           996 => x"84",
           997 => x"fc",
           998 => x"70",
           999 => x"54",
          1000 => x"25",
          1001 => x"7c",
          1002 => x"83",
          1003 => x"39",
          1004 => x"51",
          1005 => x"79",
          1006 => x"81",
          1007 => x"38",
          1008 => x"51",
          1009 => x"7a",
          1010 => x"06",
          1011 => x"2e",
          1012 => x"fa",
          1013 => x"98",
          1014 => x"31",
          1015 => x"90",
          1016 => x"80",
          1017 => x"51",
          1018 => x"90",
          1019 => x"39",
          1020 => x"51",
          1021 => x"7e",
          1022 => x"73",
          1023 => x"a2",
          1024 => x"39",
          1025 => x"98",
          1026 => x"e5",
          1027 => x"06",
          1028 => x"2e",
          1029 => x"fb",
          1030 => x"74",
          1031 => x"70",
          1032 => x"53",
          1033 => x"7c",
          1034 => x"82",
          1035 => x"39",
          1036 => x"51",
          1037 => x"ff",
          1038 => x"52",
          1039 => x"8b",
          1040 => x"8c",
          1041 => x"ff",
          1042 => x"31",
          1043 => x"5a",
          1044 => x"7a",
          1045 => x"30",
          1046 => x"bf",
          1047 => x"5b",
          1048 => x"fe",
          1049 => x"d5",
          1050 => x"75",
          1051 => x"f3",
          1052 => x"3d",
          1053 => x"3d",
          1054 => x"80",
          1055 => x"f0",
          1056 => x"33",
          1057 => x"81",
          1058 => x"06",
          1059 => x"55",
          1060 => x"72",
          1061 => x"81",
          1062 => x"38",
          1063 => x"05",
          1064 => x"72",
          1065 => x"38",
          1066 => x"08",
          1067 => x"90",
          1068 => x"72",
          1069 => x"8c",
          1070 => x"83",
          1071 => x"74",
          1072 => x"56",
          1073 => x"80",
          1074 => x"84",
          1075 => x"54",
          1076 => x"d5",
          1077 => x"84",
          1078 => x"52",
          1079 => x"14",
          1080 => x"2d",
          1081 => x"08",
          1082 => x"38",
          1083 => x"56",
          1084 => x"8c",
          1085 => x"0d",
          1086 => x"0d",
          1087 => x"54",
          1088 => x"16",
          1089 => x"2a",
          1090 => x"81",
          1091 => x"57",
          1092 => x"72",
          1093 => x"81",
          1094 => x"73",
          1095 => x"55",
          1096 => x"77",
          1097 => x"06",
          1098 => x"56",
          1099 => x"8c",
          1100 => x"0d",
          1101 => x"81",
          1102 => x"53",
          1103 => x"ea",
          1104 => x"72",
          1105 => x"08",
          1106 => x"84",
          1107 => x"80",
          1108 => x"ff",
          1109 => x"05",
          1110 => x"57",
          1111 => x"ca",
          1112 => x"0d",
          1113 => x"08",
          1114 => x"85",
          1115 => x"0d",
          1116 => x"0d",
          1117 => x"11",
          1118 => x"2a",
          1119 => x"06",
          1120 => x"57",
          1121 => x"ae",
          1122 => x"2a",
          1123 => x"73",
          1124 => x"38",
          1125 => x"53",
          1126 => x"08",
          1127 => x"74",
          1128 => x"76",
          1129 => x"81",
          1130 => x"8c",
          1131 => x"81",
          1132 => x"0c",
          1133 => x"84",
          1134 => x"88",
          1135 => x"74",
          1136 => x"ff",
          1137 => x"15",
          1138 => x"2d",
          1139 => x"ba",
          1140 => x"38",
          1141 => x"81",
          1142 => x"0c",
          1143 => x"39",
          1144 => x"77",
          1145 => x"70",
          1146 => x"70",
          1147 => x"06",
          1148 => x"56",
          1149 => x"b3",
          1150 => x"2a",
          1151 => x"71",
          1152 => x"82",
          1153 => x"52",
          1154 => x"80",
          1155 => x"08",
          1156 => x"53",
          1157 => x"80",
          1158 => x"13",
          1159 => x"16",
          1160 => x"8c",
          1161 => x"81",
          1162 => x"73",
          1163 => x"0c",
          1164 => x"04",
          1165 => x"06",
          1166 => x"17",
          1167 => x"08",
          1168 => x"17",
          1169 => x"33",
          1170 => x"0c",
          1171 => x"04",
          1172 => x"16",
          1173 => x"2d",
          1174 => x"08",
          1175 => x"8c",
          1176 => x"ff",
          1177 => x"16",
          1178 => x"07",
          1179 => x"ba",
          1180 => x"2e",
          1181 => x"a0",
          1182 => x"85",
          1183 => x"54",
          1184 => x"8c",
          1185 => x"0d",
          1186 => x"07",
          1187 => x"17",
          1188 => x"ec",
          1189 => x"0d",
          1190 => x"54",
          1191 => x"70",
          1192 => x"33",
          1193 => x"38",
          1194 => x"72",
          1195 => x"54",
          1196 => x"72",
          1197 => x"54",
          1198 => x"38",
          1199 => x"8c",
          1200 => x"0d",
          1201 => x"0d",
          1202 => x"7a",
          1203 => x"54",
          1204 => x"9d",
          1205 => x"27",
          1206 => x"80",
          1207 => x"71",
          1208 => x"53",
          1209 => x"81",
          1210 => x"ff",
          1211 => x"ef",
          1212 => x"ba",
          1213 => x"3d",
          1214 => x"12",
          1215 => x"27",
          1216 => x"14",
          1217 => x"ff",
          1218 => x"53",
          1219 => x"73",
          1220 => x"51",
          1221 => x"d9",
          1222 => x"ff",
          1223 => x"71",
          1224 => x"ff",
          1225 => x"df",
          1226 => x"fe",
          1227 => x"70",
          1228 => x"70",
          1229 => x"33",
          1230 => x"38",
          1231 => x"74",
          1232 => x"8c",
          1233 => x"3d",
          1234 => x"3d",
          1235 => x"71",
          1236 => x"72",
          1237 => x"54",
          1238 => x"72",
          1239 => x"54",
          1240 => x"38",
          1241 => x"8c",
          1242 => x"0d",
          1243 => x"0d",
          1244 => x"79",
          1245 => x"54",
          1246 => x"93",
          1247 => x"81",
          1248 => x"73",
          1249 => x"55",
          1250 => x"51",
          1251 => x"73",
          1252 => x"0c",
          1253 => x"04",
          1254 => x"76",
          1255 => x"56",
          1256 => x"2e",
          1257 => x"33",
          1258 => x"05",
          1259 => x"52",
          1260 => x"09",
          1261 => x"38",
          1262 => x"71",
          1263 => x"38",
          1264 => x"72",
          1265 => x"51",
          1266 => x"8c",
          1267 => x"0d",
          1268 => x"2e",
          1269 => x"33",
          1270 => x"72",
          1271 => x"38",
          1272 => x"52",
          1273 => x"80",
          1274 => x"72",
          1275 => x"ba",
          1276 => x"3d",
          1277 => x"84",
          1278 => x"86",
          1279 => x"fb",
          1280 => x"79",
          1281 => x"56",
          1282 => x"84",
          1283 => x"84",
          1284 => x"81",
          1285 => x"81",
          1286 => x"84",
          1287 => x"54",
          1288 => x"08",
          1289 => x"38",
          1290 => x"08",
          1291 => x"74",
          1292 => x"75",
          1293 => x"8c",
          1294 => x"b1",
          1295 => x"8c",
          1296 => x"84",
          1297 => x"87",
          1298 => x"fd",
          1299 => x"77",
          1300 => x"55",
          1301 => x"80",
          1302 => x"72",
          1303 => x"54",
          1304 => x"80",
          1305 => x"ff",
          1306 => x"ff",
          1307 => x"06",
          1308 => x"13",
          1309 => x"52",
          1310 => x"ba",
          1311 => x"3d",
          1312 => x"3d",
          1313 => x"79",
          1314 => x"54",
          1315 => x"2e",
          1316 => x"72",
          1317 => x"54",
          1318 => x"51",
          1319 => x"73",
          1320 => x"0c",
          1321 => x"04",
          1322 => x"78",
          1323 => x"a0",
          1324 => x"2e",
          1325 => x"51",
          1326 => x"84",
          1327 => x"52",
          1328 => x"73",
          1329 => x"38",
          1330 => x"e3",
          1331 => x"ba",
          1332 => x"53",
          1333 => x"9f",
          1334 => x"38",
          1335 => x"9f",
          1336 => x"38",
          1337 => x"71",
          1338 => x"31",
          1339 => x"57",
          1340 => x"80",
          1341 => x"2e",
          1342 => x"10",
          1343 => x"07",
          1344 => x"07",
          1345 => x"ff",
          1346 => x"70",
          1347 => x"72",
          1348 => x"31",
          1349 => x"56",
          1350 => x"58",
          1351 => x"da",
          1352 => x"76",
          1353 => x"84",
          1354 => x"88",
          1355 => x"fc",
          1356 => x"70",
          1357 => x"06",
          1358 => x"72",
          1359 => x"70",
          1360 => x"71",
          1361 => x"2a",
          1362 => x"80",
          1363 => x"70",
          1364 => x"2b",
          1365 => x"74",
          1366 => x"81",
          1367 => x"30",
          1368 => x"82",
          1369 => x"31",
          1370 => x"55",
          1371 => x"05",
          1372 => x"70",
          1373 => x"25",
          1374 => x"31",
          1375 => x"70",
          1376 => x"32",
          1377 => x"70",
          1378 => x"31",
          1379 => x"05",
          1380 => x"0c",
          1381 => x"55",
          1382 => x"5a",
          1383 => x"55",
          1384 => x"56",
          1385 => x"56",
          1386 => x"3d",
          1387 => x"3d",
          1388 => x"70",
          1389 => x"54",
          1390 => x"3f",
          1391 => x"08",
          1392 => x"71",
          1393 => x"8c",
          1394 => x"3d",
          1395 => x"3d",
          1396 => x"58",
          1397 => x"76",
          1398 => x"38",
          1399 => x"cf",
          1400 => x"8c",
          1401 => x"13",
          1402 => x"2e",
          1403 => x"51",
          1404 => x"72",
          1405 => x"08",
          1406 => x"53",
          1407 => x"80",
          1408 => x"53",
          1409 => x"be",
          1410 => x"74",
          1411 => x"72",
          1412 => x"2b",
          1413 => x"55",
          1414 => x"76",
          1415 => x"72",
          1416 => x"2a",
          1417 => x"77",
          1418 => x"31",
          1419 => x"2c",
          1420 => x"7b",
          1421 => x"71",
          1422 => x"5c",
          1423 => x"55",
          1424 => x"74",
          1425 => x"84",
          1426 => x"88",
          1427 => x"fa",
          1428 => x"9f",
          1429 => x"2c",
          1430 => x"7b",
          1431 => x"2c",
          1432 => x"73",
          1433 => x"31",
          1434 => x"31",
          1435 => x"59",
          1436 => x"b4",
          1437 => x"8c",
          1438 => x"75",
          1439 => x"8c",
          1440 => x"0d",
          1441 => x"0d",
          1442 => x"57",
          1443 => x"0c",
          1444 => x"33",
          1445 => x"73",
          1446 => x"81",
          1447 => x"81",
          1448 => x"0c",
          1449 => x"55",
          1450 => x"f3",
          1451 => x"2e",
          1452 => x"73",
          1453 => x"83",
          1454 => x"58",
          1455 => x"89",
          1456 => x"38",
          1457 => x"56",
          1458 => x"80",
          1459 => x"e0",
          1460 => x"38",
          1461 => x"81",
          1462 => x"53",
          1463 => x"81",
          1464 => x"53",
          1465 => x"8f",
          1466 => x"70",
          1467 => x"54",
          1468 => x"27",
          1469 => x"72",
          1470 => x"83",
          1471 => x"29",
          1472 => x"70",
          1473 => x"33",
          1474 => x"73",
          1475 => x"be",
          1476 => x"2e",
          1477 => x"30",
          1478 => x"0c",
          1479 => x"84",
          1480 => x"8b",
          1481 => x"81",
          1482 => x"79",
          1483 => x"56",
          1484 => x"b0",
          1485 => x"06",
          1486 => x"81",
          1487 => x"0c",
          1488 => x"55",
          1489 => x"2e",
          1490 => x"58",
          1491 => x"2e",
          1492 => x"56",
          1493 => x"c6",
          1494 => x"53",
          1495 => x"58",
          1496 => x"fe",
          1497 => x"84",
          1498 => x"8b",
          1499 => x"82",
          1500 => x"70",
          1501 => x"33",
          1502 => x"56",
          1503 => x"80",
          1504 => x"8c",
          1505 => x"0d",
          1506 => x"0d",
          1507 => x"57",
          1508 => x"0c",
          1509 => x"33",
          1510 => x"73",
          1511 => x"81",
          1512 => x"81",
          1513 => x"0c",
          1514 => x"55",
          1515 => x"f3",
          1516 => x"2e",
          1517 => x"73",
          1518 => x"83",
          1519 => x"58",
          1520 => x"89",
          1521 => x"38",
          1522 => x"56",
          1523 => x"80",
          1524 => x"e0",
          1525 => x"38",
          1526 => x"81",
          1527 => x"53",
          1528 => x"81",
          1529 => x"53",
          1530 => x"8f",
          1531 => x"70",
          1532 => x"54",
          1533 => x"27",
          1534 => x"72",
          1535 => x"83",
          1536 => x"29",
          1537 => x"70",
          1538 => x"33",
          1539 => x"73",
          1540 => x"be",
          1541 => x"2e",
          1542 => x"30",
          1543 => x"0c",
          1544 => x"84",
          1545 => x"8b",
          1546 => x"81",
          1547 => x"79",
          1548 => x"56",
          1549 => x"b0",
          1550 => x"06",
          1551 => x"81",
          1552 => x"0c",
          1553 => x"55",
          1554 => x"2e",
          1555 => x"58",
          1556 => x"2e",
          1557 => x"56",
          1558 => x"c6",
          1559 => x"53",
          1560 => x"58",
          1561 => x"fe",
          1562 => x"84",
          1563 => x"8b",
          1564 => x"82",
          1565 => x"70",
          1566 => x"33",
          1567 => x"56",
          1568 => x"80",
          1569 => x"8c",
          1570 => x"0d",
          1571 => x"dc",
          1572 => x"8c",
          1573 => x"06",
          1574 => x"0c",
          1575 => x"0d",
          1576 => x"93",
          1577 => x"71",
          1578 => x"be",
          1579 => x"71",
          1580 => x"ce",
          1581 => x"be",
          1582 => x"0d",
          1583 => x"f4",
          1584 => x"3f",
          1585 => x"04",
          1586 => x"51",
          1587 => x"83",
          1588 => x"83",
          1589 => x"ef",
          1590 => x"3d",
          1591 => x"cf",
          1592 => x"92",
          1593 => x"0d",
          1594 => x"cc",
          1595 => x"3f",
          1596 => x"04",
          1597 => x"51",
          1598 => x"83",
          1599 => x"83",
          1600 => x"ee",
          1601 => x"3d",
          1602 => x"d0",
          1603 => x"e6",
          1604 => x"0d",
          1605 => x"b8",
          1606 => x"3f",
          1607 => x"04",
          1608 => x"51",
          1609 => x"83",
          1610 => x"83",
          1611 => x"ee",
          1612 => x"3d",
          1613 => x"d1",
          1614 => x"ba",
          1615 => x"0d",
          1616 => x"9c",
          1617 => x"3f",
          1618 => x"04",
          1619 => x"51",
          1620 => x"83",
          1621 => x"83",
          1622 => x"ee",
          1623 => x"3d",
          1624 => x"d1",
          1625 => x"8e",
          1626 => x"0d",
          1627 => x"e0",
          1628 => x"3f",
          1629 => x"04",
          1630 => x"51",
          1631 => x"83",
          1632 => x"83",
          1633 => x"ed",
          1634 => x"3d",
          1635 => x"d2",
          1636 => x"e2",
          1637 => x"0d",
          1638 => x"0d",
          1639 => x"05",
          1640 => x"33",
          1641 => x"68",
          1642 => x"7b",
          1643 => x"51",
          1644 => x"78",
          1645 => x"ff",
          1646 => x"81",
          1647 => x"07",
          1648 => x"06",
          1649 => x"57",
          1650 => x"38",
          1651 => x"52",
          1652 => x"52",
          1653 => x"a2",
          1654 => x"8c",
          1655 => x"ba",
          1656 => x"2e",
          1657 => x"77",
          1658 => x"e0",
          1659 => x"70",
          1660 => x"25",
          1661 => x"9f",
          1662 => x"53",
          1663 => x"77",
          1664 => x"38",
          1665 => x"88",
          1666 => x"87",
          1667 => x"e0",
          1668 => x"78",
          1669 => x"51",
          1670 => x"84",
          1671 => x"54",
          1672 => x"53",
          1673 => x"d2",
          1674 => x"df",
          1675 => x"ba",
          1676 => x"3d",
          1677 => x"ba",
          1678 => x"c0",
          1679 => x"84",
          1680 => x"59",
          1681 => x"05",
          1682 => x"53",
          1683 => x"51",
          1684 => x"3f",
          1685 => x"08",
          1686 => x"8c",
          1687 => x"38",
          1688 => x"80",
          1689 => x"38",
          1690 => x"17",
          1691 => x"39",
          1692 => x"74",
          1693 => x"3f",
          1694 => x"08",
          1695 => x"f4",
          1696 => x"ba",
          1697 => x"83",
          1698 => x"78",
          1699 => x"98",
          1700 => x"3f",
          1701 => x"f8",
          1702 => x"02",
          1703 => x"05",
          1704 => x"ff",
          1705 => x"7b",
          1706 => x"fd",
          1707 => x"ba",
          1708 => x"38",
          1709 => x"91",
          1710 => x"2e",
          1711 => x"84",
          1712 => x"8a",
          1713 => x"78",
          1714 => x"ec",
          1715 => x"60",
          1716 => x"8c",
          1717 => x"7e",
          1718 => x"84",
          1719 => x"84",
          1720 => x"8a",
          1721 => x"f3",
          1722 => x"61",
          1723 => x"05",
          1724 => x"33",
          1725 => x"68",
          1726 => x"5c",
          1727 => x"78",
          1728 => x"82",
          1729 => x"83",
          1730 => x"dd",
          1731 => x"d2",
          1732 => x"f7",
          1733 => x"73",
          1734 => x"38",
          1735 => x"81",
          1736 => x"a0",
          1737 => x"38",
          1738 => x"72",
          1739 => x"a7",
          1740 => x"52",
          1741 => x"51",
          1742 => x"81",
          1743 => x"f0",
          1744 => x"a0",
          1745 => x"3f",
          1746 => x"dc",
          1747 => x"d8",
          1748 => x"3f",
          1749 => x"79",
          1750 => x"38",
          1751 => x"33",
          1752 => x"55",
          1753 => x"83",
          1754 => x"80",
          1755 => x"27",
          1756 => x"53",
          1757 => x"70",
          1758 => x"56",
          1759 => x"2e",
          1760 => x"fe",
          1761 => x"ee",
          1762 => x"f0",
          1763 => x"51",
          1764 => x"81",
          1765 => x"76",
          1766 => x"83",
          1767 => x"e9",
          1768 => x"18",
          1769 => x"58",
          1770 => x"b2",
          1771 => x"8c",
          1772 => x"70",
          1773 => x"54",
          1774 => x"81",
          1775 => x"9b",
          1776 => x"38",
          1777 => x"76",
          1778 => x"b9",
          1779 => x"84",
          1780 => x"8f",
          1781 => x"83",
          1782 => x"dc",
          1783 => x"14",
          1784 => x"08",
          1785 => x"51",
          1786 => x"78",
          1787 => x"b8",
          1788 => x"39",
          1789 => x"51",
          1790 => x"82",
          1791 => x"f0",
          1792 => x"a0",
          1793 => x"3f",
          1794 => x"fe",
          1795 => x"18",
          1796 => x"27",
          1797 => x"22",
          1798 => x"e4",
          1799 => x"3f",
          1800 => x"d5",
          1801 => x"54",
          1802 => x"c5",
          1803 => x"26",
          1804 => x"99",
          1805 => x"ec",
          1806 => x"3f",
          1807 => x"d5",
          1808 => x"54",
          1809 => x"a9",
          1810 => x"27",
          1811 => x"73",
          1812 => x"7a",
          1813 => x"72",
          1814 => x"d2",
          1815 => x"ab",
          1816 => x"84",
          1817 => x"53",
          1818 => x"ea",
          1819 => x"74",
          1820 => x"fd",
          1821 => x"d5",
          1822 => x"73",
          1823 => x"3f",
          1824 => x"fe",
          1825 => x"ce",
          1826 => x"ba",
          1827 => x"ff",
          1828 => x"59",
          1829 => x"fc",
          1830 => x"59",
          1831 => x"2e",
          1832 => x"fc",
          1833 => x"59",
          1834 => x"80",
          1835 => x"3f",
          1836 => x"08",
          1837 => x"98",
          1838 => x"32",
          1839 => x"9b",
          1840 => x"70",
          1841 => x"75",
          1842 => x"55",
          1843 => x"58",
          1844 => x"25",
          1845 => x"80",
          1846 => x"3f",
          1847 => x"08",
          1848 => x"98",
          1849 => x"32",
          1850 => x"9b",
          1851 => x"70",
          1852 => x"75",
          1853 => x"55",
          1854 => x"58",
          1855 => x"24",
          1856 => x"fd",
          1857 => x"0b",
          1858 => x"0c",
          1859 => x"04",
          1860 => x"87",
          1861 => x"08",
          1862 => x"3f",
          1863 => x"f7",
          1864 => x"b4",
          1865 => x"3f",
          1866 => x"eb",
          1867 => x"2a",
          1868 => x"51",
          1869 => x"b7",
          1870 => x"2a",
          1871 => x"51",
          1872 => x"89",
          1873 => x"2a",
          1874 => x"51",
          1875 => x"db",
          1876 => x"2a",
          1877 => x"51",
          1878 => x"ad",
          1879 => x"2a",
          1880 => x"51",
          1881 => x"ff",
          1882 => x"2a",
          1883 => x"51",
          1884 => x"d2",
          1885 => x"2a",
          1886 => x"51",
          1887 => x"38",
          1888 => x"81",
          1889 => x"88",
          1890 => x"3f",
          1891 => x"04",
          1892 => x"83",
          1893 => x"cc",
          1894 => x"3f",
          1895 => x"f7",
          1896 => x"3f",
          1897 => x"04",
          1898 => x"eb",
          1899 => x"e0",
          1900 => x"3f",
          1901 => x"df",
          1902 => x"2a",
          1903 => x"72",
          1904 => x"38",
          1905 => x"51",
          1906 => x"83",
          1907 => x"9b",
          1908 => x"51",
          1909 => x"72",
          1910 => x"81",
          1911 => x"71",
          1912 => x"9c",
          1913 => x"81",
          1914 => x"3f",
          1915 => x"51",
          1916 => x"80",
          1917 => x"3f",
          1918 => x"70",
          1919 => x"52",
          1920 => x"fe",
          1921 => x"be",
          1922 => x"9b",
          1923 => x"d4",
          1924 => x"9b",
          1925 => x"9a",
          1926 => x"85",
          1927 => x"06",
          1928 => x"80",
          1929 => x"38",
          1930 => x"81",
          1931 => x"3f",
          1932 => x"51",
          1933 => x"80",
          1934 => x"3f",
          1935 => x"70",
          1936 => x"52",
          1937 => x"fe",
          1938 => x"bd",
          1939 => x"9a",
          1940 => x"d4",
          1941 => x"d7",
          1942 => x"9a",
          1943 => x"83",
          1944 => x"06",
          1945 => x"80",
          1946 => x"38",
          1947 => x"81",
          1948 => x"3f",
          1949 => x"51",
          1950 => x"80",
          1951 => x"3f",
          1952 => x"70",
          1953 => x"52",
          1954 => x"fd",
          1955 => x"bd",
          1956 => x"0d",
          1957 => x"41",
          1958 => x"d1",
          1959 => x"81",
          1960 => x"81",
          1961 => x"84",
          1962 => x"81",
          1963 => x"3d",
          1964 => x"61",
          1965 => x"38",
          1966 => x"51",
          1967 => x"98",
          1968 => x"d5",
          1969 => x"c3",
          1970 => x"80",
          1971 => x"52",
          1972 => x"ae",
          1973 => x"83",
          1974 => x"70",
          1975 => x"5b",
          1976 => x"2e",
          1977 => x"79",
          1978 => x"88",
          1979 => x"ff",
          1980 => x"82",
          1981 => x"38",
          1982 => x"5a",
          1983 => x"83",
          1984 => x"33",
          1985 => x"2e",
          1986 => x"8c",
          1987 => x"70",
          1988 => x"7b",
          1989 => x"38",
          1990 => x"9b",
          1991 => x"7b",
          1992 => x"ef",
          1993 => x"08",
          1994 => x"ff",
          1995 => x"8c",
          1996 => x"8c",
          1997 => x"53",
          1998 => x"5d",
          1999 => x"84",
          2000 => x"8b",
          2001 => x"33",
          2002 => x"2e",
          2003 => x"81",
          2004 => x"ff",
          2005 => x"9b",
          2006 => x"38",
          2007 => x"5c",
          2008 => x"fe",
          2009 => x"f8",
          2010 => x"e9",
          2011 => x"ba",
          2012 => x"84",
          2013 => x"80",
          2014 => x"38",
          2015 => x"08",
          2016 => x"ff",
          2017 => x"91",
          2018 => x"ba",
          2019 => x"62",
          2020 => x"7a",
          2021 => x"84",
          2022 => x"8c",
          2023 => x"8b",
          2024 => x"8c",
          2025 => x"80",
          2026 => x"0b",
          2027 => x"5b",
          2028 => x"8d",
          2029 => x"82",
          2030 => x"38",
          2031 => x"82",
          2032 => x"54",
          2033 => x"d5",
          2034 => x"51",
          2035 => x"83",
          2036 => x"84",
          2037 => x"7d",
          2038 => x"80",
          2039 => x"0a",
          2040 => x"0a",
          2041 => x"f5",
          2042 => x"ba",
          2043 => x"ba",
          2044 => x"70",
          2045 => x"07",
          2046 => x"5b",
          2047 => x"5a",
          2048 => x"83",
          2049 => x"78",
          2050 => x"78",
          2051 => x"38",
          2052 => x"81",
          2053 => x"5a",
          2054 => x"38",
          2055 => x"61",
          2056 => x"5d",
          2057 => x"38",
          2058 => x"81",
          2059 => x"51",
          2060 => x"3f",
          2061 => x"51",
          2062 => x"7e",
          2063 => x"53",
          2064 => x"51",
          2065 => x"0b",
          2066 => x"80",
          2067 => x"ff",
          2068 => x"79",
          2069 => x"81",
          2070 => x"8c",
          2071 => x"9c",
          2072 => x"96",
          2073 => x"8c",
          2074 => x"38",
          2075 => x"0b",
          2076 => x"34",
          2077 => x"53",
          2078 => x"7e",
          2079 => x"91",
          2080 => x"8c",
          2081 => x"a0",
          2082 => x"8c",
          2083 => x"e6",
          2084 => x"83",
          2085 => x"70",
          2086 => x"5f",
          2087 => x"2e",
          2088 => x"fc",
          2089 => x"39",
          2090 => x"51",
          2091 => x"3f",
          2092 => x"0b",
          2093 => x"34",
          2094 => x"53",
          2095 => x"7e",
          2096 => x"3f",
          2097 => x"5a",
          2098 => x"38",
          2099 => x"1a",
          2100 => x"1b",
          2101 => x"81",
          2102 => x"80",
          2103 => x"10",
          2104 => x"05",
          2105 => x"04",
          2106 => x"51",
          2107 => x"9a",
          2108 => x"53",
          2109 => x"52",
          2110 => x"f1",
          2111 => x"7e",
          2112 => x"b8",
          2113 => x"c3",
          2114 => x"8c",
          2115 => x"09",
          2116 => x"a4",
          2117 => x"9a",
          2118 => x"41",
          2119 => x"83",
          2120 => x"de",
          2121 => x"51",
          2122 => x"3f",
          2123 => x"83",
          2124 => x"7b",
          2125 => x"98",
          2126 => x"83",
          2127 => x"7c",
          2128 => x"3f",
          2129 => x"81",
          2130 => x"fa",
          2131 => x"dd",
          2132 => x"39",
          2133 => x"51",
          2134 => x"fa",
          2135 => x"8e",
          2136 => x"de",
          2137 => x"ac",
          2138 => x"3f",
          2139 => x"04",
          2140 => x"51",
          2141 => x"d0",
          2142 => x"c6",
          2143 => x"ff",
          2144 => x"ff",
          2145 => x"ec",
          2146 => x"ba",
          2147 => x"2e",
          2148 => x"68",
          2149 => x"dc",
          2150 => x"3f",
          2151 => x"2d",
          2152 => x"08",
          2153 => x"9a",
          2154 => x"8c",
          2155 => x"d6",
          2156 => x"d7",
          2157 => x"39",
          2158 => x"84",
          2159 => x"80",
          2160 => x"c5",
          2161 => x"8c",
          2162 => x"f9",
          2163 => x"52",
          2164 => x"51",
          2165 => x"68",
          2166 => x"b8",
          2167 => x"11",
          2168 => x"05",
          2169 => x"3f",
          2170 => x"08",
          2171 => x"d2",
          2172 => x"fe",
          2173 => x"ff",
          2174 => x"e9",
          2175 => x"ba",
          2176 => x"d0",
          2177 => x"78",
          2178 => x"52",
          2179 => x"51",
          2180 => x"84",
          2181 => x"53",
          2182 => x"7e",
          2183 => x"3f",
          2184 => x"33",
          2185 => x"2e",
          2186 => x"78",
          2187 => x"d3",
          2188 => x"05",
          2189 => x"cf",
          2190 => x"fe",
          2191 => x"ff",
          2192 => x"e8",
          2193 => x"ba",
          2194 => x"2e",
          2195 => x"b8",
          2196 => x"11",
          2197 => x"05",
          2198 => x"3f",
          2199 => x"08",
          2200 => x"64",
          2201 => x"53",
          2202 => x"d7",
          2203 => x"9b",
          2204 => x"ec",
          2205 => x"f8",
          2206 => x"cf",
          2207 => x"48",
          2208 => x"78",
          2209 => x"ba",
          2210 => x"26",
          2211 => x"64",
          2212 => x"46",
          2213 => x"b8",
          2214 => x"11",
          2215 => x"05",
          2216 => x"3f",
          2217 => x"08",
          2218 => x"96",
          2219 => x"fe",
          2220 => x"ff",
          2221 => x"e9",
          2222 => x"ba",
          2223 => x"2e",
          2224 => x"b8",
          2225 => x"11",
          2226 => x"05",
          2227 => x"3f",
          2228 => x"08",
          2229 => x"ea",
          2230 => x"cc",
          2231 => x"3f",
          2232 => x"59",
          2233 => x"83",
          2234 => x"70",
          2235 => x"5f",
          2236 => x"7d",
          2237 => x"7a",
          2238 => x"78",
          2239 => x"52",
          2240 => x"51",
          2241 => x"66",
          2242 => x"81",
          2243 => x"47",
          2244 => x"b8",
          2245 => x"11",
          2246 => x"05",
          2247 => x"3f",
          2248 => x"08",
          2249 => x"9a",
          2250 => x"fe",
          2251 => x"ff",
          2252 => x"e8",
          2253 => x"ba",
          2254 => x"2e",
          2255 => x"b8",
          2256 => x"11",
          2257 => x"05",
          2258 => x"3f",
          2259 => x"08",
          2260 => x"ee",
          2261 => x"f8",
          2262 => x"3f",
          2263 => x"67",
          2264 => x"38",
          2265 => x"70",
          2266 => x"33",
          2267 => x"81",
          2268 => x"39",
          2269 => x"84",
          2270 => x"80",
          2271 => x"89",
          2272 => x"8c",
          2273 => x"f6",
          2274 => x"3d",
          2275 => x"53",
          2276 => x"51",
          2277 => x"84",
          2278 => x"b1",
          2279 => x"33",
          2280 => x"d8",
          2281 => x"e3",
          2282 => x"ec",
          2283 => x"f8",
          2284 => x"cc",
          2285 => x"48",
          2286 => x"78",
          2287 => x"82",
          2288 => x"26",
          2289 => x"68",
          2290 => x"d1",
          2291 => x"02",
          2292 => x"33",
          2293 => x"81",
          2294 => x"3d",
          2295 => x"53",
          2296 => x"51",
          2297 => x"84",
          2298 => x"80",
          2299 => x"38",
          2300 => x"80",
          2301 => x"79",
          2302 => x"05",
          2303 => x"fe",
          2304 => x"ff",
          2305 => x"e7",
          2306 => x"ba",
          2307 => x"bd",
          2308 => x"39",
          2309 => x"84",
          2310 => x"80",
          2311 => x"e9",
          2312 => x"8c",
          2313 => x"f5",
          2314 => x"3d",
          2315 => x"53",
          2316 => x"51",
          2317 => x"84",
          2318 => x"80",
          2319 => x"38",
          2320 => x"f8",
          2321 => x"80",
          2322 => x"bd",
          2323 => x"8c",
          2324 => x"84",
          2325 => x"46",
          2326 => x"51",
          2327 => x"68",
          2328 => x"78",
          2329 => x"38",
          2330 => x"79",
          2331 => x"5b",
          2332 => x"26",
          2333 => x"51",
          2334 => x"f4",
          2335 => x"3d",
          2336 => x"51",
          2337 => x"84",
          2338 => x"b9",
          2339 => x"05",
          2340 => x"d8",
          2341 => x"84",
          2342 => x"52",
          2343 => x"f9",
          2344 => x"8c",
          2345 => x"f4",
          2346 => x"ba",
          2347 => x"e7",
          2348 => x"8e",
          2349 => x"ff",
          2350 => x"ff",
          2351 => x"e5",
          2352 => x"ba",
          2353 => x"38",
          2354 => x"33",
          2355 => x"2e",
          2356 => x"83",
          2357 => x"49",
          2358 => x"fc",
          2359 => x"80",
          2360 => x"a5",
          2361 => x"8c",
          2362 => x"83",
          2363 => x"5a",
          2364 => x"83",
          2365 => x"f2",
          2366 => x"b8",
          2367 => x"11",
          2368 => x"05",
          2369 => x"3f",
          2370 => x"08",
          2371 => x"38",
          2372 => x"5c",
          2373 => x"83",
          2374 => x"7a",
          2375 => x"30",
          2376 => x"9f",
          2377 => x"5c",
          2378 => x"80",
          2379 => x"7a",
          2380 => x"38",
          2381 => x"d8",
          2382 => x"ba",
          2383 => x"68",
          2384 => x"66",
          2385 => x"eb",
          2386 => x"d8",
          2387 => x"a6",
          2388 => x"39",
          2389 => x"0c",
          2390 => x"05",
          2391 => x"fe",
          2392 => x"ff",
          2393 => x"e2",
          2394 => x"ba",
          2395 => x"2e",
          2396 => x"64",
          2397 => x"59",
          2398 => x"45",
          2399 => x"f0",
          2400 => x"80",
          2401 => x"fd",
          2402 => x"8c",
          2403 => x"f2",
          2404 => x"5e",
          2405 => x"05",
          2406 => x"82",
          2407 => x"7d",
          2408 => x"fe",
          2409 => x"ff",
          2410 => x"e1",
          2411 => x"ba",
          2412 => x"2e",
          2413 => x"64",
          2414 => x"ce",
          2415 => x"70",
          2416 => x"23",
          2417 => x"3d",
          2418 => x"53",
          2419 => x"51",
          2420 => x"84",
          2421 => x"ff",
          2422 => x"e6",
          2423 => x"fe",
          2424 => x"ff",
          2425 => x"e3",
          2426 => x"ba",
          2427 => x"2e",
          2428 => x"68",
          2429 => x"db",
          2430 => x"34",
          2431 => x"49",
          2432 => x"b8",
          2433 => x"11",
          2434 => x"05",
          2435 => x"3f",
          2436 => x"08",
          2437 => x"98",
          2438 => x"71",
          2439 => x"84",
          2440 => x"59",
          2441 => x"7a",
          2442 => x"81",
          2443 => x"38",
          2444 => x"d6",
          2445 => x"53",
          2446 => x"52",
          2447 => x"eb",
          2448 => x"39",
          2449 => x"51",
          2450 => x"f3",
          2451 => x"d8",
          2452 => x"a2",
          2453 => x"39",
          2454 => x"f0",
          2455 => x"80",
          2456 => x"a1",
          2457 => x"8c",
          2458 => x"b8",
          2459 => x"02",
          2460 => x"22",
          2461 => x"05",
          2462 => x"45",
          2463 => x"83",
          2464 => x"5c",
          2465 => x"80",
          2466 => x"f2",
          2467 => x"fc",
          2468 => x"f3",
          2469 => x"7b",
          2470 => x"38",
          2471 => x"08",
          2472 => x"39",
          2473 => x"51",
          2474 => x"64",
          2475 => x"39",
          2476 => x"51",
          2477 => x"64",
          2478 => x"39",
          2479 => x"33",
          2480 => x"2e",
          2481 => x"f2",
          2482 => x"fc",
          2483 => x"d8",
          2484 => x"a2",
          2485 => x"39",
          2486 => x"33",
          2487 => x"2e",
          2488 => x"f2",
          2489 => x"fc",
          2490 => x"f3",
          2491 => x"7d",
          2492 => x"38",
          2493 => x"08",
          2494 => x"39",
          2495 => x"33",
          2496 => x"2e",
          2497 => x"f2",
          2498 => x"fb",
          2499 => x"f3",
          2500 => x"7c",
          2501 => x"38",
          2502 => x"08",
          2503 => x"39",
          2504 => x"33",
          2505 => x"2e",
          2506 => x"f2",
          2507 => x"fb",
          2508 => x"f2",
          2509 => x"80",
          2510 => x"9c",
          2511 => x"f8",
          2512 => x"47",
          2513 => x"f3",
          2514 => x"0b",
          2515 => x"34",
          2516 => x"8c",
          2517 => x"57",
          2518 => x"52",
          2519 => x"c8",
          2520 => x"8c",
          2521 => x"77",
          2522 => x"87",
          2523 => x"75",
          2524 => x"3f",
          2525 => x"8c",
          2526 => x"0c",
          2527 => x"9c",
          2528 => x"57",
          2529 => x"52",
          2530 => x"9c",
          2531 => x"8c",
          2532 => x"77",
          2533 => x"87",
          2534 => x"75",
          2535 => x"3f",
          2536 => x"8c",
          2537 => x"0c",
          2538 => x"0b",
          2539 => x"84",
          2540 => x"83",
          2541 => x"94",
          2542 => x"bc",
          2543 => x"c7",
          2544 => x"02",
          2545 => x"05",
          2546 => x"84",
          2547 => x"89",
          2548 => x"13",
          2549 => x"0c",
          2550 => x"0c",
          2551 => x"3f",
          2552 => x"95",
          2553 => x"8d",
          2554 => x"3f",
          2555 => x"52",
          2556 => x"51",
          2557 => x"83",
          2558 => x"22",
          2559 => x"87",
          2560 => x"84",
          2561 => x"90",
          2562 => x"33",
          2563 => x"98",
          2564 => x"3f",
          2565 => x"ec",
          2566 => x"04",
          2567 => x"77",
          2568 => x"56",
          2569 => x"53",
          2570 => x"81",
          2571 => x"33",
          2572 => x"06",
          2573 => x"a0",
          2574 => x"06",
          2575 => x"15",
          2576 => x"81",
          2577 => x"53",
          2578 => x"2e",
          2579 => x"81",
          2580 => x"73",
          2581 => x"82",
          2582 => x"72",
          2583 => x"e7",
          2584 => x"33",
          2585 => x"06",
          2586 => x"70",
          2587 => x"38",
          2588 => x"80",
          2589 => x"73",
          2590 => x"38",
          2591 => x"e1",
          2592 => x"81",
          2593 => x"54",
          2594 => x"09",
          2595 => x"38",
          2596 => x"a2",
          2597 => x"70",
          2598 => x"07",
          2599 => x"72",
          2600 => x"38",
          2601 => x"81",
          2602 => x"71",
          2603 => x"51",
          2604 => x"8c",
          2605 => x"0d",
          2606 => x"2e",
          2607 => x"80",
          2608 => x"38",
          2609 => x"80",
          2610 => x"81",
          2611 => x"54",
          2612 => x"2e",
          2613 => x"54",
          2614 => x"15",
          2615 => x"53",
          2616 => x"2e",
          2617 => x"fe",
          2618 => x"39",
          2619 => x"76",
          2620 => x"8b",
          2621 => x"84",
          2622 => x"86",
          2623 => x"86",
          2624 => x"52",
          2625 => x"fd",
          2626 => x"8c",
          2627 => x"e5",
          2628 => x"ba",
          2629 => x"3d",
          2630 => x"3d",
          2631 => x"11",
          2632 => x"52",
          2633 => x"70",
          2634 => x"98",
          2635 => x"33",
          2636 => x"82",
          2637 => x"26",
          2638 => x"84",
          2639 => x"83",
          2640 => x"26",
          2641 => x"85",
          2642 => x"84",
          2643 => x"26",
          2644 => x"86",
          2645 => x"85",
          2646 => x"26",
          2647 => x"88",
          2648 => x"86",
          2649 => x"e7",
          2650 => x"38",
          2651 => x"54",
          2652 => x"87",
          2653 => x"cc",
          2654 => x"87",
          2655 => x"0c",
          2656 => x"c0",
          2657 => x"82",
          2658 => x"c0",
          2659 => x"83",
          2660 => x"c0",
          2661 => x"84",
          2662 => x"c0",
          2663 => x"85",
          2664 => x"c0",
          2665 => x"86",
          2666 => x"c0",
          2667 => x"74",
          2668 => x"a4",
          2669 => x"c0",
          2670 => x"80",
          2671 => x"98",
          2672 => x"52",
          2673 => x"8c",
          2674 => x"0d",
          2675 => x"0d",
          2676 => x"c0",
          2677 => x"81",
          2678 => x"c0",
          2679 => x"5e",
          2680 => x"87",
          2681 => x"08",
          2682 => x"1c",
          2683 => x"98",
          2684 => x"79",
          2685 => x"87",
          2686 => x"08",
          2687 => x"1c",
          2688 => x"98",
          2689 => x"79",
          2690 => x"87",
          2691 => x"08",
          2692 => x"1c",
          2693 => x"98",
          2694 => x"7b",
          2695 => x"87",
          2696 => x"08",
          2697 => x"1c",
          2698 => x"0c",
          2699 => x"ff",
          2700 => x"83",
          2701 => x"58",
          2702 => x"57",
          2703 => x"56",
          2704 => x"55",
          2705 => x"54",
          2706 => x"53",
          2707 => x"ff",
          2708 => x"d8",
          2709 => x"bf",
          2710 => x"3d",
          2711 => x"3d",
          2712 => x"05",
          2713 => x"81",
          2714 => x"72",
          2715 => x"b1",
          2716 => x"8c",
          2717 => x"70",
          2718 => x"52",
          2719 => x"09",
          2720 => x"38",
          2721 => x"e3",
          2722 => x"ba",
          2723 => x"3d",
          2724 => x"51",
          2725 => x"3f",
          2726 => x"08",
          2727 => x"98",
          2728 => x"71",
          2729 => x"81",
          2730 => x"72",
          2731 => x"f1",
          2732 => x"8c",
          2733 => x"70",
          2734 => x"52",
          2735 => x"d2",
          2736 => x"fd",
          2737 => x"70",
          2738 => x"88",
          2739 => x"51",
          2740 => x"3f",
          2741 => x"08",
          2742 => x"98",
          2743 => x"71",
          2744 => x"38",
          2745 => x"81",
          2746 => x"83",
          2747 => x"38",
          2748 => x"8c",
          2749 => x"0d",
          2750 => x"0d",
          2751 => x"33",
          2752 => x"33",
          2753 => x"06",
          2754 => x"70",
          2755 => x"f4",
          2756 => x"94",
          2757 => x"96",
          2758 => x"06",
          2759 => x"70",
          2760 => x"38",
          2761 => x"70",
          2762 => x"51",
          2763 => x"72",
          2764 => x"06",
          2765 => x"2e",
          2766 => x"93",
          2767 => x"52",
          2768 => x"73",
          2769 => x"51",
          2770 => x"80",
          2771 => x"2e",
          2772 => x"c0",
          2773 => x"74",
          2774 => x"84",
          2775 => x"86",
          2776 => x"71",
          2777 => x"81",
          2778 => x"70",
          2779 => x"81",
          2780 => x"53",
          2781 => x"cb",
          2782 => x"2a",
          2783 => x"71",
          2784 => x"38",
          2785 => x"84",
          2786 => x"2a",
          2787 => x"53",
          2788 => x"cf",
          2789 => x"ff",
          2790 => x"8f",
          2791 => x"30",
          2792 => x"51",
          2793 => x"83",
          2794 => x"83",
          2795 => x"fa",
          2796 => x"55",
          2797 => x"70",
          2798 => x"70",
          2799 => x"e7",
          2800 => x"83",
          2801 => x"70",
          2802 => x"54",
          2803 => x"80",
          2804 => x"38",
          2805 => x"94",
          2806 => x"2a",
          2807 => x"53",
          2808 => x"80",
          2809 => x"71",
          2810 => x"81",
          2811 => x"70",
          2812 => x"81",
          2813 => x"53",
          2814 => x"8a",
          2815 => x"2a",
          2816 => x"71",
          2817 => x"81",
          2818 => x"87",
          2819 => x"52",
          2820 => x"86",
          2821 => x"94",
          2822 => x"72",
          2823 => x"75",
          2824 => x"73",
          2825 => x"76",
          2826 => x"0c",
          2827 => x"04",
          2828 => x"70",
          2829 => x"51",
          2830 => x"72",
          2831 => x"06",
          2832 => x"2e",
          2833 => x"93",
          2834 => x"52",
          2835 => x"ff",
          2836 => x"c0",
          2837 => x"70",
          2838 => x"81",
          2839 => x"52",
          2840 => x"d7",
          2841 => x"0d",
          2842 => x"80",
          2843 => x"2a",
          2844 => x"52",
          2845 => x"84",
          2846 => x"c0",
          2847 => x"83",
          2848 => x"87",
          2849 => x"08",
          2850 => x"0c",
          2851 => x"94",
          2852 => x"d0",
          2853 => x"9e",
          2854 => x"f2",
          2855 => x"c0",
          2856 => x"83",
          2857 => x"87",
          2858 => x"08",
          2859 => x"0c",
          2860 => x"ac",
          2861 => x"e0",
          2862 => x"9e",
          2863 => x"f2",
          2864 => x"c0",
          2865 => x"83",
          2866 => x"87",
          2867 => x"08",
          2868 => x"0c",
          2869 => x"bc",
          2870 => x"f0",
          2871 => x"9e",
          2872 => x"f2",
          2873 => x"c0",
          2874 => x"83",
          2875 => x"87",
          2876 => x"08",
          2877 => x"f2",
          2878 => x"c0",
          2879 => x"83",
          2880 => x"87",
          2881 => x"08",
          2882 => x"0c",
          2883 => x"8c",
          2884 => x"88",
          2885 => x"83",
          2886 => x"80",
          2887 => x"9e",
          2888 => x"84",
          2889 => x"51",
          2890 => x"82",
          2891 => x"83",
          2892 => x"80",
          2893 => x"9e",
          2894 => x"88",
          2895 => x"51",
          2896 => x"80",
          2897 => x"81",
          2898 => x"f3",
          2899 => x"0b",
          2900 => x"90",
          2901 => x"80",
          2902 => x"52",
          2903 => x"2e",
          2904 => x"52",
          2905 => x"8f",
          2906 => x"87",
          2907 => x"08",
          2908 => x"80",
          2909 => x"52",
          2910 => x"83",
          2911 => x"71",
          2912 => x"34",
          2913 => x"c0",
          2914 => x"70",
          2915 => x"06",
          2916 => x"70",
          2917 => x"38",
          2918 => x"83",
          2919 => x"80",
          2920 => x"9e",
          2921 => x"90",
          2922 => x"51",
          2923 => x"80",
          2924 => x"81",
          2925 => x"f3",
          2926 => x"0b",
          2927 => x"90",
          2928 => x"80",
          2929 => x"52",
          2930 => x"2e",
          2931 => x"52",
          2932 => x"93",
          2933 => x"87",
          2934 => x"08",
          2935 => x"80",
          2936 => x"52",
          2937 => x"83",
          2938 => x"71",
          2939 => x"34",
          2940 => x"c0",
          2941 => x"70",
          2942 => x"06",
          2943 => x"70",
          2944 => x"38",
          2945 => x"83",
          2946 => x"80",
          2947 => x"9e",
          2948 => x"80",
          2949 => x"51",
          2950 => x"80",
          2951 => x"81",
          2952 => x"f3",
          2953 => x"0b",
          2954 => x"90",
          2955 => x"80",
          2956 => x"52",
          2957 => x"83",
          2958 => x"71",
          2959 => x"34",
          2960 => x"90",
          2961 => x"06",
          2962 => x"53",
          2963 => x"f3",
          2964 => x"0b",
          2965 => x"90",
          2966 => x"80",
          2967 => x"52",
          2968 => x"83",
          2969 => x"71",
          2970 => x"34",
          2971 => x"90",
          2972 => x"06",
          2973 => x"53",
          2974 => x"f3",
          2975 => x"0b",
          2976 => x"90",
          2977 => x"06",
          2978 => x"70",
          2979 => x"38",
          2980 => x"83",
          2981 => x"87",
          2982 => x"08",
          2983 => x"70",
          2984 => x"34",
          2985 => x"04",
          2986 => x"82",
          2987 => x"0d",
          2988 => x"51",
          2989 => x"3f",
          2990 => x"33",
          2991 => x"aa",
          2992 => x"a0",
          2993 => x"3f",
          2994 => x"33",
          2995 => x"fa",
          2996 => x"93",
          2997 => x"85",
          2998 => x"f3",
          2999 => x"75",
          3000 => x"83",
          3001 => x"55",
          3002 => x"38",
          3003 => x"33",
          3004 => x"d6",
          3005 => x"97",
          3006 => x"84",
          3007 => x"f3",
          3008 => x"73",
          3009 => x"83",
          3010 => x"55",
          3011 => x"38",
          3012 => x"33",
          3013 => x"cf",
          3014 => x"8f",
          3015 => x"83",
          3016 => x"f3",
          3017 => x"74",
          3018 => x"83",
          3019 => x"56",
          3020 => x"38",
          3021 => x"33",
          3022 => x"ec",
          3023 => x"b8",
          3024 => x"3f",
          3025 => x"08",
          3026 => x"c4",
          3027 => x"bb",
          3028 => x"f4",
          3029 => x"d9",
          3030 => x"b5",
          3031 => x"f2",
          3032 => x"83",
          3033 => x"ff",
          3034 => x"83",
          3035 => x"c2",
          3036 => x"f2",
          3037 => x"83",
          3038 => x"ff",
          3039 => x"83",
          3040 => x"56",
          3041 => x"52",
          3042 => x"9c",
          3043 => x"8c",
          3044 => x"c0",
          3045 => x"31",
          3046 => x"ba",
          3047 => x"83",
          3048 => x"ff",
          3049 => x"83",
          3050 => x"55",
          3051 => x"38",
          3052 => x"33",
          3053 => x"38",
          3054 => x"a5",
          3055 => x"0d",
          3056 => x"88",
          3057 => x"84",
          3058 => x"51",
          3059 => x"84",
          3060 => x"bd",
          3061 => x"76",
          3062 => x"54",
          3063 => x"08",
          3064 => x"98",
          3065 => x"a3",
          3066 => x"c2",
          3067 => x"3d",
          3068 => x"f3",
          3069 => x"bd",
          3070 => x"75",
          3071 => x"3f",
          3072 => x"08",
          3073 => x"29",
          3074 => x"54",
          3075 => x"8c",
          3076 => x"db",
          3077 => x"b3",
          3078 => x"f3",
          3079 => x"74",
          3080 => x"94",
          3081 => x"39",
          3082 => x"51",
          3083 => x"83",
          3084 => x"c0",
          3085 => x"f2",
          3086 => x"83",
          3087 => x"ff",
          3088 => x"83",
          3089 => x"52",
          3090 => x"51",
          3091 => x"3f",
          3092 => x"08",
          3093 => x"94",
          3094 => x"af",
          3095 => x"bc",
          3096 => x"3f",
          3097 => x"22",
          3098 => x"c4",
          3099 => x"9b",
          3100 => x"80",
          3101 => x"84",
          3102 => x"51",
          3103 => x"84",
          3104 => x"bd",
          3105 => x"76",
          3106 => x"54",
          3107 => x"08",
          3108 => x"ec",
          3109 => x"f3",
          3110 => x"93",
          3111 => x"80",
          3112 => x"38",
          3113 => x"83",
          3114 => x"ff",
          3115 => x"83",
          3116 => x"54",
          3117 => x"fd",
          3118 => x"ec",
          3119 => x"80",
          3120 => x"b2",
          3121 => x"95",
          3122 => x"80",
          3123 => x"38",
          3124 => x"dc",
          3125 => x"bf",
          3126 => x"f3",
          3127 => x"74",
          3128 => x"c7",
          3129 => x"83",
          3130 => x"ff",
          3131 => x"83",
          3132 => x"54",
          3133 => x"fc",
          3134 => x"39",
          3135 => x"33",
          3136 => x"ac",
          3137 => x"83",
          3138 => x"8d",
          3139 => x"80",
          3140 => x"38",
          3141 => x"f3",
          3142 => x"83",
          3143 => x"ff",
          3144 => x"83",
          3145 => x"55",
          3146 => x"fb",
          3147 => x"39",
          3148 => x"33",
          3149 => x"ec",
          3150 => x"cf",
          3151 => x"9b",
          3152 => x"80",
          3153 => x"38",
          3154 => x"f2",
          3155 => x"f2",
          3156 => x"54",
          3157 => x"8c",
          3158 => x"af",
          3159 => x"97",
          3160 => x"80",
          3161 => x"38",
          3162 => x"f2",
          3163 => x"f2",
          3164 => x"54",
          3165 => x"a8",
          3166 => x"8f",
          3167 => x"92",
          3168 => x"80",
          3169 => x"38",
          3170 => x"f2",
          3171 => x"f2",
          3172 => x"54",
          3173 => x"c4",
          3174 => x"ef",
          3175 => x"91",
          3176 => x"80",
          3177 => x"38",
          3178 => x"f2",
          3179 => x"f2",
          3180 => x"54",
          3181 => x"e0",
          3182 => x"cf",
          3183 => x"90",
          3184 => x"80",
          3185 => x"38",
          3186 => x"f2",
          3187 => x"f2",
          3188 => x"54",
          3189 => x"fc",
          3190 => x"af",
          3191 => x"93",
          3192 => x"80",
          3193 => x"38",
          3194 => x"de",
          3195 => x"b0",
          3196 => x"d9",
          3197 => x"bc",
          3198 => x"f3",
          3199 => x"74",
          3200 => x"cd",
          3201 => x"ff",
          3202 => x"8e",
          3203 => x"71",
          3204 => x"38",
          3205 => x"83",
          3206 => x"52",
          3207 => x"83",
          3208 => x"ff",
          3209 => x"83",
          3210 => x"83",
          3211 => x"ff",
          3212 => x"83",
          3213 => x"83",
          3214 => x"ff",
          3215 => x"83",
          3216 => x"83",
          3217 => x"ff",
          3218 => x"83",
          3219 => x"83",
          3220 => x"ff",
          3221 => x"83",
          3222 => x"83",
          3223 => x"ff",
          3224 => x"83",
          3225 => x"71",
          3226 => x"04",
          3227 => x"c0",
          3228 => x"04",
          3229 => x"08",
          3230 => x"84",
          3231 => x"3d",
          3232 => x"08",
          3233 => x"5a",
          3234 => x"57",
          3235 => x"83",
          3236 => x"51",
          3237 => x"3f",
          3238 => x"08",
          3239 => x"8b",
          3240 => x"0b",
          3241 => x"08",
          3242 => x"f8",
          3243 => x"82",
          3244 => x"84",
          3245 => x"80",
          3246 => x"76",
          3247 => x"3f",
          3248 => x"08",
          3249 => x"55",
          3250 => x"ba",
          3251 => x"8e",
          3252 => x"8c",
          3253 => x"70",
          3254 => x"80",
          3255 => x"09",
          3256 => x"72",
          3257 => x"51",
          3258 => x"76",
          3259 => x"73",
          3260 => x"83",
          3261 => x"8c",
          3262 => x"51",
          3263 => x"3f",
          3264 => x"08",
          3265 => x"76",
          3266 => x"77",
          3267 => x"0c",
          3268 => x"04",
          3269 => x"51",
          3270 => x"3f",
          3271 => x"09",
          3272 => x"38",
          3273 => x"51",
          3274 => x"79",
          3275 => x"fb",
          3276 => x"08",
          3277 => x"8c",
          3278 => x"76",
          3279 => x"b0",
          3280 => x"c7",
          3281 => x"84",
          3282 => x"a9",
          3283 => x"d8",
          3284 => x"3d",
          3285 => x"08",
          3286 => x"72",
          3287 => x"5a",
          3288 => x"2e",
          3289 => x"80",
          3290 => x"59",
          3291 => x"10",
          3292 => x"80",
          3293 => x"52",
          3294 => x"af",
          3295 => x"8c",
          3296 => x"52",
          3297 => x"c0",
          3298 => x"ba",
          3299 => x"38",
          3300 => x"54",
          3301 => x"81",
          3302 => x"82",
          3303 => x"81",
          3304 => x"ff",
          3305 => x"82",
          3306 => x"38",
          3307 => x"84",
          3308 => x"aa",
          3309 => x"81",
          3310 => x"3d",
          3311 => x"53",
          3312 => x"51",
          3313 => x"84",
          3314 => x"80",
          3315 => x"ff",
          3316 => x"52",
          3317 => x"a6",
          3318 => x"8c",
          3319 => x"06",
          3320 => x"2e",
          3321 => x"16",
          3322 => x"06",
          3323 => x"76",
          3324 => x"38",
          3325 => x"78",
          3326 => x"56",
          3327 => x"fe",
          3328 => x"15",
          3329 => x"33",
          3330 => x"a0",
          3331 => x"06",
          3332 => x"75",
          3333 => x"38",
          3334 => x"3d",
          3335 => x"cd",
          3336 => x"ba",
          3337 => x"83",
          3338 => x"52",
          3339 => x"b9",
          3340 => x"8c",
          3341 => x"38",
          3342 => x"08",
          3343 => x"52",
          3344 => x"cf",
          3345 => x"ba",
          3346 => x"2e",
          3347 => x"51",
          3348 => x"3f",
          3349 => x"08",
          3350 => x"84",
          3351 => x"25",
          3352 => x"ba",
          3353 => x"05",
          3354 => x"55",
          3355 => x"77",
          3356 => x"81",
          3357 => x"f8",
          3358 => x"ab",
          3359 => x"ff",
          3360 => x"06",
          3361 => x"81",
          3362 => x"8c",
          3363 => x"0d",
          3364 => x"0d",
          3365 => x"b7",
          3366 => x"3d",
          3367 => x"5c",
          3368 => x"3d",
          3369 => x"fc",
          3370 => x"f8",
          3371 => x"74",
          3372 => x"83",
          3373 => x"56",
          3374 => x"2e",
          3375 => x"77",
          3376 => x"8d",
          3377 => x"77",
          3378 => x"78",
          3379 => x"77",
          3380 => x"fd",
          3381 => x"b4",
          3382 => x"80",
          3383 => x"3f",
          3384 => x"08",
          3385 => x"98",
          3386 => x"79",
          3387 => x"38",
          3388 => x"06",
          3389 => x"33",
          3390 => x"70",
          3391 => x"d1",
          3392 => x"98",
          3393 => x"2c",
          3394 => x"05",
          3395 => x"83",
          3396 => x"70",
          3397 => x"33",
          3398 => x"5d",
          3399 => x"58",
          3400 => x"57",
          3401 => x"80",
          3402 => x"75",
          3403 => x"38",
          3404 => x"0a",
          3405 => x"0a",
          3406 => x"2c",
          3407 => x"76",
          3408 => x"38",
          3409 => x"70",
          3410 => x"57",
          3411 => x"de",
          3412 => x"42",
          3413 => x"25",
          3414 => x"de",
          3415 => x"18",
          3416 => x"41",
          3417 => x"81",
          3418 => x"80",
          3419 => x"75",
          3420 => x"34",
          3421 => x"80",
          3422 => x"38",
          3423 => x"98",
          3424 => x"2c",
          3425 => x"33",
          3426 => x"70",
          3427 => x"98",
          3428 => x"82",
          3429 => x"dc",
          3430 => x"53",
          3431 => x"5d",
          3432 => x"78",
          3433 => x"38",
          3434 => x"c8",
          3435 => x"39",
          3436 => x"ff",
          3437 => x"81",
          3438 => x"81",
          3439 => x"70",
          3440 => x"81",
          3441 => x"57",
          3442 => x"26",
          3443 => x"75",
          3444 => x"82",
          3445 => x"80",
          3446 => x"dc",
          3447 => x"57",
          3448 => x"ce",
          3449 => x"d8",
          3450 => x"70",
          3451 => x"78",
          3452 => x"bc",
          3453 => x"2e",
          3454 => x"fe",
          3455 => x"57",
          3456 => x"fe",
          3457 => x"e7",
          3458 => x"fd",
          3459 => x"57",
          3460 => x"38",
          3461 => x"c8",
          3462 => x"d1",
          3463 => x"7e",
          3464 => x"0c",
          3465 => x"95",
          3466 => x"38",
          3467 => x"83",
          3468 => x"57",
          3469 => x"83",
          3470 => x"08",
          3471 => x"0b",
          3472 => x"34",
          3473 => x"d1",
          3474 => x"39",
          3475 => x"33",
          3476 => x"2e",
          3477 => x"84",
          3478 => x"52",
          3479 => x"b6",
          3480 => x"d1",
          3481 => x"05",
          3482 => x"d1",
          3483 => x"eb",
          3484 => x"d0",
          3485 => x"ff",
          3486 => x"cc",
          3487 => x"55",
          3488 => x"fc",
          3489 => x"d5",
          3490 => x"81",
          3491 => x"84",
          3492 => x"7b",
          3493 => x"52",
          3494 => x"d5",
          3495 => x"39",
          3496 => x"8b",
          3497 => x"10",
          3498 => x"a8",
          3499 => x"57",
          3500 => x"83",
          3501 => x"d1",
          3502 => x"7c",
          3503 => x"cc",
          3504 => x"d0",
          3505 => x"74",
          3506 => x"38",
          3507 => x"08",
          3508 => x"ff",
          3509 => x"84",
          3510 => x"52",
          3511 => x"b5",
          3512 => x"d5",
          3513 => x"88",
          3514 => x"85",
          3515 => x"d0",
          3516 => x"5b",
          3517 => x"d0",
          3518 => x"ff",
          3519 => x"cc",
          3520 => x"ff",
          3521 => x"75",
          3522 => x"34",
          3523 => x"7c",
          3524 => x"f3",
          3525 => x"75",
          3526 => x"7c",
          3527 => x"f3",
          3528 => x"11",
          3529 => x"75",
          3530 => x"74",
          3531 => x"80",
          3532 => x"38",
          3533 => x"b7",
          3534 => x"ba",
          3535 => x"d1",
          3536 => x"ba",
          3537 => x"ff",
          3538 => x"53",
          3539 => x"51",
          3540 => x"3f",
          3541 => x"33",
          3542 => x"33",
          3543 => x"80",
          3544 => x"38",
          3545 => x"08",
          3546 => x"ff",
          3547 => x"84",
          3548 => x"52",
          3549 => x"b3",
          3550 => x"d5",
          3551 => x"88",
          3552 => x"ed",
          3553 => x"d0",
          3554 => x"55",
          3555 => x"d0",
          3556 => x"ff",
          3557 => x"39",
          3558 => x"33",
          3559 => x"06",
          3560 => x"33",
          3561 => x"75",
          3562 => x"af",
          3563 => x"f0",
          3564 => x"15",
          3565 => x"d1",
          3566 => x"16",
          3567 => x"55",
          3568 => x"3f",
          3569 => x"33",
          3570 => x"06",
          3571 => x"33",
          3572 => x"75",
          3573 => x"83",
          3574 => x"f0",
          3575 => x"15",
          3576 => x"d1",
          3577 => x"16",
          3578 => x"55",
          3579 => x"3f",
          3580 => x"33",
          3581 => x"06",
          3582 => x"33",
          3583 => x"77",
          3584 => x"a9",
          3585 => x"39",
          3586 => x"33",
          3587 => x"33",
          3588 => x"76",
          3589 => x"38",
          3590 => x"7a",
          3591 => x"34",
          3592 => x"70",
          3593 => x"81",
          3594 => x"57",
          3595 => x"24",
          3596 => x"84",
          3597 => x"52",
          3598 => x"b2",
          3599 => x"d1",
          3600 => x"98",
          3601 => x"2c",
          3602 => x"33",
          3603 => x"41",
          3604 => x"f9",
          3605 => x"d5",
          3606 => x"88",
          3607 => x"91",
          3608 => x"80",
          3609 => x"80",
          3610 => x"98",
          3611 => x"cc",
          3612 => x"5a",
          3613 => x"f8",
          3614 => x"d5",
          3615 => x"88",
          3616 => x"ed",
          3617 => x"80",
          3618 => x"80",
          3619 => x"98",
          3620 => x"cc",
          3621 => x"5a",
          3622 => x"ff",
          3623 => x"bb",
          3624 => x"58",
          3625 => x"78",
          3626 => x"f0",
          3627 => x"33",
          3628 => x"bd",
          3629 => x"80",
          3630 => x"80",
          3631 => x"98",
          3632 => x"cc",
          3633 => x"55",
          3634 => x"fe",
          3635 => x"16",
          3636 => x"33",
          3637 => x"d5",
          3638 => x"77",
          3639 => x"b1",
          3640 => x"81",
          3641 => x"81",
          3642 => x"70",
          3643 => x"d1",
          3644 => x"57",
          3645 => x"24",
          3646 => x"fe",
          3647 => x"d1",
          3648 => x"74",
          3649 => x"d3",
          3650 => x"f0",
          3651 => x"51",
          3652 => x"3f",
          3653 => x"33",
          3654 => x"76",
          3655 => x"34",
          3656 => x"06",
          3657 => x"84",
          3658 => x"7c",
          3659 => x"7f",
          3660 => x"f0",
          3661 => x"51",
          3662 => x"3f",
          3663 => x"52",
          3664 => x"8b",
          3665 => x"8c",
          3666 => x"06",
          3667 => x"cf",
          3668 => x"cc",
          3669 => x"80",
          3670 => x"38",
          3671 => x"33",
          3672 => x"83",
          3673 => x"70",
          3674 => x"56",
          3675 => x"38",
          3676 => x"87",
          3677 => x"f3",
          3678 => x"18",
          3679 => x"5b",
          3680 => x"3f",
          3681 => x"08",
          3682 => x"f3",
          3683 => x"10",
          3684 => x"a4",
          3685 => x"57",
          3686 => x"8b",
          3687 => x"f3",
          3688 => x"75",
          3689 => x"38",
          3690 => x"33",
          3691 => x"2e",
          3692 => x"80",
          3693 => x"d0",
          3694 => x"84",
          3695 => x"7b",
          3696 => x"0c",
          3697 => x"04",
          3698 => x"33",
          3699 => x"2e",
          3700 => x"d5",
          3701 => x"88",
          3702 => x"95",
          3703 => x"f0",
          3704 => x"51",
          3705 => x"3f",
          3706 => x"08",
          3707 => x"ff",
          3708 => x"84",
          3709 => x"ff",
          3710 => x"84",
          3711 => x"75",
          3712 => x"55",
          3713 => x"83",
          3714 => x"ff",
          3715 => x"80",
          3716 => x"d0",
          3717 => x"84",
          3718 => x"f5",
          3719 => x"7c",
          3720 => x"81",
          3721 => x"d1",
          3722 => x"74",
          3723 => x"38",
          3724 => x"08",
          3725 => x"ff",
          3726 => x"84",
          3727 => x"52",
          3728 => x"ae",
          3729 => x"d5",
          3730 => x"88",
          3731 => x"a1",
          3732 => x"d0",
          3733 => x"5d",
          3734 => x"d0",
          3735 => x"ff",
          3736 => x"cc",
          3737 => x"b8",
          3738 => x"9f",
          3739 => x"84",
          3740 => x"80",
          3741 => x"cc",
          3742 => x"ba",
          3743 => x"3d",
          3744 => x"d1",
          3745 => x"81",
          3746 => x"56",
          3747 => x"f4",
          3748 => x"d1",
          3749 => x"05",
          3750 => x"d1",
          3751 => x"16",
          3752 => x"d1",
          3753 => x"d5",
          3754 => x"88",
          3755 => x"c1",
          3756 => x"d0",
          3757 => x"2b",
          3758 => x"84",
          3759 => x"5a",
          3760 => x"76",
          3761 => x"ef",
          3762 => x"f0",
          3763 => x"51",
          3764 => x"3f",
          3765 => x"33",
          3766 => x"70",
          3767 => x"d1",
          3768 => x"57",
          3769 => x"7a",
          3770 => x"38",
          3771 => x"08",
          3772 => x"ff",
          3773 => x"74",
          3774 => x"29",
          3775 => x"05",
          3776 => x"84",
          3777 => x"5b",
          3778 => x"79",
          3779 => x"38",
          3780 => x"08",
          3781 => x"ff",
          3782 => x"74",
          3783 => x"29",
          3784 => x"05",
          3785 => x"84",
          3786 => x"5b",
          3787 => x"75",
          3788 => x"38",
          3789 => x"7b",
          3790 => x"17",
          3791 => x"84",
          3792 => x"52",
          3793 => x"ff",
          3794 => x"75",
          3795 => x"29",
          3796 => x"05",
          3797 => x"84",
          3798 => x"43",
          3799 => x"61",
          3800 => x"38",
          3801 => x"81",
          3802 => x"34",
          3803 => x"08",
          3804 => x"51",
          3805 => x"3f",
          3806 => x"0a",
          3807 => x"0a",
          3808 => x"2c",
          3809 => x"33",
          3810 => x"60",
          3811 => x"a7",
          3812 => x"39",
          3813 => x"33",
          3814 => x"06",
          3815 => x"60",
          3816 => x"38",
          3817 => x"33",
          3818 => x"27",
          3819 => x"98",
          3820 => x"2c",
          3821 => x"76",
          3822 => x"7b",
          3823 => x"33",
          3824 => x"75",
          3825 => x"29",
          3826 => x"05",
          3827 => x"84",
          3828 => x"52",
          3829 => x"78",
          3830 => x"81",
          3831 => x"84",
          3832 => x"77",
          3833 => x"7c",
          3834 => x"3d",
          3835 => x"84",
          3836 => x"57",
          3837 => x"8b",
          3838 => x"56",
          3839 => x"cc",
          3840 => x"84",
          3841 => x"70",
          3842 => x"29",
          3843 => x"05",
          3844 => x"79",
          3845 => x"44",
          3846 => x"60",
          3847 => x"ef",
          3848 => x"2b",
          3849 => x"78",
          3850 => x"5c",
          3851 => x"7a",
          3852 => x"38",
          3853 => x"08",
          3854 => x"ff",
          3855 => x"75",
          3856 => x"29",
          3857 => x"05",
          3858 => x"84",
          3859 => x"57",
          3860 => x"75",
          3861 => x"38",
          3862 => x"08",
          3863 => x"ff",
          3864 => x"75",
          3865 => x"29",
          3866 => x"05",
          3867 => x"84",
          3868 => x"57",
          3869 => x"76",
          3870 => x"38",
          3871 => x"83",
          3872 => x"56",
          3873 => x"f4",
          3874 => x"51",
          3875 => x"3f",
          3876 => x"08",
          3877 => x"34",
          3878 => x"08",
          3879 => x"81",
          3880 => x"52",
          3881 => x"ad",
          3882 => x"d1",
          3883 => x"d1",
          3884 => x"56",
          3885 => x"f4",
          3886 => x"d5",
          3887 => x"88",
          3888 => x"ad",
          3889 => x"f0",
          3890 => x"51",
          3891 => x"3f",
          3892 => x"08",
          3893 => x"ff",
          3894 => x"84",
          3895 => x"ff",
          3896 => x"84",
          3897 => x"7a",
          3898 => x"55",
          3899 => x"51",
          3900 => x"3f",
          3901 => x"08",
          3902 => x"0c",
          3903 => x"08",
          3904 => x"76",
          3905 => x"34",
          3906 => x"38",
          3907 => x"84",
          3908 => x"52",
          3909 => x"33",
          3910 => x"a8",
          3911 => x"81",
          3912 => x"81",
          3913 => x"70",
          3914 => x"d1",
          3915 => x"57",
          3916 => x"24",
          3917 => x"d1",
          3918 => x"98",
          3919 => x"2c",
          3920 => x"06",
          3921 => x"58",
          3922 => x"ef",
          3923 => x"e4",
          3924 => x"f8",
          3925 => x"ee",
          3926 => x"f3",
          3927 => x"56",
          3928 => x"74",
          3929 => x"16",
          3930 => x"56",
          3931 => x"f0",
          3932 => x"83",
          3933 => x"83",
          3934 => x"55",
          3935 => x"ee",
          3936 => x"51",
          3937 => x"3f",
          3938 => x"08",
          3939 => x"cd",
          3940 => x"83",
          3941 => x"93",
          3942 => x"5f",
          3943 => x"39",
          3944 => x"da",
          3945 => x"77",
          3946 => x"84",
          3947 => x"75",
          3948 => x"ac",
          3949 => x"39",
          3950 => x"aa",
          3951 => x"ba",
          3952 => x"d1",
          3953 => x"ba",
          3954 => x"ff",
          3955 => x"53",
          3956 => x"51",
          3957 => x"3f",
          3958 => x"d1",
          3959 => x"d1",
          3960 => x"57",
          3961 => x"2e",
          3962 => x"84",
          3963 => x"52",
          3964 => x"a6",
          3965 => x"d5",
          3966 => x"a0",
          3967 => x"f1",
          3968 => x"f0",
          3969 => x"51",
          3970 => x"3f",
          3971 => x"33",
          3972 => x"79",
          3973 => x"34",
          3974 => x"06",
          3975 => x"80",
          3976 => x"0b",
          3977 => x"34",
          3978 => x"d1",
          3979 => x"84",
          3980 => x"b4",
          3981 => x"75",
          3982 => x"ef",
          3983 => x"8c",
          3984 => x"cc",
          3985 => x"8c",
          3986 => x"06",
          3987 => x"75",
          3988 => x"ff",
          3989 => x"81",
          3990 => x"ff",
          3991 => x"cc",
          3992 => x"d0",
          3993 => x"5e",
          3994 => x"2e",
          3995 => x"84",
          3996 => x"52",
          3997 => x"a5",
          3998 => x"d5",
          3999 => x"a0",
          4000 => x"ed",
          4001 => x"f0",
          4002 => x"51",
          4003 => x"3f",
          4004 => x"33",
          4005 => x"76",
          4006 => x"34",
          4007 => x"06",
          4008 => x"75",
          4009 => x"83",
          4010 => x"8c",
          4011 => x"cc",
          4012 => x"8c",
          4013 => x"06",
          4014 => x"75",
          4015 => x"ff",
          4016 => x"ff",
          4017 => x"ff",
          4018 => x"cc",
          4019 => x"d0",
          4020 => x"5e",
          4021 => x"2e",
          4022 => x"84",
          4023 => x"52",
          4024 => x"a5",
          4025 => x"d5",
          4026 => x"a0",
          4027 => x"81",
          4028 => x"f0",
          4029 => x"51",
          4030 => x"3f",
          4031 => x"33",
          4032 => x"60",
          4033 => x"34",
          4034 => x"06",
          4035 => x"74",
          4036 => x"c9",
          4037 => x"fc",
          4038 => x"2b",
          4039 => x"83",
          4040 => x"81",
          4041 => x"52",
          4042 => x"dd",
          4043 => x"ba",
          4044 => x"0c",
          4045 => x"33",
          4046 => x"83",
          4047 => x"70",
          4048 => x"41",
          4049 => x"f4",
          4050 => x"53",
          4051 => x"51",
          4052 => x"3f",
          4053 => x"33",
          4054 => x"81",
          4055 => x"56",
          4056 => x"82",
          4057 => x"83",
          4058 => x"f4",
          4059 => x"3d",
          4060 => x"54",
          4061 => x"52",
          4062 => x"d9",
          4063 => x"f3",
          4064 => x"8a",
          4065 => x"d7",
          4066 => x"f8",
          4067 => x"e0",
          4068 => x"0b",
          4069 => x"34",
          4070 => x"d1",
          4071 => x"84",
          4072 => x"b4",
          4073 => x"93",
          4074 => x"84",
          4075 => x"51",
          4076 => x"3f",
          4077 => x"08",
          4078 => x"84",
          4079 => x"96",
          4080 => x"83",
          4081 => x"53",
          4082 => x"7a",
          4083 => x"c1",
          4084 => x"8c",
          4085 => x"ba",
          4086 => x"2e",
          4087 => x"e9",
          4088 => x"ba",
          4089 => x"ff",
          4090 => x"84",
          4091 => x"56",
          4092 => x"ba",
          4093 => x"80",
          4094 => x"ba",
          4095 => x"05",
          4096 => x"56",
          4097 => x"75",
          4098 => x"83",
          4099 => x"70",
          4100 => x"f3",
          4101 => x"08",
          4102 => x"59",
          4103 => x"38",
          4104 => x"87",
          4105 => x"f3",
          4106 => x"1a",
          4107 => x"55",
          4108 => x"3f",
          4109 => x"08",
          4110 => x"f3",
          4111 => x"10",
          4112 => x"a4",
          4113 => x"57",
          4114 => x"a0",
          4115 => x"70",
          4116 => x"5e",
          4117 => x"27",
          4118 => x"5d",
          4119 => x"09",
          4120 => x"df",
          4121 => x"ed",
          4122 => x"39",
          4123 => x"52",
          4124 => x"a5",
          4125 => x"f3",
          4126 => x"05",
          4127 => x"06",
          4128 => x"7a",
          4129 => x"38",
          4130 => x"f3",
          4131 => x"bd",
          4132 => x"80",
          4133 => x"83",
          4134 => x"70",
          4135 => x"fc",
          4136 => x"a4",
          4137 => x"70",
          4138 => x"57",
          4139 => x"3f",
          4140 => x"08",
          4141 => x"f3",
          4142 => x"10",
          4143 => x"a4",
          4144 => x"57",
          4145 => x"80",
          4146 => x"38",
          4147 => x"76",
          4148 => x"34",
          4149 => x"75",
          4150 => x"34",
          4151 => x"83",
          4152 => x"ff",
          4153 => x"77",
          4154 => x"f8",
          4155 => x"3d",
          4156 => x"c3",
          4157 => x"84",
          4158 => x"05",
          4159 => x"72",
          4160 => x"8d",
          4161 => x"2e",
          4162 => x"81",
          4163 => x"9e",
          4164 => x"2e",
          4165 => x"87",
          4166 => x"59",
          4167 => x"80",
          4168 => x"80",
          4169 => x"58",
          4170 => x"90",
          4171 => x"f9",
          4172 => x"83",
          4173 => x"75",
          4174 => x"23",
          4175 => x"33",
          4176 => x"71",
          4177 => x"71",
          4178 => x"71",
          4179 => x"56",
          4180 => x"78",
          4181 => x"38",
          4182 => x"84",
          4183 => x"74",
          4184 => x"05",
          4185 => x"74",
          4186 => x"75",
          4187 => x"38",
          4188 => x"33",
          4189 => x"17",
          4190 => x"55",
          4191 => x"0b",
          4192 => x"34",
          4193 => x"81",
          4194 => x"ff",
          4195 => x"ee",
          4196 => x"0d",
          4197 => x"a0",
          4198 => x"f9",
          4199 => x"10",
          4200 => x"f9",
          4201 => x"90",
          4202 => x"05",
          4203 => x"40",
          4204 => x"b0",
          4205 => x"b8",
          4206 => x"81",
          4207 => x"b7",
          4208 => x"81",
          4209 => x"f9",
          4210 => x"83",
          4211 => x"70",
          4212 => x"59",
          4213 => x"57",
          4214 => x"73",
          4215 => x"72",
          4216 => x"29",
          4217 => x"ff",
          4218 => x"ff",
          4219 => x"ff",
          4220 => x"ff",
          4221 => x"81",
          4222 => x"75",
          4223 => x"42",
          4224 => x"5c",
          4225 => x"8f",
          4226 => x"bc",
          4227 => x"31",
          4228 => x"29",
          4229 => x"76",
          4230 => x"7b",
          4231 => x"9c",
          4232 => x"55",
          4233 => x"26",
          4234 => x"80",
          4235 => x"05",
          4236 => x"f9",
          4237 => x"70",
          4238 => x"34",
          4239 => x"a3",
          4240 => x"87",
          4241 => x"70",
          4242 => x"33",
          4243 => x"06",
          4244 => x"33",
          4245 => x"06",
          4246 => x"22",
          4247 => x"5d",
          4248 => x"5e",
          4249 => x"74",
          4250 => x"df",
          4251 => x"ff",
          4252 => x"ff",
          4253 => x"29",
          4254 => x"54",
          4255 => x"fd",
          4256 => x"0b",
          4257 => x"34",
          4258 => x"f9",
          4259 => x"f9",
          4260 => x"98",
          4261 => x"2b",
          4262 => x"2b",
          4263 => x"7a",
          4264 => x"56",
          4265 => x"26",
          4266 => x"fd",
          4267 => x"fc",
          4268 => x"f9",
          4269 => x"81",
          4270 => x"10",
          4271 => x"f9",
          4272 => x"90",
          4273 => x"a3",
          4274 => x"5e",
          4275 => x"56",
          4276 => x"b0",
          4277 => x"84",
          4278 => x"70",
          4279 => x"84",
          4280 => x"70",
          4281 => x"83",
          4282 => x"70",
          4283 => x"06",
          4284 => x"60",
          4285 => x"41",
          4286 => x"40",
          4287 => x"73",
          4288 => x"72",
          4289 => x"70",
          4290 => x"57",
          4291 => x"ff",
          4292 => x"ff",
          4293 => x"29",
          4294 => x"ff",
          4295 => x"ff",
          4296 => x"29",
          4297 => x"5c",
          4298 => x"78",
          4299 => x"77",
          4300 => x"79",
          4301 => x"79",
          4302 => x"58",
          4303 => x"38",
          4304 => x"5c",
          4305 => x"38",
          4306 => x"74",
          4307 => x"29",
          4308 => x"39",
          4309 => x"86",
          4310 => x"54",
          4311 => x"34",
          4312 => x"34",
          4313 => x"98",
          4314 => x"34",
          4315 => x"86",
          4316 => x"56",
          4317 => x"80",
          4318 => x"80",
          4319 => x"ee",
          4320 => x"ff",
          4321 => x"87",
          4322 => x"75",
          4323 => x"34",
          4324 => x"51",
          4325 => x"87",
          4326 => x"70",
          4327 => x"81",
          4328 => x"8c",
          4329 => x"77",
          4330 => x"54",
          4331 => x"34",
          4332 => x"80",
          4333 => x"c0",
          4334 => x"72",
          4335 => x"90",
          4336 => x"70",
          4337 => x"07",
          4338 => x"87",
          4339 => x"34",
          4340 => x"f7",
          4341 => x"53",
          4342 => x"80",
          4343 => x"b8",
          4344 => x"0b",
          4345 => x"0c",
          4346 => x"04",
          4347 => x"33",
          4348 => x"0c",
          4349 => x"0d",
          4350 => x"33",
          4351 => x"b3",
          4352 => x"b7",
          4353 => x"59",
          4354 => x"75",
          4355 => x"da",
          4356 => x"80",
          4357 => x"bd",
          4358 => x"bc",
          4359 => x"29",
          4360 => x"a0",
          4361 => x"f9",
          4362 => x"51",
          4363 => x"7c",
          4364 => x"83",
          4365 => x"83",
          4366 => x"53",
          4367 => x"72",
          4368 => x"c4",
          4369 => x"ba",
          4370 => x"55",
          4371 => x"ba",
          4372 => x"bc",
          4373 => x"70",
          4374 => x"7a",
          4375 => x"55",
          4376 => x"7a",
          4377 => x"38",
          4378 => x"72",
          4379 => x"34",
          4380 => x"22",
          4381 => x"ff",
          4382 => x"fe",
          4383 => x"57",
          4384 => x"82",
          4385 => x"b8",
          4386 => x"71",
          4387 => x"80",
          4388 => x"9f",
          4389 => x"84",
          4390 => x"14",
          4391 => x"e0",
          4392 => x"e0",
          4393 => x"70",
          4394 => x"33",
          4395 => x"05",
          4396 => x"14",
          4397 => x"fd",
          4398 => x"38",
          4399 => x"26",
          4400 => x"f9",
          4401 => x"98",
          4402 => x"55",
          4403 => x"e0",
          4404 => x"73",
          4405 => x"55",
          4406 => x"54",
          4407 => x"27",
          4408 => x"b7",
          4409 => x"05",
          4410 => x"f9",
          4411 => x"57",
          4412 => x"06",
          4413 => x"ff",
          4414 => x"73",
          4415 => x"fd",
          4416 => x"31",
          4417 => x"b8",
          4418 => x"71",
          4419 => x"57",
          4420 => x"a3",
          4421 => x"87",
          4422 => x"79",
          4423 => x"75",
          4424 => x"71",
          4425 => x"5c",
          4426 => x"75",
          4427 => x"38",
          4428 => x"16",
          4429 => x"14",
          4430 => x"b8",
          4431 => x"78",
          4432 => x"5a",
          4433 => x"81",
          4434 => x"77",
          4435 => x"59",
          4436 => x"84",
          4437 => x"84",
          4438 => x"71",
          4439 => x"56",
          4440 => x"72",
          4441 => x"38",
          4442 => x"84",
          4443 => x"8b",
          4444 => x"74",
          4445 => x"34",
          4446 => x"22",
          4447 => x"ff",
          4448 => x"fe",
          4449 => x"57",
          4450 => x"fd",
          4451 => x"80",
          4452 => x"38",
          4453 => x"06",
          4454 => x"f9",
          4455 => x"53",
          4456 => x"09",
          4457 => x"c8",
          4458 => x"31",
          4459 => x"b8",
          4460 => x"71",
          4461 => x"29",
          4462 => x"59",
          4463 => x"27",
          4464 => x"83",
          4465 => x"84",
          4466 => x"74",
          4467 => x"56",
          4468 => x"e0",
          4469 => x"75",
          4470 => x"05",
          4471 => x"13",
          4472 => x"2e",
          4473 => x"a0",
          4474 => x"16",
          4475 => x"70",
          4476 => x"34",
          4477 => x"72",
          4478 => x"f4",
          4479 => x"84",
          4480 => x"55",
          4481 => x"39",
          4482 => x"15",
          4483 => x"b8",
          4484 => x"74",
          4485 => x"ff",
          4486 => x"a9",
          4487 => x"0d",
          4488 => x"05",
          4489 => x"53",
          4490 => x"26",
          4491 => x"10",
          4492 => x"b4",
          4493 => x"08",
          4494 => x"80",
          4495 => x"71",
          4496 => x"71",
          4497 => x"34",
          4498 => x"ba",
          4499 => x"3d",
          4500 => x"0b",
          4501 => x"34",
          4502 => x"33",
          4503 => x"06",
          4504 => x"80",
          4505 => x"ff",
          4506 => x"83",
          4507 => x"80",
          4508 => x"8c",
          4509 => x"0d",
          4510 => x"bc",
          4511 => x"31",
          4512 => x"9f",
          4513 => x"54",
          4514 => x"70",
          4515 => x"34",
          4516 => x"f9",
          4517 => x"05",
          4518 => x"33",
          4519 => x"56",
          4520 => x"25",
          4521 => x"53",
          4522 => x"bc",
          4523 => x"84",
          4524 => x"86",
          4525 => x"83",
          4526 => x"70",
          4527 => x"09",
          4528 => x"72",
          4529 => x"53",
          4530 => x"f9",
          4531 => x"0b",
          4532 => x"0c",
          4533 => x"04",
          4534 => x"33",
          4535 => x"b8",
          4536 => x"11",
          4537 => x"70",
          4538 => x"38",
          4539 => x"83",
          4540 => x"80",
          4541 => x"8c",
          4542 => x"0d",
          4543 => x"83",
          4544 => x"83",
          4545 => x"84",
          4546 => x"ff",
          4547 => x"71",
          4548 => x"b4",
          4549 => x"51",
          4550 => x"bc",
          4551 => x"39",
          4552 => x"02",
          4553 => x"51",
          4554 => x"b3",
          4555 => x"10",
          4556 => x"05",
          4557 => x"04",
          4558 => x"33",
          4559 => x"06",
          4560 => x"80",
          4561 => x"72",
          4562 => x"51",
          4563 => x"71",
          4564 => x"09",
          4565 => x"38",
          4566 => x"83",
          4567 => x"80",
          4568 => x"8c",
          4569 => x"0d",
          4570 => x"b8",
          4571 => x"06",
          4572 => x"70",
          4573 => x"34",
          4574 => x"ba",
          4575 => x"3d",
          4576 => x"f9",
          4577 => x"f0",
          4578 => x"83",
          4579 => x"e8",
          4580 => x"b8",
          4581 => x"06",
          4582 => x"70",
          4583 => x"34",
          4584 => x"f1",
          4585 => x"b8",
          4586 => x"84",
          4587 => x"83",
          4588 => x"83",
          4589 => x"81",
          4590 => x"07",
          4591 => x"f9",
          4592 => x"b4",
          4593 => x"b8",
          4594 => x"51",
          4595 => x"b8",
          4596 => x"39",
          4597 => x"33",
          4598 => x"85",
          4599 => x"83",
          4600 => x"ff",
          4601 => x"f9",
          4602 => x"fb",
          4603 => x"51",
          4604 => x"b8",
          4605 => x"39",
          4606 => x"33",
          4607 => x"81",
          4608 => x"83",
          4609 => x"fe",
          4610 => x"f9",
          4611 => x"f8",
          4612 => x"83",
          4613 => x"fe",
          4614 => x"f9",
          4615 => x"df",
          4616 => x"07",
          4617 => x"f9",
          4618 => x"cc",
          4619 => x"b8",
          4620 => x"06",
          4621 => x"70",
          4622 => x"34",
          4623 => x"83",
          4624 => x"81",
          4625 => x"e0",
          4626 => x"83",
          4627 => x"fe",
          4628 => x"f9",
          4629 => x"cf",
          4630 => x"07",
          4631 => x"f9",
          4632 => x"94",
          4633 => x"b8",
          4634 => x"06",
          4635 => x"70",
          4636 => x"34",
          4637 => x"83",
          4638 => x"81",
          4639 => x"70",
          4640 => x"34",
          4641 => x"83",
          4642 => x"81",
          4643 => x"07",
          4644 => x"f9",
          4645 => x"e0",
          4646 => x"0d",
          4647 => x"33",
          4648 => x"80",
          4649 => x"83",
          4650 => x"83",
          4651 => x"83",
          4652 => x"84",
          4653 => x"43",
          4654 => x"5b",
          4655 => x"2e",
          4656 => x"78",
          4657 => x"38",
          4658 => x"81",
          4659 => x"84",
          4660 => x"80",
          4661 => x"84",
          4662 => x"f9",
          4663 => x"83",
          4664 => x"7c",
          4665 => x"34",
          4666 => x"04",
          4667 => x"09",
          4668 => x"38",
          4669 => x"b8",
          4670 => x"0b",
          4671 => x"34",
          4672 => x"f9",
          4673 => x"0b",
          4674 => x"34",
          4675 => x"f9",
          4676 => x"58",
          4677 => x"33",
          4678 => x"ff",
          4679 => x"b7",
          4680 => x"7b",
          4681 => x"7a",
          4682 => x"c4",
          4683 => x"db",
          4684 => x"b8",
          4685 => x"0b",
          4686 => x"34",
          4687 => x"bc",
          4688 => x"f9",
          4689 => x"83",
          4690 => x"8f",
          4691 => x"80",
          4692 => x"82",
          4693 => x"84",
          4694 => x"80",
          4695 => x"bc",
          4696 => x"83",
          4697 => x"80",
          4698 => x"ba",
          4699 => x"8f",
          4700 => x"b9",
          4701 => x"84",
          4702 => x"56",
          4703 => x"54",
          4704 => x"52",
          4705 => x"51",
          4706 => x"3f",
          4707 => x"b9",
          4708 => x"5a",
          4709 => x"a5",
          4710 => x"84",
          4711 => x"70",
          4712 => x"83",
          4713 => x"ff",
          4714 => x"81",
          4715 => x"ff",
          4716 => x"8d",
          4717 => x"59",
          4718 => x"dd",
          4719 => x"ec",
          4720 => x"c7",
          4721 => x"b8",
          4722 => x"0b",
          4723 => x"34",
          4724 => x"bc",
          4725 => x"f9",
          4726 => x"83",
          4727 => x"8f",
          4728 => x"80",
          4729 => x"82",
          4730 => x"84",
          4731 => x"81",
          4732 => x"bc",
          4733 => x"83",
          4734 => x"81",
          4735 => x"ba",
          4736 => x"f0",
          4737 => x"a3",
          4738 => x"8c",
          4739 => x"e3",
          4740 => x"ff",
          4741 => x"59",
          4742 => x"51",
          4743 => x"3f",
          4744 => x"8c",
          4745 => x"a6",
          4746 => x"f0",
          4747 => x"83",
          4748 => x"fe",
          4749 => x"81",
          4750 => x"ff",
          4751 => x"d8",
          4752 => x"0d",
          4753 => x"05",
          4754 => x"84",
          4755 => x"83",
          4756 => x"83",
          4757 => x"72",
          4758 => x"87",
          4759 => x"11",
          4760 => x"22",
          4761 => x"5c",
          4762 => x"05",
          4763 => x"ff",
          4764 => x"92",
          4765 => x"51",
          4766 => x"72",
          4767 => x"e9",
          4768 => x"2e",
          4769 => x"75",
          4770 => x"b9",
          4771 => x"2e",
          4772 => x"75",
          4773 => x"d5",
          4774 => x"80",
          4775 => x"bc",
          4776 => x"bd",
          4777 => x"29",
          4778 => x"54",
          4779 => x"16",
          4780 => x"a0",
          4781 => x"84",
          4782 => x"83",
          4783 => x"83",
          4784 => x"72",
          4785 => x"5a",
          4786 => x"75",
          4787 => x"18",
          4788 => x"bc",
          4789 => x"29",
          4790 => x"83",
          4791 => x"87",
          4792 => x"18",
          4793 => x"80",
          4794 => x"ff",
          4795 => x"ba",
          4796 => x"bd",
          4797 => x"29",
          4798 => x"57",
          4799 => x"f9",
          4800 => x"98",
          4801 => x"81",
          4802 => x"ff",
          4803 => x"73",
          4804 => x"99",
          4805 => x"81",
          4806 => x"81",
          4807 => x"17",
          4808 => x"f9",
          4809 => x"b8",
          4810 => x"72",
          4811 => x"38",
          4812 => x"33",
          4813 => x"2e",
          4814 => x"80",
          4815 => x"8c",
          4816 => x"0d",
          4817 => x"2e",
          4818 => x"8d",
          4819 => x"38",
          4820 => x"09",
          4821 => x"c1",
          4822 => x"81",
          4823 => x"3f",
          4824 => x"f9",
          4825 => x"be",
          4826 => x"be",
          4827 => x"84",
          4828 => x"33",
          4829 => x"89",
          4830 => x"06",
          4831 => x"80",
          4832 => x"a0",
          4833 => x"3f",
          4834 => x"81",
          4835 => x"54",
          4836 => x"ff",
          4837 => x"52",
          4838 => x"a5",
          4839 => x"70",
          4840 => x"54",
          4841 => x"27",
          4842 => x"fa",
          4843 => x"f9",
          4844 => x"f2",
          4845 => x"83",
          4846 => x"3f",
          4847 => x"ba",
          4848 => x"3d",
          4849 => x"80",
          4850 => x"81",
          4851 => x"38",
          4852 => x"33",
          4853 => x"06",
          4854 => x"53",
          4855 => x"73",
          4856 => x"f9",
          4857 => x"52",
          4858 => x"d5",
          4859 => x"bd",
          4860 => x"ff",
          4861 => x"05",
          4862 => x"a5",
          4863 => x"72",
          4864 => x"34",
          4865 => x"80",
          4866 => x"bd",
          4867 => x"81",
          4868 => x"3f",
          4869 => x"80",
          4870 => x"ef",
          4871 => x"86",
          4872 => x"0d",
          4873 => x"05",
          4874 => x"88",
          4875 => x"75",
          4876 => x"b8",
          4877 => x"2e",
          4878 => x"78",
          4879 => x"b5",
          4880 => x"24",
          4881 => x"78",
          4882 => x"b9",
          4883 => x"2e",
          4884 => x"84",
          4885 => x"83",
          4886 => x"83",
          4887 => x"72",
          4888 => x"58",
          4889 => x"b8",
          4890 => x"87",
          4891 => x"17",
          4892 => x"80",
          4893 => x"bd",
          4894 => x"ba",
          4895 => x"29",
          4896 => x"42",
          4897 => x"f9",
          4898 => x"83",
          4899 => x"60",
          4900 => x"05",
          4901 => x"f9",
          4902 => x"87",
          4903 => x"05",
          4904 => x"80",
          4905 => x"ff",
          4906 => x"ba",
          4907 => x"bd",
          4908 => x"29",
          4909 => x"5d",
          4910 => x"f9",
          4911 => x"98",
          4912 => x"81",
          4913 => x"ff",
          4914 => x"76",
          4915 => x"b8",
          4916 => x"81",
          4917 => x"86",
          4918 => x"19",
          4919 => x"f9",
          4920 => x"0b",
          4921 => x"0c",
          4922 => x"04",
          4923 => x"84",
          4924 => x"79",
          4925 => x"38",
          4926 => x"9b",
          4927 => x"80",
          4928 => x"cc",
          4929 => x"84",
          4930 => x"84",
          4931 => x"83",
          4932 => x"83",
          4933 => x"72",
          4934 => x"5e",
          4935 => x"b8",
          4936 => x"87",
          4937 => x"1d",
          4938 => x"80",
          4939 => x"bd",
          4940 => x"ba",
          4941 => x"29",
          4942 => x"59",
          4943 => x"f9",
          4944 => x"83",
          4945 => x"76",
          4946 => x"5b",
          4947 => x"b8",
          4948 => x"b0",
          4949 => x"84",
          4950 => x"70",
          4951 => x"83",
          4952 => x"83",
          4953 => x"72",
          4954 => x"44",
          4955 => x"59",
          4956 => x"33",
          4957 => x"de",
          4958 => x"1f",
          4959 => x"ff",
          4960 => x"77",
          4961 => x"38",
          4962 => x"bd",
          4963 => x"84",
          4964 => x"9c",
          4965 => x"78",
          4966 => x"b7",
          4967 => x"24",
          4968 => x"78",
          4969 => x"81",
          4970 => x"38",
          4971 => x"f9",
          4972 => x"0b",
          4973 => x"0c",
          4974 => x"04",
          4975 => x"82",
          4976 => x"19",
          4977 => x"26",
          4978 => x"84",
          4979 => x"81",
          4980 => x"77",
          4981 => x"34",
          4982 => x"90",
          4983 => x"81",
          4984 => x"80",
          4985 => x"90",
          4986 => x"0b",
          4987 => x"0c",
          4988 => x"04",
          4989 => x"fd",
          4990 => x"0b",
          4991 => x"0c",
          4992 => x"33",
          4993 => x"33",
          4994 => x"33",
          4995 => x"05",
          4996 => x"84",
          4997 => x"33",
          4998 => x"80",
          4999 => x"b8",
          5000 => x"f9",
          5001 => x"f9",
          5002 => x"71",
          5003 => x"5f",
          5004 => x"83",
          5005 => x"34",
          5006 => x"33",
          5007 => x"19",
          5008 => x"f9",
          5009 => x"a3",
          5010 => x"34",
          5011 => x"33",
          5012 => x"06",
          5013 => x"22",
          5014 => x"33",
          5015 => x"11",
          5016 => x"58",
          5017 => x"b8",
          5018 => x"98",
          5019 => x"81",
          5020 => x"89",
          5021 => x"81",
          5022 => x"3f",
          5023 => x"f9",
          5024 => x"ae",
          5025 => x"80",
          5026 => x"bd",
          5027 => x"ff",
          5028 => x"bc",
          5029 => x"29",
          5030 => x"a0",
          5031 => x"f9",
          5032 => x"51",
          5033 => x"29",
          5034 => x"ff",
          5035 => x"f8",
          5036 => x"51",
          5037 => x"75",
          5038 => x"a4",
          5039 => x"ff",
          5040 => x"57",
          5041 => x"95",
          5042 => x"75",
          5043 => x"34",
          5044 => x"80",
          5045 => x"8c",
          5046 => x"84",
          5047 => x"80",
          5048 => x"8e",
          5049 => x"84",
          5050 => x"81",
          5051 => x"88",
          5052 => x"84",
          5053 => x"9c",
          5054 => x"83",
          5055 => x"84",
          5056 => x"83",
          5057 => x"84",
          5058 => x"83",
          5059 => x"84",
          5060 => x"80",
          5061 => x"88",
          5062 => x"84",
          5063 => x"9c",
          5064 => x"78",
          5065 => x"09",
          5066 => x"a7",
          5067 => x"bc",
          5068 => x"80",
          5069 => x"ff",
          5070 => x"bd",
          5071 => x"ff",
          5072 => x"29",
          5073 => x"a0",
          5074 => x"f9",
          5075 => x"40",
          5076 => x"05",
          5077 => x"ff",
          5078 => x"92",
          5079 => x"43",
          5080 => x"5c",
          5081 => x"85",
          5082 => x"81",
          5083 => x"1a",
          5084 => x"83",
          5085 => x"76",
          5086 => x"34",
          5087 => x"06",
          5088 => x"06",
          5089 => x"06",
          5090 => x"05",
          5091 => x"84",
          5092 => x"87",
          5093 => x"1e",
          5094 => x"80",
          5095 => x"bd",
          5096 => x"ba",
          5097 => x"29",
          5098 => x"42",
          5099 => x"83",
          5100 => x"34",
          5101 => x"33",
          5102 => x"62",
          5103 => x"83",
          5104 => x"87",
          5105 => x"1a",
          5106 => x"80",
          5107 => x"ff",
          5108 => x"ba",
          5109 => x"bd",
          5110 => x"29",
          5111 => x"5a",
          5112 => x"f9",
          5113 => x"84",
          5114 => x"34",
          5115 => x"81",
          5116 => x"58",
          5117 => x"95",
          5118 => x"b8",
          5119 => x"79",
          5120 => x"ff",
          5121 => x"83",
          5122 => x"83",
          5123 => x"70",
          5124 => x"58",
          5125 => x"fd",
          5126 => x"bb",
          5127 => x"38",
          5128 => x"83",
          5129 => x"bf",
          5130 => x"38",
          5131 => x"33",
          5132 => x"f9",
          5133 => x"19",
          5134 => x"26",
          5135 => x"75",
          5136 => x"c6",
          5137 => x"77",
          5138 => x"0b",
          5139 => x"34",
          5140 => x"51",
          5141 => x"80",
          5142 => x"8c",
          5143 => x"0d",
          5144 => x"bc",
          5145 => x"80",
          5146 => x"ff",
          5147 => x"bd",
          5148 => x"ff",
          5149 => x"29",
          5150 => x"a0",
          5151 => x"f9",
          5152 => x"41",
          5153 => x"05",
          5154 => x"ff",
          5155 => x"92",
          5156 => x"45",
          5157 => x"5b",
          5158 => x"82",
          5159 => x"5c",
          5160 => x"06",
          5161 => x"06",
          5162 => x"06",
          5163 => x"05",
          5164 => x"84",
          5165 => x"87",
          5166 => x"1b",
          5167 => x"80",
          5168 => x"bd",
          5169 => x"ba",
          5170 => x"29",
          5171 => x"5e",
          5172 => x"83",
          5173 => x"34",
          5174 => x"33",
          5175 => x"1e",
          5176 => x"f9",
          5177 => x"a3",
          5178 => x"34",
          5179 => x"33",
          5180 => x"06",
          5181 => x"22",
          5182 => x"33",
          5183 => x"11",
          5184 => x"40",
          5185 => x"b8",
          5186 => x"de",
          5187 => x"81",
          5188 => x"ff",
          5189 => x"7e",
          5190 => x"ac",
          5191 => x"81",
          5192 => x"92",
          5193 => x"19",
          5194 => x"f9",
          5195 => x"1c",
          5196 => x"06",
          5197 => x"83",
          5198 => x"38",
          5199 => x"33",
          5200 => x"33",
          5201 => x"33",
          5202 => x"06",
          5203 => x"06",
          5204 => x"06",
          5205 => x"05",
          5206 => x"5b",
          5207 => x"b8",
          5208 => x"a3",
          5209 => x"34",
          5210 => x"33",
          5211 => x"33",
          5212 => x"22",
          5213 => x"12",
          5214 => x"56",
          5215 => x"f9",
          5216 => x"83",
          5217 => x"76",
          5218 => x"5a",
          5219 => x"b8",
          5220 => x"b0",
          5221 => x"84",
          5222 => x"70",
          5223 => x"83",
          5224 => x"83",
          5225 => x"72",
          5226 => x"5b",
          5227 => x"59",
          5228 => x"33",
          5229 => x"18",
          5230 => x"05",
          5231 => x"06",
          5232 => x"7f",
          5233 => x"38",
          5234 => x"bd",
          5235 => x"39",
          5236 => x"b9",
          5237 => x"0b",
          5238 => x"0c",
          5239 => x"04",
          5240 => x"17",
          5241 => x"b8",
          5242 => x"7a",
          5243 => x"bd",
          5244 => x"ff",
          5245 => x"05",
          5246 => x"39",
          5247 => x"b9",
          5248 => x"0b",
          5249 => x"0c",
          5250 => x"04",
          5251 => x"17",
          5252 => x"b8",
          5253 => x"7c",
          5254 => x"bc",
          5255 => x"80",
          5256 => x"bd",
          5257 => x"5b",
          5258 => x"f4",
          5259 => x"90",
          5260 => x"dc",
          5261 => x"05",
          5262 => x"cd",
          5263 => x"8c",
          5264 => x"fb",
          5265 => x"b9",
          5266 => x"11",
          5267 => x"84",
          5268 => x"79",
          5269 => x"06",
          5270 => x"ca",
          5271 => x"84",
          5272 => x"23",
          5273 => x"83",
          5274 => x"33",
          5275 => x"88",
          5276 => x"34",
          5277 => x"33",
          5278 => x"33",
          5279 => x"33",
          5280 => x"f9",
          5281 => x"b8",
          5282 => x"f9",
          5283 => x"f9",
          5284 => x"72",
          5285 => x"5d",
          5286 => x"88",
          5287 => x"87",
          5288 => x"05",
          5289 => x"80",
          5290 => x"bd",
          5291 => x"ba",
          5292 => x"29",
          5293 => x"5b",
          5294 => x"f9",
          5295 => x"83",
          5296 => x"76",
          5297 => x"41",
          5298 => x"b8",
          5299 => x"a3",
          5300 => x"34",
          5301 => x"33",
          5302 => x"06",
          5303 => x"22",
          5304 => x"33",
          5305 => x"11",
          5306 => x"42",
          5307 => x"b8",
          5308 => x"de",
          5309 => x"1c",
          5310 => x"06",
          5311 => x"7b",
          5312 => x"38",
          5313 => x"33",
          5314 => x"e2",
          5315 => x"56",
          5316 => x"bd",
          5317 => x"84",
          5318 => x"84",
          5319 => x"40",
          5320 => x"f3",
          5321 => x"b8",
          5322 => x"75",
          5323 => x"78",
          5324 => x"ea",
          5325 => x"0b",
          5326 => x"0c",
          5327 => x"04",
          5328 => x"33",
          5329 => x"34",
          5330 => x"33",
          5331 => x"34",
          5332 => x"33",
          5333 => x"f9",
          5334 => x"b9",
          5335 => x"bc",
          5336 => x"f4",
          5337 => x"bd",
          5338 => x"f5",
          5339 => x"bb",
          5340 => x"f6",
          5341 => x"39",
          5342 => x"33",
          5343 => x"2e",
          5344 => x"84",
          5345 => x"5d",
          5346 => x"09",
          5347 => x"85",
          5348 => x"bd",
          5349 => x"55",
          5350 => x"33",
          5351 => x"9b",
          5352 => x"8c",
          5353 => x"70",
          5354 => x"ed",
          5355 => x"51",
          5356 => x"3f",
          5357 => x"08",
          5358 => x"83",
          5359 => x"57",
          5360 => x"60",
          5361 => x"cd",
          5362 => x"83",
          5363 => x"fe",
          5364 => x"fe",
          5365 => x"0b",
          5366 => x"33",
          5367 => x"81",
          5368 => x"77",
          5369 => x"ad",
          5370 => x"84",
          5371 => x"81",
          5372 => x"41",
          5373 => x"8a",
          5374 => x"10",
          5375 => x"ec",
          5376 => x"08",
          5377 => x"8d",
          5378 => x"80",
          5379 => x"38",
          5380 => x"33",
          5381 => x"33",
          5382 => x"70",
          5383 => x"2c",
          5384 => x"42",
          5385 => x"75",
          5386 => x"34",
          5387 => x"84",
          5388 => x"56",
          5389 => x"8e",
          5390 => x"b9",
          5391 => x"05",
          5392 => x"06",
          5393 => x"33",
          5394 => x"75",
          5395 => x"c5",
          5396 => x"f9",
          5397 => x"bd",
          5398 => x"83",
          5399 => x"83",
          5400 => x"70",
          5401 => x"5d",
          5402 => x"2e",
          5403 => x"ff",
          5404 => x"83",
          5405 => x"fd",
          5406 => x"0b",
          5407 => x"34",
          5408 => x"33",
          5409 => x"33",
          5410 => x"57",
          5411 => x"fd",
          5412 => x"17",
          5413 => x"f9",
          5414 => x"f9",
          5415 => x"8d",
          5416 => x"80",
          5417 => x"38",
          5418 => x"33",
          5419 => x"33",
          5420 => x"70",
          5421 => x"2c",
          5422 => x"41",
          5423 => x"75",
          5424 => x"34",
          5425 => x"84",
          5426 => x"5b",
          5427 => x"fc",
          5428 => x"b9",
          5429 => x"60",
          5430 => x"81",
          5431 => x"38",
          5432 => x"33",
          5433 => x"33",
          5434 => x"33",
          5435 => x"12",
          5436 => x"80",
          5437 => x"ba",
          5438 => x"5a",
          5439 => x"29",
          5440 => x"ff",
          5441 => x"f8",
          5442 => x"ff",
          5443 => x"42",
          5444 => x"7e",
          5445 => x"2e",
          5446 => x"80",
          5447 => x"91",
          5448 => x"39",
          5449 => x"33",
          5450 => x"2e",
          5451 => x"84",
          5452 => x"58",
          5453 => x"09",
          5454 => x"d9",
          5455 => x"83",
          5456 => x"fb",
          5457 => x"b9",
          5458 => x"75",
          5459 => x"be",
          5460 => x"e1",
          5461 => x"bd",
          5462 => x"05",
          5463 => x"33",
          5464 => x"5e",
          5465 => x"25",
          5466 => x"57",
          5467 => x"bd",
          5468 => x"39",
          5469 => x"33",
          5470 => x"2e",
          5471 => x"84",
          5472 => x"83",
          5473 => x"42",
          5474 => x"b7",
          5475 => x"11",
          5476 => x"75",
          5477 => x"38",
          5478 => x"83",
          5479 => x"fa",
          5480 => x"e4",
          5481 => x"e8",
          5482 => x"0b",
          5483 => x"33",
          5484 => x"76",
          5485 => x"38",
          5486 => x"b9",
          5487 => x"22",
          5488 => x"e3",
          5489 => x"e8",
          5490 => x"17",
          5491 => x"06",
          5492 => x"33",
          5493 => x"da",
          5494 => x"84",
          5495 => x"5f",
          5496 => x"2e",
          5497 => x"b9",
          5498 => x"75",
          5499 => x"38",
          5500 => x"52",
          5501 => x"06",
          5502 => x"3f",
          5503 => x"84",
          5504 => x"57",
          5505 => x"8e",
          5506 => x"b9",
          5507 => x"05",
          5508 => x"06",
          5509 => x"33",
          5510 => x"81",
          5511 => x"b7",
          5512 => x"81",
          5513 => x"11",
          5514 => x"5b",
          5515 => x"77",
          5516 => x"38",
          5517 => x"83",
          5518 => x"76",
          5519 => x"ff",
          5520 => x"77",
          5521 => x"38",
          5522 => x"83",
          5523 => x"84",
          5524 => x"ff",
          5525 => x"7a",
          5526 => x"b4",
          5527 => x"75",
          5528 => x"34",
          5529 => x"84",
          5530 => x"5f",
          5531 => x"8a",
          5532 => x"b9",
          5533 => x"b7",
          5534 => x"5b",
          5535 => x"f9",
          5536 => x"f9",
          5537 => x"b8",
          5538 => x"81",
          5539 => x"f9",
          5540 => x"74",
          5541 => x"a3",
          5542 => x"83",
          5543 => x"5f",
          5544 => x"29",
          5545 => x"ff",
          5546 => x"f8",
          5547 => x"52",
          5548 => x"5d",
          5549 => x"84",
          5550 => x"83",
          5551 => x"70",
          5552 => x"57",
          5553 => x"8e",
          5554 => x"b7",
          5555 => x"76",
          5556 => x"d6",
          5557 => x"56",
          5558 => x"ba",
          5559 => x"ff",
          5560 => x"31",
          5561 => x"60",
          5562 => x"38",
          5563 => x"33",
          5564 => x"27",
          5565 => x"ff",
          5566 => x"83",
          5567 => x"7e",
          5568 => x"83",
          5569 => x"57",
          5570 => x"76",
          5571 => x"38",
          5572 => x"81",
          5573 => x"ff",
          5574 => x"29",
          5575 => x"79",
          5576 => x"a0",
          5577 => x"a3",
          5578 => x"81",
          5579 => x"81",
          5580 => x"71",
          5581 => x"58",
          5582 => x"7f",
          5583 => x"38",
          5584 => x"1a",
          5585 => x"17",
          5586 => x"b8",
          5587 => x"7b",
          5588 => x"5d",
          5589 => x"81",
          5590 => x"7c",
          5591 => x"5e",
          5592 => x"84",
          5593 => x"84",
          5594 => x"71",
          5595 => x"43",
          5596 => x"77",
          5597 => x"9d",
          5598 => x"17",
          5599 => x"b8",
          5600 => x"7b",
          5601 => x"5d",
          5602 => x"81",
          5603 => x"7c",
          5604 => x"5e",
          5605 => x"84",
          5606 => x"84",
          5607 => x"71",
          5608 => x"43",
          5609 => x"7f",
          5610 => x"99",
          5611 => x"39",
          5612 => x"33",
          5613 => x"2e",
          5614 => x"80",
          5615 => x"e1",
          5616 => x"b1",
          5617 => x"39",
          5618 => x"b8",
          5619 => x"11",
          5620 => x"33",
          5621 => x"58",
          5622 => x"94",
          5623 => x"e0",
          5624 => x"78",
          5625 => x"06",
          5626 => x"83",
          5627 => x"58",
          5628 => x"06",
          5629 => x"33",
          5630 => x"5c",
          5631 => x"81",
          5632 => x"b7",
          5633 => x"7a",
          5634 => x"89",
          5635 => x"ff",
          5636 => x"76",
          5637 => x"38",
          5638 => x"61",
          5639 => x"57",
          5640 => x"38",
          5641 => x"1b",
          5642 => x"62",
          5643 => x"a0",
          5644 => x"1f",
          5645 => x"a3",
          5646 => x"79",
          5647 => x"51",
          5648 => x"ac",
          5649 => x"06",
          5650 => x"a4",
          5651 => x"b8",
          5652 => x"2b",
          5653 => x"07",
          5654 => x"07",
          5655 => x"7f",
          5656 => x"57",
          5657 => x"9e",
          5658 => x"70",
          5659 => x"0c",
          5660 => x"84",
          5661 => x"79",
          5662 => x"38",
          5663 => x"33",
          5664 => x"33",
          5665 => x"81",
          5666 => x"81",
          5667 => x"f9",
          5668 => x"73",
          5669 => x"59",
          5670 => x"77",
          5671 => x"38",
          5672 => x"1b",
          5673 => x"62",
          5674 => x"75",
          5675 => x"57",
          5676 => x"f4",
          5677 => x"f9",
          5678 => x"98",
          5679 => x"5a",
          5680 => x"e0",
          5681 => x"78",
          5682 => x"5a",
          5683 => x"57",
          5684 => x"f4",
          5685 => x"0b",
          5686 => x"34",
          5687 => x"81",
          5688 => x"81",
          5689 => x"77",
          5690 => x"f4",
          5691 => x"1f",
          5692 => x"06",
          5693 => x"8a",
          5694 => x"b8",
          5695 => x"f0",
          5696 => x"2b",
          5697 => x"71",
          5698 => x"58",
          5699 => x"80",
          5700 => x"81",
          5701 => x"80",
          5702 => x"f9",
          5703 => x"18",
          5704 => x"06",
          5705 => x"b6",
          5706 => x"be",
          5707 => x"84",
          5708 => x"33",
          5709 => x"f9",
          5710 => x"b8",
          5711 => x"f9",
          5712 => x"b7",
          5713 => x"5c",
          5714 => x"ee",
          5715 => x"b8",
          5716 => x"56",
          5717 => x"b8",
          5718 => x"70",
          5719 => x"59",
          5720 => x"39",
          5721 => x"33",
          5722 => x"85",
          5723 => x"83",
          5724 => x"e5",
          5725 => x"b8",
          5726 => x"06",
          5727 => x"75",
          5728 => x"34",
          5729 => x"f9",
          5730 => x"f9",
          5731 => x"56",
          5732 => x"b8",
          5733 => x"83",
          5734 => x"81",
          5735 => x"07",
          5736 => x"f9",
          5737 => x"b1",
          5738 => x"0b",
          5739 => x"34",
          5740 => x"81",
          5741 => x"56",
          5742 => x"83",
          5743 => x"81",
          5744 => x"75",
          5745 => x"34",
          5746 => x"83",
          5747 => x"81",
          5748 => x"07",
          5749 => x"f9",
          5750 => x"fd",
          5751 => x"b8",
          5752 => x"06",
          5753 => x"56",
          5754 => x"b8",
          5755 => x"39",
          5756 => x"33",
          5757 => x"80",
          5758 => x"75",
          5759 => x"34",
          5760 => x"83",
          5761 => x"81",
          5762 => x"07",
          5763 => x"f9",
          5764 => x"c5",
          5765 => x"b8",
          5766 => x"06",
          5767 => x"75",
          5768 => x"34",
          5769 => x"83",
          5770 => x"81",
          5771 => x"07",
          5772 => x"f9",
          5773 => x"a1",
          5774 => x"b8",
          5775 => x"06",
          5776 => x"75",
          5777 => x"34",
          5778 => x"83",
          5779 => x"81",
          5780 => x"75",
          5781 => x"34",
          5782 => x"83",
          5783 => x"80",
          5784 => x"75",
          5785 => x"34",
          5786 => x"83",
          5787 => x"80",
          5788 => x"75",
          5789 => x"34",
          5790 => x"83",
          5791 => x"81",
          5792 => x"d0",
          5793 => x"83",
          5794 => x"fd",
          5795 => x"f9",
          5796 => x"bf",
          5797 => x"56",
          5798 => x"b8",
          5799 => x"39",
          5800 => x"f9",
          5801 => x"52",
          5802 => x"c9",
          5803 => x"39",
          5804 => x"33",
          5805 => x"34",
          5806 => x"33",
          5807 => x"34",
          5808 => x"33",
          5809 => x"f9",
          5810 => x"0b",
          5811 => x"0c",
          5812 => x"81",
          5813 => x"8f",
          5814 => x"84",
          5815 => x"9c",
          5816 => x"77",
          5817 => x"34",
          5818 => x"33",
          5819 => x"06",
          5820 => x"56",
          5821 => x"84",
          5822 => x"9c",
          5823 => x"53",
          5824 => x"fe",
          5825 => x"84",
          5826 => x"a1",
          5827 => x"8c",
          5828 => x"88",
          5829 => x"84",
          5830 => x"80",
          5831 => x"8c",
          5832 => x"0d",
          5833 => x"f9",
          5834 => x"e9",
          5835 => x"8d",
          5836 => x"5c",
          5837 => x"b9",
          5838 => x"10",
          5839 => x"5d",
          5840 => x"05",
          5841 => x"e0",
          5842 => x"0b",
          5843 => x"34",
          5844 => x"0b",
          5845 => x"34",
          5846 => x"51",
          5847 => x"83",
          5848 => x"70",
          5849 => x"58",
          5850 => x"e6",
          5851 => x"0b",
          5852 => x"34",
          5853 => x"51",
          5854 => x"ef",
          5855 => x"51",
          5856 => x"3f",
          5857 => x"83",
          5858 => x"ff",
          5859 => x"70",
          5860 => x"06",
          5861 => x"f2",
          5862 => x"52",
          5863 => x"39",
          5864 => x"33",
          5865 => x"27",
          5866 => x"75",
          5867 => x"34",
          5868 => x"83",
          5869 => x"ff",
          5870 => x"70",
          5871 => x"06",
          5872 => x"f0",
          5873 => x"f9",
          5874 => x"05",
          5875 => x"33",
          5876 => x"59",
          5877 => x"25",
          5878 => x"75",
          5879 => x"39",
          5880 => x"33",
          5881 => x"06",
          5882 => x"77",
          5883 => x"38",
          5884 => x"33",
          5885 => x"33",
          5886 => x"06",
          5887 => x"33",
          5888 => x"11",
          5889 => x"80",
          5890 => x"ba",
          5891 => x"71",
          5892 => x"70",
          5893 => x"06",
          5894 => x"33",
          5895 => x"42",
          5896 => x"81",
          5897 => x"38",
          5898 => x"ff",
          5899 => x"5c",
          5900 => x"24",
          5901 => x"84",
          5902 => x"56",
          5903 => x"83",
          5904 => x"16",
          5905 => x"f9",
          5906 => x"81",
          5907 => x"11",
          5908 => x"76",
          5909 => x"38",
          5910 => x"33",
          5911 => x"27",
          5912 => x"ff",
          5913 => x"83",
          5914 => x"7b",
          5915 => x"83",
          5916 => x"57",
          5917 => x"76",
          5918 => x"38",
          5919 => x"81",
          5920 => x"ff",
          5921 => x"29",
          5922 => x"79",
          5923 => x"a0",
          5924 => x"a3",
          5925 => x"81",
          5926 => x"81",
          5927 => x"71",
          5928 => x"42",
          5929 => x"7e",
          5930 => x"38",
          5931 => x"1a",
          5932 => x"17",
          5933 => x"b8",
          5934 => x"7b",
          5935 => x"5d",
          5936 => x"81",
          5937 => x"7d",
          5938 => x"5f",
          5939 => x"84",
          5940 => x"84",
          5941 => x"71",
          5942 => x"59",
          5943 => x"77",
          5944 => x"b1",
          5945 => x"17",
          5946 => x"b8",
          5947 => x"7b",
          5948 => x"5d",
          5949 => x"81",
          5950 => x"7d",
          5951 => x"5f",
          5952 => x"84",
          5953 => x"84",
          5954 => x"71",
          5955 => x"59",
          5956 => x"75",
          5957 => x"99",
          5958 => x"39",
          5959 => x"17",
          5960 => x"b8",
          5961 => x"7b",
          5962 => x"bc",
          5963 => x"80",
          5964 => x"ba",
          5965 => x"ff",
          5966 => x"5f",
          5967 => x"39",
          5968 => x"38",
          5969 => x"33",
          5970 => x"06",
          5971 => x"42",
          5972 => x"27",
          5973 => x"5a",
          5974 => x"ba",
          5975 => x"ff",
          5976 => x"58",
          5977 => x"27",
          5978 => x"57",
          5979 => x"bc",
          5980 => x"80",
          5981 => x"ff",
          5982 => x"52",
          5983 => x"78",
          5984 => x"38",
          5985 => x"83",
          5986 => x"eb",
          5987 => x"f9",
          5988 => x"05",
          5989 => x"33",
          5990 => x"40",
          5991 => x"25",
          5992 => x"75",
          5993 => x"39",
          5994 => x"09",
          5995 => x"c0",
          5996 => x"bd",
          5997 => x"ff",
          5998 => x"bc",
          5999 => x"5d",
          6000 => x"ff",
          6001 => x"06",
          6002 => x"f6",
          6003 => x"1d",
          6004 => x"f9",
          6005 => x"93",
          6006 => x"56",
          6007 => x"ba",
          6008 => x"39",
          6009 => x"56",
          6010 => x"bc",
          6011 => x"39",
          6012 => x"56",
          6013 => x"f5",
          6014 => x"76",
          6015 => x"58",
          6016 => x"b8",
          6017 => x"81",
          6018 => x"75",
          6019 => x"ec",
          6020 => x"70",
          6021 => x"34",
          6022 => x"33",
          6023 => x"05",
          6024 => x"76",
          6025 => x"f4",
          6026 => x"7b",
          6027 => x"83",
          6028 => x"f1",
          6029 => x"0b",
          6030 => x"34",
          6031 => x"7e",
          6032 => x"23",
          6033 => x"80",
          6034 => x"ba",
          6035 => x"39",
          6036 => x"f9",
          6037 => x"a7",
          6038 => x"be",
          6039 => x"84",
          6040 => x"33",
          6041 => x"0b",
          6042 => x"34",
          6043 => x"fd",
          6044 => x"97",
          6045 => x"b8",
          6046 => x"54",
          6047 => x"90",
          6048 => x"db",
          6049 => x"0b",
          6050 => x"0c",
          6051 => x"04",
          6052 => x"51",
          6053 => x"80",
          6054 => x"8c",
          6055 => x"0d",
          6056 => x"0d",
          6057 => x"33",
          6058 => x"83",
          6059 => x"70",
          6060 => x"83",
          6061 => x"33",
          6062 => x"59",
          6063 => x"80",
          6064 => x"14",
          6065 => x"f8",
          6066 => x"59",
          6067 => x"8c",
          6068 => x"0d",
          6069 => x"ec",
          6070 => x"53",
          6071 => x"91",
          6072 => x"32",
          6073 => x"07",
          6074 => x"9f",
          6075 => x"5e",
          6076 => x"f7",
          6077 => x"59",
          6078 => x"81",
          6079 => x"06",
          6080 => x"54",
          6081 => x"70",
          6082 => x"25",
          6083 => x"5c",
          6084 => x"2e",
          6085 => x"84",
          6086 => x"83",
          6087 => x"83",
          6088 => x"72",
          6089 => x"87",
          6090 => x"05",
          6091 => x"22",
          6092 => x"71",
          6093 => x"70",
          6094 => x"06",
          6095 => x"33",
          6096 => x"58",
          6097 => x"83",
          6098 => x"f0",
          6099 => x"ee",
          6100 => x"80",
          6101 => x"98",
          6102 => x"c0",
          6103 => x"56",
          6104 => x"f6",
          6105 => x"80",
          6106 => x"76",
          6107 => x"15",
          6108 => x"70",
          6109 => x"55",
          6110 => x"74",
          6111 => x"80",
          6112 => x"ac",
          6113 => x"81",
          6114 => x"f7",
          6115 => x"58",
          6116 => x"76",
          6117 => x"38",
          6118 => x"2e",
          6119 => x"74",
          6120 => x"15",
          6121 => x"ff",
          6122 => x"81",
          6123 => x"cd",
          6124 => x"f7",
          6125 => x"83",
          6126 => x"33",
          6127 => x"15",
          6128 => x"70",
          6129 => x"55",
          6130 => x"27",
          6131 => x"83",
          6132 => x"70",
          6133 => x"80",
          6134 => x"54",
          6135 => x"e4",
          6136 => x"ff",
          6137 => x"2a",
          6138 => x"81",
          6139 => x"58",
          6140 => x"85",
          6141 => x"0b",
          6142 => x"34",
          6143 => x"06",
          6144 => x"2e",
          6145 => x"81",
          6146 => x"e6",
          6147 => x"83",
          6148 => x"83",
          6149 => x"83",
          6150 => x"70",
          6151 => x"33",
          6152 => x"33",
          6153 => x"5e",
          6154 => x"83",
          6155 => x"33",
          6156 => x"ff",
          6157 => x"83",
          6158 => x"33",
          6159 => x"2e",
          6160 => x"83",
          6161 => x"33",
          6162 => x"ff",
          6163 => x"83",
          6164 => x"33",
          6165 => x"ec",
          6166 => x"ff",
          6167 => x"81",
          6168 => x"38",
          6169 => x"16",
          6170 => x"81",
          6171 => x"38",
          6172 => x"06",
          6173 => x"ff",
          6174 => x"38",
          6175 => x"16",
          6176 => x"74",
          6177 => x"38",
          6178 => x"08",
          6179 => x"87",
          6180 => x"08",
          6181 => x"73",
          6182 => x"38",
          6183 => x"c0",
          6184 => x"83",
          6185 => x"58",
          6186 => x"81",
          6187 => x"54",
          6188 => x"fe",
          6189 => x"83",
          6190 => x"77",
          6191 => x"34",
          6192 => x"53",
          6193 => x"82",
          6194 => x"10",
          6195 => x"b4",
          6196 => x"08",
          6197 => x"94",
          6198 => x"80",
          6199 => x"83",
          6200 => x"c0",
          6201 => x"5e",
          6202 => x"27",
          6203 => x"80",
          6204 => x"92",
          6205 => x"72",
          6206 => x"38",
          6207 => x"83",
          6208 => x"87",
          6209 => x"08",
          6210 => x"0c",
          6211 => x"06",
          6212 => x"2e",
          6213 => x"f9",
          6214 => x"54",
          6215 => x"14",
          6216 => x"81",
          6217 => x"a5",
          6218 => x"ec",
          6219 => x"80",
          6220 => x"38",
          6221 => x"83",
          6222 => x"c3",
          6223 => x"f0",
          6224 => x"39",
          6225 => x"e0",
          6226 => x"56",
          6227 => x"7c",
          6228 => x"38",
          6229 => x"09",
          6230 => x"b4",
          6231 => x"2e",
          6232 => x"79",
          6233 => x"d7",
          6234 => x"ff",
          6235 => x"77",
          6236 => x"2b",
          6237 => x"80",
          6238 => x"73",
          6239 => x"38",
          6240 => x"81",
          6241 => x"10",
          6242 => x"87",
          6243 => x"98",
          6244 => x"57",
          6245 => x"73",
          6246 => x"78",
          6247 => x"79",
          6248 => x"11",
          6249 => x"05",
          6250 => x"05",
          6251 => x"56",
          6252 => x"c0",
          6253 => x"83",
          6254 => x"57",
          6255 => x"80",
          6256 => x"2e",
          6257 => x"79",
          6258 => x"59",
          6259 => x"82",
          6260 => x"39",
          6261 => x"fa",
          6262 => x"0b",
          6263 => x"33",
          6264 => x"81",
          6265 => x"38",
          6266 => x"70",
          6267 => x"25",
          6268 => x"59",
          6269 => x"38",
          6270 => x"09",
          6271 => x"cc",
          6272 => x"2e",
          6273 => x"80",
          6274 => x"10",
          6275 => x"98",
          6276 => x"5d",
          6277 => x"2e",
          6278 => x"81",
          6279 => x"ff",
          6280 => x"93",
          6281 => x"38",
          6282 => x"33",
          6283 => x"2e",
          6284 => x"84",
          6285 => x"55",
          6286 => x"38",
          6287 => x"06",
          6288 => x"cc",
          6289 => x"84",
          6290 => x"8f",
          6291 => x"be",
          6292 => x"f0",
          6293 => x"39",
          6294 => x"2e",
          6295 => x"f7",
          6296 => x"81",
          6297 => x"83",
          6298 => x"34",
          6299 => x"80",
          6300 => x"d4",
          6301 => x"0b",
          6302 => x"15",
          6303 => x"83",
          6304 => x"34",
          6305 => x"74",
          6306 => x"53",
          6307 => x"2e",
          6308 => x"83",
          6309 => x"33",
          6310 => x"27",
          6311 => x"77",
          6312 => x"54",
          6313 => x"09",
          6314 => x"fc",
          6315 => x"e0",
          6316 => x"05",
          6317 => x"9c",
          6318 => x"74",
          6319 => x"e8",
          6320 => x"98",
          6321 => x"f7",
          6322 => x"81",
          6323 => x"fb",
          6324 => x"0b",
          6325 => x"15",
          6326 => x"39",
          6327 => x"e5",
          6328 => x"81",
          6329 => x"fa",
          6330 => x"83",
          6331 => x"80",
          6332 => x"e5",
          6333 => x"ec",
          6334 => x"e6",
          6335 => x"f7",
          6336 => x"f7",
          6337 => x"5d",
          6338 => x"5e",
          6339 => x"39",
          6340 => x"09",
          6341 => x"cb",
          6342 => x"7a",
          6343 => x"ce",
          6344 => x"2e",
          6345 => x"fc",
          6346 => x"93",
          6347 => x"34",
          6348 => x"f8",
          6349 => x"0b",
          6350 => x"33",
          6351 => x"83",
          6352 => x"73",
          6353 => x"34",
          6354 => x"ac",
          6355 => x"84",
          6356 => x"58",
          6357 => x"38",
          6358 => x"84",
          6359 => x"ff",
          6360 => x"39",
          6361 => x"f7",
          6362 => x"2e",
          6363 => x"84",
          6364 => x"ec",
          6365 => x"39",
          6366 => x"33",
          6367 => x"06",
          6368 => x"5a",
          6369 => x"27",
          6370 => x"55",
          6371 => x"ba",
          6372 => x"ff",
          6373 => x"55",
          6374 => x"27",
          6375 => x"54",
          6376 => x"bc",
          6377 => x"80",
          6378 => x"ff",
          6379 => x"05",
          6380 => x"27",
          6381 => x"53",
          6382 => x"bd",
          6383 => x"f6",
          6384 => x"52",
          6385 => x"ba",
          6386 => x"59",
          6387 => x"72",
          6388 => x"39",
          6389 => x"52",
          6390 => x"51",
          6391 => x"3f",
          6392 => x"f8",
          6393 => x"f7",
          6394 => x"fc",
          6395 => x"3d",
          6396 => x"f5",
          6397 => x"3d",
          6398 => x"3d",
          6399 => x"83",
          6400 => x"54",
          6401 => x"05",
          6402 => x"34",
          6403 => x"08",
          6404 => x"72",
          6405 => x"83",
          6406 => x"56",
          6407 => x"81",
          6408 => x"0b",
          6409 => x"e8",
          6410 => x"98",
          6411 => x"f4",
          6412 => x"80",
          6413 => x"54",
          6414 => x"9c",
          6415 => x"c0",
          6416 => x"52",
          6417 => x"f6",
          6418 => x"33",
          6419 => x"9c",
          6420 => x"75",
          6421 => x"38",
          6422 => x"2e",
          6423 => x"c0",
          6424 => x"52",
          6425 => x"74",
          6426 => x"38",
          6427 => x"ff",
          6428 => x"38",
          6429 => x"9c",
          6430 => x"90",
          6431 => x"c0",
          6432 => x"53",
          6433 => x"9c",
          6434 => x"73",
          6435 => x"81",
          6436 => x"c0",
          6437 => x"53",
          6438 => x"27",
          6439 => x"81",
          6440 => x"38",
          6441 => x"a4",
          6442 => x"56",
          6443 => x"a4",
          6444 => x"72",
          6445 => x"38",
          6446 => x"a3",
          6447 => x"ff",
          6448 => x"fe",
          6449 => x"ff",
          6450 => x"77",
          6451 => x"0c",
          6452 => x"04",
          6453 => x"81",
          6454 => x"54",
          6455 => x"81",
          6456 => x"d4",
          6457 => x"d7",
          6458 => x"84",
          6459 => x"89",
          6460 => x"f9",
          6461 => x"02",
          6462 => x"05",
          6463 => x"80",
          6464 => x"98",
          6465 => x"2b",
          6466 => x"80",
          6467 => x"98",
          6468 => x"56",
          6469 => x"83",
          6470 => x"90",
          6471 => x"84",
          6472 => x"90",
          6473 => x"85",
          6474 => x"86",
          6475 => x"f4",
          6476 => x"75",
          6477 => x"83",
          6478 => x"52",
          6479 => x"34",
          6480 => x"f4",
          6481 => x"57",
          6482 => x"16",
          6483 => x"86",
          6484 => x"34",
          6485 => x"9c",
          6486 => x"98",
          6487 => x"ce",
          6488 => x"87",
          6489 => x"08",
          6490 => x"98",
          6491 => x"71",
          6492 => x"38",
          6493 => x"87",
          6494 => x"08",
          6495 => x"74",
          6496 => x"72",
          6497 => x"db",
          6498 => x"98",
          6499 => x"ff",
          6500 => x"27",
          6501 => x"72",
          6502 => x"2e",
          6503 => x"87",
          6504 => x"08",
          6505 => x"05",
          6506 => x"98",
          6507 => x"87",
          6508 => x"08",
          6509 => x"2e",
          6510 => x"15",
          6511 => x"98",
          6512 => x"53",
          6513 => x"87",
          6514 => x"ff",
          6515 => x"87",
          6516 => x"08",
          6517 => x"71",
          6518 => x"df",
          6519 => x"72",
          6520 => x"d7",
          6521 => x"2e",
          6522 => x"75",
          6523 => x"53",
          6524 => x"38",
          6525 => x"81",
          6526 => x"76",
          6527 => x"c6",
          6528 => x"80",
          6529 => x"53",
          6530 => x"92",
          6531 => x"81",
          6532 => x"72",
          6533 => x"54",
          6534 => x"26",
          6535 => x"84",
          6536 => x"89",
          6537 => x"81",
          6538 => x"e8",
          6539 => x"d4",
          6540 => x"84",
          6541 => x"89",
          6542 => x"ff",
          6543 => x"ff",
          6544 => x"76",
          6545 => x"ff",
          6546 => x"39",
          6547 => x"7a",
          6548 => x"a7",
          6549 => x"57",
          6550 => x"f4",
          6551 => x"88",
          6552 => x"80",
          6553 => x"7a",
          6554 => x"51",
          6555 => x"76",
          6556 => x"73",
          6557 => x"71",
          6558 => x"76",
          6559 => x"72",
          6560 => x"73",
          6561 => x"7b",
          6562 => x"08",
          6563 => x"84",
          6564 => x"55",
          6565 => x"74",
          6566 => x"71",
          6567 => x"53",
          6568 => x"81",
          6569 => x"73",
          6570 => x"38",
          6571 => x"08",
          6572 => x"16",
          6573 => x"98",
          6574 => x"e2",
          6575 => x"0b",
          6576 => x"08",
          6577 => x"0b",
          6578 => x"80",
          6579 => x"80",
          6580 => x"c0",
          6581 => x"83",
          6582 => x"56",
          6583 => x"05",
          6584 => x"98",
          6585 => x"87",
          6586 => x"08",
          6587 => x"2e",
          6588 => x"15",
          6589 => x"98",
          6590 => x"53",
          6591 => x"87",
          6592 => x"fe",
          6593 => x"87",
          6594 => x"08",
          6595 => x"71",
          6596 => x"cd",
          6597 => x"72",
          6598 => x"c5",
          6599 => x"98",
          6600 => x"ce",
          6601 => x"87",
          6602 => x"08",
          6603 => x"98",
          6604 => x"75",
          6605 => x"38",
          6606 => x"87",
          6607 => x"08",
          6608 => x"74",
          6609 => x"72",
          6610 => x"db",
          6611 => x"98",
          6612 => x"ff",
          6613 => x"27",
          6614 => x"56",
          6615 => x"a2",
          6616 => x"2e",
          6617 => x"81",
          6618 => x"72",
          6619 => x"75",
          6620 => x"06",
          6621 => x"a1",
          6622 => x"ba",
          6623 => x"3d",
          6624 => x"17",
          6625 => x"06",
          6626 => x"da",
          6627 => x"81",
          6628 => x"52",
          6629 => x"e1",
          6630 => x"83",
          6631 => x"58",
          6632 => x"3f",
          6633 => x"8c",
          6634 => x"0d",
          6635 => x"0d",
          6636 => x"08",
          6637 => x"71",
          6638 => x"83",
          6639 => x"56",
          6640 => x"81",
          6641 => x"0b",
          6642 => x"e8",
          6643 => x"98",
          6644 => x"f4",
          6645 => x"80",
          6646 => x"54",
          6647 => x"9c",
          6648 => x"c0",
          6649 => x"53",
          6650 => x"f6",
          6651 => x"33",
          6652 => x"9c",
          6653 => x"70",
          6654 => x"38",
          6655 => x"2e",
          6656 => x"c0",
          6657 => x"51",
          6658 => x"74",
          6659 => x"38",
          6660 => x"ff",
          6661 => x"38",
          6662 => x"9c",
          6663 => x"90",
          6664 => x"c0",
          6665 => x"52",
          6666 => x"9c",
          6667 => x"72",
          6668 => x"81",
          6669 => x"c0",
          6670 => x"52",
          6671 => x"27",
          6672 => x"81",
          6673 => x"38",
          6674 => x"a4",
          6675 => x"53",
          6676 => x"98",
          6677 => x"71",
          6678 => x"38",
          6679 => x"8a",
          6680 => x"ff",
          6681 => x"fe",
          6682 => x"39",
          6683 => x"81",
          6684 => x"54",
          6685 => x"3d",
          6686 => x"90",
          6687 => x"f6",
          6688 => x"0d",
          6689 => x"0d",
          6690 => x"08",
          6691 => x"83",
          6692 => x"ff",
          6693 => x"83",
          6694 => x"70",
          6695 => x"33",
          6696 => x"71",
          6697 => x"77",
          6698 => x"81",
          6699 => x"98",
          6700 => x"2b",
          6701 => x"41",
          6702 => x"57",
          6703 => x"57",
          6704 => x"24",
          6705 => x"72",
          6706 => x"33",
          6707 => x"71",
          6708 => x"83",
          6709 => x"05",
          6710 => x"12",
          6711 => x"2b",
          6712 => x"07",
          6713 => x"52",
          6714 => x"80",
          6715 => x"9e",
          6716 => x"33",
          6717 => x"71",
          6718 => x"83",
          6719 => x"05",
          6720 => x"52",
          6721 => x"74",
          6722 => x"73",
          6723 => x"54",
          6724 => x"34",
          6725 => x"08",
          6726 => x"12",
          6727 => x"33",
          6728 => x"07",
          6729 => x"5c",
          6730 => x"51",
          6731 => x"34",
          6732 => x"34",
          6733 => x"08",
          6734 => x"0b",
          6735 => x"80",
          6736 => x"34",
          6737 => x"08",
          6738 => x"14",
          6739 => x"14",
          6740 => x"fc",
          6741 => x"33",
          6742 => x"71",
          6743 => x"82",
          6744 => x"70",
          6745 => x"58",
          6746 => x"72",
          6747 => x"13",
          6748 => x"0d",
          6749 => x"33",
          6750 => x"71",
          6751 => x"83",
          6752 => x"11",
          6753 => x"85",
          6754 => x"88",
          6755 => x"88",
          6756 => x"54",
          6757 => x"58",
          6758 => x"34",
          6759 => x"34",
          6760 => x"08",
          6761 => x"11",
          6762 => x"33",
          6763 => x"71",
          6764 => x"56",
          6765 => x"72",
          6766 => x"33",
          6767 => x"71",
          6768 => x"70",
          6769 => x"55",
          6770 => x"86",
          6771 => x"87",
          6772 => x"b9",
          6773 => x"70",
          6774 => x"33",
          6775 => x"07",
          6776 => x"06",
          6777 => x"5a",
          6778 => x"76",
          6779 => x"81",
          6780 => x"b9",
          6781 => x"17",
          6782 => x"12",
          6783 => x"2b",
          6784 => x"07",
          6785 => x"33",
          6786 => x"71",
          6787 => x"70",
          6788 => x"ff",
          6789 => x"05",
          6790 => x"54",
          6791 => x"5c",
          6792 => x"52",
          6793 => x"34",
          6794 => x"34",
          6795 => x"08",
          6796 => x"33",
          6797 => x"71",
          6798 => x"83",
          6799 => x"05",
          6800 => x"12",
          6801 => x"2b",
          6802 => x"ff",
          6803 => x"2a",
          6804 => x"55",
          6805 => x"52",
          6806 => x"70",
          6807 => x"84",
          6808 => x"70",
          6809 => x"33",
          6810 => x"71",
          6811 => x"83",
          6812 => x"05",
          6813 => x"12",
          6814 => x"2b",
          6815 => x"07",
          6816 => x"52",
          6817 => x"53",
          6818 => x"fc",
          6819 => x"33",
          6820 => x"71",
          6821 => x"82",
          6822 => x"70",
          6823 => x"59",
          6824 => x"34",
          6825 => x"34",
          6826 => x"08",
          6827 => x"33",
          6828 => x"71",
          6829 => x"83",
          6830 => x"05",
          6831 => x"83",
          6832 => x"88",
          6833 => x"88",
          6834 => x"5c",
          6835 => x"52",
          6836 => x"15",
          6837 => x"15",
          6838 => x"0d",
          6839 => x"0d",
          6840 => x"fc",
          6841 => x"76",
          6842 => x"38",
          6843 => x"86",
          6844 => x"fb",
          6845 => x"3d",
          6846 => x"ff",
          6847 => x"b9",
          6848 => x"80",
          6849 => x"f8",
          6850 => x"80",
          6851 => x"84",
          6852 => x"fe",
          6853 => x"84",
          6854 => x"55",
          6855 => x"81",
          6856 => x"34",
          6857 => x"08",
          6858 => x"15",
          6859 => x"85",
          6860 => x"b9",
          6861 => x"76",
          6862 => x"81",
          6863 => x"34",
          6864 => x"08",
          6865 => x"22",
          6866 => x"80",
          6867 => x"83",
          6868 => x"70",
          6869 => x"51",
          6870 => x"88",
          6871 => x"89",
          6872 => x"b9",
          6873 => x"10",
          6874 => x"b9",
          6875 => x"f8",
          6876 => x"76",
          6877 => x"81",
          6878 => x"34",
          6879 => x"f7",
          6880 => x"52",
          6881 => x"51",
          6882 => x"8e",
          6883 => x"83",
          6884 => x"70",
          6885 => x"06",
          6886 => x"83",
          6887 => x"84",
          6888 => x"84",
          6889 => x"12",
          6890 => x"2b",
          6891 => x"59",
          6892 => x"81",
          6893 => x"75",
          6894 => x"cc",
          6895 => x"10",
          6896 => x"33",
          6897 => x"71",
          6898 => x"70",
          6899 => x"06",
          6900 => x"83",
          6901 => x"70",
          6902 => x"53",
          6903 => x"52",
          6904 => x"8a",
          6905 => x"2e",
          6906 => x"73",
          6907 => x"12",
          6908 => x"33",
          6909 => x"07",
          6910 => x"c1",
          6911 => x"ff",
          6912 => x"38",
          6913 => x"56",
          6914 => x"2b",
          6915 => x"33",
          6916 => x"71",
          6917 => x"70",
          6918 => x"06",
          6919 => x"56",
          6920 => x"79",
          6921 => x"81",
          6922 => x"74",
          6923 => x"8d",
          6924 => x"78",
          6925 => x"85",
          6926 => x"2e",
          6927 => x"74",
          6928 => x"2b",
          6929 => x"82",
          6930 => x"70",
          6931 => x"5c",
          6932 => x"76",
          6933 => x"81",
          6934 => x"b9",
          6935 => x"76",
          6936 => x"53",
          6937 => x"34",
          6938 => x"34",
          6939 => x"08",
          6940 => x"33",
          6941 => x"71",
          6942 => x"70",
          6943 => x"ff",
          6944 => x"05",
          6945 => x"ff",
          6946 => x"2a",
          6947 => x"57",
          6948 => x"75",
          6949 => x"72",
          6950 => x"53",
          6951 => x"34",
          6952 => x"08",
          6953 => x"74",
          6954 => x"15",
          6955 => x"fc",
          6956 => x"86",
          6957 => x"12",
          6958 => x"2b",
          6959 => x"07",
          6960 => x"5c",
          6961 => x"75",
          6962 => x"72",
          6963 => x"84",
          6964 => x"70",
          6965 => x"05",
          6966 => x"87",
          6967 => x"88",
          6968 => x"88",
          6969 => x"58",
          6970 => x"15",
          6971 => x"15",
          6972 => x"fc",
          6973 => x"84",
          6974 => x"12",
          6975 => x"2b",
          6976 => x"07",
          6977 => x"5a",
          6978 => x"75",
          6979 => x"72",
          6980 => x"84",
          6981 => x"70",
          6982 => x"05",
          6983 => x"85",
          6984 => x"88",
          6985 => x"88",
          6986 => x"57",
          6987 => x"15",
          6988 => x"15",
          6989 => x"fc",
          6990 => x"05",
          6991 => x"ba",
          6992 => x"3d",
          6993 => x"14",
          6994 => x"33",
          6995 => x"71",
          6996 => x"79",
          6997 => x"33",
          6998 => x"71",
          6999 => x"70",
          7000 => x"5b",
          7001 => x"52",
          7002 => x"34",
          7003 => x"34",
          7004 => x"08",
          7005 => x"11",
          7006 => x"33",
          7007 => x"71",
          7008 => x"74",
          7009 => x"33",
          7010 => x"71",
          7011 => x"70",
          7012 => x"5d",
          7013 => x"5b",
          7014 => x"86",
          7015 => x"87",
          7016 => x"b9",
          7017 => x"70",
          7018 => x"33",
          7019 => x"07",
          7020 => x"06",
          7021 => x"59",
          7022 => x"75",
          7023 => x"81",
          7024 => x"b9",
          7025 => x"84",
          7026 => x"f1",
          7027 => x"0d",
          7028 => x"fc",
          7029 => x"76",
          7030 => x"38",
          7031 => x"8a",
          7032 => x"ba",
          7033 => x"3d",
          7034 => x"51",
          7035 => x"84",
          7036 => x"84",
          7037 => x"89",
          7038 => x"84",
          7039 => x"84",
          7040 => x"a0",
          7041 => x"b9",
          7042 => x"80",
          7043 => x"52",
          7044 => x"51",
          7045 => x"3f",
          7046 => x"08",
          7047 => x"34",
          7048 => x"16",
          7049 => x"fc",
          7050 => x"84",
          7051 => x"0b",
          7052 => x"84",
          7053 => x"56",
          7054 => x"34",
          7055 => x"17",
          7056 => x"fc",
          7057 => x"f8",
          7058 => x"fe",
          7059 => x"70",
          7060 => x"06",
          7061 => x"58",
          7062 => x"74",
          7063 => x"73",
          7064 => x"84",
          7065 => x"70",
          7066 => x"84",
          7067 => x"05",
          7068 => x"55",
          7069 => x"34",
          7070 => x"15",
          7071 => x"77",
          7072 => x"dd",
          7073 => x"39",
          7074 => x"65",
          7075 => x"80",
          7076 => x"fc",
          7077 => x"41",
          7078 => x"84",
          7079 => x"80",
          7080 => x"38",
          7081 => x"88",
          7082 => x"54",
          7083 => x"8f",
          7084 => x"05",
          7085 => x"05",
          7086 => x"ff",
          7087 => x"73",
          7088 => x"06",
          7089 => x"83",
          7090 => x"ff",
          7091 => x"83",
          7092 => x"70",
          7093 => x"33",
          7094 => x"07",
          7095 => x"70",
          7096 => x"06",
          7097 => x"10",
          7098 => x"83",
          7099 => x"70",
          7100 => x"33",
          7101 => x"07",
          7102 => x"70",
          7103 => x"42",
          7104 => x"53",
          7105 => x"5c",
          7106 => x"5e",
          7107 => x"7a",
          7108 => x"38",
          7109 => x"83",
          7110 => x"88",
          7111 => x"10",
          7112 => x"70",
          7113 => x"33",
          7114 => x"71",
          7115 => x"53",
          7116 => x"56",
          7117 => x"24",
          7118 => x"7a",
          7119 => x"f6",
          7120 => x"58",
          7121 => x"87",
          7122 => x"80",
          7123 => x"38",
          7124 => x"77",
          7125 => x"be",
          7126 => x"59",
          7127 => x"92",
          7128 => x"1e",
          7129 => x"12",
          7130 => x"2b",
          7131 => x"07",
          7132 => x"33",
          7133 => x"71",
          7134 => x"90",
          7135 => x"43",
          7136 => x"57",
          7137 => x"60",
          7138 => x"38",
          7139 => x"11",
          7140 => x"33",
          7141 => x"71",
          7142 => x"7a",
          7143 => x"33",
          7144 => x"71",
          7145 => x"83",
          7146 => x"05",
          7147 => x"85",
          7148 => x"88",
          7149 => x"88",
          7150 => x"48",
          7151 => x"58",
          7152 => x"56",
          7153 => x"34",
          7154 => x"34",
          7155 => x"08",
          7156 => x"11",
          7157 => x"33",
          7158 => x"71",
          7159 => x"74",
          7160 => x"33",
          7161 => x"71",
          7162 => x"70",
          7163 => x"42",
          7164 => x"57",
          7165 => x"86",
          7166 => x"87",
          7167 => x"b9",
          7168 => x"70",
          7169 => x"33",
          7170 => x"07",
          7171 => x"06",
          7172 => x"5a",
          7173 => x"76",
          7174 => x"81",
          7175 => x"b9",
          7176 => x"1f",
          7177 => x"83",
          7178 => x"8b",
          7179 => x"2b",
          7180 => x"73",
          7181 => x"33",
          7182 => x"07",
          7183 => x"41",
          7184 => x"5f",
          7185 => x"79",
          7186 => x"81",
          7187 => x"b9",
          7188 => x"1f",
          7189 => x"12",
          7190 => x"2b",
          7191 => x"07",
          7192 => x"14",
          7193 => x"33",
          7194 => x"07",
          7195 => x"41",
          7196 => x"5f",
          7197 => x"79",
          7198 => x"75",
          7199 => x"84",
          7200 => x"70",
          7201 => x"33",
          7202 => x"71",
          7203 => x"66",
          7204 => x"70",
          7205 => x"52",
          7206 => x"05",
          7207 => x"fe",
          7208 => x"84",
          7209 => x"1e",
          7210 => x"65",
          7211 => x"83",
          7212 => x"5d",
          7213 => x"62",
          7214 => x"38",
          7215 => x"84",
          7216 => x"95",
          7217 => x"84",
          7218 => x"84",
          7219 => x"a0",
          7220 => x"b9",
          7221 => x"80",
          7222 => x"52",
          7223 => x"51",
          7224 => x"3f",
          7225 => x"08",
          7226 => x"34",
          7227 => x"1f",
          7228 => x"fc",
          7229 => x"84",
          7230 => x"0b",
          7231 => x"84",
          7232 => x"5c",
          7233 => x"34",
          7234 => x"1d",
          7235 => x"fc",
          7236 => x"f8",
          7237 => x"fe",
          7238 => x"70",
          7239 => x"06",
          7240 => x"5c",
          7241 => x"78",
          7242 => x"77",
          7243 => x"84",
          7244 => x"70",
          7245 => x"84",
          7246 => x"05",
          7247 => x"56",
          7248 => x"34",
          7249 => x"15",
          7250 => x"fc",
          7251 => x"fa",
          7252 => x"80",
          7253 => x"38",
          7254 => x"80",
          7255 => x"38",
          7256 => x"9b",
          7257 => x"8c",
          7258 => x"8c",
          7259 => x"0d",
          7260 => x"84",
          7261 => x"71",
          7262 => x"11",
          7263 => x"05",
          7264 => x"12",
          7265 => x"2b",
          7266 => x"ff",
          7267 => x"2a",
          7268 => x"5e",
          7269 => x"34",
          7270 => x"34",
          7271 => x"fc",
          7272 => x"88",
          7273 => x"75",
          7274 => x"7b",
          7275 => x"84",
          7276 => x"70",
          7277 => x"81",
          7278 => x"88",
          7279 => x"83",
          7280 => x"f8",
          7281 => x"64",
          7282 => x"06",
          7283 => x"4a",
          7284 => x"5e",
          7285 => x"63",
          7286 => x"76",
          7287 => x"41",
          7288 => x"05",
          7289 => x"fc",
          7290 => x"63",
          7291 => x"81",
          7292 => x"84",
          7293 => x"05",
          7294 => x"ed",
          7295 => x"54",
          7296 => x"7b",
          7297 => x"83",
          7298 => x"42",
          7299 => x"39",
          7300 => x"ff",
          7301 => x"70",
          7302 => x"06",
          7303 => x"83",
          7304 => x"88",
          7305 => x"10",
          7306 => x"70",
          7307 => x"33",
          7308 => x"71",
          7309 => x"53",
          7310 => x"58",
          7311 => x"73",
          7312 => x"f7",
          7313 => x"39",
          7314 => x"fa",
          7315 => x"7a",
          7316 => x"38",
          7317 => x"ff",
          7318 => x"7b",
          7319 => x"38",
          7320 => x"84",
          7321 => x"84",
          7322 => x"a0",
          7323 => x"b9",
          7324 => x"80",
          7325 => x"52",
          7326 => x"51",
          7327 => x"3f",
          7328 => x"08",
          7329 => x"34",
          7330 => x"1b",
          7331 => x"fc",
          7332 => x"84",
          7333 => x"0b",
          7334 => x"84",
          7335 => x"58",
          7336 => x"34",
          7337 => x"19",
          7338 => x"fc",
          7339 => x"f8",
          7340 => x"fe",
          7341 => x"70",
          7342 => x"06",
          7343 => x"58",
          7344 => x"74",
          7345 => x"34",
          7346 => x"05",
          7347 => x"f8",
          7348 => x"10",
          7349 => x"fc",
          7350 => x"05",
          7351 => x"61",
          7352 => x"81",
          7353 => x"34",
          7354 => x"80",
          7355 => x"de",
          7356 => x"ff",
          7357 => x"61",
          7358 => x"c0",
          7359 => x"39",
          7360 => x"82",
          7361 => x"51",
          7362 => x"7f",
          7363 => x"ba",
          7364 => x"3d",
          7365 => x"1e",
          7366 => x"83",
          7367 => x"8b",
          7368 => x"2b",
          7369 => x"86",
          7370 => x"12",
          7371 => x"2b",
          7372 => x"07",
          7373 => x"14",
          7374 => x"33",
          7375 => x"07",
          7376 => x"43",
          7377 => x"5b",
          7378 => x"5c",
          7379 => x"64",
          7380 => x"7a",
          7381 => x"34",
          7382 => x"08",
          7383 => x"11",
          7384 => x"33",
          7385 => x"71",
          7386 => x"74",
          7387 => x"33",
          7388 => x"71",
          7389 => x"70",
          7390 => x"41",
          7391 => x"59",
          7392 => x"64",
          7393 => x"7a",
          7394 => x"34",
          7395 => x"08",
          7396 => x"81",
          7397 => x"88",
          7398 => x"ff",
          7399 => x"88",
          7400 => x"5a",
          7401 => x"34",
          7402 => x"34",
          7403 => x"08",
          7404 => x"11",
          7405 => x"33",
          7406 => x"71",
          7407 => x"74",
          7408 => x"81",
          7409 => x"88",
          7410 => x"88",
          7411 => x"5e",
          7412 => x"45",
          7413 => x"34",
          7414 => x"34",
          7415 => x"08",
          7416 => x"33",
          7417 => x"71",
          7418 => x"83",
          7419 => x"05",
          7420 => x"83",
          7421 => x"88",
          7422 => x"88",
          7423 => x"40",
          7424 => x"55",
          7425 => x"18",
          7426 => x"18",
          7427 => x"fc",
          7428 => x"82",
          7429 => x"12",
          7430 => x"2b",
          7431 => x"62",
          7432 => x"2b",
          7433 => x"5d",
          7434 => x"05",
          7435 => x"95",
          7436 => x"fc",
          7437 => x"05",
          7438 => x"ff",
          7439 => x"fc",
          7440 => x"ff",
          7441 => x"b9",
          7442 => x"80",
          7443 => x"f8",
          7444 => x"80",
          7445 => x"84",
          7446 => x"fe",
          7447 => x"84",
          7448 => x"56",
          7449 => x"81",
          7450 => x"34",
          7451 => x"08",
          7452 => x"16",
          7453 => x"85",
          7454 => x"b9",
          7455 => x"7f",
          7456 => x"81",
          7457 => x"34",
          7458 => x"08",
          7459 => x"22",
          7460 => x"80",
          7461 => x"83",
          7462 => x"70",
          7463 => x"43",
          7464 => x"88",
          7465 => x"89",
          7466 => x"b9",
          7467 => x"10",
          7468 => x"b9",
          7469 => x"f8",
          7470 => x"7f",
          7471 => x"81",
          7472 => x"34",
          7473 => x"bd",
          7474 => x"fc",
          7475 => x"19",
          7476 => x"33",
          7477 => x"71",
          7478 => x"79",
          7479 => x"33",
          7480 => x"71",
          7481 => x"70",
          7482 => x"48",
          7483 => x"55",
          7484 => x"05",
          7485 => x"85",
          7486 => x"b9",
          7487 => x"1e",
          7488 => x"85",
          7489 => x"8b",
          7490 => x"2b",
          7491 => x"86",
          7492 => x"15",
          7493 => x"2b",
          7494 => x"2a",
          7495 => x"48",
          7496 => x"40",
          7497 => x"05",
          7498 => x"87",
          7499 => x"b9",
          7500 => x"70",
          7501 => x"33",
          7502 => x"07",
          7503 => x"06",
          7504 => x"59",
          7505 => x"75",
          7506 => x"81",
          7507 => x"b9",
          7508 => x"1f",
          7509 => x"12",
          7510 => x"2b",
          7511 => x"07",
          7512 => x"33",
          7513 => x"71",
          7514 => x"70",
          7515 => x"ff",
          7516 => x"05",
          7517 => x"48",
          7518 => x"5d",
          7519 => x"41",
          7520 => x"34",
          7521 => x"34",
          7522 => x"08",
          7523 => x"33",
          7524 => x"71",
          7525 => x"83",
          7526 => x"05",
          7527 => x"12",
          7528 => x"2b",
          7529 => x"ff",
          7530 => x"2a",
          7531 => x"5e",
          7532 => x"5b",
          7533 => x"76",
          7534 => x"34",
          7535 => x"ff",
          7536 => x"b3",
          7537 => x"33",
          7538 => x"71",
          7539 => x"83",
          7540 => x"05",
          7541 => x"85",
          7542 => x"88",
          7543 => x"88",
          7544 => x"5a",
          7545 => x"78",
          7546 => x"79",
          7547 => x"84",
          7548 => x"70",
          7549 => x"33",
          7550 => x"71",
          7551 => x"83",
          7552 => x"05",
          7553 => x"87",
          7554 => x"88",
          7555 => x"88",
          7556 => x"5e",
          7557 => x"55",
          7558 => x"86",
          7559 => x"60",
          7560 => x"84",
          7561 => x"18",
          7562 => x"12",
          7563 => x"2b",
          7564 => x"ff",
          7565 => x"2a",
          7566 => x"55",
          7567 => x"78",
          7568 => x"84",
          7569 => x"70",
          7570 => x"81",
          7571 => x"8b",
          7572 => x"2b",
          7573 => x"70",
          7574 => x"33",
          7575 => x"07",
          7576 => x"8f",
          7577 => x"77",
          7578 => x"2a",
          7579 => x"5f",
          7580 => x"5e",
          7581 => x"17",
          7582 => x"17",
          7583 => x"fc",
          7584 => x"70",
          7585 => x"33",
          7586 => x"71",
          7587 => x"74",
          7588 => x"81",
          7589 => x"88",
          7590 => x"ff",
          7591 => x"88",
          7592 => x"5e",
          7593 => x"5d",
          7594 => x"34",
          7595 => x"34",
          7596 => x"08",
          7597 => x"11",
          7598 => x"33",
          7599 => x"71",
          7600 => x"74",
          7601 => x"33",
          7602 => x"71",
          7603 => x"83",
          7604 => x"05",
          7605 => x"85",
          7606 => x"88",
          7607 => x"88",
          7608 => x"49",
          7609 => x"59",
          7610 => x"57",
          7611 => x"1d",
          7612 => x"1d",
          7613 => x"fc",
          7614 => x"84",
          7615 => x"12",
          7616 => x"2b",
          7617 => x"07",
          7618 => x"14",
          7619 => x"33",
          7620 => x"07",
          7621 => x"5f",
          7622 => x"40",
          7623 => x"77",
          7624 => x"7b",
          7625 => x"84",
          7626 => x"16",
          7627 => x"12",
          7628 => x"2b",
          7629 => x"ff",
          7630 => x"2a",
          7631 => x"59",
          7632 => x"79",
          7633 => x"84",
          7634 => x"70",
          7635 => x"33",
          7636 => x"71",
          7637 => x"83",
          7638 => x"05",
          7639 => x"15",
          7640 => x"2b",
          7641 => x"2a",
          7642 => x"5d",
          7643 => x"55",
          7644 => x"75",
          7645 => x"84",
          7646 => x"70",
          7647 => x"81",
          7648 => x"8b",
          7649 => x"2b",
          7650 => x"82",
          7651 => x"15",
          7652 => x"2b",
          7653 => x"2a",
          7654 => x"5d",
          7655 => x"55",
          7656 => x"34",
          7657 => x"34",
          7658 => x"08",
          7659 => x"11",
          7660 => x"33",
          7661 => x"07",
          7662 => x"56",
          7663 => x"42",
          7664 => x"7e",
          7665 => x"51",
          7666 => x"3f",
          7667 => x"08",
          7668 => x"61",
          7669 => x"70",
          7670 => x"06",
          7671 => x"f1",
          7672 => x"19",
          7673 => x"33",
          7674 => x"71",
          7675 => x"79",
          7676 => x"33",
          7677 => x"71",
          7678 => x"70",
          7679 => x"48",
          7680 => x"55",
          7681 => x"05",
          7682 => x"85",
          7683 => x"b9",
          7684 => x"1e",
          7685 => x"85",
          7686 => x"8b",
          7687 => x"2b",
          7688 => x"86",
          7689 => x"15",
          7690 => x"2b",
          7691 => x"2a",
          7692 => x"48",
          7693 => x"56",
          7694 => x"05",
          7695 => x"87",
          7696 => x"b9",
          7697 => x"70",
          7698 => x"33",
          7699 => x"07",
          7700 => x"06",
          7701 => x"5c",
          7702 => x"78",
          7703 => x"81",
          7704 => x"b9",
          7705 => x"1f",
          7706 => x"12",
          7707 => x"2b",
          7708 => x"07",
          7709 => x"33",
          7710 => x"71",
          7711 => x"70",
          7712 => x"ff",
          7713 => x"05",
          7714 => x"5d",
          7715 => x"58",
          7716 => x"40",
          7717 => x"34",
          7718 => x"34",
          7719 => x"08",
          7720 => x"33",
          7721 => x"71",
          7722 => x"83",
          7723 => x"05",
          7724 => x"12",
          7725 => x"2b",
          7726 => x"ff",
          7727 => x"2a",
          7728 => x"58",
          7729 => x"5b",
          7730 => x"78",
          7731 => x"77",
          7732 => x"06",
          7733 => x"39",
          7734 => x"54",
          7735 => x"84",
          7736 => x"5f",
          7737 => x"08",
          7738 => x"38",
          7739 => x"52",
          7740 => x"08",
          7741 => x"f5",
          7742 => x"df",
          7743 => x"5b",
          7744 => x"ef",
          7745 => x"e9",
          7746 => x"0d",
          7747 => x"84",
          7748 => x"58",
          7749 => x"2e",
          7750 => x"54",
          7751 => x"73",
          7752 => x"0c",
          7753 => x"04",
          7754 => x"d3",
          7755 => x"8c",
          7756 => x"ba",
          7757 => x"2e",
          7758 => x"53",
          7759 => x"ba",
          7760 => x"fe",
          7761 => x"73",
          7762 => x"0c",
          7763 => x"04",
          7764 => x"0b",
          7765 => x"0c",
          7766 => x"84",
          7767 => x"82",
          7768 => x"76",
          7769 => x"f4",
          7770 => x"96",
          7771 => x"fc",
          7772 => x"75",
          7773 => x"81",
          7774 => x"b9",
          7775 => x"76",
          7776 => x"81",
          7777 => x"34",
          7778 => x"08",
          7779 => x"17",
          7780 => x"87",
          7781 => x"b9",
          7782 => x"b9",
          7783 => x"05",
          7784 => x"07",
          7785 => x"ff",
          7786 => x"2a",
          7787 => x"56",
          7788 => x"34",
          7789 => x"34",
          7790 => x"22",
          7791 => x"10",
          7792 => x"08",
          7793 => x"55",
          7794 => x"15",
          7795 => x"83",
          7796 => x"54",
          7797 => x"fe",
          7798 => x"cc",
          7799 => x"0d",
          7800 => x"33",
          7801 => x"70",
          7802 => x"38",
          7803 => x"11",
          7804 => x"84",
          7805 => x"83",
          7806 => x"fe",
          7807 => x"93",
          7808 => x"83",
          7809 => x"26",
          7810 => x"51",
          7811 => x"84",
          7812 => x"81",
          7813 => x"72",
          7814 => x"84",
          7815 => x"34",
          7816 => x"12",
          7817 => x"84",
          7818 => x"84",
          7819 => x"f7",
          7820 => x"7e",
          7821 => x"05",
          7822 => x"5a",
          7823 => x"81",
          7824 => x"26",
          7825 => x"ba",
          7826 => x"54",
          7827 => x"54",
          7828 => x"bd",
          7829 => x"85",
          7830 => x"98",
          7831 => x"53",
          7832 => x"51",
          7833 => x"84",
          7834 => x"81",
          7835 => x"74",
          7836 => x"38",
          7837 => x"8c",
          7838 => x"e2",
          7839 => x"26",
          7840 => x"fc",
          7841 => x"54",
          7842 => x"83",
          7843 => x"73",
          7844 => x"ba",
          7845 => x"3d",
          7846 => x"80",
          7847 => x"70",
          7848 => x"5a",
          7849 => x"78",
          7850 => x"38",
          7851 => x"3d",
          7852 => x"60",
          7853 => x"af",
          7854 => x"5c",
          7855 => x"54",
          7856 => x"87",
          7857 => x"88",
          7858 => x"73",
          7859 => x"83",
          7860 => x"38",
          7861 => x"0b",
          7862 => x"8c",
          7863 => x"75",
          7864 => x"d6",
          7865 => x"ba",
          7866 => x"ff",
          7867 => x"80",
          7868 => x"87",
          7869 => x"08",
          7870 => x"38",
          7871 => x"d6",
          7872 => x"80",
          7873 => x"73",
          7874 => x"38",
          7875 => x"55",
          7876 => x"8c",
          7877 => x"0d",
          7878 => x"16",
          7879 => x"81",
          7880 => x"55",
          7881 => x"26",
          7882 => x"d5",
          7883 => x"0d",
          7884 => x"05",
          7885 => x"02",
          7886 => x"05",
          7887 => x"55",
          7888 => x"73",
          7889 => x"84",
          7890 => x"33",
          7891 => x"06",
          7892 => x"73",
          7893 => x"0b",
          7894 => x"8c",
          7895 => x"70",
          7896 => x"38",
          7897 => x"ad",
          7898 => x"2e",
          7899 => x"53",
          7900 => x"8c",
          7901 => x"0d",
          7902 => x"0a",
          7903 => x"84",
          7904 => x"86",
          7905 => x"81",
          7906 => x"80",
          7907 => x"8c",
          7908 => x"0d",
          7909 => x"2b",
          7910 => x"8c",
          7911 => x"70",
          7912 => x"08",
          7913 => x"81",
          7914 => x"70",
          7915 => x"38",
          7916 => x"8c",
          7917 => x"ea",
          7918 => x"98",
          7919 => x"70",
          7920 => x"72",
          7921 => x"92",
          7922 => x"71",
          7923 => x"54",
          7924 => x"ff",
          7925 => x"08",
          7926 => x"73",
          7927 => x"90",
          7928 => x"0d",
          7929 => x"0b",
          7930 => x"71",
          7931 => x"74",
          7932 => x"81",
          7933 => x"77",
          7934 => x"83",
          7935 => x"38",
          7936 => x"52",
          7937 => x"51",
          7938 => x"84",
          7939 => x"80",
          7940 => x"81",
          7941 => x"ba",
          7942 => x"3d",
          7943 => x"54",
          7944 => x"53",
          7945 => x"53",
          7946 => x"52",
          7947 => x"3f",
          7948 => x"ba",
          7949 => x"2e",
          7950 => x"d9",
          7951 => x"8c",
          7952 => x"34",
          7953 => x"70",
          7954 => x"31",
          7955 => x"84",
          7956 => x"5c",
          7957 => x"74",
          7958 => x"9b",
          7959 => x"33",
          7960 => x"2e",
          7961 => x"ff",
          7962 => x"54",
          7963 => x"79",
          7964 => x"33",
          7965 => x"3f",
          7966 => x"57",
          7967 => x"2e",
          7968 => x"fe",
          7969 => x"18",
          7970 => x"81",
          7971 => x"06",
          7972 => x"b8",
          7973 => x"80",
          7974 => x"80",
          7975 => x"05",
          7976 => x"17",
          7977 => x"38",
          7978 => x"84",
          7979 => x"ff",
          7980 => x"b7",
          7981 => x"d2",
          7982 => x"d2",
          7983 => x"34",
          7984 => x"ba",
          7985 => x"c1",
          7986 => x"34",
          7987 => x"84",
          7988 => x"80",
          7989 => x"9d",
          7990 => x"c1",
          7991 => x"19",
          7992 => x"0b",
          7993 => x"34",
          7994 => x"55",
          7995 => x"19",
          7996 => x"2a",
          7997 => x"a1",
          7998 => x"90",
          7999 => x"84",
          8000 => x"74",
          8001 => x"7a",
          8002 => x"34",
          8003 => x"5b",
          8004 => x"19",
          8005 => x"2a",
          8006 => x"a5",
          8007 => x"90",
          8008 => x"84",
          8009 => x"7a",
          8010 => x"74",
          8011 => x"34",
          8012 => x"81",
          8013 => x"1a",
          8014 => x"54",
          8015 => x"52",
          8016 => x"51",
          8017 => x"76",
          8018 => x"80",
          8019 => x"81",
          8020 => x"fb",
          8021 => x"ba",
          8022 => x"2e",
          8023 => x"fd",
          8024 => x"3d",
          8025 => x"70",
          8026 => x"56",
          8027 => x"88",
          8028 => x"08",
          8029 => x"38",
          8030 => x"84",
          8031 => x"8f",
          8032 => x"ff",
          8033 => x"58",
          8034 => x"81",
          8035 => x"82",
          8036 => x"38",
          8037 => x"09",
          8038 => x"38",
          8039 => x"16",
          8040 => x"a8",
          8041 => x"5a",
          8042 => x"b4",
          8043 => x"2e",
          8044 => x"17",
          8045 => x"7b",
          8046 => x"06",
          8047 => x"81",
          8048 => x"b8",
          8049 => x"17",
          8050 => x"e3",
          8051 => x"8c",
          8052 => x"85",
          8053 => x"81",
          8054 => x"18",
          8055 => x"9a",
          8056 => x"ff",
          8057 => x"11",
          8058 => x"70",
          8059 => x"1b",
          8060 => x"5d",
          8061 => x"17",
          8062 => x"b5",
          8063 => x"83",
          8064 => x"5c",
          8065 => x"7d",
          8066 => x"06",
          8067 => x"81",
          8068 => x"b8",
          8069 => x"17",
          8070 => x"93",
          8071 => x"8c",
          8072 => x"85",
          8073 => x"81",
          8074 => x"18",
          8075 => x"ca",
          8076 => x"ff",
          8077 => x"11",
          8078 => x"2b",
          8079 => x"81",
          8080 => x"2a",
          8081 => x"59",
          8082 => x"ae",
          8083 => x"ff",
          8084 => x"8c",
          8085 => x"0d",
          8086 => x"2a",
          8087 => x"05",
          8088 => x"08",
          8089 => x"38",
          8090 => x"18",
          8091 => x"5d",
          8092 => x"2e",
          8093 => x"81",
          8094 => x"54",
          8095 => x"17",
          8096 => x"33",
          8097 => x"3f",
          8098 => x"08",
          8099 => x"38",
          8100 => x"5a",
          8101 => x"0c",
          8102 => x"38",
          8103 => x"fe",
          8104 => x"b8",
          8105 => x"33",
          8106 => x"88",
          8107 => x"ba",
          8108 => x"5b",
          8109 => x"04",
          8110 => x"09",
          8111 => x"b8",
          8112 => x"2a",
          8113 => x"05",
          8114 => x"08",
          8115 => x"38",
          8116 => x"18",
          8117 => x"5e",
          8118 => x"2e",
          8119 => x"82",
          8120 => x"54",
          8121 => x"17",
          8122 => x"33",
          8123 => x"3f",
          8124 => x"08",
          8125 => x"38",
          8126 => x"5a",
          8127 => x"0c",
          8128 => x"38",
          8129 => x"83",
          8130 => x"05",
          8131 => x"11",
          8132 => x"33",
          8133 => x"71",
          8134 => x"81",
          8135 => x"72",
          8136 => x"75",
          8137 => x"ff",
          8138 => x"06",
          8139 => x"8c",
          8140 => x"5e",
          8141 => x"8f",
          8142 => x"81",
          8143 => x"08",
          8144 => x"70",
          8145 => x"33",
          8146 => x"e2",
          8147 => x"84",
          8148 => x"7b",
          8149 => x"06",
          8150 => x"84",
          8151 => x"83",
          8152 => x"17",
          8153 => x"08",
          8154 => x"8c",
          8155 => x"7d",
          8156 => x"27",
          8157 => x"82",
          8158 => x"74",
          8159 => x"81",
          8160 => x"38",
          8161 => x"17",
          8162 => x"08",
          8163 => x"52",
          8164 => x"51",
          8165 => x"7a",
          8166 => x"39",
          8167 => x"17",
          8168 => x"17",
          8169 => x"18",
          8170 => x"f6",
          8171 => x"ba",
          8172 => x"2e",
          8173 => x"82",
          8174 => x"ba",
          8175 => x"18",
          8176 => x"08",
          8177 => x"31",
          8178 => x"18",
          8179 => x"38",
          8180 => x"5e",
          8181 => x"81",
          8182 => x"ba",
          8183 => x"fb",
          8184 => x"54",
          8185 => x"53",
          8186 => x"53",
          8187 => x"52",
          8188 => x"3f",
          8189 => x"ba",
          8190 => x"2e",
          8191 => x"fd",
          8192 => x"ba",
          8193 => x"18",
          8194 => x"08",
          8195 => x"31",
          8196 => x"08",
          8197 => x"a0",
          8198 => x"fd",
          8199 => x"17",
          8200 => x"82",
          8201 => x"06",
          8202 => x"81",
          8203 => x"08",
          8204 => x"05",
          8205 => x"81",
          8206 => x"f4",
          8207 => x"5a",
          8208 => x"81",
          8209 => x"08",
          8210 => x"70",
          8211 => x"33",
          8212 => x"da",
          8213 => x"84",
          8214 => x"7d",
          8215 => x"06",
          8216 => x"84",
          8217 => x"83",
          8218 => x"17",
          8219 => x"08",
          8220 => x"8c",
          8221 => x"74",
          8222 => x"27",
          8223 => x"82",
          8224 => x"74",
          8225 => x"81",
          8226 => x"38",
          8227 => x"17",
          8228 => x"08",
          8229 => x"52",
          8230 => x"51",
          8231 => x"7c",
          8232 => x"39",
          8233 => x"17",
          8234 => x"08",
          8235 => x"52",
          8236 => x"51",
          8237 => x"fa",
          8238 => x"5b",
          8239 => x"38",
          8240 => x"f2",
          8241 => x"62",
          8242 => x"59",
          8243 => x"76",
          8244 => x"75",
          8245 => x"27",
          8246 => x"33",
          8247 => x"2e",
          8248 => x"78",
          8249 => x"38",
          8250 => x"82",
          8251 => x"84",
          8252 => x"90",
          8253 => x"75",
          8254 => x"1a",
          8255 => x"80",
          8256 => x"08",
          8257 => x"78",
          8258 => x"38",
          8259 => x"7c",
          8260 => x"7c",
          8261 => x"06",
          8262 => x"81",
          8263 => x"b8",
          8264 => x"19",
          8265 => x"87",
          8266 => x"8c",
          8267 => x"85",
          8268 => x"81",
          8269 => x"1a",
          8270 => x"79",
          8271 => x"75",
          8272 => x"06",
          8273 => x"83",
          8274 => x"58",
          8275 => x"1f",
          8276 => x"2a",
          8277 => x"1f",
          8278 => x"83",
          8279 => x"84",
          8280 => x"90",
          8281 => x"74",
          8282 => x"81",
          8283 => x"38",
          8284 => x"a8",
          8285 => x"58",
          8286 => x"1a",
          8287 => x"76",
          8288 => x"e1",
          8289 => x"33",
          8290 => x"7c",
          8291 => x"81",
          8292 => x"38",
          8293 => x"53",
          8294 => x"81",
          8295 => x"f1",
          8296 => x"ba",
          8297 => x"2e",
          8298 => x"58",
          8299 => x"b4",
          8300 => x"58",
          8301 => x"38",
          8302 => x"83",
          8303 => x"05",
          8304 => x"11",
          8305 => x"2b",
          8306 => x"7e",
          8307 => x"07",
          8308 => x"5c",
          8309 => x"7d",
          8310 => x"75",
          8311 => x"7d",
          8312 => x"79",
          8313 => x"7d",
          8314 => x"7a",
          8315 => x"81",
          8316 => x"34",
          8317 => x"75",
          8318 => x"70",
          8319 => x"1b",
          8320 => x"1b",
          8321 => x"5a",
          8322 => x"b7",
          8323 => x"83",
          8324 => x"5e",
          8325 => x"7d",
          8326 => x"06",
          8327 => x"81",
          8328 => x"b8",
          8329 => x"19",
          8330 => x"83",
          8331 => x"8c",
          8332 => x"85",
          8333 => x"81",
          8334 => x"1a",
          8335 => x"7b",
          8336 => x"79",
          8337 => x"19",
          8338 => x"1b",
          8339 => x"5f",
          8340 => x"55",
          8341 => x"8f",
          8342 => x"2b",
          8343 => x"77",
          8344 => x"71",
          8345 => x"74",
          8346 => x"0b",
          8347 => x"7d",
          8348 => x"1a",
          8349 => x"80",
          8350 => x"08",
          8351 => x"76",
          8352 => x"38",
          8353 => x"53",
          8354 => x"53",
          8355 => x"52",
          8356 => x"3f",
          8357 => x"ba",
          8358 => x"2e",
          8359 => x"80",
          8360 => x"ba",
          8361 => x"1a",
          8362 => x"08",
          8363 => x"08",
          8364 => x"08",
          8365 => x"08",
          8366 => x"5c",
          8367 => x"8b",
          8368 => x"33",
          8369 => x"2e",
          8370 => x"81",
          8371 => x"76",
          8372 => x"33",
          8373 => x"3f",
          8374 => x"08",
          8375 => x"38",
          8376 => x"58",
          8377 => x"0c",
          8378 => x"38",
          8379 => x"06",
          8380 => x"7b",
          8381 => x"56",
          8382 => x"7a",
          8383 => x"33",
          8384 => x"71",
          8385 => x"56",
          8386 => x"34",
          8387 => x"1a",
          8388 => x"39",
          8389 => x"53",
          8390 => x"53",
          8391 => x"52",
          8392 => x"3f",
          8393 => x"ba",
          8394 => x"2e",
          8395 => x"fc",
          8396 => x"ba",
          8397 => x"1a",
          8398 => x"08",
          8399 => x"08",
          8400 => x"08",
          8401 => x"08",
          8402 => x"5e",
          8403 => x"fb",
          8404 => x"19",
          8405 => x"82",
          8406 => x"06",
          8407 => x"81",
          8408 => x"53",
          8409 => x"19",
          8410 => x"c2",
          8411 => x"fb",
          8412 => x"54",
          8413 => x"19",
          8414 => x"1a",
          8415 => x"ee",
          8416 => x"5c",
          8417 => x"08",
          8418 => x"81",
          8419 => x"38",
          8420 => x"08",
          8421 => x"b4",
          8422 => x"a8",
          8423 => x"a0",
          8424 => x"ba",
          8425 => x"40",
          8426 => x"7e",
          8427 => x"38",
          8428 => x"55",
          8429 => x"09",
          8430 => x"e3",
          8431 => x"7d",
          8432 => x"52",
          8433 => x"51",
          8434 => x"7c",
          8435 => x"39",
          8436 => x"53",
          8437 => x"53",
          8438 => x"52",
          8439 => x"3f",
          8440 => x"ba",
          8441 => x"2e",
          8442 => x"fb",
          8443 => x"ba",
          8444 => x"1a",
          8445 => x"08",
          8446 => x"08",
          8447 => x"08",
          8448 => x"08",
          8449 => x"5e",
          8450 => x"fb",
          8451 => x"19",
          8452 => x"82",
          8453 => x"06",
          8454 => x"81",
          8455 => x"53",
          8456 => x"19",
          8457 => x"86",
          8458 => x"fa",
          8459 => x"54",
          8460 => x"76",
          8461 => x"33",
          8462 => x"3f",
          8463 => x"8b",
          8464 => x"10",
          8465 => x"7a",
          8466 => x"ff",
          8467 => x"5f",
          8468 => x"1f",
          8469 => x"2a",
          8470 => x"1f",
          8471 => x"39",
          8472 => x"88",
          8473 => x"82",
          8474 => x"06",
          8475 => x"11",
          8476 => x"70",
          8477 => x"0a",
          8478 => x"0a",
          8479 => x"58",
          8480 => x"7d",
          8481 => x"88",
          8482 => x"b9",
          8483 => x"90",
          8484 => x"ba",
          8485 => x"98",
          8486 => x"bb",
          8487 => x"cf",
          8488 => x"0d",
          8489 => x"08",
          8490 => x"7a",
          8491 => x"90",
          8492 => x"76",
          8493 => x"f4",
          8494 => x"1a",
          8495 => x"ec",
          8496 => x"08",
          8497 => x"73",
          8498 => x"d7",
          8499 => x"2e",
          8500 => x"76",
          8501 => x"56",
          8502 => x"76",
          8503 => x"82",
          8504 => x"26",
          8505 => x"75",
          8506 => x"f0",
          8507 => x"ba",
          8508 => x"2e",
          8509 => x"80",
          8510 => x"8c",
          8511 => x"b1",
          8512 => x"8c",
          8513 => x"30",
          8514 => x"80",
          8515 => x"07",
          8516 => x"55",
          8517 => x"38",
          8518 => x"09",
          8519 => x"b5",
          8520 => x"74",
          8521 => x"0c",
          8522 => x"04",
          8523 => x"91",
          8524 => x"8c",
          8525 => x"39",
          8526 => x"51",
          8527 => x"81",
          8528 => x"ba",
          8529 => x"db",
          8530 => x"8c",
          8531 => x"ba",
          8532 => x"2e",
          8533 => x"19",
          8534 => x"8c",
          8535 => x"38",
          8536 => x"dd",
          8537 => x"56",
          8538 => x"76",
          8539 => x"82",
          8540 => x"79",
          8541 => x"3f",
          8542 => x"ba",
          8543 => x"2e",
          8544 => x"84",
          8545 => x"09",
          8546 => x"72",
          8547 => x"70",
          8548 => x"ba",
          8549 => x"51",
          8550 => x"73",
          8551 => x"84",
          8552 => x"80",
          8553 => x"90",
          8554 => x"81",
          8555 => x"a3",
          8556 => x"1a",
          8557 => x"9b",
          8558 => x"57",
          8559 => x"39",
          8560 => x"fe",
          8561 => x"53",
          8562 => x"51",
          8563 => x"84",
          8564 => x"84",
          8565 => x"30",
          8566 => x"8c",
          8567 => x"25",
          8568 => x"7a",
          8569 => x"74",
          8570 => x"75",
          8571 => x"9c",
          8572 => x"05",
          8573 => x"56",
          8574 => x"26",
          8575 => x"15",
          8576 => x"84",
          8577 => x"07",
          8578 => x"1a",
          8579 => x"74",
          8580 => x"0c",
          8581 => x"04",
          8582 => x"ba",
          8583 => x"3d",
          8584 => x"ba",
          8585 => x"fe",
          8586 => x"80",
          8587 => x"38",
          8588 => x"52",
          8589 => x"8b",
          8590 => x"8c",
          8591 => x"a7",
          8592 => x"8c",
          8593 => x"8c",
          8594 => x"0d",
          8595 => x"74",
          8596 => x"b9",
          8597 => x"ff",
          8598 => x"3d",
          8599 => x"71",
          8600 => x"58",
          8601 => x"0a",
          8602 => x"38",
          8603 => x"53",
          8604 => x"38",
          8605 => x"0c",
          8606 => x"55",
          8607 => x"38",
          8608 => x"75",
          8609 => x"cc",
          8610 => x"2a",
          8611 => x"88",
          8612 => x"56",
          8613 => x"a9",
          8614 => x"08",
          8615 => x"74",
          8616 => x"98",
          8617 => x"82",
          8618 => x"2e",
          8619 => x"89",
          8620 => x"19",
          8621 => x"ff",
          8622 => x"05",
          8623 => x"80",
          8624 => x"ba",
          8625 => x"3d",
          8626 => x"0b",
          8627 => x"0c",
          8628 => x"04",
          8629 => x"55",
          8630 => x"ff",
          8631 => x"17",
          8632 => x"2b",
          8633 => x"76",
          8634 => x"9c",
          8635 => x"fe",
          8636 => x"54",
          8637 => x"75",
          8638 => x"38",
          8639 => x"76",
          8640 => x"19",
          8641 => x"53",
          8642 => x"0c",
          8643 => x"74",
          8644 => x"ec",
          8645 => x"ba",
          8646 => x"84",
          8647 => x"ff",
          8648 => x"81",
          8649 => x"8c",
          8650 => x"9e",
          8651 => x"08",
          8652 => x"8c",
          8653 => x"ff",
          8654 => x"76",
          8655 => x"76",
          8656 => x"ff",
          8657 => x"0b",
          8658 => x"0c",
          8659 => x"04",
          8660 => x"7f",
          8661 => x"12",
          8662 => x"5c",
          8663 => x"80",
          8664 => x"86",
          8665 => x"98",
          8666 => x"17",
          8667 => x"56",
          8668 => x"b2",
          8669 => x"ff",
          8670 => x"9d",
          8671 => x"94",
          8672 => x"58",
          8673 => x"79",
          8674 => x"1a",
          8675 => x"74",
          8676 => x"f5",
          8677 => x"18",
          8678 => x"18",
          8679 => x"b8",
          8680 => x"0c",
          8681 => x"84",
          8682 => x"8f",
          8683 => x"77",
          8684 => x"8a",
          8685 => x"05",
          8686 => x"06",
          8687 => x"38",
          8688 => x"51",
          8689 => x"84",
          8690 => x"5d",
          8691 => x"0b",
          8692 => x"08",
          8693 => x"81",
          8694 => x"8c",
          8695 => x"c6",
          8696 => x"08",
          8697 => x"08",
          8698 => x"38",
          8699 => x"81",
          8700 => x"17",
          8701 => x"51",
          8702 => x"84",
          8703 => x"5d",
          8704 => x"ba",
          8705 => x"2e",
          8706 => x"82",
          8707 => x"8c",
          8708 => x"ff",
          8709 => x"56",
          8710 => x"08",
          8711 => x"86",
          8712 => x"8c",
          8713 => x"33",
          8714 => x"80",
          8715 => x"18",
          8716 => x"fe",
          8717 => x"80",
          8718 => x"27",
          8719 => x"19",
          8720 => x"29",
          8721 => x"05",
          8722 => x"b4",
          8723 => x"19",
          8724 => x"78",
          8725 => x"76",
          8726 => x"58",
          8727 => x"55",
          8728 => x"74",
          8729 => x"22",
          8730 => x"27",
          8731 => x"81",
          8732 => x"53",
          8733 => x"19",
          8734 => x"b2",
          8735 => x"8c",
          8736 => x"38",
          8737 => x"dd",
          8738 => x"18",
          8739 => x"84",
          8740 => x"8f",
          8741 => x"75",
          8742 => x"08",
          8743 => x"70",
          8744 => x"33",
          8745 => x"86",
          8746 => x"8c",
          8747 => x"38",
          8748 => x"08",
          8749 => x"b4",
          8750 => x"1a",
          8751 => x"74",
          8752 => x"27",
          8753 => x"82",
          8754 => x"7b",
          8755 => x"81",
          8756 => x"38",
          8757 => x"19",
          8758 => x"08",
          8759 => x"52",
          8760 => x"51",
          8761 => x"fe",
          8762 => x"19",
          8763 => x"83",
          8764 => x"55",
          8765 => x"09",
          8766 => x"38",
          8767 => x"0c",
          8768 => x"1a",
          8769 => x"5e",
          8770 => x"75",
          8771 => x"85",
          8772 => x"22",
          8773 => x"b0",
          8774 => x"98",
          8775 => x"fc",
          8776 => x"0b",
          8777 => x"0c",
          8778 => x"04",
          8779 => x"64",
          8780 => x"84",
          8781 => x"5b",
          8782 => x"98",
          8783 => x"5e",
          8784 => x"2e",
          8785 => x"b8",
          8786 => x"5a",
          8787 => x"19",
          8788 => x"82",
          8789 => x"19",
          8790 => x"55",
          8791 => x"09",
          8792 => x"94",
          8793 => x"75",
          8794 => x"52",
          8795 => x"51",
          8796 => x"84",
          8797 => x"80",
          8798 => x"ff",
          8799 => x"79",
          8800 => x"76",
          8801 => x"90",
          8802 => x"08",
          8803 => x"58",
          8804 => x"82",
          8805 => x"18",
          8806 => x"70",
          8807 => x"5b",
          8808 => x"1d",
          8809 => x"e5",
          8810 => x"78",
          8811 => x"30",
          8812 => x"71",
          8813 => x"54",
          8814 => x"55",
          8815 => x"74",
          8816 => x"43",
          8817 => x"2e",
          8818 => x"75",
          8819 => x"86",
          8820 => x"5d",
          8821 => x"51",
          8822 => x"84",
          8823 => x"5b",
          8824 => x"08",
          8825 => x"98",
          8826 => x"75",
          8827 => x"7a",
          8828 => x"0c",
          8829 => x"04",
          8830 => x"19",
          8831 => x"52",
          8832 => x"51",
          8833 => x"81",
          8834 => x"8c",
          8835 => x"09",
          8836 => x"ef",
          8837 => x"8c",
          8838 => x"34",
          8839 => x"a8",
          8840 => x"84",
          8841 => x"58",
          8842 => x"1a",
          8843 => x"b5",
          8844 => x"33",
          8845 => x"2e",
          8846 => x"fe",
          8847 => x"54",
          8848 => x"a0",
          8849 => x"53",
          8850 => x"19",
          8851 => x"de",
          8852 => x"fe",
          8853 => x"8f",
          8854 => x"06",
          8855 => x"76",
          8856 => x"06",
          8857 => x"2e",
          8858 => x"18",
          8859 => x"bf",
          8860 => x"1f",
          8861 => x"05",
          8862 => x"5e",
          8863 => x"ab",
          8864 => x"55",
          8865 => x"cc",
          8866 => x"75",
          8867 => x"81",
          8868 => x"38",
          8869 => x"5b",
          8870 => x"1d",
          8871 => x"ba",
          8872 => x"3d",
          8873 => x"5b",
          8874 => x"8d",
          8875 => x"7d",
          8876 => x"81",
          8877 => x"8c",
          8878 => x"19",
          8879 => x"33",
          8880 => x"07",
          8881 => x"75",
          8882 => x"77",
          8883 => x"bf",
          8884 => x"f3",
          8885 => x"81",
          8886 => x"83",
          8887 => x"33",
          8888 => x"11",
          8889 => x"71",
          8890 => x"52",
          8891 => x"80",
          8892 => x"38",
          8893 => x"26",
          8894 => x"79",
          8895 => x"76",
          8896 => x"62",
          8897 => x"5a",
          8898 => x"8c",
          8899 => x"38",
          8900 => x"86",
          8901 => x"59",
          8902 => x"2e",
          8903 => x"81",
          8904 => x"dd",
          8905 => x"61",
          8906 => x"63",
          8907 => x"70",
          8908 => x"5e",
          8909 => x"39",
          8910 => x"ff",
          8911 => x"81",
          8912 => x"c0",
          8913 => x"38",
          8914 => x"57",
          8915 => x"75",
          8916 => x"05",
          8917 => x"05",
          8918 => x"7f",
          8919 => x"ff",
          8920 => x"59",
          8921 => x"e4",
          8922 => x"2e",
          8923 => x"ff",
          8924 => x"0c",
          8925 => x"8c",
          8926 => x"0d",
          8927 => x"0d",
          8928 => x"5c",
          8929 => x"7b",
          8930 => x"3f",
          8931 => x"08",
          8932 => x"8c",
          8933 => x"38",
          8934 => x"40",
          8935 => x"ac",
          8936 => x"1b",
          8937 => x"08",
          8938 => x"b4",
          8939 => x"2e",
          8940 => x"83",
          8941 => x"58",
          8942 => x"2e",
          8943 => x"81",
          8944 => x"54",
          8945 => x"1b",
          8946 => x"33",
          8947 => x"3f",
          8948 => x"08",
          8949 => x"38",
          8950 => x"57",
          8951 => x"0c",
          8952 => x"81",
          8953 => x"1c",
          8954 => x"58",
          8955 => x"2e",
          8956 => x"8b",
          8957 => x"06",
          8958 => x"06",
          8959 => x"86",
          8960 => x"81",
          8961 => x"f2",
          8962 => x"2a",
          8963 => x"75",
          8964 => x"ef",
          8965 => x"e2",
          8966 => x"2e",
          8967 => x"7c",
          8968 => x"7d",
          8969 => x"57",
          8970 => x"75",
          8971 => x"05",
          8972 => x"05",
          8973 => x"76",
          8974 => x"ff",
          8975 => x"59",
          8976 => x"e4",
          8977 => x"2e",
          8978 => x"ab",
          8979 => x"06",
          8980 => x"38",
          8981 => x"1d",
          8982 => x"70",
          8983 => x"33",
          8984 => x"05",
          8985 => x"71",
          8986 => x"5a",
          8987 => x"76",
          8988 => x"dc",
          8989 => x"2e",
          8990 => x"ff",
          8991 => x"ac",
          8992 => x"52",
          8993 => x"c8",
          8994 => x"8c",
          8995 => x"ba",
          8996 => x"2e",
          8997 => x"79",
          8998 => x"0c",
          8999 => x"04",
          9000 => x"1b",
          9001 => x"52",
          9002 => x"51",
          9003 => x"81",
          9004 => x"8c",
          9005 => x"09",
          9006 => x"a4",
          9007 => x"8c",
          9008 => x"34",
          9009 => x"a8",
          9010 => x"84",
          9011 => x"58",
          9012 => x"1c",
          9013 => x"ea",
          9014 => x"33",
          9015 => x"2e",
          9016 => x"fd",
          9017 => x"54",
          9018 => x"a0",
          9019 => x"53",
          9020 => x"1b",
          9021 => x"b6",
          9022 => x"fd",
          9023 => x"5a",
          9024 => x"ab",
          9025 => x"86",
          9026 => x"42",
          9027 => x"f2",
          9028 => x"2a",
          9029 => x"79",
          9030 => x"38",
          9031 => x"77",
          9032 => x"70",
          9033 => x"7f",
          9034 => x"59",
          9035 => x"7d",
          9036 => x"81",
          9037 => x"5d",
          9038 => x"51",
          9039 => x"84",
          9040 => x"5a",
          9041 => x"08",
          9042 => x"d9",
          9043 => x"39",
          9044 => x"fe",
          9045 => x"ff",
          9046 => x"ac",
          9047 => x"a2",
          9048 => x"33",
          9049 => x"2e",
          9050 => x"c7",
          9051 => x"08",
          9052 => x"9a",
          9053 => x"88",
          9054 => x"42",
          9055 => x"b3",
          9056 => x"70",
          9057 => x"29",
          9058 => x"55",
          9059 => x"56",
          9060 => x"18",
          9061 => x"81",
          9062 => x"33",
          9063 => x"07",
          9064 => x"75",
          9065 => x"ed",
          9066 => x"fe",
          9067 => x"38",
          9068 => x"a1",
          9069 => x"ba",
          9070 => x"10",
          9071 => x"22",
          9072 => x"1b",
          9073 => x"a0",
          9074 => x"84",
          9075 => x"2e",
          9076 => x"fe",
          9077 => x"56",
          9078 => x"8c",
          9079 => x"b0",
          9080 => x"70",
          9081 => x"06",
          9082 => x"80",
          9083 => x"74",
          9084 => x"38",
          9085 => x"05",
          9086 => x"41",
          9087 => x"38",
          9088 => x"81",
          9089 => x"5a",
          9090 => x"84",
          9091 => x"8c",
          9092 => x"0d",
          9093 => x"ff",
          9094 => x"bc",
          9095 => x"55",
          9096 => x"ea",
          9097 => x"70",
          9098 => x"13",
          9099 => x"06",
          9100 => x"5e",
          9101 => x"85",
          9102 => x"8c",
          9103 => x"22",
          9104 => x"74",
          9105 => x"38",
          9106 => x"10",
          9107 => x"51",
          9108 => x"f4",
          9109 => x"a0",
          9110 => x"8c",
          9111 => x"58",
          9112 => x"81",
          9113 => x"77",
          9114 => x"59",
          9115 => x"55",
          9116 => x"02",
          9117 => x"33",
          9118 => x"58",
          9119 => x"2e",
          9120 => x"80",
          9121 => x"1f",
          9122 => x"94",
          9123 => x"8c",
          9124 => x"58",
          9125 => x"61",
          9126 => x"77",
          9127 => x"59",
          9128 => x"81",
          9129 => x"ff",
          9130 => x"ef",
          9131 => x"27",
          9132 => x"7a",
          9133 => x"57",
          9134 => x"b8",
          9135 => x"1a",
          9136 => x"58",
          9137 => x"77",
          9138 => x"81",
          9139 => x"ff",
          9140 => x"90",
          9141 => x"44",
          9142 => x"60",
          9143 => x"38",
          9144 => x"a1",
          9145 => x"18",
          9146 => x"25",
          9147 => x"22",
          9148 => x"38",
          9149 => x"05",
          9150 => x"57",
          9151 => x"07",
          9152 => x"b9",
          9153 => x"38",
          9154 => x"74",
          9155 => x"16",
          9156 => x"84",
          9157 => x"56",
          9158 => x"77",
          9159 => x"fe",
          9160 => x"7a",
          9161 => x"78",
          9162 => x"79",
          9163 => x"a0",
          9164 => x"81",
          9165 => x"78",
          9166 => x"38",
          9167 => x"33",
          9168 => x"a0",
          9169 => x"06",
          9170 => x"16",
          9171 => x"77",
          9172 => x"38",
          9173 => x"05",
          9174 => x"19",
          9175 => x"59",
          9176 => x"34",
          9177 => x"87",
          9178 => x"51",
          9179 => x"84",
          9180 => x"8b",
          9181 => x"5b",
          9182 => x"27",
          9183 => x"87",
          9184 => x"e4",
          9185 => x"38",
          9186 => x"08",
          9187 => x"8c",
          9188 => x"09",
          9189 => x"d6",
          9190 => x"db",
          9191 => x"1f",
          9192 => x"02",
          9193 => x"db",
          9194 => x"58",
          9195 => x"81",
          9196 => x"5b",
          9197 => x"90",
          9198 => x"8c",
          9199 => x"89",
          9200 => x"ba",
          9201 => x"5b",
          9202 => x"51",
          9203 => x"84",
          9204 => x"56",
          9205 => x"08",
          9206 => x"84",
          9207 => x"b8",
          9208 => x"98",
          9209 => x"80",
          9210 => x"08",
          9211 => x"f3",
          9212 => x"33",
          9213 => x"2e",
          9214 => x"82",
          9215 => x"54",
          9216 => x"18",
          9217 => x"33",
          9218 => x"3f",
          9219 => x"08",
          9220 => x"38",
          9221 => x"57",
          9222 => x"0c",
          9223 => x"bc",
          9224 => x"08",
          9225 => x"42",
          9226 => x"2e",
          9227 => x"74",
          9228 => x"25",
          9229 => x"5f",
          9230 => x"81",
          9231 => x"19",
          9232 => x"2e",
          9233 => x"81",
          9234 => x"ee",
          9235 => x"ba",
          9236 => x"84",
          9237 => x"80",
          9238 => x"38",
          9239 => x"84",
          9240 => x"38",
          9241 => x"81",
          9242 => x"1b",
          9243 => x"f3",
          9244 => x"08",
          9245 => x"08",
          9246 => x"38",
          9247 => x"78",
          9248 => x"84",
          9249 => x"54",
          9250 => x"1c",
          9251 => x"33",
          9252 => x"3f",
          9253 => x"08",
          9254 => x"38",
          9255 => x"56",
          9256 => x"0c",
          9257 => x"80",
          9258 => x"0b",
          9259 => x"57",
          9260 => x"70",
          9261 => x"34",
          9262 => x"74",
          9263 => x"0b",
          9264 => x"7b",
          9265 => x"75",
          9266 => x"57",
          9267 => x"81",
          9268 => x"ff",
          9269 => x"ef",
          9270 => x"08",
          9271 => x"98",
          9272 => x"7c",
          9273 => x"81",
          9274 => x"34",
          9275 => x"84",
          9276 => x"98",
          9277 => x"81",
          9278 => x"80",
          9279 => x"57",
          9280 => x"fe",
          9281 => x"59",
          9282 => x"51",
          9283 => x"84",
          9284 => x"56",
          9285 => x"08",
          9286 => x"c7",
          9287 => x"39",
          9288 => x"18",
          9289 => x"52",
          9290 => x"51",
          9291 => x"84",
          9292 => x"77",
          9293 => x"06",
          9294 => x"84",
          9295 => x"83",
          9296 => x"18",
          9297 => x"08",
          9298 => x"a0",
          9299 => x"8b",
          9300 => x"33",
          9301 => x"2e",
          9302 => x"84",
          9303 => x"57",
          9304 => x"7f",
          9305 => x"1f",
          9306 => x"53",
          9307 => x"e9",
          9308 => x"ba",
          9309 => x"84",
          9310 => x"fe",
          9311 => x"84",
          9312 => x"56",
          9313 => x"74",
          9314 => x"81",
          9315 => x"78",
          9316 => x"5a",
          9317 => x"05",
          9318 => x"06",
          9319 => x"56",
          9320 => x"38",
          9321 => x"06",
          9322 => x"41",
          9323 => x"57",
          9324 => x"1c",
          9325 => x"b2",
          9326 => x"33",
          9327 => x"2e",
          9328 => x"82",
          9329 => x"54",
          9330 => x"1c",
          9331 => x"33",
          9332 => x"3f",
          9333 => x"08",
          9334 => x"38",
          9335 => x"56",
          9336 => x"0c",
          9337 => x"fe",
          9338 => x"1c",
          9339 => x"08",
          9340 => x"06",
          9341 => x"60",
          9342 => x"8f",
          9343 => x"34",
          9344 => x"34",
          9345 => x"34",
          9346 => x"34",
          9347 => x"f3",
          9348 => x"5a",
          9349 => x"83",
          9350 => x"8b",
          9351 => x"1f",
          9352 => x"1b",
          9353 => x"83",
          9354 => x"33",
          9355 => x"76",
          9356 => x"05",
          9357 => x"88",
          9358 => x"75",
          9359 => x"38",
          9360 => x"57",
          9361 => x"8c",
          9362 => x"38",
          9363 => x"ff",
          9364 => x"38",
          9365 => x"70",
          9366 => x"76",
          9367 => x"a6",
          9368 => x"34",
          9369 => x"1d",
          9370 => x"7d",
          9371 => x"3f",
          9372 => x"08",
          9373 => x"8c",
          9374 => x"38",
          9375 => x"40",
          9376 => x"38",
          9377 => x"81",
          9378 => x"08",
          9379 => x"70",
          9380 => x"33",
          9381 => x"96",
          9382 => x"84",
          9383 => x"fc",
          9384 => x"ba",
          9385 => x"1d",
          9386 => x"08",
          9387 => x"31",
          9388 => x"08",
          9389 => x"a0",
          9390 => x"fb",
          9391 => x"1c",
          9392 => x"82",
          9393 => x"06",
          9394 => x"81",
          9395 => x"08",
          9396 => x"05",
          9397 => x"81",
          9398 => x"cf",
          9399 => x"56",
          9400 => x"76",
          9401 => x"70",
          9402 => x"56",
          9403 => x"2e",
          9404 => x"fa",
          9405 => x"ff",
          9406 => x"57",
          9407 => x"2e",
          9408 => x"fa",
          9409 => x"80",
          9410 => x"fe",
          9411 => x"54",
          9412 => x"53",
          9413 => x"1c",
          9414 => x"92",
          9415 => x"8c",
          9416 => x"09",
          9417 => x"38",
          9418 => x"08",
          9419 => x"b4",
          9420 => x"1d",
          9421 => x"74",
          9422 => x"27",
          9423 => x"1c",
          9424 => x"82",
          9425 => x"84",
          9426 => x"56",
          9427 => x"75",
          9428 => x"58",
          9429 => x"fa",
          9430 => x"87",
          9431 => x"57",
          9432 => x"81",
          9433 => x"75",
          9434 => x"fe",
          9435 => x"39",
          9436 => x"1c",
          9437 => x"08",
          9438 => x"52",
          9439 => x"51",
          9440 => x"fc",
          9441 => x"54",
          9442 => x"a0",
          9443 => x"53",
          9444 => x"18",
          9445 => x"96",
          9446 => x"39",
          9447 => x"7f",
          9448 => x"40",
          9449 => x"0b",
          9450 => x"98",
          9451 => x"2e",
          9452 => x"ac",
          9453 => x"2e",
          9454 => x"80",
          9455 => x"8c",
          9456 => x"22",
          9457 => x"5c",
          9458 => x"2e",
          9459 => x"54",
          9460 => x"22",
          9461 => x"55",
          9462 => x"95",
          9463 => x"80",
          9464 => x"ff",
          9465 => x"5a",
          9466 => x"26",
          9467 => x"73",
          9468 => x"11",
          9469 => x"58",
          9470 => x"d4",
          9471 => x"70",
          9472 => x"30",
          9473 => x"5c",
          9474 => x"94",
          9475 => x"0b",
          9476 => x"80",
          9477 => x"59",
          9478 => x"1c",
          9479 => x"33",
          9480 => x"56",
          9481 => x"2e",
          9482 => x"85",
          9483 => x"38",
          9484 => x"70",
          9485 => x"07",
          9486 => x"5b",
          9487 => x"26",
          9488 => x"80",
          9489 => x"ae",
          9490 => x"05",
          9491 => x"18",
          9492 => x"70",
          9493 => x"34",
          9494 => x"8a",
          9495 => x"ba",
          9496 => x"88",
          9497 => x"0b",
          9498 => x"96",
          9499 => x"72",
          9500 => x"81",
          9501 => x"0b",
          9502 => x"81",
          9503 => x"94",
          9504 => x"0b",
          9505 => x"9c",
          9506 => x"11",
          9507 => x"73",
          9508 => x"89",
          9509 => x"1c",
          9510 => x"13",
          9511 => x"34",
          9512 => x"9c",
          9513 => x"33",
          9514 => x"71",
          9515 => x"88",
          9516 => x"14",
          9517 => x"07",
          9518 => x"33",
          9519 => x"0c",
          9520 => x"33",
          9521 => x"71",
          9522 => x"5f",
          9523 => x"5a",
          9524 => x"77",
          9525 => x"99",
          9526 => x"16",
          9527 => x"2b",
          9528 => x"7b",
          9529 => x"8f",
          9530 => x"81",
          9531 => x"c0",
          9532 => x"96",
          9533 => x"7a",
          9534 => x"57",
          9535 => x"7a",
          9536 => x"07",
          9537 => x"89",
          9538 => x"8c",
          9539 => x"ff",
          9540 => x"ff",
          9541 => x"38",
          9542 => x"81",
          9543 => x"88",
          9544 => x"7a",
          9545 => x"18",
          9546 => x"05",
          9547 => x"8c",
          9548 => x"5b",
          9549 => x"11",
          9550 => x"57",
          9551 => x"90",
          9552 => x"39",
          9553 => x"30",
          9554 => x"80",
          9555 => x"25",
          9556 => x"57",
          9557 => x"38",
          9558 => x"81",
          9559 => x"80",
          9560 => x"08",
          9561 => x"39",
          9562 => x"1f",
          9563 => x"57",
          9564 => x"fe",
          9565 => x"96",
          9566 => x"59",
          9567 => x"33",
          9568 => x"5a",
          9569 => x"26",
          9570 => x"1c",
          9571 => x"33",
          9572 => x"76",
          9573 => x"72",
          9574 => x"72",
          9575 => x"7d",
          9576 => x"38",
          9577 => x"83",
          9578 => x"55",
          9579 => x"70",
          9580 => x"34",
          9581 => x"16",
          9582 => x"89",
          9583 => x"57",
          9584 => x"79",
          9585 => x"fd",
          9586 => x"83",
          9587 => x"39",
          9588 => x"70",
          9589 => x"30",
          9590 => x"5d",
          9591 => x"a9",
          9592 => x"0d",
          9593 => x"70",
          9594 => x"80",
          9595 => x"57",
          9596 => x"af",
          9597 => x"81",
          9598 => x"dc",
          9599 => x"38",
          9600 => x"81",
          9601 => x"16",
          9602 => x"0c",
          9603 => x"3d",
          9604 => x"42",
          9605 => x"27",
          9606 => x"73",
          9607 => x"08",
          9608 => x"61",
          9609 => x"05",
          9610 => x"53",
          9611 => x"38",
          9612 => x"73",
          9613 => x"ec",
          9614 => x"ff",
          9615 => x"38",
          9616 => x"56",
          9617 => x"81",
          9618 => x"83",
          9619 => x"70",
          9620 => x"30",
          9621 => x"71",
          9622 => x"57",
          9623 => x"73",
          9624 => x"74",
          9625 => x"82",
          9626 => x"80",
          9627 => x"38",
          9628 => x"0b",
          9629 => x"33",
          9630 => x"06",
          9631 => x"73",
          9632 => x"ab",
          9633 => x"2e",
          9634 => x"16",
          9635 => x"81",
          9636 => x"54",
          9637 => x"38",
          9638 => x"06",
          9639 => x"84",
          9640 => x"fe",
          9641 => x"38",
          9642 => x"5d",
          9643 => x"81",
          9644 => x"70",
          9645 => x"33",
          9646 => x"73",
          9647 => x"f0",
          9648 => x"39",
          9649 => x"dc",
          9650 => x"70",
          9651 => x"07",
          9652 => x"55",
          9653 => x"a1",
          9654 => x"70",
          9655 => x"74",
          9656 => x"72",
          9657 => x"38",
          9658 => x"32",
          9659 => x"80",
          9660 => x"51",
          9661 => x"e1",
          9662 => x"1d",
          9663 => x"96",
          9664 => x"41",
          9665 => x"9f",
          9666 => x"38",
          9667 => x"b5",
          9668 => x"81",
          9669 => x"84",
          9670 => x"83",
          9671 => x"54",
          9672 => x"38",
          9673 => x"84",
          9674 => x"93",
          9675 => x"83",
          9676 => x"70",
          9677 => x"5c",
          9678 => x"2e",
          9679 => x"e4",
          9680 => x"0b",
          9681 => x"80",
          9682 => x"de",
          9683 => x"ba",
          9684 => x"ba",
          9685 => x"3d",
          9686 => x"73",
          9687 => x"70",
          9688 => x"25",
          9689 => x"55",
          9690 => x"80",
          9691 => x"81",
          9692 => x"62",
          9693 => x"55",
          9694 => x"2e",
          9695 => x"80",
          9696 => x"30",
          9697 => x"78",
          9698 => x"59",
          9699 => x"73",
          9700 => x"75",
          9701 => x"5a",
          9702 => x"84",
          9703 => x"82",
          9704 => x"38",
          9705 => x"76",
          9706 => x"38",
          9707 => x"11",
          9708 => x"22",
          9709 => x"70",
          9710 => x"2a",
          9711 => x"5f",
          9712 => x"ae",
          9713 => x"72",
          9714 => x"17",
          9715 => x"38",
          9716 => x"19",
          9717 => x"23",
          9718 => x"fe",
          9719 => x"78",
          9720 => x"ff",
          9721 => x"58",
          9722 => x"7a",
          9723 => x"e6",
          9724 => x"ff",
          9725 => x"72",
          9726 => x"f1",
          9727 => x"2e",
          9728 => x"19",
          9729 => x"22",
          9730 => x"ae",
          9731 => x"76",
          9732 => x"05",
          9733 => x"57",
          9734 => x"8f",
          9735 => x"70",
          9736 => x"7c",
          9737 => x"81",
          9738 => x"8b",
          9739 => x"55",
          9740 => x"70",
          9741 => x"34",
          9742 => x"72",
          9743 => x"73",
          9744 => x"78",
          9745 => x"81",
          9746 => x"54",
          9747 => x"2e",
          9748 => x"74",
          9749 => x"d0",
          9750 => x"32",
          9751 => x"80",
          9752 => x"54",
          9753 => x"85",
          9754 => x"83",
          9755 => x"59",
          9756 => x"83",
          9757 => x"75",
          9758 => x"30",
          9759 => x"80",
          9760 => x"07",
          9761 => x"54",
          9762 => x"83",
          9763 => x"8b",
          9764 => x"38",
          9765 => x"8a",
          9766 => x"07",
          9767 => x"26",
          9768 => x"56",
          9769 => x"7e",
          9770 => x"fc",
          9771 => x"57",
          9772 => x"15",
          9773 => x"18",
          9774 => x"74",
          9775 => x"a0",
          9776 => x"76",
          9777 => x"83",
          9778 => x"88",
          9779 => x"38",
          9780 => x"58",
          9781 => x"82",
          9782 => x"83",
          9783 => x"83",
          9784 => x"38",
          9785 => x"81",
          9786 => x"9d",
          9787 => x"06",
          9788 => x"2e",
          9789 => x"90",
          9790 => x"82",
          9791 => x"5e",
          9792 => x"85",
          9793 => x"07",
          9794 => x"1d",
          9795 => x"e4",
          9796 => x"ba",
          9797 => x"1d",
          9798 => x"84",
          9799 => x"80",
          9800 => x"38",
          9801 => x"08",
          9802 => x"81",
          9803 => x"38",
          9804 => x"81",
          9805 => x"80",
          9806 => x"38",
          9807 => x"81",
          9808 => x"82",
          9809 => x"08",
          9810 => x"73",
          9811 => x"08",
          9812 => x"f9",
          9813 => x"16",
          9814 => x"11",
          9815 => x"40",
          9816 => x"a0",
          9817 => x"75",
          9818 => x"85",
          9819 => x"07",
          9820 => x"39",
          9821 => x"56",
          9822 => x"09",
          9823 => x"ac",
          9824 => x"54",
          9825 => x"09",
          9826 => x"a0",
          9827 => x"18",
          9828 => x"23",
          9829 => x"1d",
          9830 => x"54",
          9831 => x"83",
          9832 => x"73",
          9833 => x"05",
          9834 => x"13",
          9835 => x"27",
          9836 => x"a0",
          9837 => x"ab",
          9838 => x"51",
          9839 => x"84",
          9840 => x"ab",
          9841 => x"54",
          9842 => x"08",
          9843 => x"74",
          9844 => x"06",
          9845 => x"ce",
          9846 => x"33",
          9847 => x"81",
          9848 => x"74",
          9849 => x"cd",
          9850 => x"08",
          9851 => x"60",
          9852 => x"11",
          9853 => x"12",
          9854 => x"2b",
          9855 => x"41",
          9856 => x"7d",
          9857 => x"d8",
          9858 => x"1d",
          9859 => x"65",
          9860 => x"b7",
          9861 => x"55",
          9862 => x"fe",
          9863 => x"17",
          9864 => x"88",
          9865 => x"39",
          9866 => x"76",
          9867 => x"fd",
          9868 => x"82",
          9869 => x"06",
          9870 => x"59",
          9871 => x"2e",
          9872 => x"fd",
          9873 => x"82",
          9874 => x"98",
          9875 => x"a0",
          9876 => x"88",
          9877 => x"06",
          9878 => x"d6",
          9879 => x"0b",
          9880 => x"80",
          9881 => x"8c",
          9882 => x"0d",
          9883 => x"ff",
          9884 => x"81",
          9885 => x"80",
          9886 => x"1d",
          9887 => x"26",
          9888 => x"79",
          9889 => x"77",
          9890 => x"5a",
          9891 => x"79",
          9892 => x"83",
          9893 => x"51",
          9894 => x"3f",
          9895 => x"08",
          9896 => x"06",
          9897 => x"81",
          9898 => x"78",
          9899 => x"38",
          9900 => x"06",
          9901 => x"11",
          9902 => x"74",
          9903 => x"ff",
          9904 => x"80",
          9905 => x"38",
          9906 => x"0b",
          9907 => x"33",
          9908 => x"06",
          9909 => x"73",
          9910 => x"e0",
          9911 => x"2e",
          9912 => x"19",
          9913 => x"81",
          9914 => x"54",
          9915 => x"38",
          9916 => x"06",
          9917 => x"d4",
          9918 => x"15",
          9919 => x"26",
          9920 => x"82",
          9921 => x"ff",
          9922 => x"ff",
          9923 => x"78",
          9924 => x"38",
          9925 => x"70",
          9926 => x"e0",
          9927 => x"ff",
          9928 => x"56",
          9929 => x"1b",
          9930 => x"74",
          9931 => x"1b",
          9932 => x"55",
          9933 => x"80",
          9934 => x"39",
          9935 => x"33",
          9936 => x"06",
          9937 => x"80",
          9938 => x"38",
          9939 => x"83",
          9940 => x"a0",
          9941 => x"55",
          9942 => x"81",
          9943 => x"39",
          9944 => x"33",
          9945 => x"33",
          9946 => x"71",
          9947 => x"77",
          9948 => x"0c",
          9949 => x"95",
          9950 => x"a0",
          9951 => x"2a",
          9952 => x"74",
          9953 => x"7c",
          9954 => x"5a",
          9955 => x"34",
          9956 => x"ff",
          9957 => x"83",
          9958 => x"33",
          9959 => x"81",
          9960 => x"81",
          9961 => x"38",
          9962 => x"74",
          9963 => x"06",
          9964 => x"f2",
          9965 => x"84",
          9966 => x"93",
          9967 => x"eb",
          9968 => x"69",
          9969 => x"80",
          9970 => x"42",
          9971 => x"61",
          9972 => x"08",
          9973 => x"42",
          9974 => x"85",
          9975 => x"70",
          9976 => x"33",
          9977 => x"56",
          9978 => x"2e",
          9979 => x"74",
          9980 => x"ba",
          9981 => x"38",
          9982 => x"33",
          9983 => x"24",
          9984 => x"75",
          9985 => x"d1",
          9986 => x"08",
          9987 => x"58",
          9988 => x"85",
          9989 => x"61",
          9990 => x"fe",
          9991 => x"5d",
          9992 => x"2e",
          9993 => x"17",
          9994 => x"bb",
          9995 => x"ba",
          9996 => x"ff",
          9997 => x"06",
          9998 => x"80",
          9999 => x"38",
         10000 => x"75",
         10001 => x"ba",
         10002 => x"81",
         10003 => x"52",
         10004 => x"51",
         10005 => x"3f",
         10006 => x"08",
         10007 => x"70",
         10008 => x"56",
         10009 => x"84",
         10010 => x"80",
         10011 => x"75",
         10012 => x"06",
         10013 => x"60",
         10014 => x"80",
         10015 => x"18",
         10016 => x"b4",
         10017 => x"7b",
         10018 => x"54",
         10019 => x"17",
         10020 => x"18",
         10021 => x"ff",
         10022 => x"84",
         10023 => x"7b",
         10024 => x"ff",
         10025 => x"74",
         10026 => x"84",
         10027 => x"38",
         10028 => x"33",
         10029 => x"33",
         10030 => x"07",
         10031 => x"56",
         10032 => x"d5",
         10033 => x"38",
         10034 => x"8b",
         10035 => x"81",
         10036 => x"61",
         10037 => x"81",
         10038 => x"2e",
         10039 => x"8d",
         10040 => x"26",
         10041 => x"80",
         10042 => x"80",
         10043 => x"71",
         10044 => x"5e",
         10045 => x"80",
         10046 => x"06",
         10047 => x"80",
         10048 => x"80",
         10049 => x"71",
         10050 => x"57",
         10051 => x"38",
         10052 => x"83",
         10053 => x"12",
         10054 => x"2b",
         10055 => x"07",
         10056 => x"70",
         10057 => x"2b",
         10058 => x"07",
         10059 => x"43",
         10060 => x"75",
         10061 => x"80",
         10062 => x"82",
         10063 => x"c8",
         10064 => x"11",
         10065 => x"06",
         10066 => x"8d",
         10067 => x"26",
         10068 => x"78",
         10069 => x"76",
         10070 => x"c5",
         10071 => x"5f",
         10072 => x"18",
         10073 => x"77",
         10074 => x"c4",
         10075 => x"78",
         10076 => x"87",
         10077 => x"ca",
         10078 => x"c9",
         10079 => x"88",
         10080 => x"40",
         10081 => x"23",
         10082 => x"06",
         10083 => x"58",
         10084 => x"38",
         10085 => x"33",
         10086 => x"33",
         10087 => x"07",
         10088 => x"a4",
         10089 => x"17",
         10090 => x"82",
         10091 => x"90",
         10092 => x"2b",
         10093 => x"33",
         10094 => x"88",
         10095 => x"71",
         10096 => x"5a",
         10097 => x"42",
         10098 => x"33",
         10099 => x"33",
         10100 => x"07",
         10101 => x"58",
         10102 => x"81",
         10103 => x"1c",
         10104 => x"05",
         10105 => x"26",
         10106 => x"78",
         10107 => x"31",
         10108 => x"b4",
         10109 => x"8c",
         10110 => x"ba",
         10111 => x"2e",
         10112 => x"84",
         10113 => x"80",
         10114 => x"f5",
         10115 => x"83",
         10116 => x"ff",
         10117 => x"38",
         10118 => x"9f",
         10119 => x"eb",
         10120 => x"82",
         10121 => x"19",
         10122 => x"19",
         10123 => x"70",
         10124 => x"7b",
         10125 => x"0c",
         10126 => x"83",
         10127 => x"38",
         10128 => x"5c",
         10129 => x"80",
         10130 => x"38",
         10131 => x"18",
         10132 => x"55",
         10133 => x"8d",
         10134 => x"19",
         10135 => x"7a",
         10136 => x"56",
         10137 => x"15",
         10138 => x"8d",
         10139 => x"18",
         10140 => x"38",
         10141 => x"18",
         10142 => x"90",
         10143 => x"80",
         10144 => x"34",
         10145 => x"86",
         10146 => x"77",
         10147 => x"e4",
         10148 => x"5d",
         10149 => x"e4",
         10150 => x"18",
         10151 => x"ec",
         10152 => x"0c",
         10153 => x"18",
         10154 => x"77",
         10155 => x"0c",
         10156 => x"04",
         10157 => x"ba",
         10158 => x"3d",
         10159 => x"33",
         10160 => x"81",
         10161 => x"57",
         10162 => x"26",
         10163 => x"17",
         10164 => x"06",
         10165 => x"59",
         10166 => x"87",
         10167 => x"7e",
         10168 => x"fc",
         10169 => x"7c",
         10170 => x"5b",
         10171 => x"05",
         10172 => x"70",
         10173 => x"33",
         10174 => x"5a",
         10175 => x"99",
         10176 => x"e0",
         10177 => x"ff",
         10178 => x"ff",
         10179 => x"77",
         10180 => x"38",
         10181 => x"81",
         10182 => x"55",
         10183 => x"9f",
         10184 => x"75",
         10185 => x"81",
         10186 => x"77",
         10187 => x"78",
         10188 => x"30",
         10189 => x"9f",
         10190 => x"5d",
         10191 => x"80",
         10192 => x"38",
         10193 => x"1e",
         10194 => x"7c",
         10195 => x"38",
         10196 => x"a9",
         10197 => x"2e",
         10198 => x"77",
         10199 => x"06",
         10200 => x"7d",
         10201 => x"80",
         10202 => x"39",
         10203 => x"57",
         10204 => x"e9",
         10205 => x"06",
         10206 => x"59",
         10207 => x"32",
         10208 => x"80",
         10209 => x"5a",
         10210 => x"83",
         10211 => x"81",
         10212 => x"a6",
         10213 => x"77",
         10214 => x"59",
         10215 => x"33",
         10216 => x"7a",
         10217 => x"38",
         10218 => x"33",
         10219 => x"33",
         10220 => x"71",
         10221 => x"83",
         10222 => x"70",
         10223 => x"2b",
         10224 => x"33",
         10225 => x"59",
         10226 => x"40",
         10227 => x"84",
         10228 => x"ff",
         10229 => x"57",
         10230 => x"25",
         10231 => x"84",
         10232 => x"33",
         10233 => x"9f",
         10234 => x"31",
         10235 => x"10",
         10236 => x"05",
         10237 => x"44",
         10238 => x"5b",
         10239 => x"5b",
         10240 => x"80",
         10241 => x"38",
         10242 => x"18",
         10243 => x"b4",
         10244 => x"55",
         10245 => x"ff",
         10246 => x"81",
         10247 => x"b8",
         10248 => x"17",
         10249 => x"b4",
         10250 => x"ba",
         10251 => x"2e",
         10252 => x"55",
         10253 => x"b4",
         10254 => x"58",
         10255 => x"81",
         10256 => x"33",
         10257 => x"07",
         10258 => x"58",
         10259 => x"d5",
         10260 => x"06",
         10261 => x"0b",
         10262 => x"57",
         10263 => x"e9",
         10264 => x"38",
         10265 => x"32",
         10266 => x"80",
         10267 => x"42",
         10268 => x"bc",
         10269 => x"e8",
         10270 => x"82",
         10271 => x"ff",
         10272 => x"0b",
         10273 => x"1e",
         10274 => x"7b",
         10275 => x"81",
         10276 => x"81",
         10277 => x"27",
         10278 => x"77",
         10279 => x"b7",
         10280 => x"84",
         10281 => x"83",
         10282 => x"d1",
         10283 => x"39",
         10284 => x"ee",
         10285 => x"bc",
         10286 => x"7b",
         10287 => x"5d",
         10288 => x"81",
         10289 => x"71",
         10290 => x"1b",
         10291 => x"56",
         10292 => x"80",
         10293 => x"80",
         10294 => x"85",
         10295 => x"18",
         10296 => x"40",
         10297 => x"70",
         10298 => x"33",
         10299 => x"05",
         10300 => x"71",
         10301 => x"5b",
         10302 => x"77",
         10303 => x"8e",
         10304 => x"2e",
         10305 => x"58",
         10306 => x"8d",
         10307 => x"93",
         10308 => x"ba",
         10309 => x"3d",
         10310 => x"58",
         10311 => x"fe",
         10312 => x"0b",
         10313 => x"83",
         10314 => x"5d",
         10315 => x"39",
         10316 => x"ba",
         10317 => x"3d",
         10318 => x"0b",
         10319 => x"83",
         10320 => x"5a",
         10321 => x"81",
         10322 => x"7a",
         10323 => x"5c",
         10324 => x"31",
         10325 => x"57",
         10326 => x"80",
         10327 => x"38",
         10328 => x"e1",
         10329 => x"81",
         10330 => x"e5",
         10331 => x"58",
         10332 => x"05",
         10333 => x"70",
         10334 => x"33",
         10335 => x"ff",
         10336 => x"42",
         10337 => x"2e",
         10338 => x"75",
         10339 => x"38",
         10340 => x"57",
         10341 => x"fc",
         10342 => x"58",
         10343 => x"80",
         10344 => x"80",
         10345 => x"71",
         10346 => x"57",
         10347 => x"2e",
         10348 => x"f9",
         10349 => x"1b",
         10350 => x"b4",
         10351 => x"2e",
         10352 => x"17",
         10353 => x"7a",
         10354 => x"06",
         10355 => x"81",
         10356 => x"b8",
         10357 => x"17",
         10358 => x"b0",
         10359 => x"ba",
         10360 => x"2e",
         10361 => x"58",
         10362 => x"b4",
         10363 => x"f9",
         10364 => x"84",
         10365 => x"b7",
         10366 => x"b6",
         10367 => x"88",
         10368 => x"5e",
         10369 => x"d5",
         10370 => x"06",
         10371 => x"b8",
         10372 => x"33",
         10373 => x"71",
         10374 => x"88",
         10375 => x"14",
         10376 => x"07",
         10377 => x"33",
         10378 => x"41",
         10379 => x"5c",
         10380 => x"8b",
         10381 => x"2e",
         10382 => x"f8",
         10383 => x"9c",
         10384 => x"33",
         10385 => x"71",
         10386 => x"88",
         10387 => x"14",
         10388 => x"07",
         10389 => x"33",
         10390 => x"44",
         10391 => x"5a",
         10392 => x"8a",
         10393 => x"2e",
         10394 => x"f8",
         10395 => x"a0",
         10396 => x"33",
         10397 => x"71",
         10398 => x"88",
         10399 => x"14",
         10400 => x"07",
         10401 => x"33",
         10402 => x"1e",
         10403 => x"a4",
         10404 => x"33",
         10405 => x"71",
         10406 => x"88",
         10407 => x"14",
         10408 => x"07",
         10409 => x"33",
         10410 => x"90",
         10411 => x"44",
         10412 => x"45",
         10413 => x"56",
         10414 => x"34",
         10415 => x"22",
         10416 => x"7c",
         10417 => x"23",
         10418 => x"23",
         10419 => x"0b",
         10420 => x"80",
         10421 => x"0c",
         10422 => x"7b",
         10423 => x"f0",
         10424 => x"7f",
         10425 => x"95",
         10426 => x"b4",
         10427 => x"b8",
         10428 => x"81",
         10429 => x"59",
         10430 => x"3f",
         10431 => x"08",
         10432 => x"81",
         10433 => x"38",
         10434 => x"08",
         10435 => x"b4",
         10436 => x"18",
         10437 => x"7f",
         10438 => x"27",
         10439 => x"17",
         10440 => x"82",
         10441 => x"38",
         10442 => x"08",
         10443 => x"39",
         10444 => x"80",
         10445 => x"38",
         10446 => x"8a",
         10447 => x"c0",
         10448 => x"fc",
         10449 => x"e3",
         10450 => x"e2",
         10451 => x"88",
         10452 => x"5a",
         10453 => x"f6",
         10454 => x"17",
         10455 => x"f6",
         10456 => x"e4",
         10457 => x"33",
         10458 => x"71",
         10459 => x"88",
         10460 => x"14",
         10461 => x"07",
         10462 => x"33",
         10463 => x"1e",
         10464 => x"82",
         10465 => x"44",
         10466 => x"f5",
         10467 => x"58",
         10468 => x"f9",
         10469 => x"58",
         10470 => x"75",
         10471 => x"a8",
         10472 => x"77",
         10473 => x"59",
         10474 => x"75",
         10475 => x"da",
         10476 => x"39",
         10477 => x"17",
         10478 => x"08",
         10479 => x"52",
         10480 => x"51",
         10481 => x"3f",
         10482 => x"f0",
         10483 => x"80",
         10484 => x"64",
         10485 => x"3d",
         10486 => x"ff",
         10487 => x"75",
         10488 => x"e9",
         10489 => x"81",
         10490 => x"70",
         10491 => x"55",
         10492 => x"80",
         10493 => x"ed",
         10494 => x"2e",
         10495 => x"84",
         10496 => x"54",
         10497 => x"80",
         10498 => x"10",
         10499 => x"d4",
         10500 => x"55",
         10501 => x"2e",
         10502 => x"74",
         10503 => x"73",
         10504 => x"38",
         10505 => x"62",
         10506 => x"0c",
         10507 => x"80",
         10508 => x"80",
         10509 => x"70",
         10510 => x"51",
         10511 => x"84",
         10512 => x"54",
         10513 => x"8c",
         10514 => x"0d",
         10515 => x"84",
         10516 => x"92",
         10517 => x"75",
         10518 => x"70",
         10519 => x"56",
         10520 => x"89",
         10521 => x"82",
         10522 => x"ff",
         10523 => x"5c",
         10524 => x"2e",
         10525 => x"80",
         10526 => x"e5",
         10527 => x"5b",
         10528 => x"59",
         10529 => x"81",
         10530 => x"78",
         10531 => x"5a",
         10532 => x"12",
         10533 => x"76",
         10534 => x"38",
         10535 => x"81",
         10536 => x"54",
         10537 => x"57",
         10538 => x"89",
         10539 => x"70",
         10540 => x"57",
         10541 => x"70",
         10542 => x"54",
         10543 => x"09",
         10544 => x"38",
         10545 => x"38",
         10546 => x"70",
         10547 => x"07",
         10548 => x"07",
         10549 => x"79",
         10550 => x"38",
         10551 => x"1d",
         10552 => x"7b",
         10553 => x"38",
         10554 => x"98",
         10555 => x"24",
         10556 => x"79",
         10557 => x"fe",
         10558 => x"3d",
         10559 => x"84",
         10560 => x"05",
         10561 => x"89",
         10562 => x"2e",
         10563 => x"bf",
         10564 => x"9d",
         10565 => x"53",
         10566 => x"05",
         10567 => x"9f",
         10568 => x"8c",
         10569 => x"ba",
         10570 => x"2e",
         10571 => x"79",
         10572 => x"75",
         10573 => x"0c",
         10574 => x"04",
         10575 => x"52",
         10576 => x"52",
         10577 => x"3f",
         10578 => x"08",
         10579 => x"8c",
         10580 => x"81",
         10581 => x"9c",
         10582 => x"80",
         10583 => x"38",
         10584 => x"83",
         10585 => x"84",
         10586 => x"38",
         10587 => x"58",
         10588 => x"38",
         10589 => x"81",
         10590 => x"80",
         10591 => x"38",
         10592 => x"33",
         10593 => x"71",
         10594 => x"61",
         10595 => x"58",
         10596 => x"7d",
         10597 => x"e9",
         10598 => x"8e",
         10599 => x"0b",
         10600 => x"a1",
         10601 => x"34",
         10602 => x"91",
         10603 => x"56",
         10604 => x"17",
         10605 => x"57",
         10606 => x"9a",
         10607 => x"0b",
         10608 => x"7d",
         10609 => x"83",
         10610 => x"38",
         10611 => x"0b",
         10612 => x"80",
         10613 => x"34",
         10614 => x"1c",
         10615 => x"9f",
         10616 => x"55",
         10617 => x"16",
         10618 => x"2e",
         10619 => x"7e",
         10620 => x"7d",
         10621 => x"57",
         10622 => x"7c",
         10623 => x"9c",
         10624 => x"26",
         10625 => x"82",
         10626 => x"0c",
         10627 => x"02",
         10628 => x"33",
         10629 => x"5d",
         10630 => x"25",
         10631 => x"86",
         10632 => x"5e",
         10633 => x"b8",
         10634 => x"82",
         10635 => x"c2",
         10636 => x"84",
         10637 => x"5d",
         10638 => x"91",
         10639 => x"2a",
         10640 => x"7d",
         10641 => x"38",
         10642 => x"5a",
         10643 => x"38",
         10644 => x"81",
         10645 => x"80",
         10646 => x"77",
         10647 => x"58",
         10648 => x"08",
         10649 => x"67",
         10650 => x"67",
         10651 => x"9a",
         10652 => x"88",
         10653 => x"33",
         10654 => x"57",
         10655 => x"2e",
         10656 => x"7a",
         10657 => x"9c",
         10658 => x"33",
         10659 => x"71",
         10660 => x"88",
         10661 => x"14",
         10662 => x"07",
         10663 => x"33",
         10664 => x"60",
         10665 => x"60",
         10666 => x"52",
         10667 => x"5d",
         10668 => x"22",
         10669 => x"77",
         10670 => x"80",
         10671 => x"34",
         10672 => x"1a",
         10673 => x"2a",
         10674 => x"74",
         10675 => x"ac",
         10676 => x"2e",
         10677 => x"75",
         10678 => x"8a",
         10679 => x"89",
         10680 => x"5b",
         10681 => x"70",
         10682 => x"25",
         10683 => x"76",
         10684 => x"38",
         10685 => x"06",
         10686 => x"80",
         10687 => x"38",
         10688 => x"51",
         10689 => x"3f",
         10690 => x"08",
         10691 => x"8c",
         10692 => x"83",
         10693 => x"84",
         10694 => x"ff",
         10695 => x"38",
         10696 => x"56",
         10697 => x"80",
         10698 => x"91",
         10699 => x"95",
         10700 => x"2a",
         10701 => x"74",
         10702 => x"b8",
         10703 => x"80",
         10704 => x"ed",
         10705 => x"80",
         10706 => x"e5",
         10707 => x"80",
         10708 => x"dd",
         10709 => x"cd",
         10710 => x"ba",
         10711 => x"88",
         10712 => x"76",
         10713 => x"fc",
         10714 => x"76",
         10715 => x"57",
         10716 => x"95",
         10717 => x"17",
         10718 => x"2b",
         10719 => x"07",
         10720 => x"5e",
         10721 => x"39",
         10722 => x"7b",
         10723 => x"38",
         10724 => x"51",
         10725 => x"3f",
         10726 => x"08",
         10727 => x"8c",
         10728 => x"81",
         10729 => x"ba",
         10730 => x"2e",
         10731 => x"84",
         10732 => x"ff",
         10733 => x"38",
         10734 => x"52",
         10735 => x"b2",
         10736 => x"ba",
         10737 => x"90",
         10738 => x"08",
         10739 => x"19",
         10740 => x"5b",
         10741 => x"ff",
         10742 => x"16",
         10743 => x"84",
         10744 => x"07",
         10745 => x"18",
         10746 => x"7a",
         10747 => x"a0",
         10748 => x"39",
         10749 => x"17",
         10750 => x"95",
         10751 => x"cc",
         10752 => x"33",
         10753 => x"71",
         10754 => x"90",
         10755 => x"07",
         10756 => x"80",
         10757 => x"34",
         10758 => x"17",
         10759 => x"90",
         10760 => x"cc",
         10761 => x"34",
         10762 => x"0b",
         10763 => x"7e",
         10764 => x"80",
         10765 => x"34",
         10766 => x"17",
         10767 => x"5d",
         10768 => x"09",
         10769 => x"84",
         10770 => x"39",
         10771 => x"72",
         10772 => x"5d",
         10773 => x"7e",
         10774 => x"83",
         10775 => x"79",
         10776 => x"81",
         10777 => x"81",
         10778 => x"b8",
         10779 => x"16",
         10780 => x"a3",
         10781 => x"ba",
         10782 => x"2e",
         10783 => x"57",
         10784 => x"b4",
         10785 => x"56",
         10786 => x"90",
         10787 => x"7a",
         10788 => x"bc",
         10789 => x"0c",
         10790 => x"81",
         10791 => x"08",
         10792 => x"70",
         10793 => x"33",
         10794 => x"a4",
         10795 => x"ba",
         10796 => x"2e",
         10797 => x"81",
         10798 => x"ba",
         10799 => x"17",
         10800 => x"08",
         10801 => x"31",
         10802 => x"08",
         10803 => x"a0",
         10804 => x"ff",
         10805 => x"16",
         10806 => x"82",
         10807 => x"06",
         10808 => x"81",
         10809 => x"08",
         10810 => x"05",
         10811 => x"81",
         10812 => x"ff",
         10813 => x"7c",
         10814 => x"39",
         10815 => x"0c",
         10816 => x"af",
         10817 => x"1a",
         10818 => x"a2",
         10819 => x"ff",
         10820 => x"80",
         10821 => x"38",
         10822 => x"9c",
         10823 => x"05",
         10824 => x"77",
         10825 => x"df",
         10826 => x"22",
         10827 => x"b0",
         10828 => x"56",
         10829 => x"2e",
         10830 => x"75",
         10831 => x"9c",
         10832 => x"56",
         10833 => x"75",
         10834 => x"76",
         10835 => x"39",
         10836 => x"79",
         10837 => x"39",
         10838 => x"08",
         10839 => x"0c",
         10840 => x"81",
         10841 => x"fe",
         10842 => x"3d",
         10843 => x"67",
         10844 => x"5d",
         10845 => x"0c",
         10846 => x"80",
         10847 => x"79",
         10848 => x"80",
         10849 => x"75",
         10850 => x"80",
         10851 => x"86",
         10852 => x"1b",
         10853 => x"78",
         10854 => x"b7",
         10855 => x"74",
         10856 => x"76",
         10857 => x"91",
         10858 => x"74",
         10859 => x"90",
         10860 => x"06",
         10861 => x"76",
         10862 => x"ed",
         10863 => x"08",
         10864 => x"71",
         10865 => x"7b",
         10866 => x"ef",
         10867 => x"2e",
         10868 => x"60",
         10869 => x"ff",
         10870 => x"81",
         10871 => x"19",
         10872 => x"76",
         10873 => x"5b",
         10874 => x"75",
         10875 => x"88",
         10876 => x"81",
         10877 => x"85",
         10878 => x"2e",
         10879 => x"74",
         10880 => x"60",
         10881 => x"08",
         10882 => x"1a",
         10883 => x"41",
         10884 => x"27",
         10885 => x"8a",
         10886 => x"78",
         10887 => x"08",
         10888 => x"74",
         10889 => x"d5",
         10890 => x"7c",
         10891 => x"57",
         10892 => x"83",
         10893 => x"1b",
         10894 => x"27",
         10895 => x"7b",
         10896 => x"54",
         10897 => x"52",
         10898 => x"51",
         10899 => x"3f",
         10900 => x"08",
         10901 => x"60",
         10902 => x"57",
         10903 => x"2e",
         10904 => x"19",
         10905 => x"56",
         10906 => x"9e",
         10907 => x"76",
         10908 => x"b8",
         10909 => x"55",
         10910 => x"05",
         10911 => x"70",
         10912 => x"34",
         10913 => x"74",
         10914 => x"89",
         10915 => x"78",
         10916 => x"19",
         10917 => x"1e",
         10918 => x"1a",
         10919 => x"1d",
         10920 => x"7b",
         10921 => x"80",
         10922 => x"ba",
         10923 => x"3d",
         10924 => x"84",
         10925 => x"92",
         10926 => x"74",
         10927 => x"39",
         10928 => x"57",
         10929 => x"06",
         10930 => x"31",
         10931 => x"78",
         10932 => x"7b",
         10933 => x"b4",
         10934 => x"2e",
         10935 => x"0b",
         10936 => x"71",
         10937 => x"7f",
         10938 => x"81",
         10939 => x"38",
         10940 => x"53",
         10941 => x"81",
         10942 => x"ff",
         10943 => x"84",
         10944 => x"80",
         10945 => x"ff",
         10946 => x"75",
         10947 => x"7a",
         10948 => x"60",
         10949 => x"83",
         10950 => x"79",
         10951 => x"b8",
         10952 => x"77",
         10953 => x"e6",
         10954 => x"81",
         10955 => x"77",
         10956 => x"59",
         10957 => x"56",
         10958 => x"fe",
         10959 => x"70",
         10960 => x"33",
         10961 => x"05",
         10962 => x"16",
         10963 => x"38",
         10964 => x"81",
         10965 => x"08",
         10966 => x"70",
         10967 => x"33",
         10968 => x"9e",
         10969 => x"5b",
         10970 => x"08",
         10971 => x"81",
         10972 => x"38",
         10973 => x"08",
         10974 => x"b4",
         10975 => x"1a",
         10976 => x"ba",
         10977 => x"55",
         10978 => x"08",
         10979 => x"38",
         10980 => x"55",
         10981 => x"09",
         10982 => x"d4",
         10983 => x"b4",
         10984 => x"1a",
         10985 => x"7f",
         10986 => x"33",
         10987 => x"fe",
         10988 => x"fe",
         10989 => x"9c",
         10990 => x"1a",
         10991 => x"84",
         10992 => x"08",
         10993 => x"ff",
         10994 => x"84",
         10995 => x"55",
         10996 => x"81",
         10997 => x"ff",
         10998 => x"84",
         10999 => x"81",
         11000 => x"fb",
         11001 => x"7a",
         11002 => x"fb",
         11003 => x"0b",
         11004 => x"81",
         11005 => x"8c",
         11006 => x"0d",
         11007 => x"91",
         11008 => x"0b",
         11009 => x"0c",
         11010 => x"04",
         11011 => x"62",
         11012 => x"40",
         11013 => x"80",
         11014 => x"57",
         11015 => x"9f",
         11016 => x"56",
         11017 => x"97",
         11018 => x"55",
         11019 => x"8f",
         11020 => x"22",
         11021 => x"59",
         11022 => x"2e",
         11023 => x"80",
         11024 => x"76",
         11025 => x"c4",
         11026 => x"33",
         11027 => x"bc",
         11028 => x"33",
         11029 => x"81",
         11030 => x"87",
         11031 => x"2e",
         11032 => x"94",
         11033 => x"11",
         11034 => x"77",
         11035 => x"76",
         11036 => x"80",
         11037 => x"38",
         11038 => x"06",
         11039 => x"a2",
         11040 => x"11",
         11041 => x"78",
         11042 => x"5a",
         11043 => x"38",
         11044 => x"38",
         11045 => x"55",
         11046 => x"84",
         11047 => x"81",
         11048 => x"38",
         11049 => x"86",
         11050 => x"98",
         11051 => x"1a",
         11052 => x"74",
         11053 => x"60",
         11054 => x"08",
         11055 => x"2e",
         11056 => x"98",
         11057 => x"05",
         11058 => x"fe",
         11059 => x"77",
         11060 => x"f0",
         11061 => x"22",
         11062 => x"b0",
         11063 => x"56",
         11064 => x"2e",
         11065 => x"78",
         11066 => x"2a",
         11067 => x"80",
         11068 => x"38",
         11069 => x"76",
         11070 => x"38",
         11071 => x"58",
         11072 => x"53",
         11073 => x"16",
         11074 => x"9b",
         11075 => x"ba",
         11076 => x"a1",
         11077 => x"11",
         11078 => x"56",
         11079 => x"27",
         11080 => x"80",
         11081 => x"76",
         11082 => x"57",
         11083 => x"70",
         11084 => x"33",
         11085 => x"05",
         11086 => x"16",
         11087 => x"38",
         11088 => x"83",
         11089 => x"89",
         11090 => x"79",
         11091 => x"1a",
         11092 => x"1e",
         11093 => x"1b",
         11094 => x"1f",
         11095 => x"08",
         11096 => x"5e",
         11097 => x"27",
         11098 => x"56",
         11099 => x"0c",
         11100 => x"38",
         11101 => x"58",
         11102 => x"07",
         11103 => x"1b",
         11104 => x"75",
         11105 => x"0c",
         11106 => x"04",
         11107 => x"8c",
         11108 => x"0d",
         11109 => x"33",
         11110 => x"c8",
         11111 => x"fe",
         11112 => x"9c",
         11113 => x"56",
         11114 => x"06",
         11115 => x"31",
         11116 => x"79",
         11117 => x"7a",
         11118 => x"b4",
         11119 => x"2e",
         11120 => x"0b",
         11121 => x"71",
         11122 => x"7f",
         11123 => x"81",
         11124 => x"38",
         11125 => x"53",
         11126 => x"81",
         11127 => x"ff",
         11128 => x"84",
         11129 => x"80",
         11130 => x"ff",
         11131 => x"76",
         11132 => x"7b",
         11133 => x"60",
         11134 => x"83",
         11135 => x"7a",
         11136 => x"7e",
         11137 => x"78",
         11138 => x"38",
         11139 => x"05",
         11140 => x"70",
         11141 => x"34",
         11142 => x"75",
         11143 => x"58",
         11144 => x"19",
         11145 => x"39",
         11146 => x"16",
         11147 => x"16",
         11148 => x"17",
         11149 => x"ff",
         11150 => x"81",
         11151 => x"8c",
         11152 => x"09",
         11153 => x"ab",
         11154 => x"8c",
         11155 => x"34",
         11156 => x"a8",
         11157 => x"84",
         11158 => x"5d",
         11159 => x"17",
         11160 => x"f0",
         11161 => x"33",
         11162 => x"2e",
         11163 => x"fe",
         11164 => x"54",
         11165 => x"a0",
         11166 => x"53",
         11167 => x"16",
         11168 => x"98",
         11169 => x"5c",
         11170 => x"94",
         11171 => x"8c",
         11172 => x"26",
         11173 => x"16",
         11174 => x"81",
         11175 => x"7c",
         11176 => x"94",
         11177 => x"56",
         11178 => x"1c",
         11179 => x"f8",
         11180 => x"08",
         11181 => x"ff",
         11182 => x"84",
         11183 => x"55",
         11184 => x"08",
         11185 => x"90",
         11186 => x"fd",
         11187 => x"52",
         11188 => x"ab",
         11189 => x"ba",
         11190 => x"84",
         11191 => x"fb",
         11192 => x"39",
         11193 => x"16",
         11194 => x"16",
         11195 => x"17",
         11196 => x"ff",
         11197 => x"84",
         11198 => x"81",
         11199 => x"ba",
         11200 => x"17",
         11201 => x"08",
         11202 => x"31",
         11203 => x"17",
         11204 => x"89",
         11205 => x"33",
         11206 => x"2e",
         11207 => x"fc",
         11208 => x"54",
         11209 => x"a0",
         11210 => x"53",
         11211 => x"16",
         11212 => x"96",
         11213 => x"56",
         11214 => x"81",
         11215 => x"ff",
         11216 => x"84",
         11217 => x"81",
         11218 => x"f9",
         11219 => x"7a",
         11220 => x"f9",
         11221 => x"54",
         11222 => x"53",
         11223 => x"53",
         11224 => x"52",
         11225 => x"c6",
         11226 => x"8c",
         11227 => x"38",
         11228 => x"08",
         11229 => x"b4",
         11230 => x"17",
         11231 => x"74",
         11232 => x"27",
         11233 => x"82",
         11234 => x"77",
         11235 => x"81",
         11236 => x"38",
         11237 => x"16",
         11238 => x"08",
         11239 => x"52",
         11240 => x"51",
         11241 => x"3f",
         11242 => x"12",
         11243 => x"08",
         11244 => x"f4",
         11245 => x"91",
         11246 => x"0b",
         11247 => x"0c",
         11248 => x"04",
         11249 => x"1b",
         11250 => x"84",
         11251 => x"92",
         11252 => x"f5",
         11253 => x"58",
         11254 => x"80",
         11255 => x"77",
         11256 => x"80",
         11257 => x"75",
         11258 => x"80",
         11259 => x"86",
         11260 => x"19",
         11261 => x"78",
         11262 => x"b5",
         11263 => x"74",
         11264 => x"79",
         11265 => x"90",
         11266 => x"86",
         11267 => x"5c",
         11268 => x"2e",
         11269 => x"7b",
         11270 => x"5a",
         11271 => x"08",
         11272 => x"38",
         11273 => x"5b",
         11274 => x"38",
         11275 => x"53",
         11276 => x"81",
         11277 => x"ff",
         11278 => x"84",
         11279 => x"80",
         11280 => x"ff",
         11281 => x"78",
         11282 => x"75",
         11283 => x"a4",
         11284 => x"11",
         11285 => x"5a",
         11286 => x"18",
         11287 => x"88",
         11288 => x"83",
         11289 => x"5d",
         11290 => x"9a",
         11291 => x"88",
         11292 => x"9b",
         11293 => x"17",
         11294 => x"19",
         11295 => x"74",
         11296 => x"c1",
         11297 => x"08",
         11298 => x"34",
         11299 => x"5b",
         11300 => x"34",
         11301 => x"56",
         11302 => x"34",
         11303 => x"59",
         11304 => x"34",
         11305 => x"80",
         11306 => x"34",
         11307 => x"18",
         11308 => x"0b",
         11309 => x"80",
         11310 => x"34",
         11311 => x"18",
         11312 => x"81",
         11313 => x"34",
         11314 => x"96",
         11315 => x"ba",
         11316 => x"19",
         11317 => x"06",
         11318 => x"90",
         11319 => x"84",
         11320 => x"8d",
         11321 => x"81",
         11322 => x"08",
         11323 => x"70",
         11324 => x"33",
         11325 => x"93",
         11326 => x"56",
         11327 => x"08",
         11328 => x"84",
         11329 => x"83",
         11330 => x"17",
         11331 => x"08",
         11332 => x"8c",
         11333 => x"74",
         11334 => x"27",
         11335 => x"82",
         11336 => x"74",
         11337 => x"81",
         11338 => x"38",
         11339 => x"17",
         11340 => x"08",
         11341 => x"52",
         11342 => x"51",
         11343 => x"3f",
         11344 => x"e8",
         11345 => x"2a",
         11346 => x"18",
         11347 => x"2a",
         11348 => x"18",
         11349 => x"08",
         11350 => x"34",
         11351 => x"5b",
         11352 => x"34",
         11353 => x"56",
         11354 => x"34",
         11355 => x"59",
         11356 => x"34",
         11357 => x"80",
         11358 => x"34",
         11359 => x"18",
         11360 => x"0b",
         11361 => x"80",
         11362 => x"34",
         11363 => x"18",
         11364 => x"81",
         11365 => x"34",
         11366 => x"94",
         11367 => x"ba",
         11368 => x"19",
         11369 => x"06",
         11370 => x"90",
         11371 => x"ae",
         11372 => x"33",
         11373 => x"a5",
         11374 => x"8c",
         11375 => x"55",
         11376 => x"38",
         11377 => x"56",
         11378 => x"39",
         11379 => x"79",
         11380 => x"fb",
         11381 => x"ba",
         11382 => x"84",
         11383 => x"b1",
         11384 => x"74",
         11385 => x"38",
         11386 => x"72",
         11387 => x"38",
         11388 => x"71",
         11389 => x"38",
         11390 => x"84",
         11391 => x"52",
         11392 => x"96",
         11393 => x"71",
         11394 => x"75",
         11395 => x"75",
         11396 => x"ba",
         11397 => x"3d",
         11398 => x"13",
         11399 => x"8f",
         11400 => x"ba",
         11401 => x"06",
         11402 => x"38",
         11403 => x"53",
         11404 => x"f6",
         11405 => x"7d",
         11406 => x"5b",
         11407 => x"b2",
         11408 => x"81",
         11409 => x"70",
         11410 => x"52",
         11411 => x"ac",
         11412 => x"38",
         11413 => x"a4",
         11414 => x"e8",
         11415 => x"71",
         11416 => x"70",
         11417 => x"34",
         11418 => x"ba",
         11419 => x"3d",
         11420 => x"0b",
         11421 => x"0c",
         11422 => x"04",
         11423 => x"11",
         11424 => x"06",
         11425 => x"70",
         11426 => x"38",
         11427 => x"81",
         11428 => x"05",
         11429 => x"76",
         11430 => x"38",
         11431 => x"e5",
         11432 => x"79",
         11433 => x"57",
         11434 => x"05",
         11435 => x"70",
         11436 => x"33",
         11437 => x"53",
         11438 => x"99",
         11439 => x"e0",
         11440 => x"ff",
         11441 => x"ff",
         11442 => x"70",
         11443 => x"38",
         11444 => x"81",
         11445 => x"54",
         11446 => x"9f",
         11447 => x"71",
         11448 => x"81",
         11449 => x"73",
         11450 => x"74",
         11451 => x"30",
         11452 => x"9f",
         11453 => x"59",
         11454 => x"80",
         11455 => x"81",
         11456 => x"5b",
         11457 => x"25",
         11458 => x"7a",
         11459 => x"39",
         11460 => x"f7",
         11461 => x"5e",
         11462 => x"39",
         11463 => x"80",
         11464 => x"cc",
         11465 => x"3d",
         11466 => x"3f",
         11467 => x"08",
         11468 => x"8c",
         11469 => x"8a",
         11470 => x"ba",
         11471 => x"3d",
         11472 => x"5c",
         11473 => x"3d",
         11474 => x"c5",
         11475 => x"ba",
         11476 => x"84",
         11477 => x"80",
         11478 => x"80",
         11479 => x"70",
         11480 => x"5a",
         11481 => x"80",
         11482 => x"b2",
         11483 => x"84",
         11484 => x"57",
         11485 => x"2e",
         11486 => x"63",
         11487 => x"9a",
         11488 => x"88",
         11489 => x"33",
         11490 => x"57",
         11491 => x"2e",
         11492 => x"98",
         11493 => x"84",
         11494 => x"98",
         11495 => x"84",
         11496 => x"84",
         11497 => x"06",
         11498 => x"85",
         11499 => x"8c",
         11500 => x"0d",
         11501 => x"33",
         11502 => x"71",
         11503 => x"90",
         11504 => x"07",
         11505 => x"5b",
         11506 => x"7a",
         11507 => x"0c",
         11508 => x"ba",
         11509 => x"3d",
         11510 => x"9e",
         11511 => x"e6",
         11512 => x"e6",
         11513 => x"40",
         11514 => x"80",
         11515 => x"3d",
         11516 => x"52",
         11517 => x"51",
         11518 => x"84",
         11519 => x"59",
         11520 => x"08",
         11521 => x"60",
         11522 => x"0c",
         11523 => x"11",
         11524 => x"3d",
         11525 => x"db",
         11526 => x"58",
         11527 => x"82",
         11528 => x"d8",
         11529 => x"40",
         11530 => x"7a",
         11531 => x"aa",
         11532 => x"8c",
         11533 => x"ba",
         11534 => x"92",
         11535 => x"df",
         11536 => x"56",
         11537 => x"77",
         11538 => x"84",
         11539 => x"83",
         11540 => x"5d",
         11541 => x"38",
         11542 => x"53",
         11543 => x"81",
         11544 => x"ff",
         11545 => x"84",
         11546 => x"80",
         11547 => x"ff",
         11548 => x"76",
         11549 => x"78",
         11550 => x"80",
         11551 => x"9b",
         11552 => x"12",
         11553 => x"2b",
         11554 => x"33",
         11555 => x"56",
         11556 => x"2e",
         11557 => x"76",
         11558 => x"0c",
         11559 => x"51",
         11560 => x"3f",
         11561 => x"08",
         11562 => x"8c",
         11563 => x"38",
         11564 => x"51",
         11565 => x"3f",
         11566 => x"08",
         11567 => x"8c",
         11568 => x"80",
         11569 => x"9b",
         11570 => x"12",
         11571 => x"2b",
         11572 => x"33",
         11573 => x"5e",
         11574 => x"2e",
         11575 => x"76",
         11576 => x"38",
         11577 => x"08",
         11578 => x"ff",
         11579 => x"84",
         11580 => x"59",
         11581 => x"08",
         11582 => x"b4",
         11583 => x"2e",
         11584 => x"78",
         11585 => x"80",
         11586 => x"b8",
         11587 => x"51",
         11588 => x"3f",
         11589 => x"05",
         11590 => x"79",
         11591 => x"38",
         11592 => x"81",
         11593 => x"70",
         11594 => x"57",
         11595 => x"81",
         11596 => x"78",
         11597 => x"38",
         11598 => x"9c",
         11599 => x"82",
         11600 => x"18",
         11601 => x"08",
         11602 => x"ff",
         11603 => x"56",
         11604 => x"75",
         11605 => x"38",
         11606 => x"e6",
         11607 => x"5f",
         11608 => x"34",
         11609 => x"08",
         11610 => x"bd",
         11611 => x"2e",
         11612 => x"80",
         11613 => x"e8",
         11614 => x"10",
         11615 => x"05",
         11616 => x"33",
         11617 => x"5e",
         11618 => x"2e",
         11619 => x"1a",
         11620 => x"33",
         11621 => x"74",
         11622 => x"1a",
         11623 => x"26",
         11624 => x"57",
         11625 => x"94",
         11626 => x"5f",
         11627 => x"70",
         11628 => x"34",
         11629 => x"79",
         11630 => x"38",
         11631 => x"81",
         11632 => x"76",
         11633 => x"81",
         11634 => x"38",
         11635 => x"7c",
         11636 => x"ba",
         11637 => x"e4",
         11638 => x"95",
         11639 => x"17",
         11640 => x"2b",
         11641 => x"07",
         11642 => x"56",
         11643 => x"39",
         11644 => x"94",
         11645 => x"98",
         11646 => x"2b",
         11647 => x"80",
         11648 => x"5a",
         11649 => x"7a",
         11650 => x"ce",
         11651 => x"8c",
         11652 => x"ba",
         11653 => x"2e",
         11654 => x"ff",
         11655 => x"54",
         11656 => x"53",
         11657 => x"53",
         11658 => x"52",
         11659 => x"fe",
         11660 => x"84",
         11661 => x"fc",
         11662 => x"ba",
         11663 => x"17",
         11664 => x"08",
         11665 => x"31",
         11666 => x"08",
         11667 => x"a0",
         11668 => x"fc",
         11669 => x"16",
         11670 => x"82",
         11671 => x"06",
         11672 => x"81",
         11673 => x"08",
         11674 => x"05",
         11675 => x"81",
         11676 => x"ff",
         11677 => x"7c",
         11678 => x"39",
         11679 => x"e6",
         11680 => x"5c",
         11681 => x"34",
         11682 => x"d1",
         11683 => x"10",
         11684 => x"fc",
         11685 => x"70",
         11686 => x"59",
         11687 => x"7a",
         11688 => x"06",
         11689 => x"fd",
         11690 => x"e5",
         11691 => x"81",
         11692 => x"79",
         11693 => x"81",
         11694 => x"77",
         11695 => x"8e",
         11696 => x"3d",
         11697 => x"19",
         11698 => x"33",
         11699 => x"05",
         11700 => x"78",
         11701 => x"fd",
         11702 => x"59",
         11703 => x"78",
         11704 => x"0c",
         11705 => x"0d",
         11706 => x"0d",
         11707 => x"55",
         11708 => x"80",
         11709 => x"74",
         11710 => x"80",
         11711 => x"73",
         11712 => x"80",
         11713 => x"86",
         11714 => x"16",
         11715 => x"78",
         11716 => x"a0",
         11717 => x"72",
         11718 => x"75",
         11719 => x"91",
         11720 => x"72",
         11721 => x"8c",
         11722 => x"76",
         11723 => x"b9",
         11724 => x"08",
         11725 => x"76",
         11726 => x"cc",
         11727 => x"11",
         11728 => x"2b",
         11729 => x"73",
         11730 => x"f7",
         11731 => x"ff",
         11732 => x"ba",
         11733 => x"ba",
         11734 => x"15",
         11735 => x"53",
         11736 => x"ba",
         11737 => x"ba",
         11738 => x"26",
         11739 => x"75",
         11740 => x"70",
         11741 => x"77",
         11742 => x"17",
         11743 => x"59",
         11744 => x"82",
         11745 => x"77",
         11746 => x"38",
         11747 => x"94",
         11748 => x"94",
         11749 => x"16",
         11750 => x"2a",
         11751 => x"5a",
         11752 => x"2e",
         11753 => x"73",
         11754 => x"ff",
         11755 => x"84",
         11756 => x"54",
         11757 => x"08",
         11758 => x"a3",
         11759 => x"2e",
         11760 => x"74",
         11761 => x"38",
         11762 => x"9c",
         11763 => x"82",
         11764 => x"98",
         11765 => x"ae",
         11766 => x"91",
         11767 => x"53",
         11768 => x"8c",
         11769 => x"0d",
         11770 => x"33",
         11771 => x"81",
         11772 => x"73",
         11773 => x"75",
         11774 => x"55",
         11775 => x"76",
         11776 => x"81",
         11777 => x"38",
         11778 => x"0c",
         11779 => x"54",
         11780 => x"90",
         11781 => x"16",
         11782 => x"33",
         11783 => x"57",
         11784 => x"34",
         11785 => x"06",
         11786 => x"2e",
         11787 => x"15",
         11788 => x"85",
         11789 => x"16",
         11790 => x"84",
         11791 => x"8b",
         11792 => x"80",
         11793 => x"0c",
         11794 => x"54",
         11795 => x"80",
         11796 => x"98",
         11797 => x"80",
         11798 => x"38",
         11799 => x"84",
         11800 => x"57",
         11801 => x"17",
         11802 => x"76",
         11803 => x"56",
         11804 => x"a9",
         11805 => x"15",
         11806 => x"fe",
         11807 => x"56",
         11808 => x"80",
         11809 => x"16",
         11810 => x"29",
         11811 => x"05",
         11812 => x"11",
         11813 => x"78",
         11814 => x"df",
         11815 => x"08",
         11816 => x"39",
         11817 => x"51",
         11818 => x"3f",
         11819 => x"08",
         11820 => x"39",
         11821 => x"51",
         11822 => x"3f",
         11823 => x"08",
         11824 => x"72",
         11825 => x"72",
         11826 => x"56",
         11827 => x"73",
         11828 => x"ff",
         11829 => x"84",
         11830 => x"54",
         11831 => x"08",
         11832 => x"38",
         11833 => x"08",
         11834 => x"ed",
         11835 => x"8c",
         11836 => x"0c",
         11837 => x"0c",
         11838 => x"82",
         11839 => x"34",
         11840 => x"ba",
         11841 => x"3d",
         11842 => x"3d",
         11843 => x"89",
         11844 => x"2e",
         11845 => x"53",
         11846 => x"05",
         11847 => x"84",
         11848 => x"9b",
         11849 => x"8c",
         11850 => x"ba",
         11851 => x"2e",
         11852 => x"76",
         11853 => x"73",
         11854 => x"0c",
         11855 => x"04",
         11856 => x"7d",
         11857 => x"ff",
         11858 => x"84",
         11859 => x"55",
         11860 => x"08",
         11861 => x"ab",
         11862 => x"98",
         11863 => x"80",
         11864 => x"38",
         11865 => x"70",
         11866 => x"06",
         11867 => x"80",
         11868 => x"38",
         11869 => x"9b",
         11870 => x"12",
         11871 => x"2b",
         11872 => x"33",
         11873 => x"55",
         11874 => x"2e",
         11875 => x"88",
         11876 => x"58",
         11877 => x"84",
         11878 => x"52",
         11879 => x"99",
         11880 => x"ba",
         11881 => x"74",
         11882 => x"38",
         11883 => x"ff",
         11884 => x"76",
         11885 => x"39",
         11886 => x"76",
         11887 => x"39",
         11888 => x"94",
         11889 => x"98",
         11890 => x"2b",
         11891 => x"88",
         11892 => x"5a",
         11893 => x"fa",
         11894 => x"55",
         11895 => x"80",
         11896 => x"74",
         11897 => x"80",
         11898 => x"72",
         11899 => x"80",
         11900 => x"86",
         11901 => x"16",
         11902 => x"71",
         11903 => x"38",
         11904 => x"57",
         11905 => x"73",
         11906 => x"84",
         11907 => x"88",
         11908 => x"81",
         11909 => x"fe",
         11910 => x"84",
         11911 => x"81",
         11912 => x"dc",
         11913 => x"08",
         11914 => x"39",
         11915 => x"7a",
         11916 => x"89",
         11917 => x"2e",
         11918 => x"08",
         11919 => x"2e",
         11920 => x"33",
         11921 => x"2e",
         11922 => x"14",
         11923 => x"22",
         11924 => x"78",
         11925 => x"38",
         11926 => x"59",
         11927 => x"80",
         11928 => x"80",
         11929 => x"38",
         11930 => x"51",
         11931 => x"3f",
         11932 => x"08",
         11933 => x"8c",
         11934 => x"b5",
         11935 => x"8c",
         11936 => x"76",
         11937 => x"ff",
         11938 => x"72",
         11939 => x"ff",
         11940 => x"84",
         11941 => x"84",
         11942 => x"70",
         11943 => x"2c",
         11944 => x"08",
         11945 => x"54",
         11946 => x"8c",
         11947 => x"0d",
         11948 => x"53",
         11949 => x"ff",
         11950 => x"72",
         11951 => x"ff",
         11952 => x"84",
         11953 => x"84",
         11954 => x"70",
         11955 => x"2c",
         11956 => x"08",
         11957 => x"54",
         11958 => x"52",
         11959 => x"96",
         11960 => x"ba",
         11961 => x"ba",
         11962 => x"3d",
         11963 => x"14",
         11964 => x"fd",
         11965 => x"ba",
         11966 => x"06",
         11967 => x"d8",
         11968 => x"08",
         11969 => x"d2",
         11970 => x"0d",
         11971 => x"53",
         11972 => x"53",
         11973 => x"56",
         11974 => x"84",
         11975 => x"55",
         11976 => x"08",
         11977 => x"38",
         11978 => x"8c",
         11979 => x"0d",
         11980 => x"75",
         11981 => x"a9",
         11982 => x"8c",
         11983 => x"ba",
         11984 => x"38",
         11985 => x"05",
         11986 => x"2b",
         11987 => x"74",
         11988 => x"76",
         11989 => x"38",
         11990 => x"51",
         11991 => x"3f",
         11992 => x"8c",
         11993 => x"0d",
         11994 => x"84",
         11995 => x"95",
         11996 => x"ed",
         11997 => x"68",
         11998 => x"53",
         11999 => x"05",
         12000 => x"51",
         12001 => x"84",
         12002 => x"5a",
         12003 => x"08",
         12004 => x"75",
         12005 => x"9c",
         12006 => x"11",
         12007 => x"59",
         12008 => x"75",
         12009 => x"38",
         12010 => x"79",
         12011 => x"0c",
         12012 => x"04",
         12013 => x"08",
         12014 => x"5b",
         12015 => x"82",
         12016 => x"a8",
         12017 => x"ba",
         12018 => x"5d",
         12019 => x"c1",
         12020 => x"1d",
         12021 => x"56",
         12022 => x"76",
         12023 => x"38",
         12024 => x"78",
         12025 => x"81",
         12026 => x"54",
         12027 => x"17",
         12028 => x"33",
         12029 => x"b7",
         12030 => x"8c",
         12031 => x"85",
         12032 => x"81",
         12033 => x"18",
         12034 => x"5b",
         12035 => x"cc",
         12036 => x"5e",
         12037 => x"82",
         12038 => x"17",
         12039 => x"11",
         12040 => x"33",
         12041 => x"71",
         12042 => x"81",
         12043 => x"72",
         12044 => x"75",
         12045 => x"ff",
         12046 => x"06",
         12047 => x"70",
         12048 => x"05",
         12049 => x"83",
         12050 => x"ff",
         12051 => x"43",
         12052 => x"53",
         12053 => x"56",
         12054 => x"38",
         12055 => x"7a",
         12056 => x"84",
         12057 => x"07",
         12058 => x"18",
         12059 => x"ba",
         12060 => x"3d",
         12061 => x"54",
         12062 => x"53",
         12063 => x"53",
         12064 => x"52",
         12065 => x"a6",
         12066 => x"84",
         12067 => x"fe",
         12068 => x"ba",
         12069 => x"18",
         12070 => x"08",
         12071 => x"31",
         12072 => x"08",
         12073 => x"a0",
         12074 => x"fe",
         12075 => x"17",
         12076 => x"82",
         12077 => x"06",
         12078 => x"81",
         12079 => x"08",
         12080 => x"05",
         12081 => x"81",
         12082 => x"fe",
         12083 => x"77",
         12084 => x"39",
         12085 => x"92",
         12086 => x"75",
         12087 => x"ff",
         12088 => x"84",
         12089 => x"ff",
         12090 => x"38",
         12091 => x"08",
         12092 => x"f7",
         12093 => x"8c",
         12094 => x"84",
         12095 => x"07",
         12096 => x"05",
         12097 => x"5a",
         12098 => x"9c",
         12099 => x"26",
         12100 => x"7f",
         12101 => x"18",
         12102 => x"33",
         12103 => x"77",
         12104 => x"fe",
         12105 => x"17",
         12106 => x"11",
         12107 => x"71",
         12108 => x"70",
         12109 => x"25",
         12110 => x"83",
         12111 => x"1f",
         12112 => x"59",
         12113 => x"78",
         12114 => x"fe",
         12115 => x"5a",
         12116 => x"81",
         12117 => x"7a",
         12118 => x"94",
         12119 => x"17",
         12120 => x"58",
         12121 => x"34",
         12122 => x"82",
         12123 => x"e7",
         12124 => x"0d",
         12125 => x"56",
         12126 => x"9f",
         12127 => x"55",
         12128 => x"97",
         12129 => x"54",
         12130 => x"8f",
         12131 => x"22",
         12132 => x"59",
         12133 => x"2e",
         12134 => x"80",
         12135 => x"75",
         12136 => x"91",
         12137 => x"75",
         12138 => x"90",
         12139 => x"81",
         12140 => x"55",
         12141 => x"73",
         12142 => x"c4",
         12143 => x"08",
         12144 => x"18",
         12145 => x"38",
         12146 => x"38",
         12147 => x"77",
         12148 => x"81",
         12149 => x"38",
         12150 => x"74",
         12151 => x"82",
         12152 => x"88",
         12153 => x"17",
         12154 => x"0c",
         12155 => x"07",
         12156 => x"18",
         12157 => x"2e",
         12158 => x"91",
         12159 => x"55",
         12160 => x"8c",
         12161 => x"0d",
         12162 => x"78",
         12163 => x"ff",
         12164 => x"76",
         12165 => x"ca",
         12166 => x"8c",
         12167 => x"ba",
         12168 => x"2e",
         12169 => x"84",
         12170 => x"81",
         12171 => x"38",
         12172 => x"08",
         12173 => x"e5",
         12174 => x"73",
         12175 => x"ff",
         12176 => x"84",
         12177 => x"82",
         12178 => x"16",
         12179 => x"94",
         12180 => x"55",
         12181 => x"27",
         12182 => x"81",
         12183 => x"0c",
         12184 => x"81",
         12185 => x"84",
         12186 => x"54",
         12187 => x"ff",
         12188 => x"39",
         12189 => x"51",
         12190 => x"3f",
         12191 => x"08",
         12192 => x"73",
         12193 => x"73",
         12194 => x"56",
         12195 => x"80",
         12196 => x"33",
         12197 => x"56",
         12198 => x"18",
         12199 => x"39",
         12200 => x"52",
         12201 => x"fd",
         12202 => x"ba",
         12203 => x"2e",
         12204 => x"84",
         12205 => x"81",
         12206 => x"38",
         12207 => x"38",
         12208 => x"ba",
         12209 => x"19",
         12210 => x"a1",
         12211 => x"8c",
         12212 => x"08",
         12213 => x"56",
         12214 => x"84",
         12215 => x"27",
         12216 => x"84",
         12217 => x"9c",
         12218 => x"81",
         12219 => x"80",
         12220 => x"ff",
         12221 => x"75",
         12222 => x"c7",
         12223 => x"8c",
         12224 => x"ba",
         12225 => x"e3",
         12226 => x"76",
         12227 => x"d2",
         12228 => x"8c",
         12229 => x"ba",
         12230 => x"2e",
         12231 => x"84",
         12232 => x"81",
         12233 => x"38",
         12234 => x"08",
         12235 => x"fe",
         12236 => x"73",
         12237 => x"ff",
         12238 => x"84",
         12239 => x"80",
         12240 => x"16",
         12241 => x"94",
         12242 => x"55",
         12243 => x"27",
         12244 => x"15",
         12245 => x"84",
         12246 => x"07",
         12247 => x"17",
         12248 => x"77",
         12249 => x"a1",
         12250 => x"74",
         12251 => x"33",
         12252 => x"39",
         12253 => x"bb",
         12254 => x"90",
         12255 => x"56",
         12256 => x"82",
         12257 => x"82",
         12258 => x"33",
         12259 => x"86",
         12260 => x"8c",
         12261 => x"33",
         12262 => x"fa",
         12263 => x"90",
         12264 => x"54",
         12265 => x"84",
         12266 => x"56",
         12267 => x"56",
         12268 => x"db",
         12269 => x"53",
         12270 => x"9c",
         12271 => x"3d",
         12272 => x"fb",
         12273 => x"8c",
         12274 => x"ba",
         12275 => x"2e",
         12276 => x"84",
         12277 => x"a7",
         12278 => x"7d",
         12279 => x"08",
         12280 => x"70",
         12281 => x"ab",
         12282 => x"ba",
         12283 => x"84",
         12284 => x"de",
         12285 => x"93",
         12286 => x"85",
         12287 => x"59",
         12288 => x"77",
         12289 => x"98",
         12290 => x"7b",
         12291 => x"02",
         12292 => x"33",
         12293 => x"5d",
         12294 => x"7b",
         12295 => x"7d",
         12296 => x"9b",
         12297 => x"12",
         12298 => x"2b",
         12299 => x"41",
         12300 => x"58",
         12301 => x"80",
         12302 => x"84",
         12303 => x"57",
         12304 => x"80",
         12305 => x"56",
         12306 => x"7b",
         12307 => x"38",
         12308 => x"41",
         12309 => x"08",
         12310 => x"70",
         12311 => x"8b",
         12312 => x"ba",
         12313 => x"84",
         12314 => x"fe",
         12315 => x"ba",
         12316 => x"74",
         12317 => x"b4",
         12318 => x"8c",
         12319 => x"ba",
         12320 => x"38",
         12321 => x"ba",
         12322 => x"3d",
         12323 => x"16",
         12324 => x"33",
         12325 => x"71",
         12326 => x"7d",
         12327 => x"5d",
         12328 => x"84",
         12329 => x"84",
         12330 => x"84",
         12331 => x"fe",
         12332 => x"08",
         12333 => x"08",
         12334 => x"74",
         12335 => x"d3",
         12336 => x"78",
         12337 => x"92",
         12338 => x"8c",
         12339 => x"ba",
         12340 => x"2e",
         12341 => x"30",
         12342 => x"80",
         12343 => x"7a",
         12344 => x"38",
         12345 => x"95",
         12346 => x"08",
         12347 => x"7b",
         12348 => x"9c",
         12349 => x"26",
         12350 => x"82",
         12351 => x"d2",
         12352 => x"fe",
         12353 => x"84",
         12354 => x"84",
         12355 => x"a7",
         12356 => x"b8",
         12357 => x"19",
         12358 => x"5a",
         12359 => x"76",
         12360 => x"38",
         12361 => x"7a",
         12362 => x"7a",
         12363 => x"06",
         12364 => x"81",
         12365 => x"b8",
         12366 => x"17",
         12367 => x"f1",
         12368 => x"ba",
         12369 => x"2e",
         12370 => x"56",
         12371 => x"b4",
         12372 => x"56",
         12373 => x"9c",
         12374 => x"e5",
         12375 => x"0b",
         12376 => x"90",
         12377 => x"27",
         12378 => x"80",
         12379 => x"ff",
         12380 => x"84",
         12381 => x"56",
         12382 => x"08",
         12383 => x"96",
         12384 => x"2e",
         12385 => x"fe",
         12386 => x"56",
         12387 => x"81",
         12388 => x"08",
         12389 => x"81",
         12390 => x"fe",
         12391 => x"81",
         12392 => x"8c",
         12393 => x"09",
         12394 => x"a6",
         12395 => x"8c",
         12396 => x"34",
         12397 => x"a8",
         12398 => x"84",
         12399 => x"59",
         12400 => x"18",
         12401 => x"eb",
         12402 => x"33",
         12403 => x"2e",
         12404 => x"fe",
         12405 => x"54",
         12406 => x"a0",
         12407 => x"53",
         12408 => x"17",
         12409 => x"f1",
         12410 => x"58",
         12411 => x"79",
         12412 => x"27",
         12413 => x"74",
         12414 => x"fe",
         12415 => x"84",
         12416 => x"5a",
         12417 => x"08",
         12418 => x"cb",
         12419 => x"8c",
         12420 => x"fd",
         12421 => x"ba",
         12422 => x"2e",
         12423 => x"80",
         12424 => x"76",
         12425 => x"9b",
         12426 => x"8c",
         12427 => x"9c",
         12428 => x"11",
         12429 => x"58",
         12430 => x"7b",
         12431 => x"38",
         12432 => x"18",
         12433 => x"33",
         12434 => x"7b",
         12435 => x"79",
         12436 => x"26",
         12437 => x"80",
         12438 => x"39",
         12439 => x"f7",
         12440 => x"8c",
         12441 => x"95",
         12442 => x"fd",
         12443 => x"3d",
         12444 => x"9f",
         12445 => x"05",
         12446 => x"51",
         12447 => x"3f",
         12448 => x"08",
         12449 => x"8c",
         12450 => x"8a",
         12451 => x"ba",
         12452 => x"3d",
         12453 => x"43",
         12454 => x"3d",
         12455 => x"ff",
         12456 => x"84",
         12457 => x"56",
         12458 => x"08",
         12459 => x"0b",
         12460 => x"0c",
         12461 => x"04",
         12462 => x"08",
         12463 => x"81",
         12464 => x"02",
         12465 => x"33",
         12466 => x"81",
         12467 => x"86",
         12468 => x"b9",
         12469 => x"74",
         12470 => x"70",
         12471 => x"83",
         12472 => x"ba",
         12473 => x"57",
         12474 => x"8c",
         12475 => x"87",
         12476 => x"8c",
         12477 => x"80",
         12478 => x"ba",
         12479 => x"2e",
         12480 => x"75",
         12481 => x"7d",
         12482 => x"08",
         12483 => x"5d",
         12484 => x"80",
         12485 => x"19",
         12486 => x"fe",
         12487 => x"80",
         12488 => x"27",
         12489 => x"17",
         12490 => x"29",
         12491 => x"05",
         12492 => x"b4",
         12493 => x"17",
         12494 => x"79",
         12495 => x"76",
         12496 => x"58",
         12497 => x"55",
         12498 => x"74",
         12499 => x"22",
         12500 => x"27",
         12501 => x"81",
         12502 => x"53",
         12503 => x"17",
         12504 => x"ee",
         12505 => x"ba",
         12506 => x"df",
         12507 => x"58",
         12508 => x"56",
         12509 => x"81",
         12510 => x"08",
         12511 => x"70",
         12512 => x"33",
         12513 => x"ee",
         12514 => x"56",
         12515 => x"08",
         12516 => x"ba",
         12517 => x"18",
         12518 => x"08",
         12519 => x"31",
         12520 => x"18",
         12521 => x"ee",
         12522 => x"33",
         12523 => x"2e",
         12524 => x"fe",
         12525 => x"54",
         12526 => x"a0",
         12527 => x"53",
         12528 => x"17",
         12529 => x"ed",
         12530 => x"ca",
         12531 => x"7b",
         12532 => x"55",
         12533 => x"fd",
         12534 => x"9c",
         12535 => x"fd",
         12536 => x"52",
         12537 => x"f2",
         12538 => x"ba",
         12539 => x"84",
         12540 => x"80",
         12541 => x"38",
         12542 => x"08",
         12543 => x"8d",
         12544 => x"8c",
         12545 => x"fd",
         12546 => x"53",
         12547 => x"51",
         12548 => x"3f",
         12549 => x"08",
         12550 => x"9c",
         12551 => x"11",
         12552 => x"5a",
         12553 => x"7b",
         12554 => x"81",
         12555 => x"0c",
         12556 => x"81",
         12557 => x"84",
         12558 => x"55",
         12559 => x"ff",
         12560 => x"84",
         12561 => x"9f",
         12562 => x"8a",
         12563 => x"74",
         12564 => x"06",
         12565 => x"76",
         12566 => x"81",
         12567 => x"38",
         12568 => x"1f",
         12569 => x"75",
         12570 => x"57",
         12571 => x"56",
         12572 => x"7d",
         12573 => x"b8",
         12574 => x"58",
         12575 => x"c3",
         12576 => x"59",
         12577 => x"1a",
         12578 => x"cf",
         12579 => x"0b",
         12580 => x"34",
         12581 => x"80",
         12582 => x"7d",
         12583 => x"ff",
         12584 => x"77",
         12585 => x"34",
         12586 => x"5b",
         12587 => x"17",
         12588 => x"55",
         12589 => x"81",
         12590 => x"59",
         12591 => x"d8",
         12592 => x"57",
         12593 => x"70",
         12594 => x"33",
         12595 => x"05",
         12596 => x"16",
         12597 => x"38",
         12598 => x"0b",
         12599 => x"34",
         12600 => x"83",
         12601 => x"5b",
         12602 => x"80",
         12603 => x"78",
         12604 => x"7a",
         12605 => x"34",
         12606 => x"74",
         12607 => x"f0",
         12608 => x"81",
         12609 => x"34",
         12610 => x"92",
         12611 => x"ba",
         12612 => x"84",
         12613 => x"fd",
         12614 => x"56",
         12615 => x"08",
         12616 => x"84",
         12617 => x"97",
         12618 => x"0b",
         12619 => x"80",
         12620 => x"17",
         12621 => x"58",
         12622 => x"18",
         12623 => x"2a",
         12624 => x"18",
         12625 => x"5a",
         12626 => x"80",
         12627 => x"55",
         12628 => x"16",
         12629 => x"81",
         12630 => x"34",
         12631 => x"ed",
         12632 => x"ba",
         12633 => x"75",
         12634 => x"0c",
         12635 => x"04",
         12636 => x"55",
         12637 => x"17",
         12638 => x"2a",
         12639 => x"ed",
         12640 => x"fd",
         12641 => x"2a",
         12642 => x"cc",
         12643 => x"88",
         12644 => x"80",
         12645 => x"7d",
         12646 => x"80",
         12647 => x"1b",
         12648 => x"fe",
         12649 => x"90",
         12650 => x"94",
         12651 => x"88",
         12652 => x"95",
         12653 => x"55",
         12654 => x"16",
         12655 => x"81",
         12656 => x"34",
         12657 => x"ec",
         12658 => x"ba",
         12659 => x"ff",
         12660 => x"3d",
         12661 => x"b4",
         12662 => x"59",
         12663 => x"80",
         12664 => x"79",
         12665 => x"5b",
         12666 => x"26",
         12667 => x"ba",
         12668 => x"38",
         12669 => x"75",
         12670 => x"af",
         12671 => x"b1",
         12672 => x"05",
         12673 => x"51",
         12674 => x"3f",
         12675 => x"08",
         12676 => x"8c",
         12677 => x"8a",
         12678 => x"ba",
         12679 => x"3d",
         12680 => x"a6",
         12681 => x"3d",
         12682 => x"3d",
         12683 => x"ff",
         12684 => x"84",
         12685 => x"56",
         12686 => x"08",
         12687 => x"81",
         12688 => x"81",
         12689 => x"86",
         12690 => x"38",
         12691 => x"3d",
         12692 => x"58",
         12693 => x"70",
         12694 => x"33",
         12695 => x"05",
         12696 => x"15",
         12697 => x"38",
         12698 => x"b0",
         12699 => x"58",
         12700 => x"81",
         12701 => x"77",
         12702 => x"59",
         12703 => x"55",
         12704 => x"b3",
         12705 => x"77",
         12706 => x"d5",
         12707 => x"8c",
         12708 => x"ba",
         12709 => x"d8",
         12710 => x"3d",
         12711 => x"cb",
         12712 => x"84",
         12713 => x"b1",
         12714 => x"76",
         12715 => x"70",
         12716 => x"57",
         12717 => x"89",
         12718 => x"82",
         12719 => x"ff",
         12720 => x"5d",
         12721 => x"2e",
         12722 => x"80",
         12723 => x"e5",
         12724 => x"72",
         12725 => x"5f",
         12726 => x"81",
         12727 => x"79",
         12728 => x"5b",
         12729 => x"12",
         12730 => x"77",
         12731 => x"38",
         12732 => x"81",
         12733 => x"55",
         12734 => x"58",
         12735 => x"89",
         12736 => x"70",
         12737 => x"58",
         12738 => x"70",
         12739 => x"55",
         12740 => x"09",
         12741 => x"38",
         12742 => x"38",
         12743 => x"70",
         12744 => x"07",
         12745 => x"07",
         12746 => x"7a",
         12747 => x"38",
         12748 => x"1e",
         12749 => x"83",
         12750 => x"38",
         12751 => x"5a",
         12752 => x"39",
         12753 => x"fd",
         12754 => x"7f",
         12755 => x"b1",
         12756 => x"05",
         12757 => x"51",
         12758 => x"3f",
         12759 => x"08",
         12760 => x"8c",
         12761 => x"38",
         12762 => x"6c",
         12763 => x"2e",
         12764 => x"fe",
         12765 => x"51",
         12766 => x"3f",
         12767 => x"08",
         12768 => x"8c",
         12769 => x"38",
         12770 => x"0b",
         12771 => x"88",
         12772 => x"05",
         12773 => x"75",
         12774 => x"57",
         12775 => x"81",
         12776 => x"ff",
         12777 => x"ef",
         12778 => x"cb",
         12779 => x"19",
         12780 => x"33",
         12781 => x"81",
         12782 => x"7e",
         12783 => x"a0",
         12784 => x"8b",
         12785 => x"5d",
         12786 => x"1e",
         12787 => x"33",
         12788 => x"81",
         12789 => x"75",
         12790 => x"c5",
         12791 => x"08",
         12792 => x"bd",
         12793 => x"19",
         12794 => x"33",
         12795 => x"07",
         12796 => x"58",
         12797 => x"83",
         12798 => x"38",
         12799 => x"18",
         12800 => x"5e",
         12801 => x"27",
         12802 => x"8a",
         12803 => x"71",
         12804 => x"08",
         12805 => x"75",
         12806 => x"b5",
         12807 => x"5d",
         12808 => x"08",
         12809 => x"38",
         12810 => x"5f",
         12811 => x"38",
         12812 => x"53",
         12813 => x"81",
         12814 => x"fe",
         12815 => x"84",
         12816 => x"80",
         12817 => x"ff",
         12818 => x"77",
         12819 => x"7f",
         12820 => x"d8",
         12821 => x"7b",
         12822 => x"81",
         12823 => x"79",
         12824 => x"81",
         12825 => x"6a",
         12826 => x"ff",
         12827 => x"7b",
         12828 => x"34",
         12829 => x"58",
         12830 => x"18",
         12831 => x"5b",
         12832 => x"09",
         12833 => x"38",
         12834 => x"5e",
         12835 => x"18",
         12836 => x"2a",
         12837 => x"ed",
         12838 => x"57",
         12839 => x"18",
         12840 => x"aa",
         12841 => x"3d",
         12842 => x"56",
         12843 => x"95",
         12844 => x"78",
         12845 => x"a2",
         12846 => x"8c",
         12847 => x"ba",
         12848 => x"f5",
         12849 => x"5c",
         12850 => x"57",
         12851 => x"16",
         12852 => x"b4",
         12853 => x"33",
         12854 => x"7e",
         12855 => x"81",
         12856 => x"38",
         12857 => x"53",
         12858 => x"81",
         12859 => x"fe",
         12860 => x"84",
         12861 => x"80",
         12862 => x"ff",
         12863 => x"76",
         12864 => x"77",
         12865 => x"38",
         12866 => x"5a",
         12867 => x"81",
         12868 => x"34",
         12869 => x"7b",
         12870 => x"80",
         12871 => x"fe",
         12872 => x"84",
         12873 => x"55",
         12874 => x"08",
         12875 => x"98",
         12876 => x"74",
         12877 => x"e1",
         12878 => x"74",
         12879 => x"7f",
         12880 => x"9d",
         12881 => x"8c",
         12882 => x"8c",
         12883 => x"0d",
         12884 => x"84",
         12885 => x"b1",
         12886 => x"95",
         12887 => x"19",
         12888 => x"2b",
         12889 => x"07",
         12890 => x"56",
         12891 => x"39",
         12892 => x"08",
         12893 => x"fe",
         12894 => x"8c",
         12895 => x"fe",
         12896 => x"84",
         12897 => x"b1",
         12898 => x"81",
         12899 => x"08",
         12900 => x"81",
         12901 => x"fe",
         12902 => x"81",
         12903 => x"8c",
         12904 => x"09",
         12905 => x"db",
         12906 => x"8c",
         12907 => x"34",
         12908 => x"a8",
         12909 => x"84",
         12910 => x"59",
         12911 => x"17",
         12912 => x"a0",
         12913 => x"33",
         12914 => x"2e",
         12915 => x"fe",
         12916 => x"54",
         12917 => x"a0",
         12918 => x"53",
         12919 => x"16",
         12920 => x"e1",
         12921 => x"58",
         12922 => x"81",
         12923 => x"08",
         12924 => x"70",
         12925 => x"33",
         12926 => x"e1",
         12927 => x"5c",
         12928 => x"08",
         12929 => x"84",
         12930 => x"83",
         12931 => x"17",
         12932 => x"08",
         12933 => x"8c",
         12934 => x"74",
         12935 => x"27",
         12936 => x"82",
         12937 => x"7c",
         12938 => x"81",
         12939 => x"38",
         12940 => x"17",
         12941 => x"08",
         12942 => x"52",
         12943 => x"51",
         12944 => x"3f",
         12945 => x"e8",
         12946 => x"0d",
         12947 => x"05",
         12948 => x"05",
         12949 => x"33",
         12950 => x"53",
         12951 => x"05",
         12952 => x"51",
         12953 => x"3f",
         12954 => x"08",
         12955 => x"8c",
         12956 => x"8a",
         12957 => x"ba",
         12958 => x"3d",
         12959 => x"5a",
         12960 => x"3d",
         12961 => x"ff",
         12962 => x"84",
         12963 => x"56",
         12964 => x"08",
         12965 => x"80",
         12966 => x"81",
         12967 => x"86",
         12968 => x"38",
         12969 => x"61",
         12970 => x"12",
         12971 => x"7a",
         12972 => x"51",
         12973 => x"73",
         12974 => x"78",
         12975 => x"83",
         12976 => x"51",
         12977 => x"3f",
         12978 => x"08",
         12979 => x"0c",
         12980 => x"04",
         12981 => x"67",
         12982 => x"96",
         12983 => x"52",
         12984 => x"ff",
         12985 => x"84",
         12986 => x"55",
         12987 => x"08",
         12988 => x"38",
         12989 => x"8c",
         12990 => x"0d",
         12991 => x"66",
         12992 => x"d0",
         12993 => x"95",
         12994 => x"ba",
         12995 => x"84",
         12996 => x"e0",
         12997 => x"cf",
         12998 => x"a0",
         12999 => x"55",
         13000 => x"60",
         13001 => x"86",
         13002 => x"90",
         13003 => x"59",
         13004 => x"17",
         13005 => x"2a",
         13006 => x"17",
         13007 => x"2a",
         13008 => x"17",
         13009 => x"2a",
         13010 => x"17",
         13011 => x"81",
         13012 => x"34",
         13013 => x"e1",
         13014 => x"ba",
         13015 => x"ba",
         13016 => x"3d",
         13017 => x"3d",
         13018 => x"5d",
         13019 => x"9a",
         13020 => x"52",
         13021 => x"ff",
         13022 => x"84",
         13023 => x"84",
         13024 => x"30",
         13025 => x"8c",
         13026 => x"25",
         13027 => x"7a",
         13028 => x"38",
         13029 => x"06",
         13030 => x"81",
         13031 => x"30",
         13032 => x"80",
         13033 => x"7b",
         13034 => x"8c",
         13035 => x"76",
         13036 => x"78",
         13037 => x"80",
         13038 => x"11",
         13039 => x"80",
         13040 => x"08",
         13041 => x"f6",
         13042 => x"33",
         13043 => x"74",
         13044 => x"81",
         13045 => x"38",
         13046 => x"53",
         13047 => x"81",
         13048 => x"fe",
         13049 => x"84",
         13050 => x"80",
         13051 => x"ff",
         13052 => x"76",
         13053 => x"78",
         13054 => x"38",
         13055 => x"56",
         13056 => x"56",
         13057 => x"8b",
         13058 => x"56",
         13059 => x"83",
         13060 => x"75",
         13061 => x"83",
         13062 => x"12",
         13063 => x"2b",
         13064 => x"07",
         13065 => x"70",
         13066 => x"2b",
         13067 => x"07",
         13068 => x"5d",
         13069 => x"56",
         13070 => x"8c",
         13071 => x"0d",
         13072 => x"80",
         13073 => x"8e",
         13074 => x"55",
         13075 => x"3f",
         13076 => x"08",
         13077 => x"8c",
         13078 => x"81",
         13079 => x"84",
         13080 => x"06",
         13081 => x"80",
         13082 => x"57",
         13083 => x"77",
         13084 => x"08",
         13085 => x"70",
         13086 => x"33",
         13087 => x"dc",
         13088 => x"59",
         13089 => x"08",
         13090 => x"81",
         13091 => x"38",
         13092 => x"08",
         13093 => x"b4",
         13094 => x"17",
         13095 => x"ba",
         13096 => x"55",
         13097 => x"08",
         13098 => x"38",
         13099 => x"55",
         13100 => x"09",
         13101 => x"a0",
         13102 => x"b4",
         13103 => x"17",
         13104 => x"7a",
         13105 => x"33",
         13106 => x"e2",
         13107 => x"81",
         13108 => x"b8",
         13109 => x"16",
         13110 => x"da",
         13111 => x"ba",
         13112 => x"2e",
         13113 => x"fe",
         13114 => x"52",
         13115 => x"f8",
         13116 => x"ba",
         13117 => x"84",
         13118 => x"fe",
         13119 => x"ba",
         13120 => x"ba",
         13121 => x"5c",
         13122 => x"18",
         13123 => x"1b",
         13124 => x"75",
         13125 => x"81",
         13126 => x"78",
         13127 => x"8b",
         13128 => x"58",
         13129 => x"77",
         13130 => x"f2",
         13131 => x"7b",
         13132 => x"5c",
         13133 => x"a0",
         13134 => x"fc",
         13135 => x"57",
         13136 => x"e1",
         13137 => x"53",
         13138 => x"b4",
         13139 => x"3d",
         13140 => x"eb",
         13141 => x"8c",
         13142 => x"ba",
         13143 => x"a6",
         13144 => x"5d",
         13145 => x"55",
         13146 => x"81",
         13147 => x"ff",
         13148 => x"f4",
         13149 => x"3d",
         13150 => x"70",
         13151 => x"5b",
         13152 => x"9f",
         13153 => x"b7",
         13154 => x"90",
         13155 => x"75",
         13156 => x"81",
         13157 => x"74",
         13158 => x"75",
         13159 => x"83",
         13160 => x"81",
         13161 => x"51",
         13162 => x"83",
         13163 => x"ba",
         13164 => x"9f",
         13165 => x"ba",
         13166 => x"ff",
         13167 => x"76",
         13168 => x"e0",
         13169 => x"9c",
         13170 => x"9c",
         13171 => x"ff",
         13172 => x"58",
         13173 => x"81",
         13174 => x"56",
         13175 => x"99",
         13176 => x"70",
         13177 => x"ff",
         13178 => x"58",
         13179 => x"89",
         13180 => x"2e",
         13181 => x"e9",
         13182 => x"ff",
         13183 => x"81",
         13184 => x"ff",
         13185 => x"f8",
         13186 => x"26",
         13187 => x"81",
         13188 => x"8f",
         13189 => x"2a",
         13190 => x"70",
         13191 => x"34",
         13192 => x"76",
         13193 => x"05",
         13194 => x"1a",
         13195 => x"70",
         13196 => x"ff",
         13197 => x"58",
         13198 => x"26",
         13199 => x"8f",
         13200 => x"86",
         13201 => x"e5",
         13202 => x"79",
         13203 => x"38",
         13204 => x"56",
         13205 => x"33",
         13206 => x"a0",
         13207 => x"06",
         13208 => x"1a",
         13209 => x"38",
         13210 => x"47",
         13211 => x"3d",
         13212 => x"fe",
         13213 => x"84",
         13214 => x"55",
         13215 => x"08",
         13216 => x"38",
         13217 => x"84",
         13218 => x"a1",
         13219 => x"83",
         13220 => x"51",
         13221 => x"84",
         13222 => x"83",
         13223 => x"55",
         13224 => x"38",
         13225 => x"84",
         13226 => x"a1",
         13227 => x"83",
         13228 => x"56",
         13229 => x"81",
         13230 => x"fe",
         13231 => x"84",
         13232 => x"55",
         13233 => x"08",
         13234 => x"79",
         13235 => x"c4",
         13236 => x"7e",
         13237 => x"76",
         13238 => x"58",
         13239 => x"81",
         13240 => x"ff",
         13241 => x"ef",
         13242 => x"81",
         13243 => x"34",
         13244 => x"d9",
         13245 => x"ba",
         13246 => x"74",
         13247 => x"39",
         13248 => x"fe",
         13249 => x"56",
         13250 => x"84",
         13251 => x"84",
         13252 => x"06",
         13253 => x"80",
         13254 => x"2e",
         13255 => x"75",
         13256 => x"76",
         13257 => x"ee",
         13258 => x"ba",
         13259 => x"84",
         13260 => x"75",
         13261 => x"06",
         13262 => x"84",
         13263 => x"b8",
         13264 => x"98",
         13265 => x"80",
         13266 => x"08",
         13267 => x"38",
         13268 => x"55",
         13269 => x"09",
         13270 => x"d7",
         13271 => x"76",
         13272 => x"52",
         13273 => x"51",
         13274 => x"3f",
         13275 => x"08",
         13276 => x"38",
         13277 => x"59",
         13278 => x"0c",
         13279 => x"be",
         13280 => x"17",
         13281 => x"57",
         13282 => x"81",
         13283 => x"9e",
         13284 => x"70",
         13285 => x"07",
         13286 => x"80",
         13287 => x"38",
         13288 => x"79",
         13289 => x"38",
         13290 => x"51",
         13291 => x"3f",
         13292 => x"08",
         13293 => x"8c",
         13294 => x"ff",
         13295 => x"55",
         13296 => x"fd",
         13297 => x"55",
         13298 => x"38",
         13299 => x"55",
         13300 => x"81",
         13301 => x"ff",
         13302 => x"f4",
         13303 => x"88",
         13304 => x"34",
         13305 => x"59",
         13306 => x"70",
         13307 => x"33",
         13308 => x"05",
         13309 => x"15",
         13310 => x"2e",
         13311 => x"76",
         13312 => x"58",
         13313 => x"81",
         13314 => x"ff",
         13315 => x"da",
         13316 => x"39",
         13317 => x"7a",
         13318 => x"81",
         13319 => x"34",
         13320 => x"d7",
         13321 => x"ba",
         13322 => x"fd",
         13323 => x"57",
         13324 => x"81",
         13325 => x"08",
         13326 => x"81",
         13327 => x"fe",
         13328 => x"84",
         13329 => x"79",
         13330 => x"06",
         13331 => x"84",
         13332 => x"83",
         13333 => x"18",
         13334 => x"08",
         13335 => x"a0",
         13336 => x"8a",
         13337 => x"33",
         13338 => x"2e",
         13339 => x"ba",
         13340 => x"fd",
         13341 => x"5a",
         13342 => x"51",
         13343 => x"3f",
         13344 => x"08",
         13345 => x"8c",
         13346 => x"fd",
         13347 => x"ae",
         13348 => x"58",
         13349 => x"2e",
         13350 => x"fe",
         13351 => x"54",
         13352 => x"a0",
         13353 => x"53",
         13354 => x"18",
         13355 => x"d3",
         13356 => x"a9",
         13357 => x"0d",
         13358 => x"88",
         13359 => x"05",
         13360 => x"57",
         13361 => x"80",
         13362 => x"76",
         13363 => x"80",
         13364 => x"74",
         13365 => x"80",
         13366 => x"86",
         13367 => x"18",
         13368 => x"78",
         13369 => x"c2",
         13370 => x"73",
         13371 => x"a5",
         13372 => x"33",
         13373 => x"9d",
         13374 => x"2e",
         13375 => x"8c",
         13376 => x"9c",
         13377 => x"33",
         13378 => x"81",
         13379 => x"74",
         13380 => x"8c",
         13381 => x"11",
         13382 => x"2b",
         13383 => x"54",
         13384 => x"fd",
         13385 => x"ff",
         13386 => x"70",
         13387 => x"07",
         13388 => x"ba",
         13389 => x"90",
         13390 => x"42",
         13391 => x"58",
         13392 => x"88",
         13393 => x"08",
         13394 => x"38",
         13395 => x"78",
         13396 => x"59",
         13397 => x"51",
         13398 => x"3f",
         13399 => x"55",
         13400 => x"08",
         13401 => x"38",
         13402 => x"ba",
         13403 => x"2e",
         13404 => x"84",
         13405 => x"ff",
         13406 => x"38",
         13407 => x"08",
         13408 => x"81",
         13409 => x"7d",
         13410 => x"74",
         13411 => x"81",
         13412 => x"87",
         13413 => x"73",
         13414 => x"0c",
         13415 => x"04",
         13416 => x"ba",
         13417 => x"3d",
         13418 => x"15",
         13419 => x"d0",
         13420 => x"ba",
         13421 => x"06",
         13422 => x"ad",
         13423 => x"08",
         13424 => x"a7",
         13425 => x"2e",
         13426 => x"7a",
         13427 => x"7c",
         13428 => x"38",
         13429 => x"74",
         13430 => x"e6",
         13431 => x"77",
         13432 => x"fe",
         13433 => x"84",
         13434 => x"56",
         13435 => x"08",
         13436 => x"77",
         13437 => x"17",
         13438 => x"74",
         13439 => x"7e",
         13440 => x"55",
         13441 => x"ff",
         13442 => x"88",
         13443 => x"8c",
         13444 => x"17",
         13445 => x"07",
         13446 => x"18",
         13447 => x"08",
         13448 => x"16",
         13449 => x"76",
         13450 => x"e9",
         13451 => x"31",
         13452 => x"84",
         13453 => x"07",
         13454 => x"16",
         13455 => x"fe",
         13456 => x"54",
         13457 => x"74",
         13458 => x"fe",
         13459 => x"54",
         13460 => x"81",
         13461 => x"39",
         13462 => x"ff",
         13463 => x"ba",
         13464 => x"3d",
         13465 => x"08",
         13466 => x"02",
         13467 => x"87",
         13468 => x"42",
         13469 => x"a2",
         13470 => x"5f",
         13471 => x"80",
         13472 => x"38",
         13473 => x"05",
         13474 => x"9f",
         13475 => x"75",
         13476 => x"9b",
         13477 => x"38",
         13478 => x"85",
         13479 => x"d1",
         13480 => x"80",
         13481 => x"e5",
         13482 => x"10",
         13483 => x"05",
         13484 => x"5a",
         13485 => x"84",
         13486 => x"34",
         13487 => x"ba",
         13488 => x"84",
         13489 => x"33",
         13490 => x"81",
         13491 => x"fe",
         13492 => x"84",
         13493 => x"81",
         13494 => x"81",
         13495 => x"83",
         13496 => x"ab",
         13497 => x"2a",
         13498 => x"8a",
         13499 => x"9f",
         13500 => x"fc",
         13501 => x"52",
         13502 => x"d0",
         13503 => x"ba",
         13504 => x"98",
         13505 => x"74",
         13506 => x"90",
         13507 => x"80",
         13508 => x"88",
         13509 => x"75",
         13510 => x"83",
         13511 => x"80",
         13512 => x"84",
         13513 => x"83",
         13514 => x"81",
         13515 => x"83",
         13516 => x"1f",
         13517 => x"74",
         13518 => x"7e",
         13519 => x"3d",
         13520 => x"70",
         13521 => x"59",
         13522 => x"60",
         13523 => x"ab",
         13524 => x"70",
         13525 => x"07",
         13526 => x"57",
         13527 => x"38",
         13528 => x"84",
         13529 => x"54",
         13530 => x"52",
         13531 => x"cd",
         13532 => x"57",
         13533 => x"08",
         13534 => x"60",
         13535 => x"33",
         13536 => x"05",
         13537 => x"2b",
         13538 => x"8e",
         13539 => x"d4",
         13540 => x"81",
         13541 => x"38",
         13542 => x"61",
         13543 => x"11",
         13544 => x"62",
         13545 => x"e7",
         13546 => x"18",
         13547 => x"82",
         13548 => x"90",
         13549 => x"2b",
         13550 => x"33",
         13551 => x"88",
         13552 => x"71",
         13553 => x"1f",
         13554 => x"82",
         13555 => x"90",
         13556 => x"2b",
         13557 => x"33",
         13558 => x"88",
         13559 => x"71",
         13560 => x"3d",
         13561 => x"3d",
         13562 => x"0c",
         13563 => x"45",
         13564 => x"5a",
         13565 => x"8e",
         13566 => x"79",
         13567 => x"38",
         13568 => x"81",
         13569 => x"87",
         13570 => x"2a",
         13571 => x"45",
         13572 => x"2e",
         13573 => x"61",
         13574 => x"64",
         13575 => x"38",
         13576 => x"47",
         13577 => x"38",
         13578 => x"30",
         13579 => x"7a",
         13580 => x"2e",
         13581 => x"7a",
         13582 => x"8c",
         13583 => x"0b",
         13584 => x"22",
         13585 => x"80",
         13586 => x"74",
         13587 => x"38",
         13588 => x"56",
         13589 => x"17",
         13590 => x"57",
         13591 => x"2e",
         13592 => x"75",
         13593 => x"77",
         13594 => x"fd",
         13595 => x"84",
         13596 => x"10",
         13597 => x"84",
         13598 => x"9f",
         13599 => x"38",
         13600 => x"ba",
         13601 => x"84",
         13602 => x"05",
         13603 => x"2a",
         13604 => x"4c",
         13605 => x"15",
         13606 => x"81",
         13607 => x"7b",
         13608 => x"68",
         13609 => x"ff",
         13610 => x"06",
         13611 => x"4e",
         13612 => x"83",
         13613 => x"38",
         13614 => x"77",
         13615 => x"70",
         13616 => x"57",
         13617 => x"82",
         13618 => x"7c",
         13619 => x"78",
         13620 => x"31",
         13621 => x"ff",
         13622 => x"ba",
         13623 => x"62",
         13624 => x"f6",
         13625 => x"2e",
         13626 => x"82",
         13627 => x"ff",
         13628 => x"ba",
         13629 => x"82",
         13630 => x"89",
         13631 => x"18",
         13632 => x"c0",
         13633 => x"38",
         13634 => x"a3",
         13635 => x"76",
         13636 => x"0c",
         13637 => x"84",
         13638 => x"04",
         13639 => x"fe",
         13640 => x"84",
         13641 => x"9f",
         13642 => x"ba",
         13643 => x"7c",
         13644 => x"70",
         13645 => x"57",
         13646 => x"89",
         13647 => x"82",
         13648 => x"ff",
         13649 => x"5d",
         13650 => x"2e",
         13651 => x"80",
         13652 => x"fc",
         13653 => x"08",
         13654 => x"7a",
         13655 => x"5c",
         13656 => x"81",
         13657 => x"ff",
         13658 => x"59",
         13659 => x"26",
         13660 => x"17",
         13661 => x"06",
         13662 => x"9f",
         13663 => x"99",
         13664 => x"e0",
         13665 => x"ff",
         13666 => x"76",
         13667 => x"2a",
         13668 => x"78",
         13669 => x"06",
         13670 => x"ff",
         13671 => x"7a",
         13672 => x"70",
         13673 => x"2a",
         13674 => x"4a",
         13675 => x"2e",
         13676 => x"81",
         13677 => x"5f",
         13678 => x"25",
         13679 => x"7f",
         13680 => x"39",
         13681 => x"05",
         13682 => x"79",
         13683 => x"dd",
         13684 => x"84",
         13685 => x"fe",
         13686 => x"83",
         13687 => x"84",
         13688 => x"40",
         13689 => x"38",
         13690 => x"55",
         13691 => x"75",
         13692 => x"38",
         13693 => x"59",
         13694 => x"81",
         13695 => x"39",
         13696 => x"ff",
         13697 => x"7a",
         13698 => x"56",
         13699 => x"61",
         13700 => x"93",
         13701 => x"2e",
         13702 => x"82",
         13703 => x"4a",
         13704 => x"8b",
         13705 => x"8c",
         13706 => x"26",
         13707 => x"8b",
         13708 => x"5b",
         13709 => x"27",
         13710 => x"8e",
         13711 => x"ba",
         13712 => x"3d",
         13713 => x"98",
         13714 => x"55",
         13715 => x"86",
         13716 => x"f5",
         13717 => x"38",
         13718 => x"5b",
         13719 => x"fd",
         13720 => x"80",
         13721 => x"80",
         13722 => x"05",
         13723 => x"15",
         13724 => x"38",
         13725 => x"e5",
         13726 => x"55",
         13727 => x"05",
         13728 => x"70",
         13729 => x"34",
         13730 => x"74",
         13731 => x"8b",
         13732 => x"65",
         13733 => x"8c",
         13734 => x"61",
         13735 => x"7b",
         13736 => x"06",
         13737 => x"8e",
         13738 => x"88",
         13739 => x"61",
         13740 => x"81",
         13741 => x"34",
         13742 => x"70",
         13743 => x"80",
         13744 => x"34",
         13745 => x"82",
         13746 => x"61",
         13747 => x"6c",
         13748 => x"ff",
         13749 => x"ad",
         13750 => x"ff",
         13751 => x"74",
         13752 => x"34",
         13753 => x"4c",
         13754 => x"05",
         13755 => x"95",
         13756 => x"61",
         13757 => x"80",
         13758 => x"34",
         13759 => x"05",
         13760 => x"9b",
         13761 => x"61",
         13762 => x"7e",
         13763 => x"67",
         13764 => x"34",
         13765 => x"4c",
         13766 => x"05",
         13767 => x"2a",
         13768 => x"0c",
         13769 => x"08",
         13770 => x"34",
         13771 => x"85",
         13772 => x"61",
         13773 => x"80",
         13774 => x"34",
         13775 => x"05",
         13776 => x"61",
         13777 => x"7c",
         13778 => x"06",
         13779 => x"96",
         13780 => x"88",
         13781 => x"61",
         13782 => x"ff",
         13783 => x"05",
         13784 => x"a6",
         13785 => x"61",
         13786 => x"e5",
         13787 => x"55",
         13788 => x"05",
         13789 => x"70",
         13790 => x"34",
         13791 => x"74",
         13792 => x"83",
         13793 => x"80",
         13794 => x"60",
         13795 => x"4b",
         13796 => x"34",
         13797 => x"53",
         13798 => x"51",
         13799 => x"3f",
         13800 => x"ba",
         13801 => x"e7",
         13802 => x"5c",
         13803 => x"87",
         13804 => x"61",
         13805 => x"76",
         13806 => x"58",
         13807 => x"55",
         13808 => x"63",
         13809 => x"62",
         13810 => x"c0",
         13811 => x"ff",
         13812 => x"81",
         13813 => x"f8",
         13814 => x"34",
         13815 => x"7c",
         13816 => x"64",
         13817 => x"46",
         13818 => x"2a",
         13819 => x"70",
         13820 => x"34",
         13821 => x"56",
         13822 => x"7c",
         13823 => x"76",
         13824 => x"38",
         13825 => x"54",
         13826 => x"52",
         13827 => x"c5",
         13828 => x"ba",
         13829 => x"e6",
         13830 => x"61",
         13831 => x"76",
         13832 => x"58",
         13833 => x"55",
         13834 => x"78",
         13835 => x"31",
         13836 => x"c9",
         13837 => x"05",
         13838 => x"2e",
         13839 => x"77",
         13840 => x"2e",
         13841 => x"56",
         13842 => x"66",
         13843 => x"75",
         13844 => x"7a",
         13845 => x"79",
         13846 => x"d2",
         13847 => x"8c",
         13848 => x"38",
         13849 => x"76",
         13850 => x"75",
         13851 => x"58",
         13852 => x"93",
         13853 => x"6c",
         13854 => x"26",
         13855 => x"58",
         13856 => x"83",
         13857 => x"7d",
         13858 => x"61",
         13859 => x"06",
         13860 => x"b3",
         13861 => x"61",
         13862 => x"75",
         13863 => x"57",
         13864 => x"59",
         13865 => x"80",
         13866 => x"ff",
         13867 => x"60",
         13868 => x"47",
         13869 => x"81",
         13870 => x"34",
         13871 => x"05",
         13872 => x"83",
         13873 => x"67",
         13874 => x"6c",
         13875 => x"c1",
         13876 => x"51",
         13877 => x"3f",
         13878 => x"05",
         13879 => x"8c",
         13880 => x"bf",
         13881 => x"67",
         13882 => x"84",
         13883 => x"67",
         13884 => x"7e",
         13885 => x"05",
         13886 => x"83",
         13887 => x"6b",
         13888 => x"05",
         13889 => x"98",
         13890 => x"c9",
         13891 => x"61",
         13892 => x"34",
         13893 => x"45",
         13894 => x"cb",
         13895 => x"90",
         13896 => x"61",
         13897 => x"34",
         13898 => x"5f",
         13899 => x"cd",
         13900 => x"54",
         13901 => x"52",
         13902 => x"c2",
         13903 => x"57",
         13904 => x"08",
         13905 => x"80",
         13906 => x"79",
         13907 => x"dd",
         13908 => x"84",
         13909 => x"f7",
         13910 => x"ba",
         13911 => x"ba",
         13912 => x"3d",
         13913 => x"98",
         13914 => x"55",
         13915 => x"74",
         13916 => x"45",
         13917 => x"39",
         13918 => x"78",
         13919 => x"81",
         13920 => x"c0",
         13921 => x"74",
         13922 => x"38",
         13923 => x"98",
         13924 => x"c0",
         13925 => x"82",
         13926 => x"57",
         13927 => x"80",
         13928 => x"76",
         13929 => x"38",
         13930 => x"51",
         13931 => x"3f",
         13932 => x"08",
         13933 => x"87",
         13934 => x"2a",
         13935 => x"5c",
         13936 => x"ba",
         13937 => x"80",
         13938 => x"47",
         13939 => x"0a",
         13940 => x"cb",
         13941 => x"f8",
         13942 => x"ba",
         13943 => x"ff",
         13944 => x"e6",
         13945 => x"d3",
         13946 => x"2a",
         13947 => x"bf",
         13948 => x"f8",
         13949 => x"81",
         13950 => x"80",
         13951 => x"38",
         13952 => x"ab",
         13953 => x"a0",
         13954 => x"88",
         13955 => x"61",
         13956 => x"75",
         13957 => x"7a",
         13958 => x"34",
         13959 => x"57",
         13960 => x"05",
         13961 => x"39",
         13962 => x"c3",
         13963 => x"61",
         13964 => x"34",
         13965 => x"c5",
         13966 => x"cc",
         13967 => x"05",
         13968 => x"a4",
         13969 => x"88",
         13970 => x"61",
         13971 => x"7c",
         13972 => x"78",
         13973 => x"34",
         13974 => x"56",
         13975 => x"05",
         13976 => x"ac",
         13977 => x"61",
         13978 => x"80",
         13979 => x"34",
         13980 => x"05",
         13981 => x"b0",
         13982 => x"61",
         13983 => x"86",
         13984 => x"34",
         13985 => x"05",
         13986 => x"61",
         13987 => x"34",
         13988 => x"c2",
         13989 => x"61",
         13990 => x"83",
         13991 => x"57",
         13992 => x"81",
         13993 => x"76",
         13994 => x"58",
         13995 => x"55",
         13996 => x"f9",
         13997 => x"70",
         13998 => x"33",
         13999 => x"05",
         14000 => x"15",
         14001 => x"38",
         14002 => x"81",
         14003 => x"60",
         14004 => x"fe",
         14005 => x"81",
         14006 => x"8c",
         14007 => x"38",
         14008 => x"61",
         14009 => x"62",
         14010 => x"34",
         14011 => x"ba",
         14012 => x"60",
         14013 => x"fe",
         14014 => x"fc",
         14015 => x"0b",
         14016 => x"0c",
         14017 => x"84",
         14018 => x"04",
         14019 => x"7b",
         14020 => x"70",
         14021 => x"34",
         14022 => x"81",
         14023 => x"ff",
         14024 => x"61",
         14025 => x"ff",
         14026 => x"34",
         14027 => x"05",
         14028 => x"87",
         14029 => x"61",
         14030 => x"ff",
         14031 => x"34",
         14032 => x"05",
         14033 => x"34",
         14034 => x"b1",
         14035 => x"86",
         14036 => x"52",
         14037 => x"be",
         14038 => x"80",
         14039 => x"80",
         14040 => x"05",
         14041 => x"17",
         14042 => x"38",
         14043 => x"d2",
         14044 => x"05",
         14045 => x"55",
         14046 => x"70",
         14047 => x"34",
         14048 => x"70",
         14049 => x"34",
         14050 => x"34",
         14051 => x"83",
         14052 => x"80",
         14053 => x"e5",
         14054 => x"c1",
         14055 => x"05",
         14056 => x"61",
         14057 => x"34",
         14058 => x"5b",
         14059 => x"e8",
         14060 => x"88",
         14061 => x"61",
         14062 => x"34",
         14063 => x"56",
         14064 => x"ea",
         14065 => x"98",
         14066 => x"61",
         14067 => x"34",
         14068 => x"ec",
         14069 => x"61",
         14070 => x"34",
         14071 => x"ee",
         14072 => x"61",
         14073 => x"34",
         14074 => x"34",
         14075 => x"34",
         14076 => x"1f",
         14077 => x"79",
         14078 => x"b2",
         14079 => x"81",
         14080 => x"52",
         14081 => x"bd",
         14082 => x"61",
         14083 => x"a6",
         14084 => x"0d",
         14085 => x"5b",
         14086 => x"ff",
         14087 => x"57",
         14088 => x"b8",
         14089 => x"59",
         14090 => x"05",
         14091 => x"78",
         14092 => x"ff",
         14093 => x"7b",
         14094 => x"81",
         14095 => x"8d",
         14096 => x"74",
         14097 => x"38",
         14098 => x"81",
         14099 => x"81",
         14100 => x"8a",
         14101 => x"77",
         14102 => x"38",
         14103 => x"7a",
         14104 => x"38",
         14105 => x"84",
         14106 => x"8e",
         14107 => x"f7",
         14108 => x"02",
         14109 => x"05",
         14110 => x"77",
         14111 => x"d5",
         14112 => x"08",
         14113 => x"24",
         14114 => x"17",
         14115 => x"8c",
         14116 => x"77",
         14117 => x"16",
         14118 => x"24",
         14119 => x"84",
         14120 => x"19",
         14121 => x"8b",
         14122 => x"8b",
         14123 => x"54",
         14124 => x"17",
         14125 => x"51",
         14126 => x"3f",
         14127 => x"70",
         14128 => x"07",
         14129 => x"30",
         14130 => x"81",
         14131 => x"0c",
         14132 => x"d3",
         14133 => x"76",
         14134 => x"3f",
         14135 => x"e3",
         14136 => x"80",
         14137 => x"8d",
         14138 => x"80",
         14139 => x"55",
         14140 => x"81",
         14141 => x"ff",
         14142 => x"f4",
         14143 => x"08",
         14144 => x"8a",
         14145 => x"38",
         14146 => x"76",
         14147 => x"38",
         14148 => x"8c",
         14149 => x"77",
         14150 => x"16",
         14151 => x"24",
         14152 => x"84",
         14153 => x"19",
         14154 => x"7c",
         14155 => x"24",
         14156 => x"3d",
         14157 => x"55",
         14158 => x"05",
         14159 => x"51",
         14160 => x"3f",
         14161 => x"08",
         14162 => x"7a",
         14163 => x"ff",
         14164 => x"8c",
         14165 => x"0d",
         14166 => x"ff",
         14167 => x"75",
         14168 => x"52",
         14169 => x"ff",
         14170 => x"74",
         14171 => x"30",
         14172 => x"9f",
         14173 => x"52",
         14174 => x"ff",
         14175 => x"52",
         14176 => x"eb",
         14177 => x"39",
         14178 => x"8c",
         14179 => x"0d",
         14180 => x"0d",
         14181 => x"05",
         14182 => x"52",
         14183 => x"72",
         14184 => x"90",
         14185 => x"ff",
         14186 => x"71",
         14187 => x"0c",
         14188 => x"04",
         14189 => x"73",
         14190 => x"83",
         14191 => x"81",
         14192 => x"73",
         14193 => x"38",
         14194 => x"22",
         14195 => x"2e",
         14196 => x"12",
         14197 => x"ff",
         14198 => x"71",
         14199 => x"8d",
         14200 => x"83",
         14201 => x"70",
         14202 => x"e1",
         14203 => x"12",
         14204 => x"06",
         14205 => x"0c",
         14206 => x"0d",
         14207 => x"0d",
         14208 => x"22",
         14209 => x"96",
         14210 => x"51",
         14211 => x"80",
         14212 => x"38",
         14213 => x"84",
         14214 => x"84",
         14215 => x"71",
         14216 => x"09",
         14217 => x"38",
         14218 => x"26",
         14219 => x"10",
         14220 => x"05",
         14221 => x"ba",
         14222 => x"84",
         14223 => x"fb",
         14224 => x"51",
         14225 => x"ff",
         14226 => x"38",
         14227 => x"ff",
         14228 => x"d0",
         14229 => x"9f",
         14230 => x"d9",
         14231 => x"82",
         14232 => x"75",
         14233 => x"80",
         14234 => x"26",
         14235 => x"53",
         14236 => x"38",
         14237 => x"05",
         14238 => x"71",
         14239 => x"56",
         14240 => x"70",
         14241 => x"70",
         14242 => x"38",
         14243 => x"73",
         14244 => x"70",
         14245 => x"22",
         14246 => x"70",
         14247 => x"79",
         14248 => x"55",
         14249 => x"2e",
         14250 => x"51",
         14251 => x"8c",
         14252 => x"0d",
         14253 => x"c4",
         14254 => x"39",
         14255 => x"ea",
         14256 => x"10",
         14257 => x"05",
         14258 => x"04",
         14259 => x"70",
         14260 => x"06",
         14261 => x"51",
         14262 => x"b0",
         14263 => x"ff",
         14264 => x"51",
         14265 => x"16",
         14266 => x"ff",
         14267 => x"e6",
         14268 => x"70",
         14269 => x"06",
         14270 => x"39",
         14271 => x"83",
         14272 => x"57",
         14273 => x"e0",
         14274 => x"ff",
         14275 => x"51",
         14276 => x"16",
         14277 => x"ff",
         14278 => x"ff",
         14279 => x"73",
         14280 => x"76",
         14281 => x"83",
         14282 => x"58",
         14283 => x"a6",
         14284 => x"31",
         14285 => x"70",
         14286 => x"fe",
         14287 => x"00",
         14288 => x"ff",
         14289 => x"ff",
         14290 => x"ff",
         14291 => x"00",
         14292 => x"00",
         14293 => x"00",
         14294 => x"00",
         14295 => x"00",
         14296 => x"00",
         14297 => x"00",
         14298 => x"00",
         14299 => x"00",
         14300 => x"00",
         14301 => x"00",
         14302 => x"00",
         14303 => x"00",
         14304 => x"00",
         14305 => x"00",
         14306 => x"00",
         14307 => x"00",
         14308 => x"00",
         14309 => x"00",
         14310 => x"00",
         14311 => x"00",
         14312 => x"00",
         14313 => x"00",
         14314 => x"00",
         14315 => x"00",
         14316 => x"00",
         14317 => x"00",
         14318 => x"00",
         14319 => x"00",
         14320 => x"00",
         14321 => x"00",
         14322 => x"00",
         14323 => x"00",
         14324 => x"00",
         14325 => x"00",
         14326 => x"00",
         14327 => x"00",
         14328 => x"00",
         14329 => x"00",
         14330 => x"00",
         14331 => x"00",
         14332 => x"00",
         14333 => x"00",
         14334 => x"00",
         14335 => x"00",
         14336 => x"00",
         14337 => x"00",
         14338 => x"00",
         14339 => x"00",
         14340 => x"00",
         14341 => x"00",
         14342 => x"00",
         14343 => x"00",
         14344 => x"00",
         14345 => x"00",
         14346 => x"00",
         14347 => x"00",
         14348 => x"00",
         14349 => x"00",
         14350 => x"00",
         14351 => x"00",
         14352 => x"00",
         14353 => x"00",
         14354 => x"00",
         14355 => x"00",
         14356 => x"00",
         14357 => x"00",
         14358 => x"00",
         14359 => x"00",
         14360 => x"00",
         14361 => x"00",
         14362 => x"00",
         14363 => x"00",
         14364 => x"00",
         14365 => x"00",
         14366 => x"00",
         14367 => x"00",
         14368 => x"00",
         14369 => x"00",
         14370 => x"00",
         14371 => x"00",
         14372 => x"00",
         14373 => x"00",
         14374 => x"00",
         14375 => x"00",
         14376 => x"00",
         14377 => x"00",
         14378 => x"00",
         14379 => x"00",
         14380 => x"00",
         14381 => x"00",
         14382 => x"00",
         14383 => x"00",
         14384 => x"00",
         14385 => x"00",
         14386 => x"00",
         14387 => x"00",
         14388 => x"00",
         14389 => x"00",
         14390 => x"00",
         14391 => x"00",
         14392 => x"00",
         14393 => x"00",
         14394 => x"00",
         14395 => x"00",
         14396 => x"00",
         14397 => x"00",
         14398 => x"00",
         14399 => x"00",
         14400 => x"00",
         14401 => x"00",
         14402 => x"00",
         14403 => x"00",
         14404 => x"00",
         14405 => x"00",
         14406 => x"00",
         14407 => x"00",
         14408 => x"00",
         14409 => x"00",
         14410 => x"00",
         14411 => x"00",
         14412 => x"00",
         14413 => x"00",
         14414 => x"00",
         14415 => x"00",
         14416 => x"00",
         14417 => x"00",
         14418 => x"00",
         14419 => x"00",
         14420 => x"00",
         14421 => x"00",
         14422 => x"00",
         14423 => x"00",
         14424 => x"00",
         14425 => x"00",
         14426 => x"00",
         14427 => x"00",
         14428 => x"00",
         14429 => x"00",
         14430 => x"00",
         14431 => x"00",
         14432 => x"00",
         14433 => x"00",
         14434 => x"00",
         14435 => x"00",
         14436 => x"00",
         14437 => x"00",
         14438 => x"00",
         14439 => x"00",
         14440 => x"00",
         14441 => x"00",
         14442 => x"00",
         14443 => x"00",
         14444 => x"00",
         14445 => x"00",
         14446 => x"00",
         14447 => x"00",
         14448 => x"00",
         14449 => x"00",
         14450 => x"00",
         14451 => x"00",
         14452 => x"00",
         14453 => x"00",
         14454 => x"00",
         14455 => x"00",
         14456 => x"00",
         14457 => x"00",
         14458 => x"00",
         14459 => x"00",
         14460 => x"00",
         14461 => x"00",
         14462 => x"00",
         14463 => x"00",
         14464 => x"00",
         14465 => x"00",
         14466 => x"00",
         14467 => x"00",
         14468 => x"00",
         14469 => x"00",
         14470 => x"00",
         14471 => x"00",
         14472 => x"00",
         14473 => x"00",
         14474 => x"00",
         14475 => x"00",
         14476 => x"00",
         14477 => x"00",
         14478 => x"00",
         14479 => x"00",
         14480 => x"00",
         14481 => x"00",
         14482 => x"00",
         14483 => x"00",
         14484 => x"00",
         14485 => x"00",
         14486 => x"00",
         14487 => x"00",
         14488 => x"00",
         14489 => x"00",
         14490 => x"00",
         14491 => x"00",
         14492 => x"00",
         14493 => x"00",
         14494 => x"00",
         14495 => x"00",
         14496 => x"00",
         14497 => x"00",
         14498 => x"00",
         14499 => x"00",
         14500 => x"00",
         14501 => x"00",
         14502 => x"00",
         14503 => x"00",
         14504 => x"00",
         14505 => x"00",
         14506 => x"00",
         14507 => x"00",
         14508 => x"00",
         14509 => x"00",
         14510 => x"00",
         14511 => x"00",
         14512 => x"00",
         14513 => x"00",
         14514 => x"00",
         14515 => x"00",
         14516 => x"00",
         14517 => x"00",
         14518 => x"00",
         14519 => x"00",
         14520 => x"00",
         14521 => x"00",
         14522 => x"00",
         14523 => x"00",
         14524 => x"00",
         14525 => x"00",
         14526 => x"00",
         14527 => x"00",
         14528 => x"00",
         14529 => x"00",
         14530 => x"00",
         14531 => x"00",
         14532 => x"00",
         14533 => x"00",
         14534 => x"00",
         14535 => x"00",
         14536 => x"00",
         14537 => x"00",
         14538 => x"00",
         14539 => x"00",
         14540 => x"00",
         14541 => x"00",
         14542 => x"00",
         14543 => x"00",
         14544 => x"00",
         14545 => x"00",
         14546 => x"00",
         14547 => x"00",
         14548 => x"00",
         14549 => x"00",
         14550 => x"00",
         14551 => x"00",
         14552 => x"00",
         14553 => x"00",
         14554 => x"00",
         14555 => x"00",
         14556 => x"00",
         14557 => x"00",
         14558 => x"00",
         14559 => x"00",
         14560 => x"00",
         14561 => x"00",
         14562 => x"00",
         14563 => x"00",
         14564 => x"00",
         14565 => x"00",
         14566 => x"00",
         14567 => x"00",
         14568 => x"00",
         14569 => x"00",
         14570 => x"00",
         14571 => x"00",
         14572 => x"00",
         14573 => x"00",
         14574 => x"00",
         14575 => x"00",
         14576 => x"00",
         14577 => x"00",
         14578 => x"00",
         14579 => x"00",
         14580 => x"00",
         14581 => x"00",
         14582 => x"00",
         14583 => x"00",
         14584 => x"00",
         14585 => x"00",
         14586 => x"00",
         14587 => x"00",
         14588 => x"00",
         14589 => x"00",
         14590 => x"00",
         14591 => x"00",
         14592 => x"00",
         14593 => x"00",
         14594 => x"00",
         14595 => x"00",
         14596 => x"00",
         14597 => x"00",
         14598 => x"00",
         14599 => x"00",
         14600 => x"00",
         14601 => x"00",
         14602 => x"00",
         14603 => x"00",
         14604 => x"00",
         14605 => x"00",
         14606 => x"00",
         14607 => x"00",
         14608 => x"00",
         14609 => x"00",
         14610 => x"00",
         14611 => x"00",
         14612 => x"00",
         14613 => x"00",
         14614 => x"00",
         14615 => x"00",
         14616 => x"00",
         14617 => x"00",
         14618 => x"00",
         14619 => x"00",
         14620 => x"00",
         14621 => x"00",
         14622 => x"00",
         14623 => x"00",
         14624 => x"00",
         14625 => x"00",
         14626 => x"00",
         14627 => x"00",
         14628 => x"00",
         14629 => x"00",
         14630 => x"00",
         14631 => x"00",
         14632 => x"00",
         14633 => x"00",
         14634 => x"00",
         14635 => x"00",
         14636 => x"00",
         14637 => x"00",
         14638 => x"00",
         14639 => x"00",
         14640 => x"00",
         14641 => x"00",
         14642 => x"00",
         14643 => x"00",
         14644 => x"00",
         14645 => x"00",
         14646 => x"00",
         14647 => x"00",
         14648 => x"00",
         14649 => x"00",
         14650 => x"00",
         14651 => x"00",
         14652 => x"00",
         14653 => x"00",
         14654 => x"00",
         14655 => x"00",
         14656 => x"00",
         14657 => x"00",
         14658 => x"00",
         14659 => x"00",
         14660 => x"00",
         14661 => x"00",
         14662 => x"00",
         14663 => x"00",
         14664 => x"00",
         14665 => x"00",
         14666 => x"00",
         14667 => x"00",
         14668 => x"00",
         14669 => x"00",
         14670 => x"00",
         14671 => x"00",
         14672 => x"00",
         14673 => x"00",
         14674 => x"00",
         14675 => x"00",
         14676 => x"00",
         14677 => x"00",
         14678 => x"00",
         14679 => x"00",
         14680 => x"00",
         14681 => x"00",
         14682 => x"00",
         14683 => x"00",
         14684 => x"00",
         14685 => x"00",
         14686 => x"00",
         14687 => x"00",
         14688 => x"00",
         14689 => x"00",
         14690 => x"00",
         14691 => x"00",
         14692 => x"00",
         14693 => x"00",
         14694 => x"00",
         14695 => x"00",
         14696 => x"00",
         14697 => x"00",
         14698 => x"00",
         14699 => x"00",
         14700 => x"00",
         14701 => x"00",
         14702 => x"00",
         14703 => x"00",
         14704 => x"00",
         14705 => x"00",
         14706 => x"00",
         14707 => x"00",
         14708 => x"00",
         14709 => x"00",
         14710 => x"00",
         14711 => x"00",
         14712 => x"00",
         14713 => x"00",
         14714 => x"00",
         14715 => x"00",
         14716 => x"00",
         14717 => x"00",
         14718 => x"00",
         14719 => x"00",
         14720 => x"00",
         14721 => x"00",
         14722 => x"00",
         14723 => x"00",
         14724 => x"00",
         14725 => x"00",
         14726 => x"00",
         14727 => x"00",
         14728 => x"00",
         14729 => x"00",
         14730 => x"00",
         14731 => x"00",
         14732 => x"00",
         14733 => x"00",
         14734 => x"00",
         14735 => x"00",
         14736 => x"00",
         14737 => x"00",
         14738 => x"00",
         14739 => x"00",
         14740 => x"00",
         14741 => x"00",
         14742 => x"00",
         14743 => x"00",
         14744 => x"00",
         14745 => x"00",
         14746 => x"00",
         14747 => x"00",
         14748 => x"00",
         14749 => x"00",
         14750 => x"00",
         14751 => x"00",
         14752 => x"00",
         14753 => x"00",
         14754 => x"00",
         14755 => x"00",
         14756 => x"00",
         14757 => x"00",
         14758 => x"00",
         14759 => x"00",
         14760 => x"00",
         14761 => x"00",
         14762 => x"00",
         14763 => x"00",
         14764 => x"64",
         14765 => x"74",
         14766 => x"64",
         14767 => x"74",
         14768 => x"66",
         14769 => x"74",
         14770 => x"66",
         14771 => x"64",
         14772 => x"66",
         14773 => x"63",
         14774 => x"6d",
         14775 => x"61",
         14776 => x"6d",
         14777 => x"79",
         14778 => x"6d",
         14779 => x"66",
         14780 => x"6d",
         14781 => x"70",
         14782 => x"6d",
         14783 => x"6d",
         14784 => x"6d",
         14785 => x"68",
         14786 => x"68",
         14787 => x"68",
         14788 => x"68",
         14789 => x"63",
         14790 => x"00",
         14791 => x"6a",
         14792 => x"72",
         14793 => x"61",
         14794 => x"72",
         14795 => x"74",
         14796 => x"69",
         14797 => x"00",
         14798 => x"74",
         14799 => x"00",
         14800 => x"63",
         14801 => x"7a",
         14802 => x"74",
         14803 => x"69",
         14804 => x"6d",
         14805 => x"69",
         14806 => x"6b",
         14807 => x"00",
         14808 => x"65",
         14809 => x"55",
         14810 => x"6f",
         14811 => x"65",
         14812 => x"72",
         14813 => x"50",
         14814 => x"6d",
         14815 => x"72",
         14816 => x"6e",
         14817 => x"72",
         14818 => x"2e",
         14819 => x"54",
         14820 => x"6d",
         14821 => x"20",
         14822 => x"6e",
         14823 => x"6c",
         14824 => x"00",
         14825 => x"49",
         14826 => x"66",
         14827 => x"69",
         14828 => x"20",
         14829 => x"6f",
         14830 => x"00",
         14831 => x"46",
         14832 => x"20",
         14833 => x"6c",
         14834 => x"65",
         14835 => x"54",
         14836 => x"6f",
         14837 => x"20",
         14838 => x"72",
         14839 => x"6f",
         14840 => x"61",
         14841 => x"6c",
         14842 => x"2e",
         14843 => x"46",
         14844 => x"61",
         14845 => x"62",
         14846 => x"65",
         14847 => x"4e",
         14848 => x"6f",
         14849 => x"74",
         14850 => x"65",
         14851 => x"6c",
         14852 => x"73",
         14853 => x"20",
         14854 => x"6e",
         14855 => x"6e",
         14856 => x"73",
         14857 => x"44",
         14858 => x"20",
         14859 => x"20",
         14860 => x"62",
         14861 => x"2e",
         14862 => x"44",
         14863 => x"65",
         14864 => x"6d",
         14865 => x"20",
         14866 => x"69",
         14867 => x"6c",
         14868 => x"00",
         14869 => x"53",
         14870 => x"73",
         14871 => x"69",
         14872 => x"70",
         14873 => x"65",
         14874 => x"64",
         14875 => x"46",
         14876 => x"20",
         14877 => x"64",
         14878 => x"69",
         14879 => x"6c",
         14880 => x"00",
         14881 => x"46",
         14882 => x"20",
         14883 => x"65",
         14884 => x"20",
         14885 => x"73",
         14886 => x"00",
         14887 => x"41",
         14888 => x"73",
         14889 => x"65",
         14890 => x"64",
         14891 => x"49",
         14892 => x"6c",
         14893 => x"66",
         14894 => x"6e",
         14895 => x"2e",
         14896 => x"4e",
         14897 => x"61",
         14898 => x"66",
         14899 => x"64",
         14900 => x"4e",
         14901 => x"69",
         14902 => x"66",
         14903 => x"64",
         14904 => x"44",
         14905 => x"20",
         14906 => x"20",
         14907 => x"64",
         14908 => x"49",
         14909 => x"72",
         14910 => x"20",
         14911 => x"6f",
         14912 => x"44",
         14913 => x"20",
         14914 => x"6f",
         14915 => x"53",
         14916 => x"65",
         14917 => x"00",
         14918 => x"0a",
         14919 => x"20",
         14920 => x"65",
         14921 => x"73",
         14922 => x"20",
         14923 => x"20",
         14924 => x"65",
         14925 => x"65",
         14926 => x"00",
         14927 => x"72",
         14928 => x"00",
         14929 => x"25",
         14930 => x"58",
         14931 => x"3a",
         14932 => x"25",
         14933 => x"00",
         14934 => x"20",
         14935 => x"7c",
         14936 => x"20",
         14937 => x"25",
         14938 => x"00",
         14939 => x"20",
         14940 => x"20",
         14941 => x"00",
         14942 => x"7a",
         14943 => x"2a",
         14944 => x"73",
         14945 => x"31",
         14946 => x"32",
         14947 => x"32",
         14948 => x"76",
         14949 => x"64",
         14950 => x"20",
         14951 => x"2c",
         14952 => x"76",
         14953 => x"32",
         14954 => x"25",
         14955 => x"73",
         14956 => x"0a",
         14957 => x"5a",
         14958 => x"49",
         14959 => x"72",
         14960 => x"74",
         14961 => x"6e",
         14962 => x"72",
         14963 => x"55",
         14964 => x"31",
         14965 => x"20",
         14966 => x"65",
         14967 => x"70",
         14968 => x"55",
         14969 => x"31",
         14970 => x"20",
         14971 => x"65",
         14972 => x"70",
         14973 => x"55",
         14974 => x"30",
         14975 => x"20",
         14976 => x"65",
         14977 => x"70",
         14978 => x"55",
         14979 => x"30",
         14980 => x"20",
         14981 => x"65",
         14982 => x"70",
         14983 => x"49",
         14984 => x"4c",
         14985 => x"20",
         14986 => x"65",
         14987 => x"70",
         14988 => x"49",
         14989 => x"4c",
         14990 => x"20",
         14991 => x"65",
         14992 => x"70",
         14993 => x"50",
         14994 => x"69",
         14995 => x"72",
         14996 => x"74",
         14997 => x"54",
         14998 => x"72",
         14999 => x"74",
         15000 => x"75",
         15001 => x"53",
         15002 => x"69",
         15003 => x"75",
         15004 => x"69",
         15005 => x"2e",
         15006 => x"45",
         15007 => x"6c",
         15008 => x"20",
         15009 => x"65",
         15010 => x"2e",
         15011 => x"61",
         15012 => x"65",
         15013 => x"2e",
         15014 => x"00",
         15015 => x"7a",
         15016 => x"7a",
         15017 => x"68",
         15018 => x"46",
         15019 => x"65",
         15020 => x"6f",
         15021 => x"69",
         15022 => x"6c",
         15023 => x"20",
         15024 => x"63",
         15025 => x"20",
         15026 => x"70",
         15027 => x"73",
         15028 => x"6e",
         15029 => x"6d",
         15030 => x"61",
         15031 => x"2e",
         15032 => x"2a",
         15033 => x"25",
         15034 => x"25",
         15035 => x"44",
         15036 => x"20",
         15037 => x"74",
         15038 => x"69",
         15039 => x"00",
         15040 => x"30",
         15041 => x"42",
         15042 => x"63",
         15043 => x"61",
         15044 => x"00",
         15045 => x"5a",
         15046 => x"62",
         15047 => x"25",
         15048 => x"25",
         15049 => x"73",
         15050 => x"00",
         15051 => x"43",
         15052 => x"20",
         15053 => x"6f",
         15054 => x"6e",
         15055 => x"2e",
         15056 => x"52",
         15057 => x"61",
         15058 => x"6e",
         15059 => x"70",
         15060 => x"63",
         15061 => x"6f",
         15062 => x"2e",
         15063 => x"43",
         15064 => x"69",
         15065 => x"63",
         15066 => x"20",
         15067 => x"30",
         15068 => x"20",
         15069 => x"0a",
         15070 => x"43",
         15071 => x"20",
         15072 => x"75",
         15073 => x"64",
         15074 => x"64",
         15075 => x"25",
         15076 => x"0a",
         15077 => x"45",
         15078 => x"75",
         15079 => x"67",
         15080 => x"64",
         15081 => x"20",
         15082 => x"6c",
         15083 => x"2e",
         15084 => x"25",
         15085 => x"58",
         15086 => x"38",
         15087 => x"00",
         15088 => x"25",
         15089 => x"58",
         15090 => x"34",
         15091 => x"43",
         15092 => x"61",
         15093 => x"67",
         15094 => x"00",
         15095 => x"25",
         15096 => x"78",
         15097 => x"38",
         15098 => x"3e",
         15099 => x"6c",
         15100 => x"30",
         15101 => x"0a",
         15102 => x"43",
         15103 => x"69",
         15104 => x"2e",
         15105 => x"25",
         15106 => x"58",
         15107 => x"32",
         15108 => x"43",
         15109 => x"72",
         15110 => x"2e",
         15111 => x"00",
         15112 => x"44",
         15113 => x"20",
         15114 => x"6f",
         15115 => x"0a",
         15116 => x"70",
         15117 => x"65",
         15118 => x"25",
         15119 => x"25",
         15120 => x"73",
         15121 => x"4d",
         15122 => x"72",
         15123 => x"78",
         15124 => x"73",
         15125 => x"2c",
         15126 => x"6e",
         15127 => x"20",
         15128 => x"63",
         15129 => x"20",
         15130 => x"6d",
         15131 => x"2e",
         15132 => x"3f",
         15133 => x"25",
         15134 => x"64",
         15135 => x"20",
         15136 => x"25",
         15137 => x"64",
         15138 => x"25",
         15139 => x"53",
         15140 => x"43",
         15141 => x"69",
         15142 => x"61",
         15143 => x"6e",
         15144 => x"3a",
         15145 => x"76",
         15146 => x"73",
         15147 => x"70",
         15148 => x"65",
         15149 => x"64",
         15150 => x"41",
         15151 => x"65",
         15152 => x"73",
         15153 => x"20",
         15154 => x"43",
         15155 => x"52",
         15156 => x"74",
         15157 => x"63",
         15158 => x"20",
         15159 => x"72",
         15160 => x"20",
         15161 => x"30",
         15162 => x"00",
         15163 => x"20",
         15164 => x"43",
         15165 => x"4d",
         15166 => x"72",
         15167 => x"74",
         15168 => x"20",
         15169 => x"72",
         15170 => x"20",
         15171 => x"30",
         15172 => x"00",
         15173 => x"20",
         15174 => x"53",
         15175 => x"6b",
         15176 => x"61",
         15177 => x"41",
         15178 => x"65",
         15179 => x"20",
         15180 => x"20",
         15181 => x"30",
         15182 => x"00",
         15183 => x"4d",
         15184 => x"3a",
         15185 => x"20",
         15186 => x"5a",
         15187 => x"49",
         15188 => x"20",
         15189 => x"20",
         15190 => x"20",
         15191 => x"20",
         15192 => x"20",
         15193 => x"30",
         15194 => x"00",
         15195 => x"20",
         15196 => x"53",
         15197 => x"65",
         15198 => x"6c",
         15199 => x"20",
         15200 => x"71",
         15201 => x"20",
         15202 => x"20",
         15203 => x"64",
         15204 => x"34",
         15205 => x"7a",
         15206 => x"20",
         15207 => x"57",
         15208 => x"62",
         15209 => x"20",
         15210 => x"41",
         15211 => x"6c",
         15212 => x"20",
         15213 => x"71",
         15214 => x"64",
         15215 => x"34",
         15216 => x"7a",
         15217 => x"20",
         15218 => x"53",
         15219 => x"4d",
         15220 => x"6f",
         15221 => x"46",
         15222 => x"20",
         15223 => x"20",
         15224 => x"20",
         15225 => x"64",
         15226 => x"34",
         15227 => x"7a",
         15228 => x"20",
         15229 => x"53",
         15230 => x"20",
         15231 => x"50",
         15232 => x"20",
         15233 => x"49",
         15234 => x"4c",
         15235 => x"20",
         15236 => x"57",
         15237 => x"32",
         15238 => x"20",
         15239 => x"57",
         15240 => x"42",
         15241 => x"20",
         15242 => x"00",
         15243 => x"20",
         15244 => x"49",
         15245 => x"20",
         15246 => x"4c",
         15247 => x"68",
         15248 => x"65",
         15249 => x"25",
         15250 => x"29",
         15251 => x"20",
         15252 => x"54",
         15253 => x"52",
         15254 => x"20",
         15255 => x"69",
         15256 => x"73",
         15257 => x"25",
         15258 => x"29",
         15259 => x"20",
         15260 => x"53",
         15261 => x"41",
         15262 => x"20",
         15263 => x"65",
         15264 => x"65",
         15265 => x"25",
         15266 => x"29",
         15267 => x"20",
         15268 => x"52",
         15269 => x"20",
         15270 => x"20",
         15271 => x"30",
         15272 => x"25",
         15273 => x"29",
         15274 => x"20",
         15275 => x"42",
         15276 => x"20",
         15277 => x"20",
         15278 => x"30",
         15279 => x"25",
         15280 => x"29",
         15281 => x"20",
         15282 => x"49",
         15283 => x"20",
         15284 => x"4d",
         15285 => x"30",
         15286 => x"25",
         15287 => x"29",
         15288 => x"20",
         15289 => x"53",
         15290 => x"4d",
         15291 => x"20",
         15292 => x"30",
         15293 => x"25",
         15294 => x"29",
         15295 => x"20",
         15296 => x"57",
         15297 => x"44",
         15298 => x"20",
         15299 => x"30",
         15300 => x"25",
         15301 => x"29",
         15302 => x"20",
         15303 => x"6f",
         15304 => x"6f",
         15305 => x"6f",
         15306 => x"67",
         15307 => x"55",
         15308 => x"6f",
         15309 => x"45",
         15310 => x"00",
         15311 => x"53",
         15312 => x"6c",
         15313 => x"4d",
         15314 => x"75",
         15315 => x"46",
         15316 => x"00",
         15317 => x"45",
         15318 => x"00",
         15319 => x"01",
         15320 => x"00",
         15321 => x"00",
         15322 => x"01",
         15323 => x"00",
         15324 => x"00",
         15325 => x"01",
         15326 => x"00",
         15327 => x"00",
         15328 => x"01",
         15329 => x"00",
         15330 => x"00",
         15331 => x"01",
         15332 => x"00",
         15333 => x"00",
         15334 => x"01",
         15335 => x"00",
         15336 => x"00",
         15337 => x"01",
         15338 => x"00",
         15339 => x"00",
         15340 => x"01",
         15341 => x"00",
         15342 => x"00",
         15343 => x"01",
         15344 => x"00",
         15345 => x"00",
         15346 => x"01",
         15347 => x"00",
         15348 => x"00",
         15349 => x"01",
         15350 => x"00",
         15351 => x"00",
         15352 => x"04",
         15353 => x"00",
         15354 => x"00",
         15355 => x"04",
         15356 => x"00",
         15357 => x"00",
         15358 => x"04",
         15359 => x"00",
         15360 => x"00",
         15361 => x"03",
         15362 => x"00",
         15363 => x"00",
         15364 => x"04",
         15365 => x"00",
         15366 => x"00",
         15367 => x"04",
         15368 => x"00",
         15369 => x"00",
         15370 => x"04",
         15371 => x"00",
         15372 => x"00",
         15373 => x"03",
         15374 => x"00",
         15375 => x"00",
         15376 => x"03",
         15377 => x"00",
         15378 => x"00",
         15379 => x"03",
         15380 => x"00",
         15381 => x"00",
         15382 => x"03",
         15383 => x"00",
         15384 => x"1b",
         15385 => x"1b",
         15386 => x"1b",
         15387 => x"1b",
         15388 => x"1b",
         15389 => x"1b",
         15390 => x"1b",
         15391 => x"1b",
         15392 => x"1b",
         15393 => x"1b",
         15394 => x"1b",
         15395 => x"10",
         15396 => x"0e",
         15397 => x"0d",
         15398 => x"0b",
         15399 => x"08",
         15400 => x"06",
         15401 => x"05",
         15402 => x"04",
         15403 => x"03",
         15404 => x"02",
         15405 => x"01",
         15406 => x"43",
         15407 => x"6f",
         15408 => x"70",
         15409 => x"63",
         15410 => x"74",
         15411 => x"69",
         15412 => x"72",
         15413 => x"69",
         15414 => x"20",
         15415 => x"61",
         15416 => x"6e",
         15417 => x"68",
         15418 => x"6f",
         15419 => x"68",
         15420 => x"00",
         15421 => x"21",
         15422 => x"25",
         15423 => x"75",
         15424 => x"73",
         15425 => x"46",
         15426 => x"65",
         15427 => x"6f",
         15428 => x"73",
         15429 => x"74",
         15430 => x"68",
         15431 => x"6f",
         15432 => x"66",
         15433 => x"20",
         15434 => x"45",
         15435 => x"00",
         15436 => x"3e",
         15437 => x"00",
         15438 => x"1b",
         15439 => x"00",
         15440 => x"1b",
         15441 => x"1b",
         15442 => x"1b",
         15443 => x"1b",
         15444 => x"1b",
         15445 => x"7e",
         15446 => x"1b",
         15447 => x"7e",
         15448 => x"1b",
         15449 => x"7e",
         15450 => x"1b",
         15451 => x"7e",
         15452 => x"1b",
         15453 => x"7e",
         15454 => x"1b",
         15455 => x"7e",
         15456 => x"1b",
         15457 => x"7e",
         15458 => x"1b",
         15459 => x"7e",
         15460 => x"1b",
         15461 => x"7e",
         15462 => x"1b",
         15463 => x"7e",
         15464 => x"1b",
         15465 => x"00",
         15466 => x"1b",
         15467 => x"00",
         15468 => x"1b",
         15469 => x"1b",
         15470 => x"00",
         15471 => x"1b",
         15472 => x"00",
         15473 => x"58",
         15474 => x"2c",
         15475 => x"25",
         15476 => x"64",
         15477 => x"2c",
         15478 => x"25",
         15479 => x"00",
         15480 => x"44",
         15481 => x"2d",
         15482 => x"25",
         15483 => x"63",
         15484 => x"2c",
         15485 => x"25",
         15486 => x"25",
         15487 => x"4b",
         15488 => x"3a",
         15489 => x"25",
         15490 => x"2c",
         15491 => x"25",
         15492 => x"64",
         15493 => x"52",
         15494 => x"52",
         15495 => x"72",
         15496 => x"75",
         15497 => x"72",
         15498 => x"55",
         15499 => x"30",
         15500 => x"25",
         15501 => x"00",
         15502 => x"44",
         15503 => x"30",
         15504 => x"25",
         15505 => x"00",
         15506 => x"48",
         15507 => x"30",
         15508 => x"00",
         15509 => x"42",
         15510 => x"65",
         15511 => x"2c",
         15512 => x"20",
         15513 => x"74",
         15514 => x"42",
         15515 => x"65",
         15516 => x"2c",
         15517 => x"20",
         15518 => x"64",
         15519 => x"42",
         15520 => x"65",
         15521 => x"2c",
         15522 => x"20",
         15523 => x"74",
         15524 => x"4e",
         15525 => x"65",
         15526 => x"64",
         15527 => x"6e",
         15528 => x"00",
         15529 => x"53",
         15530 => x"22",
         15531 => x"3e",
         15532 => x"00",
         15533 => x"2b",
         15534 => x"5b",
         15535 => x"46",
         15536 => x"46",
         15537 => x"32",
         15538 => x"eb",
         15539 => x"53",
         15540 => x"35",
         15541 => x"4e",
         15542 => x"41",
         15543 => x"20",
         15544 => x"41",
         15545 => x"20",
         15546 => x"4e",
         15547 => x"41",
         15548 => x"20",
         15549 => x"41",
         15550 => x"20",
         15551 => x"00",
         15552 => x"00",
         15553 => x"00",
         15554 => x"00",
         15555 => x"01",
         15556 => x"09",
         15557 => x"14",
         15558 => x"1e",
         15559 => x"80",
         15560 => x"8e",
         15561 => x"45",
         15562 => x"49",
         15563 => x"90",
         15564 => x"99",
         15565 => x"59",
         15566 => x"9c",
         15567 => x"41",
         15568 => x"a5",
         15569 => x"a8",
         15570 => x"ac",
         15571 => x"b0",
         15572 => x"b4",
         15573 => x"b8",
         15574 => x"bc",
         15575 => x"c0",
         15576 => x"c4",
         15577 => x"c8",
         15578 => x"cc",
         15579 => x"d0",
         15580 => x"d4",
         15581 => x"d8",
         15582 => x"dc",
         15583 => x"e0",
         15584 => x"e4",
         15585 => x"e8",
         15586 => x"ec",
         15587 => x"f0",
         15588 => x"f4",
         15589 => x"f8",
         15590 => x"fc",
         15591 => x"2b",
         15592 => x"3d",
         15593 => x"5c",
         15594 => x"3c",
         15595 => x"7f",
         15596 => x"00",
         15597 => x"00",
         15598 => x"01",
         15599 => x"00",
         15600 => x"00",
         15601 => x"00",
         15602 => x"00",
         15603 => x"00",
         15604 => x"00",
         15605 => x"00",
         15606 => x"00",
         15607 => x"00",
         15608 => x"00",
         15609 => x"00",
         15610 => x"00",
         15611 => x"00",
         15612 => x"00",
         15613 => x"00",
         15614 => x"00",
         15615 => x"00",
         15616 => x"00",
         15617 => x"00",
         15618 => x"00",
         15619 => x"20",
         15620 => x"00",
         15621 => x"00",
         15622 => x"00",
         15623 => x"00",
         15624 => x"00",
         15625 => x"00",
         15626 => x"00",
         15627 => x"00",
         15628 => x"25",
         15629 => x"25",
         15630 => x"25",
         15631 => x"25",
         15632 => x"25",
         15633 => x"25",
         15634 => x"25",
         15635 => x"25",
         15636 => x"25",
         15637 => x"25",
         15638 => x"25",
         15639 => x"25",
         15640 => x"25",
         15641 => x"25",
         15642 => x"25",
         15643 => x"25",
         15644 => x"25",
         15645 => x"25",
         15646 => x"25",
         15647 => x"25",
         15648 => x"25",
         15649 => x"25",
         15650 => x"25",
         15651 => x"25",
         15652 => x"03",
         15653 => x"03",
         15654 => x"03",
         15655 => x"00",
         15656 => x"03",
         15657 => x"03",
         15658 => x"22",
         15659 => x"03",
         15660 => x"22",
         15661 => x"22",
         15662 => x"23",
         15663 => x"00",
         15664 => x"00",
         15665 => x"00",
         15666 => x"20",
         15667 => x"25",
         15668 => x"00",
         15669 => x"00",
         15670 => x"00",
         15671 => x"00",
         15672 => x"01",
         15673 => x"01",
         15674 => x"01",
         15675 => x"01",
         15676 => x"01",
         15677 => x"01",
         15678 => x"00",
         15679 => x"01",
         15680 => x"01",
         15681 => x"01",
         15682 => x"01",
         15683 => x"01",
         15684 => x"01",
         15685 => x"01",
         15686 => x"01",
         15687 => x"01",
         15688 => x"01",
         15689 => x"01",
         15690 => x"01",
         15691 => x"01",
         15692 => x"01",
         15693 => x"01",
         15694 => x"01",
         15695 => x"01",
         15696 => x"01",
         15697 => x"01",
         15698 => x"01",
         15699 => x"01",
         15700 => x"01",
         15701 => x"01",
         15702 => x"01",
         15703 => x"01",
         15704 => x"01",
         15705 => x"01",
         15706 => x"01",
         15707 => x"01",
         15708 => x"01",
         15709 => x"01",
         15710 => x"01",
         15711 => x"01",
         15712 => x"01",
         15713 => x"01",
         15714 => x"01",
         15715 => x"01",
         15716 => x"01",
         15717 => x"01",
         15718 => x"01",
         15719 => x"01",
         15720 => x"01",
         15721 => x"00",
         15722 => x"01",
         15723 => x"01",
         15724 => x"02",
         15725 => x"02",
         15726 => x"2c",
         15727 => x"02",
         15728 => x"2c",
         15729 => x"02",
         15730 => x"02",
         15731 => x"01",
         15732 => x"00",
         15733 => x"01",
         15734 => x"01",
         15735 => x"02",
         15736 => x"02",
         15737 => x"02",
         15738 => x"02",
         15739 => x"01",
         15740 => x"02",
         15741 => x"02",
         15742 => x"02",
         15743 => x"01",
         15744 => x"02",
         15745 => x"02",
         15746 => x"02",
         15747 => x"02",
         15748 => x"01",
         15749 => x"02",
         15750 => x"02",
         15751 => x"02",
         15752 => x"02",
         15753 => x"02",
         15754 => x"02",
         15755 => x"01",
         15756 => x"02",
         15757 => x"02",
         15758 => x"02",
         15759 => x"01",
         15760 => x"01",
         15761 => x"02",
         15762 => x"02",
         15763 => x"02",
         15764 => x"01",
         15765 => x"00",
         15766 => x"03",
         15767 => x"03",
         15768 => x"03",
         15769 => x"03",
         15770 => x"03",
         15771 => x"03",
         15772 => x"03",
         15773 => x"03",
         15774 => x"03",
         15775 => x"03",
         15776 => x"03",
         15777 => x"01",
         15778 => x"00",
         15779 => x"03",
         15780 => x"03",
         15781 => x"03",
         15782 => x"03",
         15783 => x"03",
         15784 => x"03",
         15785 => x"07",
         15786 => x"01",
         15787 => x"01",
         15788 => x"01",
         15789 => x"00",
         15790 => x"04",
         15791 => x"05",
         15792 => x"00",
         15793 => x"1d",
         15794 => x"2c",
         15795 => x"01",
         15796 => x"01",
         15797 => x"06",
         15798 => x"06",
         15799 => x"06",
         15800 => x"06",
         15801 => x"06",
         15802 => x"00",
         15803 => x"1f",
         15804 => x"1f",
         15805 => x"1f",
         15806 => x"1f",
         15807 => x"1f",
         15808 => x"1f",
         15809 => x"1f",
         15810 => x"1f",
         15811 => x"1f",
         15812 => x"1f",
         15813 => x"1f",
         15814 => x"1f",
         15815 => x"1f",
         15816 => x"1f",
         15817 => x"1f",
         15818 => x"1f",
         15819 => x"1f",
         15820 => x"1f",
         15821 => x"1f",
         15822 => x"1f",
         15823 => x"06",
         15824 => x"06",
         15825 => x"00",
         15826 => x"1f",
         15827 => x"1f",
         15828 => x"00",
         15829 => x"21",
         15830 => x"21",
         15831 => x"21",
         15832 => x"05",
         15833 => x"04",
         15834 => x"01",
         15835 => x"01",
         15836 => x"01",
         15837 => x"01",
         15838 => x"08",
         15839 => x"03",
         15840 => x"00",
         15841 => x"00",
         15842 => x"01",
         15843 => x"00",
         15844 => x"00",
         15845 => x"00",
         15846 => x"01",
         15847 => x"00",
         15848 => x"00",
         15849 => x"00",
         15850 => x"01",
         15851 => x"00",
         15852 => x"00",
         15853 => x"00",
         15854 => x"01",
         15855 => x"00",
         15856 => x"00",
         15857 => x"00",
         15858 => x"01",
         15859 => x"00",
         15860 => x"00",
         15861 => x"00",
         15862 => x"01",
         15863 => x"00",
         15864 => x"00",
         15865 => x"00",
         15866 => x"01",
         15867 => x"00",
         15868 => x"00",
         15869 => x"00",
         15870 => x"01",
         15871 => x"00",
         15872 => x"00",
         15873 => x"00",
         15874 => x"01",
         15875 => x"00",
         15876 => x"00",
         15877 => x"00",
         15878 => x"01",
         15879 => x"00",
         15880 => x"00",
         15881 => x"00",
         15882 => x"01",
         15883 => x"00",
         15884 => x"00",
         15885 => x"00",
         15886 => x"01",
         15887 => x"00",
         15888 => x"00",
         15889 => x"00",
         15890 => x"01",
         15891 => x"00",
         15892 => x"00",
         15893 => x"00",
         15894 => x"01",
         15895 => x"00",
         15896 => x"00",
         15897 => x"00",
         15898 => x"01",
         15899 => x"00",
         15900 => x"00",
         15901 => x"00",
         15902 => x"01",
         15903 => x"00",
         15904 => x"00",
         15905 => x"00",
         15906 => x"01",
         15907 => x"00",
         15908 => x"00",
         15909 => x"00",
         15910 => x"01",
         15911 => x"00",
         15912 => x"00",
         15913 => x"00",
         15914 => x"01",
         15915 => x"00",
         15916 => x"00",
         15917 => x"00",
         15918 => x"01",
         15919 => x"00",
         15920 => x"00",
         15921 => x"00",
         15922 => x"01",
         15923 => x"00",
         15924 => x"00",
         15925 => x"00",
         15926 => x"01",
         15927 => x"00",
         15928 => x"00",
         15929 => x"00",
         15930 => x"01",
         15931 => x"00",
         15932 => x"00",
         15933 => x"00",
         15934 => x"01",
         15935 => x"00",
         15936 => x"00",
         15937 => x"00",
         15938 => x"01",
         15939 => x"00",
         15940 => x"00",
         15941 => x"00",
         15942 => x"01",
         15943 => x"00",
         15944 => x"00",
         15945 => x"00",
         15946 => x"01",
         15947 => x"00",
         15948 => x"00",
         15949 => x"00",
         15950 => x"01",
         15951 => x"00",
         15952 => x"00",
         15953 => x"00",
         15954 => x"00",
         15955 => x"00",
         15956 => x"00",
         15957 => x"00",
         15958 => x"00",
         15959 => x"00",
         15960 => x"00",
         15961 => x"00",
         15962 => x"01",
         15963 => x"01",
         15964 => x"00",
         15965 => x"00",
         15966 => x"00",
         15967 => x"00",
         15968 => x"05",
         15969 => x"05",
         15970 => x"05",
         15971 => x"00",
         15972 => x"01",
         15973 => x"01",
         15974 => x"01",
         15975 => x"01",
         15976 => x"00",
         15977 => x"00",
         15978 => x"00",
         15979 => x"00",
         15980 => x"00",
         15981 => x"00",
         15982 => x"00",
         15983 => x"00",
         15984 => x"00",
         15985 => x"00",
         15986 => x"00",
         15987 => x"00",
         15988 => x"00",
         15989 => x"00",
         15990 => x"00",
         15991 => x"00",
         15992 => x"00",
         15993 => x"00",
         15994 => x"00",
         15995 => x"00",
         15996 => x"00",
         15997 => x"00",
         15998 => x"00",
         15999 => x"00",
         16000 => x"00",
         16001 => x"01",
         16002 => x"00",
         16003 => x"01",
         16004 => x"00",
         16005 => x"02",
         16006 => x"00",
         16007 => x"1b",
         16008 => x"f0",
         16009 => x"79",
         16010 => x"5d",
         16011 => x"71",
         16012 => x"75",
         16013 => x"69",
         16014 => x"6d",
         16015 => x"61",
         16016 => x"65",
         16017 => x"31",
         16018 => x"35",
         16019 => x"5c",
         16020 => x"30",
         16021 => x"f6",
         16022 => x"f1",
         16023 => x"08",
         16024 => x"f0",
         16025 => x"80",
         16026 => x"84",
         16027 => x"1b",
         16028 => x"f0",
         16029 => x"59",
         16030 => x"5d",
         16031 => x"51",
         16032 => x"55",
         16033 => x"49",
         16034 => x"4d",
         16035 => x"41",
         16036 => x"45",
         16037 => x"31",
         16038 => x"35",
         16039 => x"5c",
         16040 => x"30",
         16041 => x"f6",
         16042 => x"f1",
         16043 => x"08",
         16044 => x"f0",
         16045 => x"80",
         16046 => x"84",
         16047 => x"1b",
         16048 => x"f0",
         16049 => x"59",
         16050 => x"7d",
         16051 => x"51",
         16052 => x"55",
         16053 => x"49",
         16054 => x"4d",
         16055 => x"41",
         16056 => x"45",
         16057 => x"21",
         16058 => x"25",
         16059 => x"7c",
         16060 => x"20",
         16061 => x"f7",
         16062 => x"f9",
         16063 => x"fb",
         16064 => x"f0",
         16065 => x"85",
         16066 => x"89",
         16067 => x"1b",
         16068 => x"f0",
         16069 => x"19",
         16070 => x"1d",
         16071 => x"11",
         16072 => x"15",
         16073 => x"09",
         16074 => x"0d",
         16075 => x"01",
         16076 => x"05",
         16077 => x"f0",
         16078 => x"f0",
         16079 => x"f0",
         16080 => x"f0",
         16081 => x"f0",
         16082 => x"f0",
         16083 => x"f0",
         16084 => x"f0",
         16085 => x"80",
         16086 => x"84",
         16087 => x"bf",
         16088 => x"f0",
         16089 => x"35",
         16090 => x"b7",
         16091 => x"7c",
         16092 => x"39",
         16093 => x"3d",
         16094 => x"1d",
         16095 => x"46",
         16096 => x"74",
         16097 => x"3f",
         16098 => x"7a",
         16099 => x"d3",
         16100 => x"9d",
         16101 => x"c6",
         16102 => x"c3",
         16103 => x"f0",
         16104 => x"f0",
         16105 => x"80",
         16106 => x"84",
         16107 => x"00",
         16108 => x"00",
         16109 => x"00",
         16110 => x"00",
         16111 => x"00",
         16112 => x"00",
         16113 => x"00",
         16114 => x"00",
         16115 => x"00",
         16116 => x"00",
         16117 => x"00",
         16118 => x"00",
         16119 => x"00",
         16120 => x"00",
         16121 => x"00",
         16122 => x"00",
         16123 => x"00",
         16124 => x"00",
         16125 => x"00",
         16126 => x"00",
         16127 => x"00",
         16128 => x"00",
         16129 => x"00",
         16130 => x"00",
         16131 => x"00",
         16132 => x"00",
         16133 => x"00",
         16134 => x"f8",
         16135 => x"00",
         16136 => x"f3",
         16137 => x"00",
         16138 => x"f4",
         16139 => x"00",
         16140 => x"f1",
         16141 => x"00",
         16142 => x"f2",
         16143 => x"00",
         16144 => x"80",
         16145 => x"00",
         16146 => x"81",
         16147 => x"00",
         16148 => x"82",
         16149 => x"00",
         16150 => x"83",
         16151 => x"00",
         16152 => x"84",
         16153 => x"00",
         16154 => x"85",
         16155 => x"00",
         16156 => x"86",
         16157 => x"00",
         16158 => x"87",
         16159 => x"00",
         16160 => x"88",
         16161 => x"00",
         16162 => x"89",
         16163 => x"00",
         16164 => x"f6",
         16165 => x"00",
         16166 => x"7f",
         16167 => x"00",
         16168 => x"f9",
         16169 => x"00",
         16170 => x"e0",
         16171 => x"00",
         16172 => x"e1",
         16173 => x"00",
         16174 => x"71",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"00",
         18159 => x"00",
         18160 => x"00",
         18161 => x"00",
         18162 => x"00",
         18163 => x"00",
         18164 => x"00",
         18165 => x"00",
         18166 => x"00",
         18167 => x"00",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"00",
         18176 => x"50",
         18177 => x"00",
         18178 => x"cc",
         18179 => x"ce",
         18180 => x"f8",
         18181 => x"fc",
         18182 => x"e1",
         18183 => x"c4",
         18184 => x"e3",
         18185 => x"eb",
         18186 => x"00",
         18187 => x"64",
         18188 => x"68",
         18189 => x"2f",
         18190 => x"20",
         18191 => x"24",
         18192 => x"28",
         18193 => x"51",
         18194 => x"55",
         18195 => x"04",
         18196 => x"08",
         18197 => x"0c",
         18198 => x"10",
         18199 => x"14",
         18200 => x"18",
         18201 => x"59",
         18202 => x"c7",
         18203 => x"84",
         18204 => x"88",
         18205 => x"8c",
         18206 => x"90",
         18207 => x"94",
         18208 => x"98",
         18209 => x"80",
         18210 => x"00",
         18211 => x"00",
         18212 => x"00",
         18213 => x"00",
         18214 => x"00",
         18215 => x"00",
         18216 => x"00",
         18217 => x"00",
         18218 => x"00",
         18219 => x"00",
         18220 => x"00",
         18221 => x"00",
         18222 => x"00",
         18223 => x"00",
         18224 => x"00",
         18225 => x"00",
         18226 => x"00",
         18227 => x"00",
         18228 => x"00",
         18229 => x"00",
         18230 => x"00",
         18231 => x"00",
         18232 => x"00",
         18233 => x"00",
         18234 => x"00",
         18235 => x"00",
         18236 => x"00",
         18237 => x"00",
         18238 => x"00",
         18239 => x"00",
         18240 => x"00",
         18241 => x"00",
         18242 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
