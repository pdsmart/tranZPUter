SFL_IV_inst : SFL_IV PORT MAP (
		noe_in	 => noe_in_sig
	);
