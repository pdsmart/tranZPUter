-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"800b0b0b",
             2 => x"0b8eae04",
             3 => x"ffffffff",
             4 => x"ffffffff",
             5 => x"ffffffff",
             6 => x"ffffffff",
             7 => x"ffffffff",
             8 => x"0b0b0b88",
             9 => x"80040b0b",
            10 => x"0b888404",
            11 => x"0b0b0b88",
            12 => x"94040b0b",
            13 => x"0b88a404",
            14 => x"0b0b0b88",
            15 => x"b4040b0b",
            16 => x"0b88c404",
            17 => x"0b0b0b88",
            18 => x"d4040b0b",
            19 => x"0b88e404",
            20 => x"0b0b0b88",
            21 => x"f4040b0b",
            22 => x"0b898404",
            23 => x"0b0b0b89",
            24 => x"94040b0b",
            25 => x"0b89a404",
            26 => x"0b0b0b89",
            27 => x"b4040b0b",
            28 => x"0b89c404",
            29 => x"0b0b0b89",
            30 => x"d4040b0b",
            31 => x"0b89e404",
            32 => x"0b0b0b89",
            33 => x"f4040b0b",
            34 => x"0b8a8404",
            35 => x"0b0b0b8a",
            36 => x"94040b0b",
            37 => x"0b8aa504",
            38 => x"0b0b0b8a",
            39 => x"b6040b0b",
            40 => x"0b8ac704",
            41 => x"0b0b0b8a",
            42 => x"d8040b0b",
            43 => x"0b8ae904",
            44 => x"0b0b0b8a",
            45 => x"fa040b0b",
            46 => x"0b8b8b04",
            47 => x"0b0b0b8b",
            48 => x"9c040b0b",
            49 => x"0b8bad04",
            50 => x"0b0b0b8b",
            51 => x"be040b0b",
            52 => x"0b8bcf04",
            53 => x"0b0b0b8b",
            54 => x"e0040b0b",
            55 => x"0b8bf104",
            56 => x"0b0b0b8c",
            57 => x"82040b0b",
            58 => x"0b8c9304",
            59 => x"0b0b0b8c",
            60 => x"a4040b0b",
            61 => x"0b8cb504",
            62 => x"0b0b0b8c",
            63 => x"c6040b0b",
            64 => x"0b8cd704",
            65 => x"0b0b0b8c",
            66 => x"e8040b0b",
            67 => x"0b8cf904",
            68 => x"0b0b0b8d",
            69 => x"8a040b0b",
            70 => x"0b8d9b04",
            71 => x"0b0b0b8d",
            72 => x"ac040b0b",
            73 => x"0b8dbd04",
            74 => x"0b0b0b8d",
            75 => x"cd040b0b",
            76 => x"0b8ddd04",
            77 => x"0b0b0b8d",
            78 => x"ed040b0b",
            79 => x"0b8dfd04",
            80 => x"0b0b0b8e",
            81 => x"8d040b0b",
            82 => x"0b8e9d04",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"00000000",
            89 => x"00000000",
            90 => x"00000000",
            91 => x"00000000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"00000000",
            97 => x"00000000",
            98 => x"00000000",
            99 => x"00000000",
           100 => x"00000000",
           101 => x"00000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"00000000",
           105 => x"00000000",
           106 => x"00000000",
           107 => x"00000000",
           108 => x"00000000",
           109 => x"00000000",
           110 => x"00000000",
           111 => x"00000000",
           112 => x"00000000",
           113 => x"00000000",
           114 => x"00000000",
           115 => x"00000000",
           116 => x"00000000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"00000000",
           121 => x"00000000",
           122 => x"00000000",
           123 => x"00000000",
           124 => x"00000000",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"00000000",
           129 => x"00000000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"00000000",
           137 => x"00000000",
           138 => x"00000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"00000000",
           145 => x"00000000",
           146 => x"00000000",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"00000000",
           153 => x"00000000",
           154 => x"00000000",
           155 => x"00000000",
           156 => x"00000000",
           157 => x"00000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"00000000",
           161 => x"00000000",
           162 => x"00000000",
           163 => x"00000000",
           164 => x"00000000",
           165 => x"00000000",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"00000000",
           169 => x"00000000",
           170 => x"00000000",
           171 => x"00000000",
           172 => x"00000000",
           173 => x"00000000",
           174 => x"00000000",
           175 => x"00000000",
           176 => x"00000000",
           177 => x"00000000",
           178 => x"00000000",
           179 => x"00000000",
           180 => x"00000000",
           181 => x"00000000",
           182 => x"00000000",
           183 => x"00000000",
           184 => x"00000000",
           185 => x"00000000",
           186 => x"00000000",
           187 => x"00000000",
           188 => x"00000000",
           189 => x"00000000",
           190 => x"00000000",
           191 => x"00000000",
           192 => x"00000000",
           193 => x"00000000",
           194 => x"00000000",
           195 => x"00000000",
           196 => x"00000000",
           197 => x"00000000",
           198 => x"00000000",
           199 => x"00000000",
           200 => x"00000000",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"00000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"00000000",
           217 => x"00000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"00000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"00000000",
           233 => x"00000000",
           234 => x"00000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"00000000",
           249 => x"00000000",
           250 => x"00000000",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00888004",
           257 => x"81cbe00c",
           258 => x"98f62d81",
           259 => x"cbe00888",
           260 => x"80809004",
           261 => x"81cbe00c",
           262 => x"a3a62d81",
           263 => x"cbe00888",
           264 => x"80809004",
           265 => x"81cbe00c",
           266 => x"a3e52d81",
           267 => x"cbe00888",
           268 => x"80809004",
           269 => x"81cbe00c",
           270 => x"a4832d81",
           271 => x"cbe00888",
           272 => x"80809004",
           273 => x"81cbe00c",
           274 => x"aac12d81",
           275 => x"cbe00888",
           276 => x"80809004",
           277 => x"81cbe00c",
           278 => x"abbf2d81",
           279 => x"cbe00888",
           280 => x"80809004",
           281 => x"81cbe00c",
           282 => x"a4a62d81",
           283 => x"cbe00888",
           284 => x"80809004",
           285 => x"81cbe00c",
           286 => x"abdc2d81",
           287 => x"cbe00888",
           288 => x"80809004",
           289 => x"81cbe00c",
           290 => x"adce2d81",
           291 => x"cbe00888",
           292 => x"80809004",
           293 => x"81cbe00c",
           294 => x"a9e72d81",
           295 => x"cbe00888",
           296 => x"80809004",
           297 => x"81cbe00c",
           298 => x"a9fd2d81",
           299 => x"cbe00888",
           300 => x"80809004",
           301 => x"81cbe00c",
           302 => x"aaa12d81",
           303 => x"cbe00888",
           304 => x"80809004",
           305 => x"81cbe00c",
           306 => x"9b832d81",
           307 => x"cbe00888",
           308 => x"80809004",
           309 => x"81cbe00c",
           310 => x"9bd42d81",
           311 => x"cbe00888",
           312 => x"80809004",
           313 => x"81cbe00c",
           314 => x"93f02d81",
           315 => x"cbe00888",
           316 => x"80809004",
           317 => x"81cbe00c",
           318 => x"95a52d81",
           319 => x"cbe00888",
           320 => x"80809004",
           321 => x"81cbe00c",
           322 => x"96d82d81",
           323 => x"cbe00888",
           324 => x"80809004",
           325 => x"81cbe00c",
           326 => x"80e0832d",
           327 => x"81cbe008",
           328 => x"88808090",
           329 => x"0481cbe0",
           330 => x"0c80ecf4",
           331 => x"2d81cbe0",
           332 => x"08888080",
           333 => x"900481cb",
           334 => x"e00c80e4",
           335 => x"e82d81cb",
           336 => x"e0088880",
           337 => x"80900481",
           338 => x"cbe00c80",
           339 => x"e7e52d81",
           340 => x"cbe00888",
           341 => x"80809004",
           342 => x"81cbe00c",
           343 => x"80f2832d",
           344 => x"81cbe008",
           345 => x"88808090",
           346 => x"0481cbe0",
           347 => x"0c80fae3",
           348 => x"2d81cbe0",
           349 => x"08888080",
           350 => x"900481cb",
           351 => x"e00c80eb",
           352 => x"d62d81cb",
           353 => x"e0088880",
           354 => x"80900481",
           355 => x"cbe00c80",
           356 => x"f5a22d81",
           357 => x"cbe00888",
           358 => x"80809004",
           359 => x"81cbe00c",
           360 => x"80f6c12d",
           361 => x"81cbe008",
           362 => x"88808090",
           363 => x"0481cbe0",
           364 => x"0c80f6e0",
           365 => x"2d81cbe0",
           366 => x"08888080",
           367 => x"900481cb",
           368 => x"e00c80fe",
           369 => x"ca2d81cb",
           370 => x"e0088880",
           371 => x"80900481",
           372 => x"cbe00c80",
           373 => x"fcb02d81",
           374 => x"cbe00888",
           375 => x"80809004",
           376 => x"81cbe00c",
           377 => x"81819e2d",
           378 => x"81cbe008",
           379 => x"88808090",
           380 => x"0481cbe0",
           381 => x"0c80f7e4",
           382 => x"2d81cbe0",
           383 => x"08888080",
           384 => x"900481cb",
           385 => x"e00c8184",
           386 => x"9e2d81cb",
           387 => x"e0088880",
           388 => x"80900481",
           389 => x"cbe00c81",
           390 => x"859f2d81",
           391 => x"cbe00888",
           392 => x"80809004",
           393 => x"81cbe00c",
           394 => x"80edd42d",
           395 => x"81cbe008",
           396 => x"88808090",
           397 => x"0481cbe0",
           398 => x"0c80edad",
           399 => x"2d81cbe0",
           400 => x"08888080",
           401 => x"900481cb",
           402 => x"e00c80ee",
           403 => x"d82d81cb",
           404 => x"e0088880",
           405 => x"80900481",
           406 => x"cbe00c80",
           407 => x"f8bb2d81",
           408 => x"cbe00888",
           409 => x"80809004",
           410 => x"81cbe00c",
           411 => x"8186902d",
           412 => x"81cbe008",
           413 => x"88808090",
           414 => x"0481cbe0",
           415 => x"0c81889a",
           416 => x"2d81cbe0",
           417 => x"08888080",
           418 => x"900481cb",
           419 => x"e00c818b",
           420 => x"dc2d81cb",
           421 => x"e0088880",
           422 => x"80900481",
           423 => x"cbe00c80",
           424 => x"dfa22d81",
           425 => x"cbe00888",
           426 => x"80809004",
           427 => x"81cbe00c",
           428 => x"818ec82d",
           429 => x"81cbe008",
           430 => x"88808090",
           431 => x"0481cbe0",
           432 => x"0cb0dd2d",
           433 => x"81cbe008",
           434 => x"88808090",
           435 => x"0481cbe0",
           436 => x"0cb2c72d",
           437 => x"81cbe008",
           438 => x"88808090",
           439 => x"0481cbe0",
           440 => x"0cb4ab2d",
           441 => x"81cbe008",
           442 => x"88808090",
           443 => x"0481cbe0",
           444 => x"0c94992d",
           445 => x"81cbe008",
           446 => x"88808090",
           447 => x"0481cbe0",
           448 => x"0c94fb2d",
           449 => x"81cbe008",
           450 => x"88808090",
           451 => x"0481cbe0",
           452 => x"0c97e82d",
           453 => x"81cbe008",
           454 => x"88808090",
           455 => x"0481cbe0",
           456 => x"0c819ae9",
           457 => x"2d81cbe0",
           458 => x"08888080",
           459 => x"900481cb",
           460 => x"d47081e2",
           461 => x"d8278e38",
           462 => x"80717084",
           463 => x"05530c0b",
           464 => x"0b0b8eb1",
           465 => x"04888051",
           466 => x"81b4bd04",
           467 => x"3c0481cb",
           468 => x"e0080281",
           469 => x"cbe00cfd",
           470 => x"3d0d8053",
           471 => x"81cbe008",
           472 => x"8c050852",
           473 => x"81cbe008",
           474 => x"88050851",
           475 => x"80c53f81",
           476 => x"cbd40870",
           477 => x"81cbd40c",
           478 => x"54853d0d",
           479 => x"81cbe00c",
           480 => x"0481cbe0",
           481 => x"080281cb",
           482 => x"e00cfd3d",
           483 => x"0d815381",
           484 => x"cbe0088c",
           485 => x"05085281",
           486 => x"cbe00888",
           487 => x"05085193",
           488 => x"3f81cbd4",
           489 => x"087081cb",
           490 => x"d40c5485",
           491 => x"3d0d81cb",
           492 => x"e00c0481",
           493 => x"cbe00802",
           494 => x"81cbe00c",
           495 => x"fd3d0d81",
           496 => x"0b81cbe0",
           497 => x"08fc050c",
           498 => x"800b81cb",
           499 => x"e008f805",
           500 => x"0c81cbe0",
           501 => x"088c0508",
           502 => x"81cbe008",
           503 => x"88050827",
           504 => x"b93881cb",
           505 => x"e008fc05",
           506 => x"08802eae",
           507 => x"38800b81",
           508 => x"cbe0088c",
           509 => x"050824a2",
           510 => x"3881cbe0",
           511 => x"088c0508",
           512 => x"1081cbe0",
           513 => x"088c050c",
           514 => x"81cbe008",
           515 => x"fc050810",
           516 => x"81cbe008",
           517 => x"fc050cff",
           518 => x"b83981cb",
           519 => x"e008fc05",
           520 => x"08802e80",
           521 => x"e13881cb",
           522 => x"e0088c05",
           523 => x"0881cbe0",
           524 => x"08880508",
           525 => x"26ad3881",
           526 => x"cbe00888",
           527 => x"050881cb",
           528 => x"e0088c05",
           529 => x"083181cb",
           530 => x"e0088805",
           531 => x"0c81cbe0",
           532 => x"08f80508",
           533 => x"81cbe008",
           534 => x"fc050807",
           535 => x"81cbe008",
           536 => x"f8050c81",
           537 => x"cbe008fc",
           538 => x"0508812a",
           539 => x"81cbe008",
           540 => x"fc050c81",
           541 => x"cbe0088c",
           542 => x"0508812a",
           543 => x"81cbe008",
           544 => x"8c050cff",
           545 => x"953981cb",
           546 => x"e0089005",
           547 => x"08802e93",
           548 => x"3881cbe0",
           549 => x"08880508",
           550 => x"7081cbe0",
           551 => x"08f4050c",
           552 => x"51913981",
           553 => x"cbe008f8",
           554 => x"05087081",
           555 => x"cbe008f4",
           556 => x"050c5181",
           557 => x"cbe008f4",
           558 => x"050881cb",
           559 => x"d40c853d",
           560 => x"0d81cbe0",
           561 => x"0c04fc3d",
           562 => x"0d767971",
           563 => x"028c059f",
           564 => x"05335755",
           565 => x"53558372",
           566 => x"278a3874",
           567 => x"83065170",
           568 => x"802ea438",
           569 => x"ff125271",
           570 => x"ff2e9338",
           571 => x"73737081",
           572 => x"055534ff",
           573 => x"125271ff",
           574 => x"2e098106",
           575 => x"ef387481",
           576 => x"cbd40c86",
           577 => x"3d0d0474",
           578 => x"74882b75",
           579 => x"07707190",
           580 => x"2b075154",
           581 => x"518f7227",
           582 => x"a5387271",
           583 => x"70840553",
           584 => x"0c727170",
           585 => x"8405530c",
           586 => x"72717084",
           587 => x"05530c72",
           588 => x"71708405",
           589 => x"530cf012",
           590 => x"52718f26",
           591 => x"dd388372",
           592 => x"27903872",
           593 => x"71708405",
           594 => x"530cfc12",
           595 => x"52718326",
           596 => x"f2387053",
           597 => x"ff8e39fb",
           598 => x"3d0d7779",
           599 => x"70720783",
           600 => x"06535452",
           601 => x"70933871",
           602 => x"73730854",
           603 => x"56547173",
           604 => x"082e80c6",
           605 => x"38737554",
           606 => x"52713370",
           607 => x"81ff0652",
           608 => x"5470802e",
           609 => x"9d387233",
           610 => x"5570752e",
           611 => x"09810695",
           612 => x"38811281",
           613 => x"14713370",
           614 => x"81ff0654",
           615 => x"56545270",
           616 => x"e5387233",
           617 => x"557381ff",
           618 => x"067581ff",
           619 => x"06717131",
           620 => x"81cbd40c",
           621 => x"5252873d",
           622 => x"0d047109",
           623 => x"70f7fbfd",
           624 => x"ff140670",
           625 => x"f8848281",
           626 => x"80065151",
           627 => x"51709738",
           628 => x"84148416",
           629 => x"71085456",
           630 => x"54717508",
           631 => x"2edc3873",
           632 => x"755452ff",
           633 => x"9439800b",
           634 => x"81cbd40c",
           635 => x"873d0d04",
           636 => x"fe3d0d80",
           637 => x"52835371",
           638 => x"882b5287",
           639 => x"863f81cb",
           640 => x"d40881ff",
           641 => x"067207ff",
           642 => x"14545272",
           643 => x"8025e838",
           644 => x"7181cbd4",
           645 => x"0c843d0d",
           646 => x"04fb3d0d",
           647 => x"77700870",
           648 => x"53535671",
           649 => x"802e80ca",
           650 => x"38713351",
           651 => x"70a02e09",
           652 => x"81068638",
           653 => x"811252f1",
           654 => x"39715384",
           655 => x"39811353",
           656 => x"80733370",
           657 => x"81ff0653",
           658 => x"555570a0",
           659 => x"2e833881",
           660 => x"5570802e",
           661 => x"843874e5",
           662 => x"387381ff",
           663 => x"065170a0",
           664 => x"2e098106",
           665 => x"88388073",
           666 => x"70810555",
           667 => x"3472760c",
           668 => x"71517081",
           669 => x"cbd40c87",
           670 => x"3d0d04fc",
           671 => x"3d0d7653",
           672 => x"7208802e",
           673 => x"9138863d",
           674 => x"fc055272",
           675 => x"5198bf3f",
           676 => x"81cbd408",
           677 => x"85388053",
           678 => x"83397453",
           679 => x"7281cbd4",
           680 => x"0c863d0d",
           681 => x"04fc3d0d",
           682 => x"76821133",
           683 => x"ff055253",
           684 => x"8152708b",
           685 => x"26819838",
           686 => x"831333ff",
           687 => x"05518252",
           688 => x"709e2681",
           689 => x"8a388413",
           690 => x"33518352",
           691 => x"70972680",
           692 => x"fe388513",
           693 => x"33518452",
           694 => x"70bb2680",
           695 => x"f2388613",
           696 => x"33518552",
           697 => x"70bb2680",
           698 => x"e6388813",
           699 => x"22558652",
           700 => x"7487e726",
           701 => x"80d9388a",
           702 => x"13225487",
           703 => x"527387e7",
           704 => x"2680cc38",
           705 => x"810b87c0",
           706 => x"989c0c72",
           707 => x"2287c098",
           708 => x"bc0c8213",
           709 => x"3387c098",
           710 => x"b80c8313",
           711 => x"3387c098",
           712 => x"b40c8413",
           713 => x"3387c098",
           714 => x"b00c8513",
           715 => x"3387c098",
           716 => x"ac0c8613",
           717 => x"3387c098",
           718 => x"a80c7487",
           719 => x"c098a40c",
           720 => x"7387c098",
           721 => x"a00c800b",
           722 => x"87c0989c",
           723 => x"0c805271",
           724 => x"81cbd40c",
           725 => x"863d0d04",
           726 => x"f33d0d7f",
           727 => x"5b87c098",
           728 => x"9c5d817d",
           729 => x"0c87c098",
           730 => x"bc085e7d",
           731 => x"7b2387c0",
           732 => x"98b8085a",
           733 => x"79821c34",
           734 => x"87c098b4",
           735 => x"085a7983",
           736 => x"1c3487c0",
           737 => x"98b0085a",
           738 => x"79841c34",
           739 => x"87c098ac",
           740 => x"085a7985",
           741 => x"1c3487c0",
           742 => x"98a8085a",
           743 => x"79861c34",
           744 => x"87c098a4",
           745 => x"085c7b88",
           746 => x"1c2387c0",
           747 => x"98a0085a",
           748 => x"798a1c23",
           749 => x"807d0c79",
           750 => x"83ffff06",
           751 => x"597b83ff",
           752 => x"ff065886",
           753 => x"1b335785",
           754 => x"1b335684",
           755 => x"1b335583",
           756 => x"1b335482",
           757 => x"1b33537d",
           758 => x"83ffff06",
           759 => x"5281b688",
           760 => x"5192843f",
           761 => x"8f3d0d04",
           762 => x"ff3d0d02",
           763 => x"8f053370",
           764 => x"30709f2a",
           765 => x"51525270",
           766 => x"0b0b81c8",
           767 => x"bc34833d",
           768 => x"0d04fb3d",
           769 => x"0d770b0b",
           770 => x"81c8bc33",
           771 => x"7081ff06",
           772 => x"57555687",
           773 => x"c0948451",
           774 => x"74802e86",
           775 => x"3887c094",
           776 => x"94517008",
           777 => x"70962a70",
           778 => x"81065354",
           779 => x"5270802e",
           780 => x"8c387191",
           781 => x"2a708106",
           782 => x"515170d7",
           783 => x"38728132",
           784 => x"70810651",
           785 => x"5170802e",
           786 => x"8d387193",
           787 => x"2a708106",
           788 => x"515170ff",
           789 => x"be387381",
           790 => x"ff065187",
           791 => x"c0948052",
           792 => x"70802e86",
           793 => x"3887c094",
           794 => x"90527572",
           795 => x"0c7581cb",
           796 => x"d40c873d",
           797 => x"0d04fb3d",
           798 => x"0d029f05",
           799 => x"330b0b81",
           800 => x"c8bc3370",
           801 => x"81ff0657",
           802 => x"555687c0",
           803 => x"94845174",
           804 => x"802e8638",
           805 => x"87c09494",
           806 => x"51700870",
           807 => x"962a7081",
           808 => x"06535452",
           809 => x"70802e8c",
           810 => x"3871912a",
           811 => x"70810651",
           812 => x"5170d738",
           813 => x"72813270",
           814 => x"81065151",
           815 => x"70802e8d",
           816 => x"3871932a",
           817 => x"70810651",
           818 => x"5170ffbe",
           819 => x"387381ff",
           820 => x"065187c0",
           821 => x"94805270",
           822 => x"802e8638",
           823 => x"87c09490",
           824 => x"5275720c",
           825 => x"873d0d04",
           826 => x"f93d0d79",
           827 => x"54807433",
           828 => x"7081ff06",
           829 => x"53535770",
           830 => x"772e80fe",
           831 => x"387181ff",
           832 => x"0681150b",
           833 => x"0b81c8bc",
           834 => x"337081ff",
           835 => x"06595755",
           836 => x"5887c094",
           837 => x"84517580",
           838 => x"2e863887",
           839 => x"c0949451",
           840 => x"70087096",
           841 => x"2a708106",
           842 => x"53545270",
           843 => x"802e8c38",
           844 => x"71912a70",
           845 => x"81065151",
           846 => x"70d73872",
           847 => x"81327081",
           848 => x"06515170",
           849 => x"802e8d38",
           850 => x"71932a70",
           851 => x"81065151",
           852 => x"70ffbe38",
           853 => x"7481ff06",
           854 => x"5187c094",
           855 => x"80527080",
           856 => x"2e863887",
           857 => x"c0949052",
           858 => x"77720c81",
           859 => x"17743370",
           860 => x"81ff0653",
           861 => x"535770ff",
           862 => x"84387681",
           863 => x"cbd40c89",
           864 => x"3d0d04fe",
           865 => x"3d0d0b0b",
           866 => x"81c8bc33",
           867 => x"7081ff06",
           868 => x"545287c0",
           869 => x"94845172",
           870 => x"802e8638",
           871 => x"87c09494",
           872 => x"51700870",
           873 => x"822a7081",
           874 => x"06515151",
           875 => x"70802ee2",
           876 => x"387181ff",
           877 => x"065187c0",
           878 => x"94805270",
           879 => x"802e8638",
           880 => x"87c09490",
           881 => x"52710870",
           882 => x"81ff0681",
           883 => x"cbd40c51",
           884 => x"843d0d04",
           885 => x"fe3d0d0b",
           886 => x"0b81c8bc",
           887 => x"337081ff",
           888 => x"06525387",
           889 => x"c0948452",
           890 => x"70802e86",
           891 => x"3887c094",
           892 => x"94527108",
           893 => x"70822a70",
           894 => x"81065151",
           895 => x"51ff5270",
           896 => x"802ea038",
           897 => x"7281ff06",
           898 => x"5187c094",
           899 => x"80527080",
           900 => x"2e863887",
           901 => x"c0949052",
           902 => x"71087098",
           903 => x"2b70982c",
           904 => x"51535171",
           905 => x"81cbd40c",
           906 => x"843d0d04",
           907 => x"ff3d0d87",
           908 => x"c09e8008",
           909 => x"709c2a8a",
           910 => x"06515170",
           911 => x"802e8393",
           912 => x"3887c09e",
           913 => x"9c0881c8",
           914 => x"c00c87c0",
           915 => x"9ea00881",
           916 => x"c8c40c87",
           917 => x"c09e8c08",
           918 => x"81c8c80c",
           919 => x"87c09e90",
           920 => x"0881c8cc",
           921 => x"0c87c09e",
           922 => x"940881c8",
           923 => x"d00c87c0",
           924 => x"9e980881",
           925 => x"c8d40c87",
           926 => x"c09ea408",
           927 => x"81c8d80c",
           928 => x"87c09ea8",
           929 => x"0881c8dc",
           930 => x"0c87c09e",
           931 => x"ac0881c8",
           932 => x"e00c87c0",
           933 => x"9e800851",
           934 => x"7081c8e4",
           935 => x"2387c09e",
           936 => x"840881c8",
           937 => x"e80c810b",
           938 => x"81c8ec34",
           939 => x"800b87c0",
           940 => x"9e880870",
           941 => x"a0800651",
           942 => x"52527080",
           943 => x"2e833881",
           944 => x"527181c8",
           945 => x"ed34800b",
           946 => x"87c09e88",
           947 => x"08708180",
           948 => x"80065152",
           949 => x"5270802e",
           950 => x"83388152",
           951 => x"7181c8ee",
           952 => x"34800b87",
           953 => x"c09e8808",
           954 => x"7080c080",
           955 => x"06515252",
           956 => x"70802e83",
           957 => x"38815271",
           958 => x"81c8ef34",
           959 => x"800b87c0",
           960 => x"9e880870",
           961 => x"90800651",
           962 => x"52527080",
           963 => x"2e833881",
           964 => x"527181c8",
           965 => x"f034800b",
           966 => x"87c09e88",
           967 => x"08708880",
           968 => x"06515252",
           969 => x"70802e83",
           970 => x"38815271",
           971 => x"81c8f134",
           972 => x"800b87c0",
           973 => x"9e880870",
           974 => x"84800651",
           975 => x"52527080",
           976 => x"2e833881",
           977 => x"527181c8",
           978 => x"f234800b",
           979 => x"87c09e88",
           980 => x"08708280",
           981 => x"06515252",
           982 => x"70802e83",
           983 => x"38815271",
           984 => x"81c8f334",
           985 => x"800b87c0",
           986 => x"9e880870",
           987 => x"81800651",
           988 => x"52527080",
           989 => x"2e833881",
           990 => x"527181c8",
           991 => x"f43487c0",
           992 => x"9e880870",
           993 => x"80e00670",
           994 => x"862c5151",
           995 => x"517081c8",
           996 => x"f534800b",
           997 => x"87c09e88",
           998 => x"08709006",
           999 => x"51525270",
          1000 => x"802e8338",
          1001 => x"81527181",
          1002 => x"c8f63480",
          1003 => x"0b87c09e",
          1004 => x"88087088",
          1005 => x"06515252",
          1006 => x"70802e83",
          1007 => x"38815271",
          1008 => x"81c8f734",
          1009 => x"87c09e88",
          1010 => x"08708706",
          1011 => x"51517081",
          1012 => x"c8f83483",
          1013 => x"3d0d04fd",
          1014 => x"3d0d81b6",
          1015 => x"a05184a3",
          1016 => x"3f81c8ec",
          1017 => x"33547380",
          1018 => x"2e883881",
          1019 => x"b6b45184",
          1020 => x"923f81b6",
          1021 => x"c851848b",
          1022 => x"3f81c8ed",
          1023 => x"33547380",
          1024 => x"2e923881",
          1025 => x"c8c40853",
          1026 => x"81c8c008",
          1027 => x"5281b6e0",
          1028 => x"5189d43f",
          1029 => x"81c8ee33",
          1030 => x"5473802e",
          1031 => x"923881c8",
          1032 => x"cc085381",
          1033 => x"c8c80852",
          1034 => x"81b78851",
          1035 => x"89b93f81",
          1036 => x"c8ef3354",
          1037 => x"738b3881",
          1038 => x"c8f03354",
          1039 => x"73802e92",
          1040 => x"3881c8d4",
          1041 => x"085381c8",
          1042 => x"d0085281",
          1043 => x"b7ac5189",
          1044 => x"963f81c8",
          1045 => x"f1335473",
          1046 => x"802e8838",
          1047 => x"81b7d051",
          1048 => x"83a13f81",
          1049 => x"c8f23354",
          1050 => x"73802e88",
          1051 => x"3881b7dc",
          1052 => x"5183903f",
          1053 => x"81c8f333",
          1054 => x"5473802e",
          1055 => x"883881b7",
          1056 => x"e85182ff",
          1057 => x"3f81c8f4",
          1058 => x"33547380",
          1059 => x"2e8d3881",
          1060 => x"c8f53352",
          1061 => x"81b7f451",
          1062 => x"88cd3f81",
          1063 => x"c8f63354",
          1064 => x"73802e88",
          1065 => x"3881b894",
          1066 => x"5182d83f",
          1067 => x"81c8f733",
          1068 => x"5473802e",
          1069 => x"8d3881c8",
          1070 => x"f8335281",
          1071 => x"b8b05188",
          1072 => x"a63f81b8",
          1073 => x"cc5182bb",
          1074 => x"3f81c8d8",
          1075 => x"085281b8",
          1076 => x"d8518893",
          1077 => x"3f81c8dc",
          1078 => x"085281b9",
          1079 => x"80518887",
          1080 => x"3f81c8e0",
          1081 => x"085281b9",
          1082 => x"a85187fb",
          1083 => x"3f81c8e4",
          1084 => x"225281b9",
          1085 => x"d05187ef",
          1086 => x"3f81c8e8",
          1087 => x"085281b9",
          1088 => x"f85187e3",
          1089 => x"3f853d0d",
          1090 => x"04fe3d0d",
          1091 => x"02920533",
          1092 => x"ff055271",
          1093 => x"8426ac38",
          1094 => x"7184290b",
          1095 => x"0b81b5a4",
          1096 => x"05527108",
          1097 => x"0481baa0",
          1098 => x"519d3981",
          1099 => x"baa85197",
          1100 => x"3981bab0",
          1101 => x"51913981",
          1102 => x"bab8518b",
          1103 => x"3981babc",
          1104 => x"51853981",
          1105 => x"bac451f7",
          1106 => x"9f3f843d",
          1107 => x"0d047188",
          1108 => x"800c0480",
          1109 => x"0b87c096",
          1110 => x"840c04ff",
          1111 => x"3d0d87c0",
          1112 => x"96847008",
          1113 => x"52528072",
          1114 => x"0c707407",
          1115 => x"7081c8fc",
          1116 => x"0c720c83",
          1117 => x"3d0d04ff",
          1118 => x"3d0d87c0",
          1119 => x"96847008",
          1120 => x"81c8fc0c",
          1121 => x"5280720c",
          1122 => x"73097081",
          1123 => x"c8fc0806",
          1124 => x"7081c8fc",
          1125 => x"0c730c51",
          1126 => x"833d0d04",
          1127 => x"81c8fc08",
          1128 => x"87c09684",
          1129 => x"0c04fe3d",
          1130 => x"0d029305",
          1131 => x"3353728a",
          1132 => x"2e098106",
          1133 => x"85388d51",
          1134 => x"ed3f81cb",
          1135 => x"ec085271",
          1136 => x"802e9038",
          1137 => x"72723481",
          1138 => x"cbec0881",
          1139 => x"0581cbec",
          1140 => x"0c8f3981",
          1141 => x"cbe40852",
          1142 => x"71802e85",
          1143 => x"38725171",
          1144 => x"2d843d0d",
          1145 => x"04fe3d0d",
          1146 => x"02970533",
          1147 => x"81cbe408",
          1148 => x"7681cbe4",
          1149 => x"0c5451ff",
          1150 => x"ad3f7281",
          1151 => x"cbe40c84",
          1152 => x"3d0d04fd",
          1153 => x"3d0d7554",
          1154 => x"73337081",
          1155 => x"ff065353",
          1156 => x"71802e8e",
          1157 => x"387281ff",
          1158 => x"06518114",
          1159 => x"54ff873f",
          1160 => x"e739853d",
          1161 => x"0d04fc3d",
          1162 => x"0d7781cb",
          1163 => x"e4087881",
          1164 => x"cbe40c56",
          1165 => x"54733370",
          1166 => x"81ff0653",
          1167 => x"5371802e",
          1168 => x"8e387281",
          1169 => x"ff065181",
          1170 => x"1454feda",
          1171 => x"3fe73974",
          1172 => x"81cbe40c",
          1173 => x"863d0d04",
          1174 => x"ec3d0d66",
          1175 => x"68595978",
          1176 => x"7081055a",
          1177 => x"33567580",
          1178 => x"2e84f838",
          1179 => x"75a52e09",
          1180 => x"810682de",
          1181 => x"3880707a",
          1182 => x"7081055c",
          1183 => x"33585b5b",
          1184 => x"75b02e09",
          1185 => x"81068538",
          1186 => x"815a8b39",
          1187 => x"75ad2e09",
          1188 => x"81068a38",
          1189 => x"825a7870",
          1190 => x"81055a33",
          1191 => x"5675aa2e",
          1192 => x"09810692",
          1193 => x"38778419",
          1194 => x"71087b70",
          1195 => x"81055d33",
          1196 => x"595d5953",
          1197 => x"9d39d016",
          1198 => x"53728926",
          1199 => x"95387a88",
          1200 => x"297b1005",
          1201 => x"7605d005",
          1202 => x"79708105",
          1203 => x"5b33575b",
          1204 => x"e5397580",
          1205 => x"ec327030",
          1206 => x"70720780",
          1207 => x"257880cc",
          1208 => x"32703070",
          1209 => x"72078025",
          1210 => x"73075354",
          1211 => x"58515553",
          1212 => x"73802e8c",
          1213 => x"38798407",
          1214 => x"79708105",
          1215 => x"5b33575a",
          1216 => x"75802e83",
          1217 => x"de387554",
          1218 => x"80e07627",
          1219 => x"8938e016",
          1220 => x"7081ff06",
          1221 => x"55537380",
          1222 => x"cf2e81aa",
          1223 => x"387380cf",
          1224 => x"24a23873",
          1225 => x"80c32e81",
          1226 => x"8e387380",
          1227 => x"c3248b38",
          1228 => x"7380c22e",
          1229 => x"818c3881",
          1230 => x"99397380",
          1231 => x"c42e818a",
          1232 => x"38818f39",
          1233 => x"7380d52e",
          1234 => x"81803873",
          1235 => x"80d5248a",
          1236 => x"387380d3",
          1237 => x"2e8e3880",
          1238 => x"f9397380",
          1239 => x"d82e80ee",
          1240 => x"3880ef39",
          1241 => x"77841971",
          1242 => x"08565953",
          1243 => x"80743354",
          1244 => x"5572752e",
          1245 => x"8d388115",
          1246 => x"70157033",
          1247 => x"51545572",
          1248 => x"f5387981",
          1249 => x"2a569039",
          1250 => x"74811656",
          1251 => x"53727b27",
          1252 => x"8f38a051",
          1253 => x"fc903f75",
          1254 => x"81065372",
          1255 => x"802ee938",
          1256 => x"7351fcdf",
          1257 => x"3f748116",
          1258 => x"5653727b",
          1259 => x"27fdb038",
          1260 => x"a051fbf2",
          1261 => x"3fef3977",
          1262 => x"84198312",
          1263 => x"33535953",
          1264 => x"9339825c",
          1265 => x"9539885c",
          1266 => x"91398a5c",
          1267 => x"8d39905c",
          1268 => x"89397551",
          1269 => x"fbd03ffd",
          1270 => x"86397982",
          1271 => x"2a708106",
          1272 => x"51537280",
          1273 => x"2e883877",
          1274 => x"84195953",
          1275 => x"86398418",
          1276 => x"78545872",
          1277 => x"087480c4",
          1278 => x"32703070",
          1279 => x"72078025",
          1280 => x"51555555",
          1281 => x"7480258d",
          1282 => x"3872802e",
          1283 => x"88387430",
          1284 => x"7a90075b",
          1285 => x"55800b8f",
          1286 => x"3d5e577b",
          1287 => x"527451e6",
          1288 => x"e03f81cb",
          1289 => x"d40881ff",
          1290 => x"067c5375",
          1291 => x"5254e69e",
          1292 => x"3f81cbd4",
          1293 => x"08558974",
          1294 => x"279238a7",
          1295 => x"14537580",
          1296 => x"f82e8438",
          1297 => x"87145372",
          1298 => x"81ff0654",
          1299 => x"b0145372",
          1300 => x"7d708105",
          1301 => x"5f348117",
          1302 => x"75307077",
          1303 => x"079f2a51",
          1304 => x"5457769f",
          1305 => x"26853872",
          1306 => x"ffb13879",
          1307 => x"842a7081",
          1308 => x"06515372",
          1309 => x"802e8e38",
          1310 => x"963d7705",
          1311 => x"e00553ad",
          1312 => x"73348117",
          1313 => x"57767a81",
          1314 => x"065455b0",
          1315 => x"54728338",
          1316 => x"a0547981",
          1317 => x"2a708106",
          1318 => x"5456729f",
          1319 => x"38811755",
          1320 => x"767b2797",
          1321 => x"387351f9",
          1322 => x"fd3f7581",
          1323 => x"0653728b",
          1324 => x"38748116",
          1325 => x"56537a73",
          1326 => x"26eb3896",
          1327 => x"3d7705e0",
          1328 => x"0553ff17",
          1329 => x"ff147033",
          1330 => x"535457f9",
          1331 => x"d93f76f2",
          1332 => x"38748116",
          1333 => x"5653727b",
          1334 => x"27fb8438",
          1335 => x"a051f9c6",
          1336 => x"3fef3996",
          1337 => x"3d0d04fd",
          1338 => x"3d0d863d",
          1339 => x"70708405",
          1340 => x"52085552",
          1341 => x"7351fae0",
          1342 => x"3f853d0d",
          1343 => x"04fe3d0d",
          1344 => x"7481cbec",
          1345 => x"0c853d88",
          1346 => x"05527551",
          1347 => x"faca3f81",
          1348 => x"cbec0853",
          1349 => x"80733480",
          1350 => x"0b81cbec",
          1351 => x"0c843d0d",
          1352 => x"04fd3d0d",
          1353 => x"81cbe408",
          1354 => x"7681cbe4",
          1355 => x"0c873d88",
          1356 => x"05537752",
          1357 => x"53faa13f",
          1358 => x"7281cbe4",
          1359 => x"0c853d0d",
          1360 => x"04fb3d0d",
          1361 => x"777981cb",
          1362 => x"e8087056",
          1363 => x"54575580",
          1364 => x"5471802e",
          1365 => x"80e03881",
          1366 => x"cbe80852",
          1367 => x"712d81cb",
          1368 => x"d40881ff",
          1369 => x"06537280",
          1370 => x"2e80cb38",
          1371 => x"728d2eb9",
          1372 => x"38728832",
          1373 => x"70307080",
          1374 => x"25515152",
          1375 => x"73802e8b",
          1376 => x"3871802e",
          1377 => x"8638ff14",
          1378 => x"5497399f",
          1379 => x"7325c838",
          1380 => x"ff165273",
          1381 => x"7225c038",
          1382 => x"74145272",
          1383 => x"72348114",
          1384 => x"547251f8",
          1385 => x"813fffaf",
          1386 => x"39731552",
          1387 => x"8072348a",
          1388 => x"51f7f33f",
          1389 => x"81537281",
          1390 => x"cbd40c87",
          1391 => x"3d0d04fe",
          1392 => x"3d0d81cb",
          1393 => x"e8087581",
          1394 => x"cbe80c77",
          1395 => x"53765253",
          1396 => x"feef3f72",
          1397 => x"81cbe80c",
          1398 => x"843d0d04",
          1399 => x"f83d0d7a",
          1400 => x"7c5a5680",
          1401 => x"707a0c58",
          1402 => x"75087033",
          1403 => x"555373a0",
          1404 => x"2e098106",
          1405 => x"87388113",
          1406 => x"760ced39",
          1407 => x"73ad2e09",
          1408 => x"81068e38",
          1409 => x"81760811",
          1410 => x"770c7608",
          1411 => x"70335654",
          1412 => x"5873b02e",
          1413 => x"09810680",
          1414 => x"c2387508",
          1415 => x"8105760c",
          1416 => x"75087033",
          1417 => x"55537380",
          1418 => x"e22e8b38",
          1419 => x"90577380",
          1420 => x"f82e8538",
          1421 => x"8f398257",
          1422 => x"8113760c",
          1423 => x"75087033",
          1424 => x"5553ac39",
          1425 => x"8155a074",
          1426 => x"2780fa38",
          1427 => x"d0145380",
          1428 => x"55885789",
          1429 => x"73279838",
          1430 => x"80eb39d0",
          1431 => x"14538055",
          1432 => x"72892680",
          1433 => x"e0388639",
          1434 => x"805580d9",
          1435 => x"398a5780",
          1436 => x"55a07427",
          1437 => x"80c23880",
          1438 => x"e0742789",
          1439 => x"38e01470",
          1440 => x"81ff0655",
          1441 => x"53d01470",
          1442 => x"81ff0655",
          1443 => x"53907427",
          1444 => x"8e38f914",
          1445 => x"7081ff06",
          1446 => x"55538974",
          1447 => x"27ca3873",
          1448 => x"7727c538",
          1449 => x"74772914",
          1450 => x"76088105",
          1451 => x"770c7608",
          1452 => x"70335654",
          1453 => x"55ffba39",
          1454 => x"77802e84",
          1455 => x"38743055",
          1456 => x"74790c81",
          1457 => x"557481cb",
          1458 => x"d40c8a3d",
          1459 => x"0d04f83d",
          1460 => x"0d7a7c5a",
          1461 => x"5680707a",
          1462 => x"0c587508",
          1463 => x"70335553",
          1464 => x"73a02e09",
          1465 => x"81068738",
          1466 => x"8113760c",
          1467 => x"ed3973ad",
          1468 => x"2e098106",
          1469 => x"8e388176",
          1470 => x"0811770c",
          1471 => x"76087033",
          1472 => x"56545873",
          1473 => x"b02e0981",
          1474 => x"0680c238",
          1475 => x"75088105",
          1476 => x"760c7508",
          1477 => x"70335553",
          1478 => x"7380e22e",
          1479 => x"8b389057",
          1480 => x"7380f82e",
          1481 => x"85388f39",
          1482 => x"82578113",
          1483 => x"760c7508",
          1484 => x"70335553",
          1485 => x"ac398155",
          1486 => x"a0742780",
          1487 => x"fa38d014",
          1488 => x"53805588",
          1489 => x"57897327",
          1490 => x"983880eb",
          1491 => x"39d01453",
          1492 => x"80557289",
          1493 => x"2680e038",
          1494 => x"86398055",
          1495 => x"80d9398a",
          1496 => x"578055a0",
          1497 => x"742780c2",
          1498 => x"3880e074",
          1499 => x"278938e0",
          1500 => x"147081ff",
          1501 => x"065553d0",
          1502 => x"147081ff",
          1503 => x"06555390",
          1504 => x"74278e38",
          1505 => x"f9147081",
          1506 => x"ff065553",
          1507 => x"897427ca",
          1508 => x"38737727",
          1509 => x"c5387477",
          1510 => x"29147608",
          1511 => x"8105770c",
          1512 => x"76087033",
          1513 => x"565455ff",
          1514 => x"ba397780",
          1515 => x"2e843874",
          1516 => x"30557479",
          1517 => x"0c815574",
          1518 => x"81cbd40c",
          1519 => x"8a3d0d04",
          1520 => x"ff3d0d02",
          1521 => x"8f053351",
          1522 => x"81527072",
          1523 => x"26873881",
          1524 => x"c9801133",
          1525 => x"527181cb",
          1526 => x"d40c833d",
          1527 => x"0d04fc3d",
          1528 => x"0d029b05",
          1529 => x"33028405",
          1530 => x"9f053356",
          1531 => x"53835172",
          1532 => x"812680e0",
          1533 => x"3872842b",
          1534 => x"87c0928c",
          1535 => x"11535188",
          1536 => x"5474802e",
          1537 => x"84388188",
          1538 => x"5473720c",
          1539 => x"87c0928c",
          1540 => x"11518171",
          1541 => x"0c850b87",
          1542 => x"c0988c0c",
          1543 => x"70527108",
          1544 => x"70820651",
          1545 => x"5170802e",
          1546 => x"8a3887c0",
          1547 => x"988c0851",
          1548 => x"70ec3871",
          1549 => x"08fc8080",
          1550 => x"06527192",
          1551 => x"3887c098",
          1552 => x"8c085170",
          1553 => x"802e8738",
          1554 => x"7181c980",
          1555 => x"143481c9",
          1556 => x"80133351",
          1557 => x"7081cbd4",
          1558 => x"0c863d0d",
          1559 => x"04f33d0d",
          1560 => x"60626402",
          1561 => x"8c05bf05",
          1562 => x"33574058",
          1563 => x"5b837452",
          1564 => x"5afecd3f",
          1565 => x"81cbd408",
          1566 => x"81067a54",
          1567 => x"527181be",
          1568 => x"38717275",
          1569 => x"842b87c0",
          1570 => x"92801187",
          1571 => x"c0928c12",
          1572 => x"87c09284",
          1573 => x"13415a40",
          1574 => x"575a5885",
          1575 => x"0b87c098",
          1576 => x"8c0c767d",
          1577 => x"0c84760c",
          1578 => x"75087085",
          1579 => x"2a708106",
          1580 => x"51535471",
          1581 => x"802e8e38",
          1582 => x"7b085271",
          1583 => x"7b708105",
          1584 => x"5d348119",
          1585 => x"598074a2",
          1586 => x"06535371",
          1587 => x"732e8338",
          1588 => x"81537883",
          1589 => x"ff268f38",
          1590 => x"72802e8a",
          1591 => x"3887c098",
          1592 => x"8c085271",
          1593 => x"c33887c0",
          1594 => x"988c0852",
          1595 => x"71802e87",
          1596 => x"38788480",
          1597 => x"2e993881",
          1598 => x"760c87c0",
          1599 => x"928c1553",
          1600 => x"72087082",
          1601 => x"06515271",
          1602 => x"f738ff1a",
          1603 => x"5a8d3984",
          1604 => x"80178119",
          1605 => x"7081ff06",
          1606 => x"5a535779",
          1607 => x"802e9038",
          1608 => x"73fc8080",
          1609 => x"06527187",
          1610 => x"387d7826",
          1611 => x"feed3873",
          1612 => x"fc808006",
          1613 => x"5271802e",
          1614 => x"83388152",
          1615 => x"71537281",
          1616 => x"cbd40c8f",
          1617 => x"3d0d04f3",
          1618 => x"3d0d6062",
          1619 => x"64028c05",
          1620 => x"bf053357",
          1621 => x"40585b83",
          1622 => x"59807452",
          1623 => x"58fce13f",
          1624 => x"81cbd408",
          1625 => x"81067954",
          1626 => x"5271782e",
          1627 => x"09810681",
          1628 => x"b1387774",
          1629 => x"842b87c0",
          1630 => x"92801187",
          1631 => x"c0928c12",
          1632 => x"87c09284",
          1633 => x"1340595f",
          1634 => x"565a850b",
          1635 => x"87c0988c",
          1636 => x"0c767d0c",
          1637 => x"82760c80",
          1638 => x"58750870",
          1639 => x"842a7081",
          1640 => x"06515354",
          1641 => x"71802e8c",
          1642 => x"387a7081",
          1643 => x"055c337c",
          1644 => x"0c811858",
          1645 => x"73812a70",
          1646 => x"81065152",
          1647 => x"71802e8a",
          1648 => x"3887c098",
          1649 => x"8c085271",
          1650 => x"d03887c0",
          1651 => x"988c0852",
          1652 => x"71802e87",
          1653 => x"38778480",
          1654 => x"2e993881",
          1655 => x"760c87c0",
          1656 => x"928c1553",
          1657 => x"72087082",
          1658 => x"06515271",
          1659 => x"f738ff19",
          1660 => x"598d3981",
          1661 => x"1a7081ff",
          1662 => x"06848019",
          1663 => x"595b5278",
          1664 => x"802e9038",
          1665 => x"73fc8080",
          1666 => x"06527187",
          1667 => x"387d7a26",
          1668 => x"fef83873",
          1669 => x"fc808006",
          1670 => x"5271802e",
          1671 => x"83388152",
          1672 => x"71537281",
          1673 => x"cbd40c8f",
          1674 => x"3d0d04f6",
          1675 => x"3d0d7e02",
          1676 => x"8405b305",
          1677 => x"33028805",
          1678 => x"b7053371",
          1679 => x"54545657",
          1680 => x"fafe3f81",
          1681 => x"cbd40881",
          1682 => x"06538354",
          1683 => x"7280fe38",
          1684 => x"850b87c0",
          1685 => x"988c0c81",
          1686 => x"5671762e",
          1687 => x"80dc3871",
          1688 => x"76249338",
          1689 => x"74842b87",
          1690 => x"c0928c11",
          1691 => x"54547180",
          1692 => x"2e8d3880",
          1693 => x"d4397183",
          1694 => x"2e80c638",
          1695 => x"80cb3972",
          1696 => x"0870812a",
          1697 => x"70810651",
          1698 => x"51527180",
          1699 => x"2e8a3887",
          1700 => x"c0988c08",
          1701 => x"5271e838",
          1702 => x"87c0988c",
          1703 => x"08527196",
          1704 => x"3881730c",
          1705 => x"87c0928c",
          1706 => x"14537208",
          1707 => x"70820651",
          1708 => x"5271f738",
          1709 => x"96398056",
          1710 => x"92398880",
          1711 => x"0a770c85",
          1712 => x"39818077",
          1713 => x"0c725683",
          1714 => x"39845675",
          1715 => x"547381cb",
          1716 => x"d40c8c3d",
          1717 => x"0d04fe3d",
          1718 => x"0d748111",
          1719 => x"33713371",
          1720 => x"882b0781",
          1721 => x"cbd40c53",
          1722 => x"51843d0d",
          1723 => x"04fd3d0d",
          1724 => x"75831133",
          1725 => x"82123371",
          1726 => x"902b7188",
          1727 => x"2b078114",
          1728 => x"33707207",
          1729 => x"882b7533",
          1730 => x"710781cb",
          1731 => x"d40c5253",
          1732 => x"54565452",
          1733 => x"853d0d04",
          1734 => x"ff3d0d73",
          1735 => x"02840592",
          1736 => x"05225252",
          1737 => x"70727081",
          1738 => x"05543470",
          1739 => x"882a5170",
          1740 => x"7234833d",
          1741 => x"0d04ff3d",
          1742 => x"0d737552",
          1743 => x"52707270",
          1744 => x"81055434",
          1745 => x"70882a51",
          1746 => x"70727081",
          1747 => x"05543470",
          1748 => x"882a5170",
          1749 => x"72708105",
          1750 => x"54347088",
          1751 => x"2a517072",
          1752 => x"34833d0d",
          1753 => x"04fe3d0d",
          1754 => x"76757754",
          1755 => x"54517080",
          1756 => x"2e923871",
          1757 => x"70810553",
          1758 => x"33737081",
          1759 => x"055534ff",
          1760 => x"1151eb39",
          1761 => x"843d0d04",
          1762 => x"fe3d0d75",
          1763 => x"77765452",
          1764 => x"53727270",
          1765 => x"81055434",
          1766 => x"ff115170",
          1767 => x"f438843d",
          1768 => x"0d04fc3d",
          1769 => x"0d787779",
          1770 => x"56565374",
          1771 => x"70810556",
          1772 => x"33747081",
          1773 => x"05563371",
          1774 => x"7131ff16",
          1775 => x"56525252",
          1776 => x"72802e86",
          1777 => x"3871802e",
          1778 => x"e2387181",
          1779 => x"cbd40c86",
          1780 => x"3d0d04fe",
          1781 => x"3d0d7476",
          1782 => x"54518939",
          1783 => x"71732e8a",
          1784 => x"38811151",
          1785 => x"70335271",
          1786 => x"f3387033",
          1787 => x"81cbd40c",
          1788 => x"843d0d04",
          1789 => x"800b81cb",
          1790 => x"d40c0480",
          1791 => x"0b81cbd4",
          1792 => x"0c04f73d",
          1793 => x"0d7b5680",
          1794 => x"0b831733",
          1795 => x"565a747a",
          1796 => x"2e80d638",
          1797 => x"8154b016",
          1798 => x"0853b416",
          1799 => x"70538117",
          1800 => x"335259fa",
          1801 => x"a23f81cb",
          1802 => x"d4087a2e",
          1803 => x"098106b7",
          1804 => x"3881cbd4",
          1805 => x"08831734",
          1806 => x"b0160870",
          1807 => x"a4180831",
          1808 => x"9c180859",
          1809 => x"56587477",
          1810 => x"279f3882",
          1811 => x"16335574",
          1812 => x"822e0981",
          1813 => x"06933881",
          1814 => x"54761853",
          1815 => x"78528116",
          1816 => x"3351f9e3",
          1817 => x"3f833981",
          1818 => x"5a7981cb",
          1819 => x"d40c8b3d",
          1820 => x"0d04fa3d",
          1821 => x"0d787a56",
          1822 => x"56805774",
          1823 => x"b017082e",
          1824 => x"af387551",
          1825 => x"fefc3f81",
          1826 => x"cbd40857",
          1827 => x"81cbd408",
          1828 => x"9f388154",
          1829 => x"7453b416",
          1830 => x"52811633",
          1831 => x"51f7be3f",
          1832 => x"81cbd408",
          1833 => x"802e8538",
          1834 => x"ff558157",
          1835 => x"74b0170c",
          1836 => x"7681cbd4",
          1837 => x"0c883d0d",
          1838 => x"04f83d0d",
          1839 => x"7a705257",
          1840 => x"fec03f81",
          1841 => x"cbd40858",
          1842 => x"81cbd408",
          1843 => x"81913876",
          1844 => x"33557483",
          1845 => x"2e098106",
          1846 => x"80f03884",
          1847 => x"17335978",
          1848 => x"812e0981",
          1849 => x"0680e338",
          1850 => x"84805381",
          1851 => x"cbd40852",
          1852 => x"b4177052",
          1853 => x"56fd913f",
          1854 => x"82d4d552",
          1855 => x"84b21751",
          1856 => x"fc963f84",
          1857 => x"8b85a4d2",
          1858 => x"527551fc",
          1859 => x"a93f868a",
          1860 => x"85e4f252",
          1861 => x"84981751",
          1862 => x"fc9c3f90",
          1863 => x"17085284",
          1864 => x"9c1751fc",
          1865 => x"913f8c17",
          1866 => x"085284a0",
          1867 => x"1751fc86",
          1868 => x"3fa01708",
          1869 => x"810570b0",
          1870 => x"190c7955",
          1871 => x"53755281",
          1872 => x"173351f8",
          1873 => x"823f7784",
          1874 => x"18348053",
          1875 => x"80528117",
          1876 => x"3351f9d7",
          1877 => x"3f81cbd4",
          1878 => x"08802e83",
          1879 => x"38815877",
          1880 => x"81cbd40c",
          1881 => x"8a3d0d04",
          1882 => x"fb3d0d77",
          1883 => x"fe1a9812",
          1884 => x"08fe0555",
          1885 => x"56548056",
          1886 => x"7473278d",
          1887 => x"388a1422",
          1888 => x"757129ac",
          1889 => x"16080557",
          1890 => x"537581cb",
          1891 => x"d40c873d",
          1892 => x"0d04f93d",
          1893 => x"0d7a7a70",
          1894 => x"08565457",
          1895 => x"81772781",
          1896 => x"df387698",
          1897 => x"15082781",
          1898 => x"d738ff74",
          1899 => x"33545872",
          1900 => x"822e80f5",
          1901 => x"38728224",
          1902 => x"89387281",
          1903 => x"2e8d3881",
          1904 => x"bf397283",
          1905 => x"2e818e38",
          1906 => x"81b63976",
          1907 => x"812a1770",
          1908 => x"892aa416",
          1909 => x"08055374",
          1910 => x"5255fd96",
          1911 => x"3f81cbd4",
          1912 => x"08819f38",
          1913 => x"7483ff06",
          1914 => x"14b41133",
          1915 => x"81177089",
          1916 => x"2aa41808",
          1917 => x"05557654",
          1918 => x"575753fc",
          1919 => x"f53f81cb",
          1920 => x"d40880fe",
          1921 => x"387483ff",
          1922 => x"0614b411",
          1923 => x"3370882b",
          1924 => x"78077981",
          1925 => x"0671842a",
          1926 => x"5c525851",
          1927 => x"537280e2",
          1928 => x"38759fff",
          1929 => x"065880da",
          1930 => x"3976882a",
          1931 => x"a4150805",
          1932 => x"527351fc",
          1933 => x"bd3f81cb",
          1934 => x"d40880c6",
          1935 => x"38761083",
          1936 => x"fe067405",
          1937 => x"b40551f9",
          1938 => x"8d3f81cb",
          1939 => x"d40883ff",
          1940 => x"ff0658ae",
          1941 => x"3976872a",
          1942 => x"a4150805",
          1943 => x"527351fc",
          1944 => x"913f81cb",
          1945 => x"d4089b38",
          1946 => x"76822b83",
          1947 => x"fc067405",
          1948 => x"b40551f8",
          1949 => x"f83f81cb",
          1950 => x"d408f00a",
          1951 => x"06588339",
          1952 => x"81587781",
          1953 => x"cbd40c89",
          1954 => x"3d0d04f8",
          1955 => x"3d0d7a7c",
          1956 => x"7e5a5856",
          1957 => x"82598177",
          1958 => x"27829e38",
          1959 => x"76981708",
          1960 => x"27829638",
          1961 => x"75335372",
          1962 => x"792e819d",
          1963 => x"38727924",
          1964 => x"89387281",
          1965 => x"2e8d3882",
          1966 => x"80397283",
          1967 => x"2e81b838",
          1968 => x"81f73976",
          1969 => x"812a1770",
          1970 => x"892aa418",
          1971 => x"08055376",
          1972 => x"5255fb9e",
          1973 => x"3f81cbd4",
          1974 => x"085981cb",
          1975 => x"d40881d9",
          1976 => x"387483ff",
          1977 => x"0616b405",
          1978 => x"81167881",
          1979 => x"06595654",
          1980 => x"77537680",
          1981 => x"2e8f3877",
          1982 => x"842b9ff0",
          1983 => x"0674338f",
          1984 => x"06710751",
          1985 => x"53727434",
          1986 => x"810b8317",
          1987 => x"3474892a",
          1988 => x"a4170805",
          1989 => x"527551fa",
          1990 => x"d93f81cb",
          1991 => x"d4085981",
          1992 => x"cbd40881",
          1993 => x"94387483",
          1994 => x"ff0616b4",
          1995 => x"0578842a",
          1996 => x"5454768f",
          1997 => x"3877882a",
          1998 => x"743381f0",
          1999 => x"06718f06",
          2000 => x"07515372",
          2001 => x"743480ec",
          2002 => x"3976882a",
          2003 => x"a4170805",
          2004 => x"527551fa",
          2005 => x"9d3f81cb",
          2006 => x"d4085981",
          2007 => x"cbd40880",
          2008 => x"d8387783",
          2009 => x"ffff0652",
          2010 => x"761083fe",
          2011 => x"067605b4",
          2012 => x"0551f7a4",
          2013 => x"3fbe3976",
          2014 => x"872aa417",
          2015 => x"08055275",
          2016 => x"51f9ef3f",
          2017 => x"81cbd408",
          2018 => x"5981cbd4",
          2019 => x"08ab3877",
          2020 => x"f00a0677",
          2021 => x"822b83fc",
          2022 => x"067018b4",
          2023 => x"05705451",
          2024 => x"5454f6c9",
          2025 => x"3f81cbd4",
          2026 => x"088f0a06",
          2027 => x"74075272",
          2028 => x"51f7833f",
          2029 => x"810b8317",
          2030 => x"347881cb",
          2031 => x"d40c8a3d",
          2032 => x"0d04f83d",
          2033 => x"0d7a7c7e",
          2034 => x"72085956",
          2035 => x"56598175",
          2036 => x"27a43874",
          2037 => x"98170827",
          2038 => x"9d387380",
          2039 => x"2eaa38ff",
          2040 => x"53735275",
          2041 => x"51fda43f",
          2042 => x"81cbd408",
          2043 => x"5481cbd4",
          2044 => x"0880f238",
          2045 => x"93398254",
          2046 => x"80eb3981",
          2047 => x"5480e639",
          2048 => x"81cbd408",
          2049 => x"5480de39",
          2050 => x"74527851",
          2051 => x"fb843f81",
          2052 => x"cbd40858",
          2053 => x"81cbd408",
          2054 => x"802e80c7",
          2055 => x"3881cbd4",
          2056 => x"08812ed2",
          2057 => x"3881cbd4",
          2058 => x"08ff2ecf",
          2059 => x"38805374",
          2060 => x"527551fc",
          2061 => x"d63f81cb",
          2062 => x"d408c538",
          2063 => x"981608fe",
          2064 => x"11901808",
          2065 => x"57555774",
          2066 => x"74279038",
          2067 => x"81159017",
          2068 => x"0c841633",
          2069 => x"81075473",
          2070 => x"84173477",
          2071 => x"55767826",
          2072 => x"ffa63880",
          2073 => x"547381cb",
          2074 => x"d40c8a3d",
          2075 => x"0d04f63d",
          2076 => x"0d7c7e71",
          2077 => x"08595b5b",
          2078 => x"7995388c",
          2079 => x"17085877",
          2080 => x"802e8838",
          2081 => x"98170878",
          2082 => x"26b23881",
          2083 => x"58ae3979",
          2084 => x"527a51f9",
          2085 => x"fd3f8155",
          2086 => x"7481cbd4",
          2087 => x"082782e0",
          2088 => x"3881cbd4",
          2089 => x"085581cb",
          2090 => x"d408ff2e",
          2091 => x"82d23898",
          2092 => x"170881cb",
          2093 => x"d4082682",
          2094 => x"c7387958",
          2095 => x"90170870",
          2096 => x"56547380",
          2097 => x"2e82b938",
          2098 => x"777a2e09",
          2099 => x"810680e2",
          2100 => x"38811a56",
          2101 => x"98170876",
          2102 => x"26833882",
          2103 => x"5675527a",
          2104 => x"51f9af3f",
          2105 => x"805981cb",
          2106 => x"d408812e",
          2107 => x"09810686",
          2108 => x"3881cbd4",
          2109 => x"085981cb",
          2110 => x"d4080970",
          2111 => x"30707207",
          2112 => x"8025707c",
          2113 => x"0781cbd4",
          2114 => x"08545151",
          2115 => x"55557381",
          2116 => x"ef3881cb",
          2117 => x"d408802e",
          2118 => x"95388c17",
          2119 => x"08548174",
          2120 => x"27903873",
          2121 => x"98180827",
          2122 => x"89387358",
          2123 => x"85397580",
          2124 => x"db387756",
          2125 => x"81165698",
          2126 => x"17087626",
          2127 => x"89388256",
          2128 => x"75782681",
          2129 => x"ac387552",
          2130 => x"7a51f8c6",
          2131 => x"3f81cbd4",
          2132 => x"08802eb8",
          2133 => x"38805981",
          2134 => x"cbd40881",
          2135 => x"2e098106",
          2136 => x"863881cb",
          2137 => x"d4085981",
          2138 => x"cbd40809",
          2139 => x"70307072",
          2140 => x"07802570",
          2141 => x"7c075151",
          2142 => x"55557380",
          2143 => x"f8387578",
          2144 => x"2e098106",
          2145 => x"ffae3873",
          2146 => x"5580f539",
          2147 => x"ff537552",
          2148 => x"7651f9f7",
          2149 => x"3f81cbd4",
          2150 => x"0881cbd4",
          2151 => x"08307081",
          2152 => x"cbd40807",
          2153 => x"80255155",
          2154 => x"5579802e",
          2155 => x"94387380",
          2156 => x"2e8f3875",
          2157 => x"53795276",
          2158 => x"51f9d03f",
          2159 => x"81cbd408",
          2160 => x"5574a538",
          2161 => x"758c180c",
          2162 => x"981708fe",
          2163 => x"05901808",
          2164 => x"56547474",
          2165 => x"268638ff",
          2166 => x"1590180c",
          2167 => x"84173381",
          2168 => x"07547384",
          2169 => x"18349739",
          2170 => x"ff567481",
          2171 => x"2e90388c",
          2172 => x"3980558c",
          2173 => x"3981cbd4",
          2174 => x"08558539",
          2175 => x"81567555",
          2176 => x"7481cbd4",
          2177 => x"0c8c3d0d",
          2178 => x"04f83d0d",
          2179 => x"7a705255",
          2180 => x"f3f03f81",
          2181 => x"cbd40858",
          2182 => x"815681cb",
          2183 => x"d40880d8",
          2184 => x"387b5274",
          2185 => x"51f6c13f",
          2186 => x"81cbd408",
          2187 => x"81cbd408",
          2188 => x"b0170c59",
          2189 => x"84805377",
          2190 => x"52b41570",
          2191 => x"5257f2c8",
          2192 => x"3f775684",
          2193 => x"39811656",
          2194 => x"8a152258",
          2195 => x"75782797",
          2196 => x"38815475",
          2197 => x"19537652",
          2198 => x"81153351",
          2199 => x"ede93f81",
          2200 => x"cbd40880",
          2201 => x"2edf388a",
          2202 => x"15227632",
          2203 => x"70307072",
          2204 => x"07709f2a",
          2205 => x"53515656",
          2206 => x"7581cbd4",
          2207 => x"0c8a3d0d",
          2208 => x"04f83d0d",
          2209 => x"7a7c7108",
          2210 => x"58565774",
          2211 => x"f0800a26",
          2212 => x"80f13874",
          2213 => x"9f065372",
          2214 => x"80e93874",
          2215 => x"90180c88",
          2216 => x"17085473",
          2217 => x"aa387533",
          2218 => x"53827327",
          2219 => x"8838a816",
          2220 => x"0854739b",
          2221 => x"3874852a",
          2222 => x"53820b88",
          2223 => x"17225a58",
          2224 => x"72792780",
          2225 => x"fe38a816",
          2226 => x"0898180c",
          2227 => x"80cd398a",
          2228 => x"16227089",
          2229 => x"2b545872",
          2230 => x"7526b238",
          2231 => x"73527651",
          2232 => x"f5b03f81",
          2233 => x"cbd40854",
          2234 => x"81cbd408",
          2235 => x"ff2ebd38",
          2236 => x"810b81cb",
          2237 => x"d408278b",
          2238 => x"38981608",
          2239 => x"81cbd408",
          2240 => x"26853882",
          2241 => x"58bd3974",
          2242 => x"733155cb",
          2243 => x"39735275",
          2244 => x"51f4d53f",
          2245 => x"81cbd408",
          2246 => x"98180c73",
          2247 => x"94180c98",
          2248 => x"17085382",
          2249 => x"5872802e",
          2250 => x"9a388539",
          2251 => x"81589439",
          2252 => x"74892a13",
          2253 => x"98180c74",
          2254 => x"83ff0616",
          2255 => x"b4059c18",
          2256 => x"0c805877",
          2257 => x"81cbd40c",
          2258 => x"8a3d0d04",
          2259 => x"f83d0d7a",
          2260 => x"70089012",
          2261 => x"08a00559",
          2262 => x"5754f080",
          2263 => x"0a772786",
          2264 => x"38800b98",
          2265 => x"150c9814",
          2266 => x"08538455",
          2267 => x"72802e81",
          2268 => x"cb387683",
          2269 => x"ff065877",
          2270 => x"81b53881",
          2271 => x"1398150c",
          2272 => x"94140855",
          2273 => x"74923876",
          2274 => x"852a8817",
          2275 => x"22565374",
          2276 => x"7326819b",
          2277 => x"3880c039",
          2278 => x"8a1622ff",
          2279 => x"0577892a",
          2280 => x"06537281",
          2281 => x"8a387452",
          2282 => x"7351f3e6",
          2283 => x"3f81cbd4",
          2284 => x"08538255",
          2285 => x"810b81cb",
          2286 => x"d4082780",
          2287 => x"ff388155",
          2288 => x"81cbd408",
          2289 => x"ff2e80f4",
          2290 => x"38981608",
          2291 => x"81cbd408",
          2292 => x"2680ca38",
          2293 => x"7b8a3877",
          2294 => x"98150c84",
          2295 => x"5580dd39",
          2296 => x"94140852",
          2297 => x"7351f986",
          2298 => x"3f81cbd4",
          2299 => x"08538755",
          2300 => x"81cbd408",
          2301 => x"802e80c4",
          2302 => x"38825581",
          2303 => x"cbd40881",
          2304 => x"2eba3881",
          2305 => x"5581cbd4",
          2306 => x"08ff2eb0",
          2307 => x"3881cbd4",
          2308 => x"08527551",
          2309 => x"fbf33f81",
          2310 => x"cbd408a0",
          2311 => x"38729415",
          2312 => x"0c725275",
          2313 => x"51f2c13f",
          2314 => x"81cbd408",
          2315 => x"98150c76",
          2316 => x"90150c77",
          2317 => x"16b4059c",
          2318 => x"150c8055",
          2319 => x"7481cbd4",
          2320 => x"0c8a3d0d",
          2321 => x"04f73d0d",
          2322 => x"7b7d7108",
          2323 => x"5b5b5780",
          2324 => x"527651fc",
          2325 => x"ac3f81cb",
          2326 => x"d4085481",
          2327 => x"cbd40880",
          2328 => x"ec3881cb",
          2329 => x"d4085698",
          2330 => x"17085278",
          2331 => x"51f0833f",
          2332 => x"81cbd408",
          2333 => x"5481cbd4",
          2334 => x"0880d238",
          2335 => x"81cbd408",
          2336 => x"9c180870",
          2337 => x"33515458",
          2338 => x"7281e52e",
          2339 => x"09810683",
          2340 => x"38815881",
          2341 => x"cbd40855",
          2342 => x"72833881",
          2343 => x"55777507",
          2344 => x"5372802e",
          2345 => x"8e388116",
          2346 => x"56757a2e",
          2347 => x"09810688",
          2348 => x"38a53981",
          2349 => x"cbd40856",
          2350 => x"81527651",
          2351 => x"fd8e3f81",
          2352 => x"cbd40854",
          2353 => x"81cbd408",
          2354 => x"802eff9b",
          2355 => x"3873842e",
          2356 => x"09810683",
          2357 => x"38875473",
          2358 => x"81cbd40c",
          2359 => x"8b3d0d04",
          2360 => x"fd3d0d76",
          2361 => x"9a115254",
          2362 => x"ebec3f81",
          2363 => x"cbd40883",
          2364 => x"ffff0676",
          2365 => x"70335153",
          2366 => x"5371832e",
          2367 => x"09810690",
          2368 => x"38941451",
          2369 => x"ebd03f81",
          2370 => x"cbd40890",
          2371 => x"2b730753",
          2372 => x"7281cbd4",
          2373 => x"0c853d0d",
          2374 => x"04fc3d0d",
          2375 => x"77797083",
          2376 => x"ffff0654",
          2377 => x"9a125355",
          2378 => x"55ebed3f",
          2379 => x"76703351",
          2380 => x"5372832e",
          2381 => x"0981068b",
          2382 => x"3873902a",
          2383 => x"52941551",
          2384 => x"ebd63f86",
          2385 => x"3d0d04f7",
          2386 => x"3d0d7b7d",
          2387 => x"5b558475",
          2388 => x"085a5898",
          2389 => x"1508802e",
          2390 => x"818a3898",
          2391 => x"15085278",
          2392 => x"51ee8f3f",
          2393 => x"81cbd408",
          2394 => x"5881cbd4",
          2395 => x"0880f538",
          2396 => x"9c150870",
          2397 => x"33555373",
          2398 => x"86388458",
          2399 => x"80e6398b",
          2400 => x"133370bf",
          2401 => x"067081ff",
          2402 => x"06585153",
          2403 => x"72861634",
          2404 => x"81cbd408",
          2405 => x"537381e5",
          2406 => x"2e833881",
          2407 => x"5373ae2e",
          2408 => x"a9388170",
          2409 => x"74065457",
          2410 => x"72802e9e",
          2411 => x"38758f2e",
          2412 => x"993881cb",
          2413 => x"d40876df",
          2414 => x"06545472",
          2415 => x"882e0981",
          2416 => x"06833876",
          2417 => x"54737a2e",
          2418 => x"a0388052",
          2419 => x"7451fafc",
          2420 => x"3f81cbd4",
          2421 => x"085881cb",
          2422 => x"d4088938",
          2423 => x"981508fe",
          2424 => x"fa388639",
          2425 => x"800b9816",
          2426 => x"0c7781cb",
          2427 => x"d40c8b3d",
          2428 => x"0d04fb3d",
          2429 => x"0d777008",
          2430 => x"57548152",
          2431 => x"7351fcc5",
          2432 => x"3f81cbd4",
          2433 => x"085581cb",
          2434 => x"d408b438",
          2435 => x"98140852",
          2436 => x"7551ecde",
          2437 => x"3f81cbd4",
          2438 => x"085581cb",
          2439 => x"d408a038",
          2440 => x"a05381cb",
          2441 => x"d408529c",
          2442 => x"140851ea",
          2443 => x"db3f8b53",
          2444 => x"a014529c",
          2445 => x"140851ea",
          2446 => x"ac3f810b",
          2447 => x"83173474",
          2448 => x"81cbd40c",
          2449 => x"873d0d04",
          2450 => x"fd3d0d75",
          2451 => x"70089812",
          2452 => x"08547053",
          2453 => x"5553ec9a",
          2454 => x"3f81cbd4",
          2455 => x"088d389c",
          2456 => x"130853e5",
          2457 => x"7334810b",
          2458 => x"83153485",
          2459 => x"3d0d04fa",
          2460 => x"3d0d787a",
          2461 => x"5757800b",
          2462 => x"89173498",
          2463 => x"1708802e",
          2464 => x"81823880",
          2465 => x"70891855",
          2466 => x"55559c17",
          2467 => x"08147033",
          2468 => x"81165651",
          2469 => x"5271a02e",
          2470 => x"a8387185",
          2471 => x"2e098106",
          2472 => x"843881e5",
          2473 => x"5273892e",
          2474 => x"0981068b",
          2475 => x"38ae7370",
          2476 => x"81055534",
          2477 => x"81155571",
          2478 => x"73708105",
          2479 => x"55348115",
          2480 => x"558a7427",
          2481 => x"c5387515",
          2482 => x"88055280",
          2483 => x"0b811334",
          2484 => x"9c170852",
          2485 => x"8b123388",
          2486 => x"17349c17",
          2487 => x"089c1152",
          2488 => x"52e88a3f",
          2489 => x"81cbd408",
          2490 => x"760c9612",
          2491 => x"51e7e73f",
          2492 => x"81cbd408",
          2493 => x"86172398",
          2494 => x"1251e7da",
          2495 => x"3f81cbd4",
          2496 => x"08841723",
          2497 => x"883d0d04",
          2498 => x"f33d0d7f",
          2499 => x"70085e5b",
          2500 => x"80617033",
          2501 => x"51555573",
          2502 => x"af2e8338",
          2503 => x"81557380",
          2504 => x"dc2e9138",
          2505 => x"74802e8c",
          2506 => x"38941d08",
          2507 => x"881c0caa",
          2508 => x"39811541",
          2509 => x"80617033",
          2510 => x"56565673",
          2511 => x"af2e0981",
          2512 => x"06833881",
          2513 => x"567380dc",
          2514 => x"32703070",
          2515 => x"80257807",
          2516 => x"51515473",
          2517 => x"dc387388",
          2518 => x"1c0c6070",
          2519 => x"33515473",
          2520 => x"9f269638",
          2521 => x"ff800bab",
          2522 => x"1c348052",
          2523 => x"7a51f691",
          2524 => x"3f81cbd4",
          2525 => x"08558598",
          2526 => x"39913d61",
          2527 => x"a01d5c5a",
          2528 => x"5e8b53a0",
          2529 => x"527951e7",
          2530 => x"ff3f8070",
          2531 => x"59578879",
          2532 => x"33555c73",
          2533 => x"ae2e0981",
          2534 => x"0680d438",
          2535 => x"78187033",
          2536 => x"811a71ae",
          2537 => x"32703070",
          2538 => x"9f2a7382",
          2539 => x"26075151",
          2540 => x"535a5754",
          2541 => x"738c3879",
          2542 => x"17547574",
          2543 => x"34811757",
          2544 => x"db3975af",
          2545 => x"32703070",
          2546 => x"9f2a5151",
          2547 => x"547580dc",
          2548 => x"2e8c3873",
          2549 => x"802e8738",
          2550 => x"75a02682",
          2551 => x"bd387719",
          2552 => x"7e0ca454",
          2553 => x"a0762782",
          2554 => x"bd38a054",
          2555 => x"82b83978",
          2556 => x"18703381",
          2557 => x"1a5a5754",
          2558 => x"a0762781",
          2559 => x"fc3875af",
          2560 => x"32703077",
          2561 => x"80dc3270",
          2562 => x"30728025",
          2563 => x"71802507",
          2564 => x"51515651",
          2565 => x"5573802e",
          2566 => x"ac388439",
          2567 => x"81185880",
          2568 => x"781a7033",
          2569 => x"51555573",
          2570 => x"af2e0981",
          2571 => x"06833881",
          2572 => x"557380dc",
          2573 => x"32703070",
          2574 => x"80257707",
          2575 => x"51515473",
          2576 => x"db3881b5",
          2577 => x"3975ae2e",
          2578 => x"09810683",
          2579 => x"38815476",
          2580 => x"7c277407",
          2581 => x"5473802e",
          2582 => x"a2387b8b",
          2583 => x"32703077",
          2584 => x"ae327030",
          2585 => x"72802571",
          2586 => x"9f2a0753",
          2587 => x"51565155",
          2588 => x"7481a738",
          2589 => x"88578b5c",
          2590 => x"fef53975",
          2591 => x"982b5473",
          2592 => x"80258c38",
          2593 => x"7580ff06",
          2594 => x"81bbb011",
          2595 => x"33575475",
          2596 => x"51e6e13f",
          2597 => x"81cbd408",
          2598 => x"802eb238",
          2599 => x"78187033",
          2600 => x"811a7154",
          2601 => x"5a5654e6",
          2602 => x"d23f81cb",
          2603 => x"d408802e",
          2604 => x"80e838ff",
          2605 => x"1c547674",
          2606 => x"2780df38",
          2607 => x"79175475",
          2608 => x"74348117",
          2609 => x"7a115557",
          2610 => x"747434a7",
          2611 => x"39755281",
          2612 => x"bad051e5",
          2613 => x"fe3f81cb",
          2614 => x"d408bf38",
          2615 => x"ff9f1654",
          2616 => x"73992689",
          2617 => x"38e01670",
          2618 => x"81ff0657",
          2619 => x"54791754",
          2620 => x"75743481",
          2621 => x"1757fdf7",
          2622 => x"3977197e",
          2623 => x"0c76802e",
          2624 => x"99387933",
          2625 => x"547381e5",
          2626 => x"2e098106",
          2627 => x"8438857a",
          2628 => x"348454a0",
          2629 => x"76278f38",
          2630 => x"8b398655",
          2631 => x"81f23984",
          2632 => x"5680f339",
          2633 => x"8054738b",
          2634 => x"1b34807b",
          2635 => x"0858527a",
          2636 => x"51f2ce3f",
          2637 => x"81cbd408",
          2638 => x"5681cbd4",
          2639 => x"0880d738",
          2640 => x"981b0852",
          2641 => x"7651e6aa",
          2642 => x"3f81cbd4",
          2643 => x"085681cb",
          2644 => x"d40880c2",
          2645 => x"389c1b08",
          2646 => x"70335555",
          2647 => x"73802eff",
          2648 => x"be388b15",
          2649 => x"33bf0654",
          2650 => x"73861c34",
          2651 => x"8b153370",
          2652 => x"832a7081",
          2653 => x"06515558",
          2654 => x"7392388b",
          2655 => x"53795274",
          2656 => x"51e49f3f",
          2657 => x"81cbd408",
          2658 => x"802e8b38",
          2659 => x"75527a51",
          2660 => x"f3ba3fff",
          2661 => x"9f3975ab",
          2662 => x"1c335755",
          2663 => x"74802ebb",
          2664 => x"3874842e",
          2665 => x"09810680",
          2666 => x"e7387585",
          2667 => x"2a708106",
          2668 => x"77822a58",
          2669 => x"51547380",
          2670 => x"2e963875",
          2671 => x"81065473",
          2672 => x"802efbb5",
          2673 => x"38ff800b",
          2674 => x"ab1c3480",
          2675 => x"5580c139",
          2676 => x"75810654",
          2677 => x"73ba3885",
          2678 => x"55b63975",
          2679 => x"822a7081",
          2680 => x"06515473",
          2681 => x"ab38861b",
          2682 => x"3370842a",
          2683 => x"70810651",
          2684 => x"55557380",
          2685 => x"2ee13890",
          2686 => x"1b0883ff",
          2687 => x"061db405",
          2688 => x"527c51f5",
          2689 => x"db3f81cb",
          2690 => x"d408881c",
          2691 => x"0cfaea39",
          2692 => x"7481cbd4",
          2693 => x"0c8f3d0d",
          2694 => x"04f63d0d",
          2695 => x"7c5bff7b",
          2696 => x"08707173",
          2697 => x"55595c55",
          2698 => x"5973802e",
          2699 => x"81c63875",
          2700 => x"70810557",
          2701 => x"3370a026",
          2702 => x"525271ba",
          2703 => x"2e8d3870",
          2704 => x"ee3871ba",
          2705 => x"2e098106",
          2706 => x"81a53873",
          2707 => x"33d01170",
          2708 => x"81ff0651",
          2709 => x"52537089",
          2710 => x"26913882",
          2711 => x"147381ff",
          2712 => x"06d00556",
          2713 => x"5271762e",
          2714 => x"80f73880",
          2715 => x"0b81bba0",
          2716 => x"59557708",
          2717 => x"7a555776",
          2718 => x"70810558",
          2719 => x"33747081",
          2720 => x"055633ff",
          2721 => x"9f125353",
          2722 => x"53709926",
          2723 => x"8938e013",
          2724 => x"7081ff06",
          2725 => x"5451ff9f",
          2726 => x"12517099",
          2727 => x"268938e0",
          2728 => x"127081ff",
          2729 => x"06535172",
          2730 => x"30709f2a",
          2731 => x"51517272",
          2732 => x"2e098106",
          2733 => x"853870ff",
          2734 => x"be387230",
          2735 => x"74773270",
          2736 => x"30707207",
          2737 => x"9f2a739f",
          2738 => x"2a075354",
          2739 => x"54517080",
          2740 => x"2e8f3881",
          2741 => x"15841959",
          2742 => x"55837525",
          2743 => x"ff94388b",
          2744 => x"39748324",
          2745 => x"86387476",
          2746 => x"7c0c5978",
          2747 => x"51863981",
          2748 => x"cc843351",
          2749 => x"7081cbd4",
          2750 => x"0c8c3d0d",
          2751 => x"04fa3d0d",
          2752 => x"7856800b",
          2753 => x"831734ff",
          2754 => x"0bb0170c",
          2755 => x"79527551",
          2756 => x"e2e03f84",
          2757 => x"5581cbd4",
          2758 => x"08818038",
          2759 => x"84b21651",
          2760 => x"dfb43f81",
          2761 => x"cbd40883",
          2762 => x"ffff0654",
          2763 => x"83557382",
          2764 => x"d4d52e09",
          2765 => x"810680e3",
          2766 => x"38800bb4",
          2767 => x"17335657",
          2768 => x"7481e92e",
          2769 => x"09810683",
          2770 => x"38815774",
          2771 => x"81eb3270",
          2772 => x"30708025",
          2773 => x"79075151",
          2774 => x"54738a38",
          2775 => x"7481e82e",
          2776 => x"098106b5",
          2777 => x"38835381",
          2778 => x"bae05280",
          2779 => x"ea1651e0",
          2780 => x"b13f81cb",
          2781 => x"d4085581",
          2782 => x"cbd40880",
          2783 => x"2e9d3885",
          2784 => x"5381bae4",
          2785 => x"52818616",
          2786 => x"51e0973f",
          2787 => x"81cbd408",
          2788 => x"5581cbd4",
          2789 => x"08802e83",
          2790 => x"38825574",
          2791 => x"81cbd40c",
          2792 => x"883d0d04",
          2793 => x"f23d0d61",
          2794 => x"02840580",
          2795 => x"cb053358",
          2796 => x"5580750c",
          2797 => x"6051fce1",
          2798 => x"3f81cbd4",
          2799 => x"08588b56",
          2800 => x"800b81cb",
          2801 => x"d4082486",
          2802 => x"fc3881cb",
          2803 => x"d4088429",
          2804 => x"81cbf005",
          2805 => x"70085553",
          2806 => x"8c567380",
          2807 => x"2e86e638",
          2808 => x"73750c76",
          2809 => x"81fe0674",
          2810 => x"33545772",
          2811 => x"802eae38",
          2812 => x"81143351",
          2813 => x"d7ca3f81",
          2814 => x"cbd40881",
          2815 => x"ff067081",
          2816 => x"06545572",
          2817 => x"98387680",
          2818 => x"2e86b838",
          2819 => x"74822a70",
          2820 => x"81065153",
          2821 => x"8a567286",
          2822 => x"ac3886a7",
          2823 => x"39807434",
          2824 => x"77811534",
          2825 => x"81528114",
          2826 => x"3351d7b2",
          2827 => x"3f81cbd4",
          2828 => x"0881ff06",
          2829 => x"70810654",
          2830 => x"55835672",
          2831 => x"86873876",
          2832 => x"802e8f38",
          2833 => x"74822a70",
          2834 => x"81065153",
          2835 => x"8a567285",
          2836 => x"f4388070",
          2837 => x"5374525b",
          2838 => x"fda33f81",
          2839 => x"cbd40881",
          2840 => x"ff065776",
          2841 => x"822e0981",
          2842 => x"0680e238",
          2843 => x"8c3d7456",
          2844 => x"58835683",
          2845 => x"f6153370",
          2846 => x"58537280",
          2847 => x"2e8d3883",
          2848 => x"fa1551dc",
          2849 => x"e83f81cb",
          2850 => x"d4085776",
          2851 => x"78708405",
          2852 => x"5a0cff16",
          2853 => x"90165656",
          2854 => x"758025d7",
          2855 => x"38800b8d",
          2856 => x"3d545672",
          2857 => x"70840554",
          2858 => x"085b8357",
          2859 => x"7a802e95",
          2860 => x"387a5273",
          2861 => x"51fcc63f",
          2862 => x"81cbd408",
          2863 => x"81ff0657",
          2864 => x"81772789",
          2865 => x"38811656",
          2866 => x"837627d7",
          2867 => x"38815676",
          2868 => x"842e84f1",
          2869 => x"388d5676",
          2870 => x"812684e9",
          2871 => x"38bf1451",
          2872 => x"dbf43f81",
          2873 => x"cbd40883",
          2874 => x"ffff0653",
          2875 => x"7284802e",
          2876 => x"09810684",
          2877 => x"d03880ca",
          2878 => x"1451dbda",
          2879 => x"3f81cbd4",
          2880 => x"0883ffff",
          2881 => x"0658778d",
          2882 => x"3880d814",
          2883 => x"51dbde3f",
          2884 => x"81cbd408",
          2885 => x"58779c15",
          2886 => x"0c80c414",
          2887 => x"33821534",
          2888 => x"80c41433",
          2889 => x"ff117081",
          2890 => x"ff065154",
          2891 => x"558d5672",
          2892 => x"81268491",
          2893 => x"387481ff",
          2894 => x"06787129",
          2895 => x"80c11633",
          2896 => x"52595372",
          2897 => x"8a152372",
          2898 => x"802e8b38",
          2899 => x"ff137306",
          2900 => x"5372802e",
          2901 => x"86388d56",
          2902 => x"83eb3980",
          2903 => x"c51451da",
          2904 => x"f53f81cb",
          2905 => x"d4085381",
          2906 => x"cbd40888",
          2907 => x"1523728f",
          2908 => x"06578d56",
          2909 => x"7683ce38",
          2910 => x"80c71451",
          2911 => x"dad83f81",
          2912 => x"cbd40883",
          2913 => x"ffff0655",
          2914 => x"748d3880",
          2915 => x"d41451da",
          2916 => x"dc3f81cb",
          2917 => x"d4085580",
          2918 => x"c21451da",
          2919 => x"b93f81cb",
          2920 => x"d40883ff",
          2921 => x"ff06538d",
          2922 => x"5672802e",
          2923 => x"83973888",
          2924 => x"14227814",
          2925 => x"71842a05",
          2926 => x"5a5a7875",
          2927 => x"26838638",
          2928 => x"8a142252",
          2929 => x"74793151",
          2930 => x"ffb3833f",
          2931 => x"81cbd408",
          2932 => x"5581cbd4",
          2933 => x"08802e82",
          2934 => x"ec3881cb",
          2935 => x"d40880ff",
          2936 => x"fffff526",
          2937 => x"83388357",
          2938 => x"7483fff5",
          2939 => x"26833882",
          2940 => x"57749ff5",
          2941 => x"26853881",
          2942 => x"5789398d",
          2943 => x"5676802e",
          2944 => x"82c33882",
          2945 => x"15709816",
          2946 => x"0c7ba016",
          2947 => x"0c731c70",
          2948 => x"a4170c7a",
          2949 => x"1dac170c",
          2950 => x"54557683",
          2951 => x"2e098106",
          2952 => x"af3880de",
          2953 => x"1451d9ae",
          2954 => x"3f81cbd4",
          2955 => x"0883ffff",
          2956 => x"06538d56",
          2957 => x"72828e38",
          2958 => x"79828a38",
          2959 => x"80e01451",
          2960 => x"d9ab3f81",
          2961 => x"cbd408a8",
          2962 => x"150c7482",
          2963 => x"2b53a239",
          2964 => x"8d567980",
          2965 => x"2e81ee38",
          2966 => x"7713a815",
          2967 => x"0c741553",
          2968 => x"76822e8d",
          2969 => x"38741015",
          2970 => x"70812a76",
          2971 => x"81060551",
          2972 => x"5383ff13",
          2973 => x"892a538d",
          2974 => x"56729c15",
          2975 => x"082681c5",
          2976 => x"38ff0b90",
          2977 => x"150cff0b",
          2978 => x"8c150cff",
          2979 => x"800b8415",
          2980 => x"3476832e",
          2981 => x"09810681",
          2982 => x"923880e4",
          2983 => x"1451d8b6",
          2984 => x"3f81cbd4",
          2985 => x"0883ffff",
          2986 => x"06537281",
          2987 => x"2e098106",
          2988 => x"80f93881",
          2989 => x"1b527351",
          2990 => x"dbb83f81",
          2991 => x"cbd40880",
          2992 => x"ea3881cb",
          2993 => x"d4088415",
          2994 => x"3484b214",
          2995 => x"51d8873f",
          2996 => x"81cbd408",
          2997 => x"83ffff06",
          2998 => x"537282d4",
          2999 => x"d52e0981",
          3000 => x"0680c838",
          3001 => x"b41451d8",
          3002 => x"843f81cb",
          3003 => x"d408848b",
          3004 => x"85a4d22e",
          3005 => x"098106b3",
          3006 => x"38849814",
          3007 => x"51d7ee3f",
          3008 => x"81cbd408",
          3009 => x"868a85e4",
          3010 => x"f22e0981",
          3011 => x"069d3884",
          3012 => x"9c1451d7",
          3013 => x"d83f81cb",
          3014 => x"d4089015",
          3015 => x"0c84a014",
          3016 => x"51d7ca3f",
          3017 => x"81cbd408",
          3018 => x"8c150c76",
          3019 => x"743481cc",
          3020 => x"80228105",
          3021 => x"537281cc",
          3022 => x"80237286",
          3023 => x"1523800b",
          3024 => x"94150c80",
          3025 => x"567581cb",
          3026 => x"d40c903d",
          3027 => x"0d04fb3d",
          3028 => x"0d775489",
          3029 => x"5573802e",
          3030 => x"b9387308",
          3031 => x"5372802e",
          3032 => x"b1387233",
          3033 => x"5271802e",
          3034 => x"a9388613",
          3035 => x"22841522",
          3036 => x"57527176",
          3037 => x"2e098106",
          3038 => x"99388113",
          3039 => x"3351d0c0",
          3040 => x"3f81cbd4",
          3041 => x"08810652",
          3042 => x"71883871",
          3043 => x"74085455",
          3044 => x"83398053",
          3045 => x"7873710c",
          3046 => x"527481cb",
          3047 => x"d40c873d",
          3048 => x"0d04fa3d",
          3049 => x"0d02ab05",
          3050 => x"337a5889",
          3051 => x"3dfc0552",
          3052 => x"56f4e63f",
          3053 => x"8b54800b",
          3054 => x"81cbd408",
          3055 => x"24bc3881",
          3056 => x"cbd40884",
          3057 => x"2981cbf0",
          3058 => x"05700855",
          3059 => x"5573802e",
          3060 => x"84388074",
          3061 => x"34785473",
          3062 => x"802e8438",
          3063 => x"80743478",
          3064 => x"750c7554",
          3065 => x"75802e92",
          3066 => x"38805389",
          3067 => x"3d705384",
          3068 => x"0551f7b0",
          3069 => x"3f81cbd4",
          3070 => x"08547381",
          3071 => x"cbd40c88",
          3072 => x"3d0d04eb",
          3073 => x"3d0d6702",
          3074 => x"840580e7",
          3075 => x"05335959",
          3076 => x"89547880",
          3077 => x"2e84c838",
          3078 => x"77bf0670",
          3079 => x"54983dd0",
          3080 => x"0553993d",
          3081 => x"84055258",
          3082 => x"f6fa3f81",
          3083 => x"cbd40855",
          3084 => x"81cbd408",
          3085 => x"84a4387a",
          3086 => x"5c68528c",
          3087 => x"3d705256",
          3088 => x"edc63f81",
          3089 => x"cbd40855",
          3090 => x"81cbd408",
          3091 => x"92380280",
          3092 => x"d7053370",
          3093 => x"982b5557",
          3094 => x"73802583",
          3095 => x"38865577",
          3096 => x"9c065473",
          3097 => x"802e81ab",
          3098 => x"3874802e",
          3099 => x"95387484",
          3100 => x"2e098106",
          3101 => x"aa387551",
          3102 => x"eaf83f81",
          3103 => x"cbd40855",
          3104 => x"9e3902b2",
          3105 => x"05339106",
          3106 => x"547381b8",
          3107 => x"3877822a",
          3108 => x"70810651",
          3109 => x"5473802e",
          3110 => x"8e388855",
          3111 => x"83bc3977",
          3112 => x"88075874",
          3113 => x"83b43877",
          3114 => x"832a7081",
          3115 => x"06515473",
          3116 => x"802e81af",
          3117 => x"3862527a",
          3118 => x"51e8a53f",
          3119 => x"81cbd408",
          3120 => x"568288b2",
          3121 => x"0a52628e",
          3122 => x"0551d4ea",
          3123 => x"3f6254a0",
          3124 => x"0b8b1534",
          3125 => x"80536252",
          3126 => x"7a51e8bd",
          3127 => x"3f805262",
          3128 => x"9c0551d4",
          3129 => x"d13f7a54",
          3130 => x"810b8315",
          3131 => x"3475802e",
          3132 => x"80f1387a",
          3133 => x"b0110851",
          3134 => x"54805375",
          3135 => x"52973dd4",
          3136 => x"0551ddbe",
          3137 => x"3f81cbd4",
          3138 => x"085581cb",
          3139 => x"d40882ca",
          3140 => x"38b73974",
          3141 => x"82c43802",
          3142 => x"b2053370",
          3143 => x"842a7081",
          3144 => x"06515556",
          3145 => x"73802e86",
          3146 => x"38845582",
          3147 => x"ad397781",
          3148 => x"2a708106",
          3149 => x"51547380",
          3150 => x"2ea93875",
          3151 => x"81065473",
          3152 => x"802ea038",
          3153 => x"87558292",
          3154 => x"3973527a",
          3155 => x"51d6a33f",
          3156 => x"81cbd408",
          3157 => x"7bff188c",
          3158 => x"120c5555",
          3159 => x"81cbd408",
          3160 => x"81f83877",
          3161 => x"832a7081",
          3162 => x"06515473",
          3163 => x"802e8638",
          3164 => x"7780c007",
          3165 => x"587ab011",
          3166 => x"08a01b0c",
          3167 => x"63a41b0c",
          3168 => x"63537052",
          3169 => x"57e6d93f",
          3170 => x"81cbd408",
          3171 => x"81cbd408",
          3172 => x"881b0c63",
          3173 => x"9c05525a",
          3174 => x"d2d33f81",
          3175 => x"cbd40881",
          3176 => x"cbd4088c",
          3177 => x"1b0c777a",
          3178 => x"0c568617",
          3179 => x"22841a23",
          3180 => x"77901a34",
          3181 => x"800b911a",
          3182 => x"34800b9c",
          3183 => x"1a0c800b",
          3184 => x"941a0c77",
          3185 => x"852a7081",
          3186 => x"06515473",
          3187 => x"802e818d",
          3188 => x"3881cbd4",
          3189 => x"08802e81",
          3190 => x"843881cb",
          3191 => x"d408941a",
          3192 => x"0c8a1722",
          3193 => x"70892b7b",
          3194 => x"525957a8",
          3195 => x"39765278",
          3196 => x"51d79f3f",
          3197 => x"81cbd408",
          3198 => x"5781cbd4",
          3199 => x"08812683",
          3200 => x"38825581",
          3201 => x"cbd408ff",
          3202 => x"2e098106",
          3203 => x"83387955",
          3204 => x"75783156",
          3205 => x"74307076",
          3206 => x"07802551",
          3207 => x"54777627",
          3208 => x"8a388170",
          3209 => x"7506555a",
          3210 => x"73c33876",
          3211 => x"981a0c74",
          3212 => x"a9387583",
          3213 => x"ff065473",
          3214 => x"802ea238",
          3215 => x"76527a51",
          3216 => x"d6a63f81",
          3217 => x"cbd40885",
          3218 => x"3882558e",
          3219 => x"3975892a",
          3220 => x"81cbd408",
          3221 => x"059c1a0c",
          3222 => x"84398079",
          3223 => x"0c745473",
          3224 => x"81cbd40c",
          3225 => x"973d0d04",
          3226 => x"f23d0d60",
          3227 => x"63656440",
          3228 => x"405d5980",
          3229 => x"7e0c903d",
          3230 => x"fc055278",
          3231 => x"51f9cf3f",
          3232 => x"81cbd408",
          3233 => x"5581cbd4",
          3234 => x"088a3891",
          3235 => x"19335574",
          3236 => x"802e8638",
          3237 => x"745682c4",
          3238 => x"39901933",
          3239 => x"81065587",
          3240 => x"5674802e",
          3241 => x"82b63895",
          3242 => x"39820b91",
          3243 => x"1a348256",
          3244 => x"82aa3981",
          3245 => x"0b911a34",
          3246 => x"815682a0",
          3247 => x"398c1908",
          3248 => x"941a0831",
          3249 => x"55747c27",
          3250 => x"8338745c",
          3251 => x"7b802e82",
          3252 => x"89389419",
          3253 => x"087083ff",
          3254 => x"06565674",
          3255 => x"81b2387e",
          3256 => x"8a1122ff",
          3257 => x"0577892a",
          3258 => x"065b5579",
          3259 => x"a8387587",
          3260 => x"38881908",
          3261 => x"558f3998",
          3262 => x"19085278",
          3263 => x"51d5933f",
          3264 => x"81cbd408",
          3265 => x"55817527",
          3266 => x"ff9f3874",
          3267 => x"ff2effa3",
          3268 => x"3874981a",
          3269 => x"0c981908",
          3270 => x"527e51d4",
          3271 => x"cb3f81cb",
          3272 => x"d408802e",
          3273 => x"ff833881",
          3274 => x"cbd4081a",
          3275 => x"7c892a59",
          3276 => x"5777802e",
          3277 => x"80d63877",
          3278 => x"1a7f8a11",
          3279 => x"22585c55",
          3280 => x"75752785",
          3281 => x"38757a31",
          3282 => x"58775476",
          3283 => x"537c5281",
          3284 => x"1b3351ca",
          3285 => x"883f81cb",
          3286 => x"d408fed7",
          3287 => x"387e8311",
          3288 => x"33565674",
          3289 => x"802e9f38",
          3290 => x"b0160877",
          3291 => x"31557478",
          3292 => x"27943884",
          3293 => x"8053b416",
          3294 => x"52b01608",
          3295 => x"7731892b",
          3296 => x"7d0551cf",
          3297 => x"e03f7789",
          3298 => x"2b56b939",
          3299 => x"769c1a0c",
          3300 => x"94190883",
          3301 => x"ff068480",
          3302 => x"71315755",
          3303 => x"7b762783",
          3304 => x"387b569c",
          3305 => x"1908527e",
          3306 => x"51d1c73f",
          3307 => x"81cbd408",
          3308 => x"fe813875",
          3309 => x"53941908",
          3310 => x"83ff061f",
          3311 => x"b405527c",
          3312 => x"51cfa23f",
          3313 => x"7b76317e",
          3314 => x"08177f0c",
          3315 => x"761e941b",
          3316 => x"0818941c",
          3317 => x"0c5e5cfd",
          3318 => x"f3398056",
          3319 => x"7581cbd4",
          3320 => x"0c903d0d",
          3321 => x"04f23d0d",
          3322 => x"60636564",
          3323 => x"40405d58",
          3324 => x"807e0c90",
          3325 => x"3dfc0552",
          3326 => x"7751f6d2",
          3327 => x"3f81cbd4",
          3328 => x"085581cb",
          3329 => x"d4088a38",
          3330 => x"91183355",
          3331 => x"74802e86",
          3332 => x"38745683",
          3333 => x"b8399018",
          3334 => x"3370812a",
          3335 => x"70810651",
          3336 => x"56568756",
          3337 => x"74802e83",
          3338 => x"a4389539",
          3339 => x"820b9119",
          3340 => x"34825683",
          3341 => x"9839810b",
          3342 => x"91193481",
          3343 => x"56838e39",
          3344 => x"9418087c",
          3345 => x"11565674",
          3346 => x"76278438",
          3347 => x"75095c7b",
          3348 => x"802e82ec",
          3349 => x"38941808",
          3350 => x"7083ff06",
          3351 => x"56567481",
          3352 => x"fd387e8a",
          3353 => x"1122ff05",
          3354 => x"77892a06",
          3355 => x"5c557abf",
          3356 => x"38758c38",
          3357 => x"88180855",
          3358 => x"749c387a",
          3359 => x"52853998",
          3360 => x"18085277",
          3361 => x"51d7e73f",
          3362 => x"81cbd408",
          3363 => x"5581cbd4",
          3364 => x"08802e82",
          3365 => x"ab387481",
          3366 => x"2eff9138",
          3367 => x"74ff2eff",
          3368 => x"95387498",
          3369 => x"190c8818",
          3370 => x"08853874",
          3371 => x"88190c7e",
          3372 => x"55b01508",
          3373 => x"9c19082e",
          3374 => x"0981068d",
          3375 => x"387451ce",
          3376 => x"c13f81cb",
          3377 => x"d408feee",
          3378 => x"38981808",
          3379 => x"527e51d1",
          3380 => x"973f81cb",
          3381 => x"d408802e",
          3382 => x"fed23881",
          3383 => x"cbd4081b",
          3384 => x"7c892a5a",
          3385 => x"5778802e",
          3386 => x"80d53878",
          3387 => x"1b7f8a11",
          3388 => x"22585b55",
          3389 => x"75752785",
          3390 => x"38757b31",
          3391 => x"59785476",
          3392 => x"537c5281",
          3393 => x"1a3351c8",
          3394 => x"be3f81cb",
          3395 => x"d408fea6",
          3396 => x"387eb011",
          3397 => x"08783156",
          3398 => x"56747927",
          3399 => x"9b388480",
          3400 => x"53b01608",
          3401 => x"7731892b",
          3402 => x"7d0552b4",
          3403 => x"1651ccb5",
          3404 => x"3f7e5580",
          3405 => x"0b831634",
          3406 => x"78892b56",
          3407 => x"80db398c",
          3408 => x"18089419",
          3409 => x"08269338",
          3410 => x"7e51cdb6",
          3411 => x"3f81cbd4",
          3412 => x"08fde338",
          3413 => x"7e77b012",
          3414 => x"0c55769c",
          3415 => x"190c9418",
          3416 => x"0883ff06",
          3417 => x"84807131",
          3418 => x"57557b76",
          3419 => x"2783387b",
          3420 => x"569c1808",
          3421 => x"527e51cd",
          3422 => x"f93f81cb",
          3423 => x"d408fdb6",
          3424 => x"3875537c",
          3425 => x"52941808",
          3426 => x"83ff061f",
          3427 => x"b40551cb",
          3428 => x"d43f7e55",
          3429 => x"810b8316",
          3430 => x"347b7631",
          3431 => x"7e08177f",
          3432 => x"0c761e94",
          3433 => x"1a081870",
          3434 => x"941c0c8c",
          3435 => x"1b085858",
          3436 => x"5e5c7476",
          3437 => x"27833875",
          3438 => x"55748c19",
          3439 => x"0cfd9039",
          3440 => x"90183380",
          3441 => x"c0075574",
          3442 => x"90193480",
          3443 => x"567581cb",
          3444 => x"d40c903d",
          3445 => x"0d04f83d",
          3446 => x"0d7a8b3d",
          3447 => x"fc055370",
          3448 => x"5256f2ea",
          3449 => x"3f81cbd4",
          3450 => x"085781cb",
          3451 => x"d40880fb",
          3452 => x"38901633",
          3453 => x"70862a70",
          3454 => x"81065155",
          3455 => x"5573802e",
          3456 => x"80e938a0",
          3457 => x"16085278",
          3458 => x"51cce73f",
          3459 => x"81cbd408",
          3460 => x"5781cbd4",
          3461 => x"0880d438",
          3462 => x"a416088b",
          3463 => x"1133a007",
          3464 => x"5555738b",
          3465 => x"16348816",
          3466 => x"08537452",
          3467 => x"750851dd",
          3468 => x"e83f8c16",
          3469 => x"08529c15",
          3470 => x"51c9fb3f",
          3471 => x"8288b20a",
          3472 => x"52961551",
          3473 => x"c9f03f76",
          3474 => x"52921551",
          3475 => x"c9ca3f78",
          3476 => x"54810b83",
          3477 => x"15347851",
          3478 => x"ccdf3f81",
          3479 => x"cbd40890",
          3480 => x"173381bf",
          3481 => x"06555773",
          3482 => x"90173476",
          3483 => x"81cbd40c",
          3484 => x"8a3d0d04",
          3485 => x"fc3d0d76",
          3486 => x"705254fe",
          3487 => x"d93f81cb",
          3488 => x"d4085381",
          3489 => x"cbd4089c",
          3490 => x"38863dfc",
          3491 => x"05527351",
          3492 => x"f1bc3f81",
          3493 => x"cbd40853",
          3494 => x"81cbd408",
          3495 => x"873881cb",
          3496 => x"d408740c",
          3497 => x"7281cbd4",
          3498 => x"0c863d0d",
          3499 => x"04ff3d0d",
          3500 => x"843d51e6",
          3501 => x"e43f8b52",
          3502 => x"800b81cb",
          3503 => x"d408248b",
          3504 => x"3881cbd4",
          3505 => x"0881cc84",
          3506 => x"34805271",
          3507 => x"81cbd40c",
          3508 => x"833d0d04",
          3509 => x"ef3d0d80",
          3510 => x"53933dd0",
          3511 => x"0552943d",
          3512 => x"51e9c13f",
          3513 => x"81cbd408",
          3514 => x"5581cbd4",
          3515 => x"0880e038",
          3516 => x"76586352",
          3517 => x"933dd405",
          3518 => x"51e08d3f",
          3519 => x"81cbd408",
          3520 => x"5581cbd4",
          3521 => x"08bc3802",
          3522 => x"80c70533",
          3523 => x"70982b55",
          3524 => x"56738025",
          3525 => x"8938767a",
          3526 => x"94120c54",
          3527 => x"b23902a2",
          3528 => x"05337084",
          3529 => x"2a708106",
          3530 => x"51555673",
          3531 => x"802e9e38",
          3532 => x"767f5370",
          3533 => x"5254dba8",
          3534 => x"3f81cbd4",
          3535 => x"0894150c",
          3536 => x"8e3981cb",
          3537 => x"d408842e",
          3538 => x"09810683",
          3539 => x"38855574",
          3540 => x"81cbd40c",
          3541 => x"933d0d04",
          3542 => x"e43d0d6f",
          3543 => x"6f5b5b80",
          3544 => x"7a348053",
          3545 => x"9e3dffb8",
          3546 => x"05529f3d",
          3547 => x"51e8b53f",
          3548 => x"81cbd408",
          3549 => x"5781cbd4",
          3550 => x"0882fc38",
          3551 => x"7b437a7c",
          3552 => x"94110847",
          3553 => x"55586454",
          3554 => x"73802e81",
          3555 => x"ed38a052",
          3556 => x"933d7052",
          3557 => x"55d5ea3f",
          3558 => x"81cbd408",
          3559 => x"5781cbd4",
          3560 => x"0882d438",
          3561 => x"68527b51",
          3562 => x"c9c83f81",
          3563 => x"cbd40857",
          3564 => x"81cbd408",
          3565 => x"82c13869",
          3566 => x"527b51da",
          3567 => x"a33f81cb",
          3568 => x"d4084576",
          3569 => x"527451d5",
          3570 => x"b83f81cb",
          3571 => x"d4085781",
          3572 => x"cbd40882",
          3573 => x"a2388052",
          3574 => x"7451daeb",
          3575 => x"3f81cbd4",
          3576 => x"085781cb",
          3577 => x"d408a438",
          3578 => x"69527b51",
          3579 => x"d9f23f73",
          3580 => x"81cbd408",
          3581 => x"2ea63876",
          3582 => x"527451d6",
          3583 => x"cf3f81cb",
          3584 => x"d4085781",
          3585 => x"cbd40880",
          3586 => x"2ecc3876",
          3587 => x"842e0981",
          3588 => x"06863882",
          3589 => x"5781e039",
          3590 => x"7681dc38",
          3591 => x"9e3dffbc",
          3592 => x"05527451",
          3593 => x"dcc93f76",
          3594 => x"903d7811",
          3595 => x"81113351",
          3596 => x"565a5673",
          3597 => x"802e9138",
          3598 => x"02b90555",
          3599 => x"81168116",
          3600 => x"70335656",
          3601 => x"5673f538",
          3602 => x"81165473",
          3603 => x"78268190",
          3604 => x"3875802e",
          3605 => x"99387816",
          3606 => x"810555ff",
          3607 => x"186f11ff",
          3608 => x"18ff1858",
          3609 => x"58555874",
          3610 => x"33743475",
          3611 => x"ee38ff18",
          3612 => x"6f115558",
          3613 => x"af7434fe",
          3614 => x"8d39777b",
          3615 => x"2e098106",
          3616 => x"8a38ff18",
          3617 => x"6f115558",
          3618 => x"af743480",
          3619 => x"0b81cc84",
          3620 => x"33708429",
          3621 => x"81bba005",
          3622 => x"70087033",
          3623 => x"525c5656",
          3624 => x"5673762e",
          3625 => x"8d388116",
          3626 => x"701a7033",
          3627 => x"51555673",
          3628 => x"f5388216",
          3629 => x"54737826",
          3630 => x"a7388055",
          3631 => x"74762791",
          3632 => x"38741954",
          3633 => x"73337a70",
          3634 => x"81055c34",
          3635 => x"811555ec",
          3636 => x"39ba7a70",
          3637 => x"81055c34",
          3638 => x"74ff2e09",
          3639 => x"81068538",
          3640 => x"91579439",
          3641 => x"6e188119",
          3642 => x"59547333",
          3643 => x"7a708105",
          3644 => x"5c347a78",
          3645 => x"26ee3880",
          3646 => x"7a347681",
          3647 => x"cbd40c9e",
          3648 => x"3d0d04f7",
          3649 => x"3d0d7b7d",
          3650 => x"8d3dfc05",
          3651 => x"54715357",
          3652 => x"55ecbb3f",
          3653 => x"81cbd408",
          3654 => x"5381cbd4",
          3655 => x"0882fa38",
          3656 => x"91153353",
          3657 => x"7282f238",
          3658 => x"8c150854",
          3659 => x"73762792",
          3660 => x"38901533",
          3661 => x"70812a70",
          3662 => x"81065154",
          3663 => x"57728338",
          3664 => x"73569415",
          3665 => x"08548070",
          3666 => x"94170c58",
          3667 => x"75782e82",
          3668 => x"9738798a",
          3669 => x"11227089",
          3670 => x"2b595153",
          3671 => x"73782eb7",
          3672 => x"387652ff",
          3673 => x"1651ff9b",
          3674 => x"e53f81cb",
          3675 => x"d408ff15",
          3676 => x"78547053",
          3677 => x"5553ff9b",
          3678 => x"d53f81cb",
          3679 => x"d4087326",
          3680 => x"96387630",
          3681 => x"70750670",
          3682 => x"94180c77",
          3683 => x"71319818",
          3684 => x"08575851",
          3685 => x"53b13988",
          3686 => x"15085473",
          3687 => x"a6387352",
          3688 => x"7451cdca",
          3689 => x"3f81cbd4",
          3690 => x"085481cb",
          3691 => x"d408812e",
          3692 => x"819a3881",
          3693 => x"cbd408ff",
          3694 => x"2e819b38",
          3695 => x"81cbd408",
          3696 => x"88160c73",
          3697 => x"98160c73",
          3698 => x"802e819c",
          3699 => x"38767627",
          3700 => x"80dc3875",
          3701 => x"77319416",
          3702 => x"08189417",
          3703 => x"0c901633",
          3704 => x"70812a70",
          3705 => x"81065155",
          3706 => x"5a567280",
          3707 => x"2e9a3873",
          3708 => x"527451cc",
          3709 => x"f93f81cb",
          3710 => x"d4085481",
          3711 => x"cbd40894",
          3712 => x"3881cbd4",
          3713 => x"0856a739",
          3714 => x"73527451",
          3715 => x"c7843f81",
          3716 => x"cbd40854",
          3717 => x"73ff2ebe",
          3718 => x"38817427",
          3719 => x"af387953",
          3720 => x"73981408",
          3721 => x"27a63873",
          3722 => x"98160cff",
          3723 => x"a0399415",
          3724 => x"08169416",
          3725 => x"0c7583ff",
          3726 => x"06537280",
          3727 => x"2eaa3873",
          3728 => x"527951c6",
          3729 => x"a33f81cb",
          3730 => x"d4089438",
          3731 => x"820b9116",
          3732 => x"34825380",
          3733 => x"c439810b",
          3734 => x"91163481",
          3735 => x"53bb3975",
          3736 => x"892a81cb",
          3737 => x"d4080558",
          3738 => x"94150854",
          3739 => x"8c150874",
          3740 => x"27903873",
          3741 => x"8c160c90",
          3742 => x"153380c0",
          3743 => x"07537290",
          3744 => x"16347383",
          3745 => x"ff065372",
          3746 => x"802e8c38",
          3747 => x"779c1608",
          3748 => x"2e853877",
          3749 => x"9c160c80",
          3750 => x"537281cb",
          3751 => x"d40c8b3d",
          3752 => x"0d04f93d",
          3753 => x"0d795689",
          3754 => x"5475802e",
          3755 => x"818a3880",
          3756 => x"53893dfc",
          3757 => x"05528a3d",
          3758 => x"840551e1",
          3759 => x"e73f81cb",
          3760 => x"d4085581",
          3761 => x"cbd40880",
          3762 => x"ea387776",
          3763 => x"0c7a5275",
          3764 => x"51d8b53f",
          3765 => x"81cbd408",
          3766 => x"5581cbd4",
          3767 => x"0880c338",
          3768 => x"ab163370",
          3769 => x"982b5557",
          3770 => x"807424a2",
          3771 => x"38861633",
          3772 => x"70842a70",
          3773 => x"81065155",
          3774 => x"5773802e",
          3775 => x"ad389c16",
          3776 => x"08527751",
          3777 => x"d3da3f81",
          3778 => x"cbd40888",
          3779 => x"170c7754",
          3780 => x"86142284",
          3781 => x"17237452",
          3782 => x"7551cee5",
          3783 => x"3f81cbd4",
          3784 => x"08557484",
          3785 => x"2e098106",
          3786 => x"85388555",
          3787 => x"86397480",
          3788 => x"2e843880",
          3789 => x"760c7454",
          3790 => x"7381cbd4",
          3791 => x"0c893d0d",
          3792 => x"04fc3d0d",
          3793 => x"76873dfc",
          3794 => x"05537052",
          3795 => x"53e7ff3f",
          3796 => x"81cbd408",
          3797 => x"873881cb",
          3798 => x"d408730c",
          3799 => x"863d0d04",
          3800 => x"fb3d0d77",
          3801 => x"79893dfc",
          3802 => x"05547153",
          3803 => x"5654e7de",
          3804 => x"3f81cbd4",
          3805 => x"085381cb",
          3806 => x"d40880df",
          3807 => x"38749338",
          3808 => x"81cbd408",
          3809 => x"527351cd",
          3810 => x"f83f81cb",
          3811 => x"d4085380",
          3812 => x"ca3981cb",
          3813 => x"d4085273",
          3814 => x"51d3ac3f",
          3815 => x"81cbd408",
          3816 => x"5381cbd4",
          3817 => x"08842e09",
          3818 => x"81068538",
          3819 => x"80538739",
          3820 => x"81cbd408",
          3821 => x"a6387452",
          3822 => x"7351d5b3",
          3823 => x"3f725273",
          3824 => x"51cf893f",
          3825 => x"81cbd408",
          3826 => x"84327030",
          3827 => x"7072079f",
          3828 => x"2c7081cb",
          3829 => x"d4080651",
          3830 => x"51545472",
          3831 => x"81cbd40c",
          3832 => x"873d0d04",
          3833 => x"ee3d0d65",
          3834 => x"57805389",
          3835 => x"3d705396",
          3836 => x"3d5256df",
          3837 => x"af3f81cb",
          3838 => x"d4085581",
          3839 => x"cbd408b2",
          3840 => x"38645275",
          3841 => x"51d6813f",
          3842 => x"81cbd408",
          3843 => x"5581cbd4",
          3844 => x"08a03802",
          3845 => x"80cb0533",
          3846 => x"70982b55",
          3847 => x"58738025",
          3848 => x"85388655",
          3849 => x"8d397680",
          3850 => x"2e883876",
          3851 => x"527551d4",
          3852 => x"be3f7481",
          3853 => x"cbd40c94",
          3854 => x"3d0d04f0",
          3855 => x"3d0d6365",
          3856 => x"555c8053",
          3857 => x"923dec05",
          3858 => x"52933d51",
          3859 => x"ded63f81",
          3860 => x"cbd4085b",
          3861 => x"81cbd408",
          3862 => x"8280387c",
          3863 => x"740c7308",
          3864 => x"981108fe",
          3865 => x"11901308",
          3866 => x"59565855",
          3867 => x"75742691",
          3868 => x"38757c0c",
          3869 => x"81e43981",
          3870 => x"5b81cc39",
          3871 => x"825b81c7",
          3872 => x"3981cbd4",
          3873 => x"08753355",
          3874 => x"5973812e",
          3875 => x"098106bf",
          3876 => x"3882755f",
          3877 => x"57765292",
          3878 => x"3df00551",
          3879 => x"c1f43f81",
          3880 => x"cbd408ff",
          3881 => x"2ed13881",
          3882 => x"cbd40881",
          3883 => x"2ece3881",
          3884 => x"cbd40830",
          3885 => x"7081cbd4",
          3886 => x"08078025",
          3887 => x"7a058119",
          3888 => x"7f53595a",
          3889 => x"54981408",
          3890 => x"7726ca38",
          3891 => x"80f939a4",
          3892 => x"150881cb",
          3893 => x"d4085758",
          3894 => x"75983877",
          3895 => x"5281187d",
          3896 => x"5258ffbf",
          3897 => x"8d3f81cb",
          3898 => x"d4085b81",
          3899 => x"cbd40880",
          3900 => x"d6387c70",
          3901 => x"337712ff",
          3902 => x"1a5d5256",
          3903 => x"5474822e",
          3904 => x"0981069e",
          3905 => x"38b41451",
          3906 => x"ffbbcb3f",
          3907 => x"81cbd408",
          3908 => x"83ffff06",
          3909 => x"70307080",
          3910 => x"251b8219",
          3911 => x"595b5154",
          3912 => x"9b39b414",
          3913 => x"51ffbbc5",
          3914 => x"3f81cbd4",
          3915 => x"08f00a06",
          3916 => x"70307080",
          3917 => x"251b8419",
          3918 => x"595b5154",
          3919 => x"7583ff06",
          3920 => x"7a585679",
          3921 => x"ff923878",
          3922 => x"7c0c7c79",
          3923 => x"90120c84",
          3924 => x"11338107",
          3925 => x"56547484",
          3926 => x"15347a81",
          3927 => x"cbd40c92",
          3928 => x"3d0d04f9",
          3929 => x"3d0d798a",
          3930 => x"3dfc0553",
          3931 => x"705257e3",
          3932 => x"dd3f81cb",
          3933 => x"d4085681",
          3934 => x"cbd40881",
          3935 => x"a8389117",
          3936 => x"33567581",
          3937 => x"a0389017",
          3938 => x"3370812a",
          3939 => x"70810651",
          3940 => x"55558755",
          3941 => x"73802e81",
          3942 => x"8e389417",
          3943 => x"0854738c",
          3944 => x"18082781",
          3945 => x"8038739b",
          3946 => x"3881cbd4",
          3947 => x"08538817",
          3948 => x"08527651",
          3949 => x"c48c3f81",
          3950 => x"cbd40874",
          3951 => x"88190c56",
          3952 => x"80c93998",
          3953 => x"17085276",
          3954 => x"51ffbfc6",
          3955 => x"3f81cbd4",
          3956 => x"08ff2e09",
          3957 => x"81068338",
          3958 => x"815681cb",
          3959 => x"d408812e",
          3960 => x"09810685",
          3961 => x"388256a3",
          3962 => x"3975a038",
          3963 => x"775481cb",
          3964 => x"d4089815",
          3965 => x"08279438",
          3966 => x"98170853",
          3967 => x"81cbd408",
          3968 => x"527651c3",
          3969 => x"bd3f81cb",
          3970 => x"d4085694",
          3971 => x"17088c18",
          3972 => x"0c901733",
          3973 => x"80c00754",
          3974 => x"73901834",
          3975 => x"75802e85",
          3976 => x"38759118",
          3977 => x"34755574",
          3978 => x"81cbd40c",
          3979 => x"893d0d04",
          3980 => x"e23d0d82",
          3981 => x"53a03dff",
          3982 => x"a40552a1",
          3983 => x"3d51dae4",
          3984 => x"3f81cbd4",
          3985 => x"085581cb",
          3986 => x"d40881f5",
          3987 => x"387845a1",
          3988 => x"3d085295",
          3989 => x"3d705258",
          3990 => x"d1ae3f81",
          3991 => x"cbd40855",
          3992 => x"81cbd408",
          3993 => x"81db3802",
          3994 => x"80fb0533",
          3995 => x"70852a70",
          3996 => x"81065155",
          3997 => x"56865573",
          3998 => x"81c73875",
          3999 => x"982b5480",
          4000 => x"742481bd",
          4001 => x"380280d6",
          4002 => x"05337081",
          4003 => x"06585487",
          4004 => x"557681ad",
          4005 => x"386b5278",
          4006 => x"51ccc53f",
          4007 => x"81cbd408",
          4008 => x"74842a70",
          4009 => x"81065155",
          4010 => x"5673802e",
          4011 => x"80d43878",
          4012 => x"5481cbd4",
          4013 => x"08941508",
          4014 => x"2e818638",
          4015 => x"735a81cb",
          4016 => x"d4085c76",
          4017 => x"528a3d70",
          4018 => x"5254c7b5",
          4019 => x"3f81cbd4",
          4020 => x"085581cb",
          4021 => x"d40880e9",
          4022 => x"3881cbd4",
          4023 => x"08527351",
          4024 => x"cce53f81",
          4025 => x"cbd40855",
          4026 => x"81cbd408",
          4027 => x"86388755",
          4028 => x"80cf3981",
          4029 => x"cbd40884",
          4030 => x"2e883881",
          4031 => x"cbd40880",
          4032 => x"c0387751",
          4033 => x"cec23f81",
          4034 => x"cbd40881",
          4035 => x"cbd40830",
          4036 => x"7081cbd4",
          4037 => x"08078025",
          4038 => x"51555575",
          4039 => x"802e9438",
          4040 => x"73802e8f",
          4041 => x"38805375",
          4042 => x"527751c1",
          4043 => x"953f81cb",
          4044 => x"d4085574",
          4045 => x"8c387851",
          4046 => x"ffbafe3f",
          4047 => x"81cbd408",
          4048 => x"557481cb",
          4049 => x"d40ca03d",
          4050 => x"0d04e93d",
          4051 => x"0d825399",
          4052 => x"3dc00552",
          4053 => x"9a3d51d8",
          4054 => x"cb3f81cb",
          4055 => x"d4085481",
          4056 => x"cbd40882",
          4057 => x"b038785e",
          4058 => x"69528e3d",
          4059 => x"705258cf",
          4060 => x"973f81cb",
          4061 => x"d4085481",
          4062 => x"cbd40886",
          4063 => x"38885482",
          4064 => x"943981cb",
          4065 => x"d408842e",
          4066 => x"09810682",
          4067 => x"88380280",
          4068 => x"df053370",
          4069 => x"852a8106",
          4070 => x"51558654",
          4071 => x"7481f638",
          4072 => x"785a7452",
          4073 => x"8a3d7052",
          4074 => x"57c1c33f",
          4075 => x"81cbd408",
          4076 => x"75555681",
          4077 => x"cbd40883",
          4078 => x"38875481",
          4079 => x"cbd40881",
          4080 => x"2e098106",
          4081 => x"83388254",
          4082 => x"81cbd408",
          4083 => x"ff2e0981",
          4084 => x"06863881",
          4085 => x"5481b439",
          4086 => x"7381b038",
          4087 => x"81cbd408",
          4088 => x"527851c4",
          4089 => x"a43f81cb",
          4090 => x"d4085481",
          4091 => x"cbd40881",
          4092 => x"9a388b53",
          4093 => x"a052b419",
          4094 => x"51ffb78c",
          4095 => x"3f7854ae",
          4096 => x"0bb41534",
          4097 => x"7854900b",
          4098 => x"bf153482",
          4099 => x"88b20a52",
          4100 => x"80ca1951",
          4101 => x"ffb69f3f",
          4102 => x"755378b4",
          4103 => x"115351c9",
          4104 => x"f83fa053",
          4105 => x"78b41153",
          4106 => x"80d40551",
          4107 => x"ffb6b63f",
          4108 => x"7854ae0b",
          4109 => x"80d51534",
          4110 => x"7f537880",
          4111 => x"d4115351",
          4112 => x"c9d73f78",
          4113 => x"54810b83",
          4114 => x"15347751",
          4115 => x"cba43f81",
          4116 => x"cbd40854",
          4117 => x"81cbd408",
          4118 => x"b2388288",
          4119 => x"b20a5264",
          4120 => x"960551ff",
          4121 => x"b5d03f75",
          4122 => x"53645278",
          4123 => x"51c9aa3f",
          4124 => x"6454900b",
          4125 => x"8b153478",
          4126 => x"54810b83",
          4127 => x"15347851",
          4128 => x"ffb8b63f",
          4129 => x"81cbd408",
          4130 => x"548b3980",
          4131 => x"53755276",
          4132 => x"51ffbeae",
          4133 => x"3f7381cb",
          4134 => x"d40c993d",
          4135 => x"0d04da3d",
          4136 => x"0da93d84",
          4137 => x"0551d2f1",
          4138 => x"3f8253a8",
          4139 => x"3dff8405",
          4140 => x"52a93d51",
          4141 => x"d5ee3f81",
          4142 => x"cbd40855",
          4143 => x"81cbd408",
          4144 => x"82d33878",
          4145 => x"4da93d08",
          4146 => x"529d3d70",
          4147 => x"5258ccb8",
          4148 => x"3f81cbd4",
          4149 => x"085581cb",
          4150 => x"d40882b9",
          4151 => x"3802819b",
          4152 => x"053381a0",
          4153 => x"06548655",
          4154 => x"7382aa38",
          4155 => x"a053a43d",
          4156 => x"0852a83d",
          4157 => x"ff880551",
          4158 => x"ffb4ea3f",
          4159 => x"ac537752",
          4160 => x"923d7052",
          4161 => x"54ffb4dd",
          4162 => x"3faa3d08",
          4163 => x"527351cb",
          4164 => x"f73f81cb",
          4165 => x"d4085581",
          4166 => x"cbd40895",
          4167 => x"38636f2e",
          4168 => x"09810688",
          4169 => x"3865a23d",
          4170 => x"082e9238",
          4171 => x"885581e5",
          4172 => x"3981cbd4",
          4173 => x"08842e09",
          4174 => x"810681b8",
          4175 => x"387351c9",
          4176 => x"b13f81cb",
          4177 => x"d4085581",
          4178 => x"cbd40881",
          4179 => x"c8386856",
          4180 => x"9353a83d",
          4181 => x"ff950552",
          4182 => x"8d1651ff",
          4183 => x"b4873f02",
          4184 => x"af05338b",
          4185 => x"17348b16",
          4186 => x"3370842a",
          4187 => x"70810651",
          4188 => x"55557389",
          4189 => x"3874a007",
          4190 => x"54738b17",
          4191 => x"34785481",
          4192 => x"0b831534",
          4193 => x"8b163370",
          4194 => x"842a7081",
          4195 => x"06515555",
          4196 => x"73802e80",
          4197 => x"e5386e64",
          4198 => x"2e80df38",
          4199 => x"75527851",
          4200 => x"c6be3f81",
          4201 => x"cbd40852",
          4202 => x"7851ffb7",
          4203 => x"bb3f8255",
          4204 => x"81cbd408",
          4205 => x"802e80dd",
          4206 => x"3881cbd4",
          4207 => x"08527851",
          4208 => x"ffb5af3f",
          4209 => x"81cbd408",
          4210 => x"7980d411",
          4211 => x"58585581",
          4212 => x"cbd40880",
          4213 => x"c0388116",
          4214 => x"335473ae",
          4215 => x"2e098106",
          4216 => x"99386353",
          4217 => x"75527651",
          4218 => x"c6af3f78",
          4219 => x"54810b83",
          4220 => x"15348739",
          4221 => x"81cbd408",
          4222 => x"9c387751",
          4223 => x"c8ca3f81",
          4224 => x"cbd40855",
          4225 => x"81cbd408",
          4226 => x"8c387851",
          4227 => x"ffb5aa3f",
          4228 => x"81cbd408",
          4229 => x"557481cb",
          4230 => x"d40ca83d",
          4231 => x"0d04ed3d",
          4232 => x"0d0280db",
          4233 => x"05330284",
          4234 => x"0580df05",
          4235 => x"33575782",
          4236 => x"53953dd0",
          4237 => x"0552963d",
          4238 => x"51d2e93f",
          4239 => x"81cbd408",
          4240 => x"5581cbd4",
          4241 => x"0880cf38",
          4242 => x"785a6552",
          4243 => x"953dd405",
          4244 => x"51c9b53f",
          4245 => x"81cbd408",
          4246 => x"5581cbd4",
          4247 => x"08b83802",
          4248 => x"80cf0533",
          4249 => x"81a00654",
          4250 => x"865573aa",
          4251 => x"3875a706",
          4252 => x"6171098b",
          4253 => x"12337106",
          4254 => x"7a740607",
          4255 => x"51575556",
          4256 => x"748b1534",
          4257 => x"7854810b",
          4258 => x"83153478",
          4259 => x"51ffb4a9",
          4260 => x"3f81cbd4",
          4261 => x"08557481",
          4262 => x"cbd40c95",
          4263 => x"3d0d04ef",
          4264 => x"3d0d6456",
          4265 => x"8253933d",
          4266 => x"d0055294",
          4267 => x"3d51d1f4",
          4268 => x"3f81cbd4",
          4269 => x"085581cb",
          4270 => x"d40880cb",
          4271 => x"38765863",
          4272 => x"52933dd4",
          4273 => x"0551c8c0",
          4274 => x"3f81cbd4",
          4275 => x"085581cb",
          4276 => x"d408b438",
          4277 => x"0280c705",
          4278 => x"3381a006",
          4279 => x"54865573",
          4280 => x"a6388416",
          4281 => x"22861722",
          4282 => x"71902b07",
          4283 => x"5354961f",
          4284 => x"51ffb0c2",
          4285 => x"3f765481",
          4286 => x"0b831534",
          4287 => x"7651ffb3",
          4288 => x"b83f81cb",
          4289 => x"d4085574",
          4290 => x"81cbd40c",
          4291 => x"933d0d04",
          4292 => x"ea3d0d69",
          4293 => x"6b5c5a80",
          4294 => x"53983dd0",
          4295 => x"0552993d",
          4296 => x"51d1813f",
          4297 => x"81cbd408",
          4298 => x"81cbd408",
          4299 => x"307081cb",
          4300 => x"d4080780",
          4301 => x"25515557",
          4302 => x"79802e81",
          4303 => x"85388170",
          4304 => x"75065555",
          4305 => x"73802e80",
          4306 => x"f9387b5d",
          4307 => x"805f8052",
          4308 => x"8d3d7052",
          4309 => x"54ffbea9",
          4310 => x"3f81cbd4",
          4311 => x"085781cb",
          4312 => x"d40880d1",
          4313 => x"38745273",
          4314 => x"51c3dc3f",
          4315 => x"81cbd408",
          4316 => x"5781cbd4",
          4317 => x"08bf3881",
          4318 => x"cbd40881",
          4319 => x"cbd40865",
          4320 => x"5b595678",
          4321 => x"1881197b",
          4322 => x"18565955",
          4323 => x"74337434",
          4324 => x"8116568a",
          4325 => x"7827ec38",
          4326 => x"8b56751a",
          4327 => x"54807434",
          4328 => x"75802e9e",
          4329 => x"38ff1670",
          4330 => x"1b703351",
          4331 => x"555673a0",
          4332 => x"2ee8388e",
          4333 => x"3976842e",
          4334 => x"09810686",
          4335 => x"38807a34",
          4336 => x"80577630",
          4337 => x"70780780",
          4338 => x"2551547a",
          4339 => x"802e80c1",
          4340 => x"3873802e",
          4341 => x"bc387ba0",
          4342 => x"11085351",
          4343 => x"ffb1933f",
          4344 => x"81cbd408",
          4345 => x"5781cbd4",
          4346 => x"08a7387b",
          4347 => x"70335555",
          4348 => x"80c35673",
          4349 => x"832e8b38",
          4350 => x"80e45673",
          4351 => x"842e8338",
          4352 => x"a7567515",
          4353 => x"b40551ff",
          4354 => x"ade33f81",
          4355 => x"cbd4087b",
          4356 => x"0c7681cb",
          4357 => x"d40c983d",
          4358 => x"0d04e63d",
          4359 => x"0d82539c",
          4360 => x"3dffb805",
          4361 => x"529d3d51",
          4362 => x"cefa3f81",
          4363 => x"cbd40881",
          4364 => x"cbd40856",
          4365 => x"5481cbd4",
          4366 => x"08839838",
          4367 => x"8b53a052",
          4368 => x"8b3d7052",
          4369 => x"59ffaec0",
          4370 => x"3f736d70",
          4371 => x"337081ff",
          4372 => x"06525755",
          4373 => x"579f7427",
          4374 => x"81bc3878",
          4375 => x"587481ff",
          4376 => x"066d8105",
          4377 => x"4e705255",
          4378 => x"ffaf893f",
          4379 => x"81cbd408",
          4380 => x"802ea538",
          4381 => x"6c703370",
          4382 => x"535754ff",
          4383 => x"aefd3f81",
          4384 => x"cbd40880",
          4385 => x"2e8d3874",
          4386 => x"882b7607",
          4387 => x"6d81054e",
          4388 => x"55863981",
          4389 => x"cbd40855",
          4390 => x"ff9f1570",
          4391 => x"83ffff06",
          4392 => x"51547399",
          4393 => x"268a38e0",
          4394 => x"157083ff",
          4395 => x"ff065654",
          4396 => x"80ff7527",
          4397 => x"873881ba",
          4398 => x"b0153355",
          4399 => x"74802ea3",
          4400 => x"38745281",
          4401 => x"bcb051ff",
          4402 => x"ae893f81",
          4403 => x"cbd40893",
          4404 => x"3881ff75",
          4405 => x"27883876",
          4406 => x"89268838",
          4407 => x"8b398a77",
          4408 => x"27863886",
          4409 => x"5581ec39",
          4410 => x"81ff7527",
          4411 => x"8f387488",
          4412 => x"2a547378",
          4413 => x"7081055a",
          4414 => x"34811757",
          4415 => x"74787081",
          4416 => x"055a3481",
          4417 => x"176d7033",
          4418 => x"7081ff06",
          4419 => x"52575557",
          4420 => x"739f26fe",
          4421 => x"c8388b3d",
          4422 => x"33548655",
          4423 => x"7381e52e",
          4424 => x"81b13876",
          4425 => x"802e9938",
          4426 => x"02a70555",
          4427 => x"76157033",
          4428 => x"515473a0",
          4429 => x"2e098106",
          4430 => x"8738ff17",
          4431 => x"5776ed38",
          4432 => x"79418043",
          4433 => x"8052913d",
          4434 => x"705255ff",
          4435 => x"bab33f81",
          4436 => x"cbd40854",
          4437 => x"81cbd408",
          4438 => x"80f73881",
          4439 => x"527451ff",
          4440 => x"bfe53f81",
          4441 => x"cbd40854",
          4442 => x"81cbd408",
          4443 => x"8d387680",
          4444 => x"c4386754",
          4445 => x"e5743480",
          4446 => x"c63981cb",
          4447 => x"d408842e",
          4448 => x"09810680",
          4449 => x"cc388054",
          4450 => x"76742e80",
          4451 => x"c4388152",
          4452 => x"7451ffbd",
          4453 => x"b03f81cb",
          4454 => x"d4085481",
          4455 => x"cbd408b1",
          4456 => x"38a05381",
          4457 => x"cbd40852",
          4458 => x"6751ffab",
          4459 => x"db3f6754",
          4460 => x"880b8b15",
          4461 => x"348b5378",
          4462 => x"526751ff",
          4463 => x"aba73f79",
          4464 => x"54810b83",
          4465 => x"15347951",
          4466 => x"ffadee3f",
          4467 => x"81cbd408",
          4468 => x"54735574",
          4469 => x"81cbd40c",
          4470 => x"9c3d0d04",
          4471 => x"f23d0d60",
          4472 => x"62028805",
          4473 => x"80cb0533",
          4474 => x"933dfc05",
          4475 => x"55725440",
          4476 => x"5e5ad2da",
          4477 => x"3f81cbd4",
          4478 => x"085881cb",
          4479 => x"d40882bd",
          4480 => x"38911a33",
          4481 => x"587782b5",
          4482 => x"387c802e",
          4483 => x"97388c1a",
          4484 => x"08597890",
          4485 => x"38901a33",
          4486 => x"70812a70",
          4487 => x"81065155",
          4488 => x"55739038",
          4489 => x"87548297",
          4490 => x"39825882",
          4491 => x"90398158",
          4492 => x"828b397e",
          4493 => x"8a112270",
          4494 => x"892b7055",
          4495 => x"7f545656",
          4496 => x"56ff828a",
          4497 => x"3fff147d",
          4498 => x"06703070",
          4499 => x"72079f2a",
          4500 => x"81cbd408",
          4501 => x"058c1908",
          4502 => x"7c405a5d",
          4503 => x"55558177",
          4504 => x"27883898",
          4505 => x"16087726",
          4506 => x"83388257",
          4507 => x"76775659",
          4508 => x"80567452",
          4509 => x"7951ffae",
          4510 => x"993f8115",
          4511 => x"7f555598",
          4512 => x"14087526",
          4513 => x"83388255",
          4514 => x"81cbd408",
          4515 => x"812eff99",
          4516 => x"3881cbd4",
          4517 => x"08ff2eff",
          4518 => x"953881cb",
          4519 => x"d4088e38",
          4520 => x"81165675",
          4521 => x"7b2e0981",
          4522 => x"06873893",
          4523 => x"39745980",
          4524 => x"5674772e",
          4525 => x"098106ff",
          4526 => x"b9388758",
          4527 => x"80ff397d",
          4528 => x"802eba38",
          4529 => x"787b5555",
          4530 => x"7a802eb4",
          4531 => x"38811556",
          4532 => x"73812e09",
          4533 => x"81068338",
          4534 => x"ff567553",
          4535 => x"74527e51",
          4536 => x"ffafa83f",
          4537 => x"81cbd408",
          4538 => x"5881cbd4",
          4539 => x"0880ce38",
          4540 => x"748116ff",
          4541 => x"1656565c",
          4542 => x"73d33884",
          4543 => x"39ff195c",
          4544 => x"7e7c8c12",
          4545 => x"0c557d80",
          4546 => x"2eb33878",
          4547 => x"881b0c7c",
          4548 => x"8c1b0c90",
          4549 => x"1a3380c0",
          4550 => x"07547390",
          4551 => x"1b349815",
          4552 => x"08fe0590",
          4553 => x"16085754",
          4554 => x"75742691",
          4555 => x"38757b31",
          4556 => x"90160c84",
          4557 => x"15338107",
          4558 => x"54738416",
          4559 => x"34775473",
          4560 => x"81cbd40c",
          4561 => x"903d0d04",
          4562 => x"e93d0d6b",
          4563 => x"6d028805",
          4564 => x"80eb0533",
          4565 => x"9d3d545a",
          4566 => x"5c59c5bd",
          4567 => x"3f8b5680",
          4568 => x"0b81cbd4",
          4569 => x"08248bf8",
          4570 => x"3881cbd4",
          4571 => x"08842981",
          4572 => x"cbf00570",
          4573 => x"08515574",
          4574 => x"802e8438",
          4575 => x"80753481",
          4576 => x"cbd40881",
          4577 => x"ff065f81",
          4578 => x"527e51ff",
          4579 => x"a0d03f81",
          4580 => x"cbd40881",
          4581 => x"ff067081",
          4582 => x"06565783",
          4583 => x"56748bc0",
          4584 => x"3876822a",
          4585 => x"70810651",
          4586 => x"558a5674",
          4587 => x"8bb23899",
          4588 => x"3dfc0553",
          4589 => x"83527e51",
          4590 => x"ffa4f03f",
          4591 => x"81cbd408",
          4592 => x"99386755",
          4593 => x"74802e92",
          4594 => x"38748280",
          4595 => x"80268b38",
          4596 => x"ff157506",
          4597 => x"5574802e",
          4598 => x"83388148",
          4599 => x"78802e87",
          4600 => x"38848079",
          4601 => x"26923878",
          4602 => x"81800a26",
          4603 => x"8b38ff19",
          4604 => x"79065574",
          4605 => x"802e8638",
          4606 => x"93568ae4",
          4607 => x"3978892a",
          4608 => x"6e892a70",
          4609 => x"892b7759",
          4610 => x"4843597a",
          4611 => x"83388156",
          4612 => x"61307080",
          4613 => x"25770751",
          4614 => x"55915674",
          4615 => x"8ac23899",
          4616 => x"3df80553",
          4617 => x"81527e51",
          4618 => x"ffa4803f",
          4619 => x"815681cb",
          4620 => x"d4088aac",
          4621 => x"3877832a",
          4622 => x"70770681",
          4623 => x"cbd40843",
          4624 => x"56457483",
          4625 => x"38bf4166",
          4626 => x"558e5660",
          4627 => x"75268a90",
          4628 => x"38746131",
          4629 => x"70485580",
          4630 => x"ff75278a",
          4631 => x"83389356",
          4632 => x"78818026",
          4633 => x"89fa3877",
          4634 => x"812a7081",
          4635 => x"06564374",
          4636 => x"802e9538",
          4637 => x"77870655",
          4638 => x"74822e83",
          4639 => x"8d387781",
          4640 => x"06557480",
          4641 => x"2e838338",
          4642 => x"77810655",
          4643 => x"9356825e",
          4644 => x"74802e89",
          4645 => x"cb38785a",
          4646 => x"7d832e09",
          4647 => x"810680e1",
          4648 => x"3878ae38",
          4649 => x"66912a57",
          4650 => x"810b81bc",
          4651 => x"d422565a",
          4652 => x"74802e9d",
          4653 => x"38747726",
          4654 => x"983881bc",
          4655 => x"d4567910",
          4656 => x"82177022",
          4657 => x"57575a74",
          4658 => x"802e8638",
          4659 => x"767527ee",
          4660 => x"38795266",
          4661 => x"51fefcf6",
          4662 => x"3f81cbd4",
          4663 => x"08842984",
          4664 => x"87057089",
          4665 => x"2a5e55a0",
          4666 => x"5c800b81",
          4667 => x"cbd408fc",
          4668 => x"808a0556",
          4669 => x"44fdfff0",
          4670 => x"0a752780",
          4671 => x"ec3888d3",
          4672 => x"3978ae38",
          4673 => x"668c2a57",
          4674 => x"810b81bc",
          4675 => x"c422565a",
          4676 => x"74802e9d",
          4677 => x"38747726",
          4678 => x"983881bc",
          4679 => x"c4567910",
          4680 => x"82177022",
          4681 => x"57575a74",
          4682 => x"802e8638",
          4683 => x"767527ee",
          4684 => x"38795266",
          4685 => x"51fefc96",
          4686 => x"3f81cbd4",
          4687 => x"08108405",
          4688 => x"5781cbd4",
          4689 => x"089ff526",
          4690 => x"9638810b",
          4691 => x"81cbd408",
          4692 => x"1081cbd4",
          4693 => x"08057111",
          4694 => x"722a8305",
          4695 => x"59565e83",
          4696 => x"ff17892a",
          4697 => x"5d815ca0",
          4698 => x"44601c7d",
          4699 => x"11650569",
          4700 => x"7012ff05",
          4701 => x"71307072",
          4702 => x"0674315c",
          4703 => x"52595759",
          4704 => x"407d832e",
          4705 => x"09810689",
          4706 => x"38761c60",
          4707 => x"18415c84",
          4708 => x"39761d5d",
          4709 => x"79902918",
          4710 => x"70623168",
          4711 => x"58515574",
          4712 => x"762687af",
          4713 => x"38757c31",
          4714 => x"7d317a53",
          4715 => x"70653152",
          4716 => x"55fefb9a",
          4717 => x"3f81cbd4",
          4718 => x"08587d83",
          4719 => x"2e098106",
          4720 => x"9b3881cb",
          4721 => x"d40883ff",
          4722 => x"f52680dd",
          4723 => x"38788783",
          4724 => x"3879812a",
          4725 => x"5978fdbe",
          4726 => x"3886f839",
          4727 => x"7d822e09",
          4728 => x"810680c5",
          4729 => x"3883fff5",
          4730 => x"0b81cbd4",
          4731 => x"0827a038",
          4732 => x"788f3879",
          4733 => x"1a557480",
          4734 => x"c0268638",
          4735 => x"7459fd96",
          4736 => x"39628106",
          4737 => x"5574802e",
          4738 => x"8f38835e",
          4739 => x"fd883981",
          4740 => x"cbd4089f",
          4741 => x"f5269238",
          4742 => x"7886b838",
          4743 => x"791a5981",
          4744 => x"807927fc",
          4745 => x"f13886ab",
          4746 => x"3980557d",
          4747 => x"812e0981",
          4748 => x"0683387d",
          4749 => x"559ff578",
          4750 => x"278b3874",
          4751 => x"8106558e",
          4752 => x"5674869c",
          4753 => x"38848053",
          4754 => x"80527a51",
          4755 => x"ffa2b93f",
          4756 => x"8b5381ba",
          4757 => x"ec527a51",
          4758 => x"ffa28a3f",
          4759 => x"8480528b",
          4760 => x"1b51ffa1",
          4761 => x"b33f798d",
          4762 => x"1c347b83",
          4763 => x"ffff0652",
          4764 => x"8e1b51ff",
          4765 => x"a1a23f81",
          4766 => x"0b901c34",
          4767 => x"7d833270",
          4768 => x"3070962a",
          4769 => x"84800654",
          4770 => x"5155911b",
          4771 => x"51ffa188",
          4772 => x"3f665574",
          4773 => x"83ffff26",
          4774 => x"90387483",
          4775 => x"ffff0652",
          4776 => x"931b51ff",
          4777 => x"a0f23f8a",
          4778 => x"397452a0",
          4779 => x"1b51ffa1",
          4780 => x"853ff80b",
          4781 => x"951c34bf",
          4782 => x"52981b51",
          4783 => x"ffa0d93f",
          4784 => x"81ff529a",
          4785 => x"1b51ffa0",
          4786 => x"cf3f6052",
          4787 => x"9c1b51ff",
          4788 => x"a0e43f7d",
          4789 => x"832e0981",
          4790 => x"0680cb38",
          4791 => x"8288b20a",
          4792 => x"5280c31b",
          4793 => x"51ffa0ce",
          4794 => x"3f7c52a4",
          4795 => x"1b51ffa0",
          4796 => x"c53f8252",
          4797 => x"ac1b51ff",
          4798 => x"a0bc3f81",
          4799 => x"52b01b51",
          4800 => x"ffa0953f",
          4801 => x"8652b21b",
          4802 => x"51ffa08c",
          4803 => x"3fff800b",
          4804 => x"80c01c34",
          4805 => x"a90b80c2",
          4806 => x"1c349353",
          4807 => x"81baf852",
          4808 => x"80c71b51",
          4809 => x"ae398288",
          4810 => x"b20a52a7",
          4811 => x"1b51ffa0",
          4812 => x"853f7c83",
          4813 => x"ffff0652",
          4814 => x"961b51ff",
          4815 => x"9fda3fff",
          4816 => x"800ba41c",
          4817 => x"34a90ba6",
          4818 => x"1c349353",
          4819 => x"81bb8c52",
          4820 => x"ab1b51ff",
          4821 => x"a08f3f82",
          4822 => x"d4d55283",
          4823 => x"fe1b7052",
          4824 => x"59ff9fb4",
          4825 => x"3f815460",
          4826 => x"537a527e",
          4827 => x"51ff9bd7",
          4828 => x"3f815681",
          4829 => x"cbd40883",
          4830 => x"e7387d83",
          4831 => x"2e098106",
          4832 => x"80ee3875",
          4833 => x"54608605",
          4834 => x"537a527e",
          4835 => x"51ff9bb7",
          4836 => x"3f848053",
          4837 => x"80527a51",
          4838 => x"ff9fed3f",
          4839 => x"848b85a4",
          4840 => x"d2527a51",
          4841 => x"ff9f8f3f",
          4842 => x"868a85e4",
          4843 => x"f25283e4",
          4844 => x"1b51ff9f",
          4845 => x"813fff18",
          4846 => x"5283e81b",
          4847 => x"51ff9ef6",
          4848 => x"3f825283",
          4849 => x"ec1b51ff",
          4850 => x"9eec3f82",
          4851 => x"d4d55278",
          4852 => x"51ff9ec4",
          4853 => x"3f755460",
          4854 => x"8705537a",
          4855 => x"527e51ff",
          4856 => x"9ae53f75",
          4857 => x"54601653",
          4858 => x"7a527e51",
          4859 => x"ff9ad83f",
          4860 => x"65538052",
          4861 => x"7a51ff9f",
          4862 => x"8f3f7f56",
          4863 => x"80587d83",
          4864 => x"2e098106",
          4865 => x"9a38f852",
          4866 => x"7a51ff9e",
          4867 => x"a93fff52",
          4868 => x"841b51ff",
          4869 => x"9ea03ff0",
          4870 => x"0a52881b",
          4871 => x"51913987",
          4872 => x"fffff855",
          4873 => x"7d812e83",
          4874 => x"38f85574",
          4875 => x"527a51ff",
          4876 => x"9e843f7c",
          4877 => x"55615774",
          4878 => x"62268338",
          4879 => x"74577654",
          4880 => x"75537a52",
          4881 => x"7e51ff99",
          4882 => x"fe3f81cb",
          4883 => x"d4088287",
          4884 => x"38848053",
          4885 => x"81cbd408",
          4886 => x"527a51ff",
          4887 => x"9eaa3f76",
          4888 => x"16757831",
          4889 => x"565674cd",
          4890 => x"38811858",
          4891 => x"77802eff",
          4892 => x"8d387955",
          4893 => x"7d832e83",
          4894 => x"38635561",
          4895 => x"57746226",
          4896 => x"83387457",
          4897 => x"76547553",
          4898 => x"7a527e51",
          4899 => x"ff99b83f",
          4900 => x"81cbd408",
          4901 => x"81c13876",
          4902 => x"16757831",
          4903 => x"565674db",
          4904 => x"388c567d",
          4905 => x"832e9338",
          4906 => x"86566683",
          4907 => x"ffff268a",
          4908 => x"3884567d",
          4909 => x"822e8338",
          4910 => x"81566481",
          4911 => x"06587780",
          4912 => x"fe388480",
          4913 => x"5377527a",
          4914 => x"51ff9dbc",
          4915 => x"3f82d4d5",
          4916 => x"527851ff",
          4917 => x"9cc23f83",
          4918 => x"be1b5577",
          4919 => x"7534810b",
          4920 => x"81163481",
          4921 => x"0b821634",
          4922 => x"77831634",
          4923 => x"75841634",
          4924 => x"60670556",
          4925 => x"80fdc152",
          4926 => x"7551fef4",
          4927 => x"d13ffe0b",
          4928 => x"85163481",
          4929 => x"cbd40882",
          4930 => x"2abf0756",
          4931 => x"75861634",
          4932 => x"81cbd408",
          4933 => x"87163460",
          4934 => x"5283c61b",
          4935 => x"51ff9c96",
          4936 => x"3f665283",
          4937 => x"ca1b51ff",
          4938 => x"9c8c3f81",
          4939 => x"5477537a",
          4940 => x"527e51ff",
          4941 => x"98913f81",
          4942 => x"5681cbd4",
          4943 => x"08a23880",
          4944 => x"5380527e",
          4945 => x"51ff99e3",
          4946 => x"3f815681",
          4947 => x"cbd40890",
          4948 => x"3889398e",
          4949 => x"568a3981",
          4950 => x"56863981",
          4951 => x"cbd40856",
          4952 => x"7581cbd4",
          4953 => x"0c993d0d",
          4954 => x"04ff3d0d",
          4955 => x"73527193",
          4956 => x"26818e38",
          4957 => x"71842981",
          4958 => x"b5b80552",
          4959 => x"71080481",
          4960 => x"bdec5181",
          4961 => x"803981bd",
          4962 => x"f85180f9",
          4963 => x"3981be8c",
          4964 => x"5180f239",
          4965 => x"81bea051",
          4966 => x"80eb3981",
          4967 => x"beb05180",
          4968 => x"e43981be",
          4969 => x"c05180dd",
          4970 => x"3981bed4",
          4971 => x"5180d639",
          4972 => x"81bee451",
          4973 => x"80cf3981",
          4974 => x"befc5180",
          4975 => x"c83981bf",
          4976 => x"945180c1",
          4977 => x"3981bfac",
          4978 => x"51bb3981",
          4979 => x"bfc851b5",
          4980 => x"3981bfdc",
          4981 => x"51af3981",
          4982 => x"c08851a9",
          4983 => x"3981c09c",
          4984 => x"51a33981",
          4985 => x"c0bc519d",
          4986 => x"3981c0d0",
          4987 => x"51973981",
          4988 => x"c0e85191",
          4989 => x"3981c180",
          4990 => x"518b3981",
          4991 => x"c1985185",
          4992 => x"3981c1a4",
          4993 => x"51ff87fb",
          4994 => x"3f833d0d",
          4995 => x"04fb3d0d",
          4996 => x"77795656",
          4997 => x"7487e726",
          4998 => x"8a387452",
          4999 => x"7587e829",
          5000 => x"51913987",
          5001 => x"e8527451",
          5002 => x"fef2a33f",
          5003 => x"81cbd408",
          5004 => x"527551fe",
          5005 => x"f2983f81",
          5006 => x"cbd40854",
          5007 => x"79537552",
          5008 => x"81c1b451",
          5009 => x"ff8da03f",
          5010 => x"873d0d04",
          5011 => x"f53d0d7d",
          5012 => x"7f61028c",
          5013 => x"0580c705",
          5014 => x"33737315",
          5015 => x"665f5d5a",
          5016 => x"5a5c5c5c",
          5017 => x"785281c1",
          5018 => x"d851ff8c",
          5019 => x"fa3f81c1",
          5020 => x"e051ff87",
          5021 => x"8e3f8055",
          5022 => x"74772780",
          5023 => x"fc387990",
          5024 => x"2e893879",
          5025 => x"a02ea738",
          5026 => x"80c63974",
          5027 => x"16537278",
          5028 => x"278e3872",
          5029 => x"225281c1",
          5030 => x"e451ff8c",
          5031 => x"ca3f8939",
          5032 => x"81c1f051",
          5033 => x"ff86dc3f",
          5034 => x"82155580",
          5035 => x"c3397416",
          5036 => x"53727827",
          5037 => x"8e387208",
          5038 => x"5281c1d8",
          5039 => x"51ff8ca7",
          5040 => x"3f893981",
          5041 => x"c1ec51ff",
          5042 => x"86b93f84",
          5043 => x"1555a139",
          5044 => x"74165372",
          5045 => x"78278e38",
          5046 => x"72335281",
          5047 => x"c1f851ff",
          5048 => x"8c853f89",
          5049 => x"3981c280",
          5050 => x"51ff8697",
          5051 => x"3f811555",
          5052 => x"a051fefa",
          5053 => x"8d3fff80",
          5054 => x"3981c284",
          5055 => x"51ff8683",
          5056 => x"3f805574",
          5057 => x"7727aa38",
          5058 => x"74167033",
          5059 => x"79722652",
          5060 => x"55539f74",
          5061 => x"27903872",
          5062 => x"802e8b38",
          5063 => x"7380fe26",
          5064 => x"85387351",
          5065 => x"8339a051",
          5066 => x"fef9d73f",
          5067 => x"811555d3",
          5068 => x"3981c288",
          5069 => x"51ff85cb",
          5070 => x"3f761677",
          5071 => x"1a5a56fe",
          5072 => x"fd923f81",
          5073 => x"cbd40898",
          5074 => x"2b70982c",
          5075 => x"515574a0",
          5076 => x"2e098106",
          5077 => x"a538fefc",
          5078 => x"fb3f81cb",
          5079 => x"d408982b",
          5080 => x"70982c70",
          5081 => x"a0327030",
          5082 => x"7072079f",
          5083 => x"2a515656",
          5084 => x"5155749b",
          5085 => x"2e8c3872",
          5086 => x"dd38749b",
          5087 => x"2e098106",
          5088 => x"85388053",
          5089 => x"8c397a1c",
          5090 => x"53727626",
          5091 => x"fdd638ff",
          5092 => x"537281cb",
          5093 => x"d40c8d3d",
          5094 => x"0d04ec3d",
          5095 => x"0d660284",
          5096 => x"0580e305",
          5097 => x"33697230",
          5098 => x"70740780",
          5099 => x"257087ff",
          5100 => x"74270751",
          5101 => x"51585a5b",
          5102 => x"56935774",
          5103 => x"80fb3881",
          5104 => x"5375528c",
          5105 => x"3d705257",
          5106 => x"c0b93f81",
          5107 => x"cbd40856",
          5108 => x"81cbd408",
          5109 => x"b83881cb",
          5110 => x"d40887c0",
          5111 => x"98880c81",
          5112 => x"cbd40859",
          5113 => x"963dd405",
          5114 => x"54848053",
          5115 => x"77527651",
          5116 => x"c4f63f81",
          5117 => x"cbd40856",
          5118 => x"81cbd408",
          5119 => x"90387a55",
          5120 => x"74802e89",
          5121 => x"38741975",
          5122 => x"195959d8",
          5123 => x"39963dd8",
          5124 => x"0551cce0",
          5125 => x"3f753070",
          5126 => x"77078025",
          5127 => x"51557980",
          5128 => x"2e953874",
          5129 => x"802e9038",
          5130 => x"81c28c53",
          5131 => x"87c09888",
          5132 => x"08527851",
          5133 => x"fbd73f75",
          5134 => x"577681cb",
          5135 => x"d40c963d",
          5136 => x"0d04f93d",
          5137 => x"0d7b0284",
          5138 => x"05b30533",
          5139 => x"5758ff57",
          5140 => x"80537a52",
          5141 => x"7951fec2",
          5142 => x"3f81cbd4",
          5143 => x"08a43875",
          5144 => x"802e8838",
          5145 => x"75812e98",
          5146 => x"38983960",
          5147 => x"557f5481",
          5148 => x"cbd4537e",
          5149 => x"527d5177",
          5150 => x"2d81cbd4",
          5151 => x"08578339",
          5152 => x"77047681",
          5153 => x"cbd40c89",
          5154 => x"3d0d04fc",
          5155 => x"3d0d029b",
          5156 => x"053381c2",
          5157 => x"945381c2",
          5158 => x"9c5255ff",
          5159 => x"88c93f81",
          5160 => x"c8e42251",
          5161 => x"ff80e23f",
          5162 => x"81c2a854",
          5163 => x"81c2b453",
          5164 => x"81c8e533",
          5165 => x"5281c2bc",
          5166 => x"51ff88ab",
          5167 => x"3f74802e",
          5168 => x"8538fefe",
          5169 => x"923f863d",
          5170 => x"0d04fe3d",
          5171 => x"0d87c096",
          5172 => x"800853ff",
          5173 => x"80fd3f81",
          5174 => x"51fef68c",
          5175 => x"3f81c2d8",
          5176 => x"51fef884",
          5177 => x"3f8051fe",
          5178 => x"f5fe3f72",
          5179 => x"812a7081",
          5180 => x"06515271",
          5181 => x"802e9538",
          5182 => x"8151fef5",
          5183 => x"eb3f81c2",
          5184 => x"f451fef7",
          5185 => x"e33f8051",
          5186 => x"fef5dd3f",
          5187 => x"72822a70",
          5188 => x"81065152",
          5189 => x"71802e95",
          5190 => x"388151fe",
          5191 => x"f5ca3f81",
          5192 => x"c38851fe",
          5193 => x"f7c23f80",
          5194 => x"51fef5bc",
          5195 => x"3f72832a",
          5196 => x"70810651",
          5197 => x"5271802e",
          5198 => x"95388151",
          5199 => x"fef5a93f",
          5200 => x"81c39851",
          5201 => x"fef7a13f",
          5202 => x"8051fef5",
          5203 => x"9b3f7284",
          5204 => x"2a708106",
          5205 => x"51527180",
          5206 => x"2e953881",
          5207 => x"51fef588",
          5208 => x"3f81c3ac",
          5209 => x"51fef780",
          5210 => x"3f8051fe",
          5211 => x"f4fa3f72",
          5212 => x"852a7081",
          5213 => x"06515271",
          5214 => x"802e9538",
          5215 => x"8151fef4",
          5216 => x"e73f81c3",
          5217 => x"c051fef6",
          5218 => x"df3f8051",
          5219 => x"fef4d93f",
          5220 => x"72862a70",
          5221 => x"81065152",
          5222 => x"71802e95",
          5223 => x"388151fe",
          5224 => x"f4c63f81",
          5225 => x"c3d451fe",
          5226 => x"f6be3f80",
          5227 => x"51fef4b8",
          5228 => x"3f72872a",
          5229 => x"70810651",
          5230 => x"5271802e",
          5231 => x"95388151",
          5232 => x"fef4a53f",
          5233 => x"81c3e851",
          5234 => x"fef69d3f",
          5235 => x"8051fef4",
          5236 => x"973f7288",
          5237 => x"2a708106",
          5238 => x"51527180",
          5239 => x"2e953881",
          5240 => x"51fef484",
          5241 => x"3f81c3fc",
          5242 => x"51fef5fc",
          5243 => x"3f8051fe",
          5244 => x"f3f63ffe",
          5245 => x"ffa63f84",
          5246 => x"3d0d04fa",
          5247 => x"3d0d7870",
          5248 => x"08705555",
          5249 => x"5773802e",
          5250 => x"80f0388e",
          5251 => x"3973770c",
          5252 => x"85153353",
          5253 => x"80e43981",
          5254 => x"14548074",
          5255 => x"337081ff",
          5256 => x"06575753",
          5257 => x"74a02e83",
          5258 => x"38815374",
          5259 => x"802e8438",
          5260 => x"72e53875",
          5261 => x"81ff0653",
          5262 => x"72a02e09",
          5263 => x"81068838",
          5264 => x"80747081",
          5265 => x"05563480",
          5266 => x"56759029",
          5267 => x"81c98405",
          5268 => x"77085370",
          5269 => x"085255fe",
          5270 => x"edfd3f81",
          5271 => x"cbd4088b",
          5272 => x"38841533",
          5273 => x"5372812e",
          5274 => x"ffa33881",
          5275 => x"167081ff",
          5276 => x"06575394",
          5277 => x"7627d238",
          5278 => x"ff537281",
          5279 => x"cbd40c88",
          5280 => x"3d0d04cb",
          5281 => x"3d0d8070",
          5282 => x"7181e2d4",
          5283 => x"0c5e5c81",
          5284 => x"527b51ff",
          5285 => x"8ac83f81",
          5286 => x"cbd40881",
          5287 => x"ff065978",
          5288 => x"7c2e0981",
          5289 => x"06a23881",
          5290 => x"c4bc5299",
          5291 => x"3d705259",
          5292 => x"ff84ca3f",
          5293 => x"7b537852",
          5294 => x"81cd8451",
          5295 => x"ffb9e33f",
          5296 => x"81cbd408",
          5297 => x"7c2e8838",
          5298 => x"81c4c051",
          5299 => x"8ee83981",
          5300 => x"705e5c81",
          5301 => x"c4f851fe",
          5302 => x"fea93f99",
          5303 => x"3d70465a",
          5304 => x"80f85380",
          5305 => x"527951fe",
          5306 => x"ebdc3f80",
          5307 => x"f8526451",
          5308 => x"ff84ce3f",
          5309 => x"b73dfef8",
          5310 => x"0551fdff",
          5311 => x"3f81cbd4",
          5312 => x"08902b70",
          5313 => x"902c5159",
          5314 => x"7880c32e",
          5315 => x"8a9b3878",
          5316 => x"80c32480",
          5317 => x"dc3878ab",
          5318 => x"2e83bc38",
          5319 => x"78ab24a4",
          5320 => x"3878822e",
          5321 => x"81af3878",
          5322 => x"82248a38",
          5323 => x"78802eff",
          5324 => x"a2388d88",
          5325 => x"3978842e",
          5326 => x"82823878",
          5327 => x"942e82ad",
          5328 => x"388cf939",
          5329 => x"7880c02e",
          5330 => x"858a3878",
          5331 => x"80c02490",
          5332 => x"3878b02e",
          5333 => x"83a93878",
          5334 => x"bc2e848b",
          5335 => x"388cdd39",
          5336 => x"7880c12e",
          5337 => x"86eb3878",
          5338 => x"80c22e88",
          5339 => x"8c388ccc",
          5340 => x"397880f8",
          5341 => x"2e8bba38",
          5342 => x"7880f824",
          5343 => x"a9387880",
          5344 => x"d12e8ae2",
          5345 => x"387880d1",
          5346 => x"248b3878",
          5347 => x"80d02e8a",
          5348 => x"c4388ca8",
          5349 => x"397880d4",
          5350 => x"2e8adc38",
          5351 => x"7880d52e",
          5352 => x"8af2388c",
          5353 => x"97397881",
          5354 => x"832e8bfc",
          5355 => x"38788183",
          5356 => x"24923878",
          5357 => x"80f92e8b",
          5358 => x"9d387881",
          5359 => x"822e8bd9",
          5360 => x"388bf939",
          5361 => x"7881852e",
          5362 => x"8beb3878",
          5363 => x"81872efe",
          5364 => x"82388be8",
          5365 => x"39b73dfe",
          5366 => x"f41153fe",
          5367 => x"f80551ff",
          5368 => x"83fa3f81",
          5369 => x"cbd40888",
          5370 => x"3881c4fc",
          5371 => x"518cc739",
          5372 => x"b73dfef0",
          5373 => x"1153fef8",
          5374 => x"0551ff83",
          5375 => x"df3f81cb",
          5376 => x"d408802e",
          5377 => x"88388163",
          5378 => x"25833880",
          5379 => x"430280cb",
          5380 => x"05335202",
          5381 => x"80cf0533",
          5382 => x"51ff87c2",
          5383 => x"3f81cbd4",
          5384 => x"0881ff06",
          5385 => x"59788e38",
          5386 => x"81c58c51",
          5387 => x"fefbd43f",
          5388 => x"815dfd9f",
          5389 => x"3981c59c",
          5390 => x"5189d239",
          5391 => x"b73dfef4",
          5392 => x"1153fef8",
          5393 => x"0551ff83",
          5394 => x"933f81cb",
          5395 => x"d408802e",
          5396 => x"fd813880",
          5397 => x"53805202",
          5398 => x"80cf0533",
          5399 => x"51ff8bcb",
          5400 => x"3f81cbd4",
          5401 => x"085281c5",
          5402 => x"b4518aa6",
          5403 => x"39b73dfe",
          5404 => x"f41153fe",
          5405 => x"f80551ff",
          5406 => x"82e23f81",
          5407 => x"cbd40880",
          5408 => x"2e873863",
          5409 => x"8926fccb",
          5410 => x"38b73dfe",
          5411 => x"f01153fe",
          5412 => x"f80551ff",
          5413 => x"82c63f81",
          5414 => x"cbd40886",
          5415 => x"3881cbd4",
          5416 => x"08436353",
          5417 => x"81c5bc52",
          5418 => x"7951ff80",
          5419 => x"d03f0280",
          5420 => x"cb053353",
          5421 => x"79526384",
          5422 => x"b42981cd",
          5423 => x"840551ff",
          5424 => x"b5e03f81",
          5425 => x"cbd40881",
          5426 => x"933881c5",
          5427 => x"8c51fefa",
          5428 => x"b23f815c",
          5429 => x"fbfd39b7",
          5430 => x"3dfef805",
          5431 => x"51feeab9",
          5432 => x"3f81cbd4",
          5433 => x"08b83dfe",
          5434 => x"f805525b",
          5435 => x"feeb8c3f",
          5436 => x"815381cb",
          5437 => x"d408527a",
          5438 => x"51f59f3f",
          5439 => x"80d539b7",
          5440 => x"3dfef805",
          5441 => x"51feea91",
          5442 => x"3f81cbd4",
          5443 => x"08b83dfe",
          5444 => x"f805525b",
          5445 => x"feeae43f",
          5446 => x"81cbd408",
          5447 => x"b83dfef8",
          5448 => x"05525afe",
          5449 => x"ead53f81",
          5450 => x"cbd408b8",
          5451 => x"3dfef805",
          5452 => x"5259feea",
          5453 => x"c63f81c8",
          5454 => x"c05881cc",
          5455 => x"88578056",
          5456 => x"805581cb",
          5457 => x"d40881ff",
          5458 => x"06547853",
          5459 => x"79527a51",
          5460 => x"f5f03f81",
          5461 => x"cbd40880",
          5462 => x"2efaf838",
          5463 => x"81cbd408",
          5464 => x"51f0863f",
          5465 => x"faed39b7",
          5466 => x"3dfef411",
          5467 => x"53fef805",
          5468 => x"51ff80e8",
          5469 => x"3f81cbd4",
          5470 => x"08802efa",
          5471 => x"d638b73d",
          5472 => x"fef01153",
          5473 => x"fef80551",
          5474 => x"ff80d13f",
          5475 => x"81cbd408",
          5476 => x"802efabf",
          5477 => x"38b73dfe",
          5478 => x"ec1153fe",
          5479 => x"f80551ff",
          5480 => x"80ba3f81",
          5481 => x"cbd40886",
          5482 => x"3881cbd4",
          5483 => x"084281c5",
          5484 => x"c051fef8",
          5485 => x"ce3f6363",
          5486 => x"5c5a797b",
          5487 => x"278f3861",
          5488 => x"59787a70",
          5489 => x"84055c0c",
          5490 => x"7a7a26f5",
          5491 => x"3881c588",
          5492 => x"5186ba39",
          5493 => x"b73dfef4",
          5494 => x"1153fef8",
          5495 => x"0551feff",
          5496 => x"fb3f81cb",
          5497 => x"d40880c4",
          5498 => x"3881c8ed",
          5499 => x"33597880",
          5500 => x"2e883881",
          5501 => x"c8c00844",
          5502 => x"b33981c8",
          5503 => x"ee335978",
          5504 => x"802e8838",
          5505 => x"81c8c808",
          5506 => x"44a23981",
          5507 => x"c8ef3359",
          5508 => x"788b3881",
          5509 => x"c8f03359",
          5510 => x"78802e88",
          5511 => x"3881c8d0",
          5512 => x"08448939",
          5513 => x"81c8e008",
          5514 => x"fc800544",
          5515 => x"b73dfef0",
          5516 => x"1153fef8",
          5517 => x"0551feff",
          5518 => x"a33f81cb",
          5519 => x"d40880c3",
          5520 => x"3881c8ed",
          5521 => x"33597880",
          5522 => x"2e883881",
          5523 => x"c8c40843",
          5524 => x"b23981c8",
          5525 => x"ee335978",
          5526 => x"802e8838",
          5527 => x"81c8cc08",
          5528 => x"43a13981",
          5529 => x"c8ef3359",
          5530 => x"788b3881",
          5531 => x"c8f03359",
          5532 => x"78802e88",
          5533 => x"3881c8d4",
          5534 => x"08438839",
          5535 => x"81c8e008",
          5536 => x"880543b7",
          5537 => x"3dfeec11",
          5538 => x"53fef805",
          5539 => x"51fefecc",
          5540 => x"3f81cbd4",
          5541 => x"08802e9b",
          5542 => x"3880625b",
          5543 => x"5979882e",
          5544 => x"83388159",
          5545 => x"79902e8d",
          5546 => x"3878802e",
          5547 => x"883879a0",
          5548 => x"2e833888",
          5549 => x"4281c5cc",
          5550 => x"51fef6c7",
          5551 => x"3fa05563",
          5552 => x"54615362",
          5553 => x"526351ef",
          5554 => x"833f81c5",
          5555 => x"dc5184bd",
          5556 => x"39b73dfe",
          5557 => x"f41153fe",
          5558 => x"f80551fe",
          5559 => x"fdfe3f81",
          5560 => x"cbd40880",
          5561 => x"2ef7ec38",
          5562 => x"b73dfef0",
          5563 => x"1153fef8",
          5564 => x"0551fefd",
          5565 => x"e73f81cb",
          5566 => x"d408802e",
          5567 => x"a5386359",
          5568 => x"0280cb05",
          5569 => x"33793463",
          5570 => x"810544b7",
          5571 => x"3dfef011",
          5572 => x"53fef805",
          5573 => x"51fefdc4",
          5574 => x"3f81cbd4",
          5575 => x"08e038f7",
          5576 => x"b2396370",
          5577 => x"33545281",
          5578 => x"c5e851fe",
          5579 => x"fbb93f80",
          5580 => x"f8527951",
          5581 => x"fefc8a3f",
          5582 => x"79457933",
          5583 => x"5978ae2e",
          5584 => x"f791389f",
          5585 => x"7927a038",
          5586 => x"b73dfef0",
          5587 => x"1153fef8",
          5588 => x"0551fefd",
          5589 => x"873f81cb",
          5590 => x"d408802e",
          5591 => x"91386359",
          5592 => x"0280cb05",
          5593 => x"33793463",
          5594 => x"810544ff",
          5595 => x"b53981c5",
          5596 => x"f451fef5",
          5597 => x"8e3fffaa",
          5598 => x"39b73dfe",
          5599 => x"e81153fe",
          5600 => x"f80551fe",
          5601 => x"fec83f81",
          5602 => x"cbd40880",
          5603 => x"2ef6c438",
          5604 => x"b73dfee4",
          5605 => x"1153fef8",
          5606 => x"0551fefe",
          5607 => x"b13f81cb",
          5608 => x"d408802e",
          5609 => x"a6386059",
          5610 => x"02be0522",
          5611 => x"79708205",
          5612 => x"5b237841",
          5613 => x"b73dfee4",
          5614 => x"1153fef8",
          5615 => x"0551fefe",
          5616 => x"8d3f81cb",
          5617 => x"d408df38",
          5618 => x"f6893960",
          5619 => x"70225452",
          5620 => x"81c5fc51",
          5621 => x"fefa903f",
          5622 => x"80f85279",
          5623 => x"51fefae1",
          5624 => x"3f794579",
          5625 => x"335978ae",
          5626 => x"2ef5e838",
          5627 => x"789f2687",
          5628 => x"38608405",
          5629 => x"41d539b7",
          5630 => x"3dfee411",
          5631 => x"53fef805",
          5632 => x"51fefdca",
          5633 => x"3f81cbd4",
          5634 => x"08802e92",
          5635 => x"38605902",
          5636 => x"be052279",
          5637 => x"7082055b",
          5638 => x"237841ff",
          5639 => x"ae3981c5",
          5640 => x"f451fef3",
          5641 => x"de3fffa3",
          5642 => x"39b73dfe",
          5643 => x"e81153fe",
          5644 => x"f80551fe",
          5645 => x"fd983f81",
          5646 => x"cbd40880",
          5647 => x"2ef59438",
          5648 => x"b73dfee4",
          5649 => x"1153fef8",
          5650 => x"0551fefd",
          5651 => x"813f81cb",
          5652 => x"d408802e",
          5653 => x"a1386060",
          5654 => x"710c5960",
          5655 => x"840541b7",
          5656 => x"3dfee411",
          5657 => x"53fef805",
          5658 => x"51fefce2",
          5659 => x"3f81cbd4",
          5660 => x"08e438f4",
          5661 => x"de396070",
          5662 => x"08545281",
          5663 => x"c68851fe",
          5664 => x"f8e53f80",
          5665 => x"f8527951",
          5666 => x"fef9b63f",
          5667 => x"79457933",
          5668 => x"5978ae2e",
          5669 => x"f4bd389f",
          5670 => x"7927a838",
          5671 => x"b73dfee4",
          5672 => x"1153fef8",
          5673 => x"0551fefc",
          5674 => x"a53f81cb",
          5675 => x"d408802e",
          5676 => x"99387f53",
          5677 => x"605281c6",
          5678 => x"8851fef8",
          5679 => x"aa3f6060",
          5680 => x"710c5960",
          5681 => x"840541ff",
          5682 => x"ad3981c5",
          5683 => x"f451fef2",
          5684 => x"b23fffa2",
          5685 => x"3981c694",
          5686 => x"51fef2a7",
          5687 => x"3f8251fe",
          5688 => x"f1953ff3",
          5689 => x"ee3981c6",
          5690 => x"ac51fef2",
          5691 => x"963fa251",
          5692 => x"fef0e83f",
          5693 => x"f3dd3984",
          5694 => x"80810b87",
          5695 => x"c094840c",
          5696 => x"8480810b",
          5697 => x"87c09494",
          5698 => x"0c81c6c4",
          5699 => x"51fef1f3",
          5700 => x"3ff3c039",
          5701 => x"81c6d851",
          5702 => x"fef1e83f",
          5703 => x"8c80830b",
          5704 => x"87c09484",
          5705 => x"0c8c8083",
          5706 => x"0b87c094",
          5707 => x"940cf3a3",
          5708 => x"39b73dfe",
          5709 => x"f41153fe",
          5710 => x"f80551fe",
          5711 => x"f99e3f81",
          5712 => x"cbd40880",
          5713 => x"2ef38c38",
          5714 => x"635281c6",
          5715 => x"ec51fef7",
          5716 => x"963f6359",
          5717 => x"7804b73d",
          5718 => x"fef41153",
          5719 => x"fef80551",
          5720 => x"fef8f93f",
          5721 => x"81cbd408",
          5722 => x"802ef2e7",
          5723 => x"38635281",
          5724 => x"c78851fe",
          5725 => x"f6f13f63",
          5726 => x"59782d81",
          5727 => x"cbd4085e",
          5728 => x"81cbd408",
          5729 => x"802ef2cb",
          5730 => x"3881cbd4",
          5731 => x"085281c7",
          5732 => x"a451fef6",
          5733 => x"d23ff2bb",
          5734 => x"3981c7c0",
          5735 => x"51fef0e3",
          5736 => x"3ffeccdc",
          5737 => x"3ff2ac39",
          5738 => x"81c7dc51",
          5739 => x"fef0d43f",
          5740 => x"8059ffa0",
          5741 => x"39feec9f",
          5742 => x"3ff29839",
          5743 => x"64703351",
          5744 => x"5978802e",
          5745 => x"f28d387b",
          5746 => x"802e80d2",
          5747 => x"387c802e",
          5748 => x"80cc38b7",
          5749 => x"3dfef805",
          5750 => x"51fee0bd",
          5751 => x"3f81c7f0",
          5752 => x"5681cbd4",
          5753 => x"085581c7",
          5754 => x"f4548053",
          5755 => x"81c7f852",
          5756 => x"a33d7052",
          5757 => x"5afef685",
          5758 => x"3f81c8c0",
          5759 => x"5881cc88",
          5760 => x"57805664",
          5761 => x"81114681",
          5762 => x"05558054",
          5763 => x"81800a53",
          5764 => x"81800a52",
          5765 => x"7951ecaa",
          5766 => x"3f81cbd4",
          5767 => x"085e7c81",
          5768 => x"327c8132",
          5769 => x"0759788a",
          5770 => x"387dff2e",
          5771 => x"098106f1",
          5772 => x"a23881c8",
          5773 => x"8851fef5",
          5774 => x"ae3ff197",
          5775 => x"39803d0d",
          5776 => x"800b81cc",
          5777 => x"88349b90",
          5778 => x"86e40b87",
          5779 => x"c0948c0c",
          5780 => x"9b9086e4",
          5781 => x"0b87c094",
          5782 => x"9c0c8c80",
          5783 => x"830b87c0",
          5784 => x"94840c8c",
          5785 => x"80830b87",
          5786 => x"c094940c",
          5787 => x"98820b81",
          5788 => x"cbe40c9b",
          5789 => x"830b81cb",
          5790 => x"e80cfee7",
          5791 => x"af3ffeed",
          5792 => x"d23f81c8",
          5793 => x"9851fee4",
          5794 => x"df3f81c8",
          5795 => x"a451feee",
          5796 => x"f23f81a1",
          5797 => x"ca51feed",
          5798 => x"b53f8151",
          5799 => x"ebed3fef",
          5800 => x"e23f8004",
          5801 => x"00001125",
          5802 => x"0000112b",
          5803 => x"00001131",
          5804 => x"00001137",
          5805 => x"0000113d",
          5806 => x"00004dfb",
          5807 => x"00004d7f",
          5808 => x"00004d86",
          5809 => x"00004d8d",
          5810 => x"00004d94",
          5811 => x"00004d9b",
          5812 => x"00004da2",
          5813 => x"00004da9",
          5814 => x"00004db0",
          5815 => x"00004db7",
          5816 => x"00004dbe",
          5817 => x"00004dc5",
          5818 => x"00004dcb",
          5819 => x"00004dd1",
          5820 => x"00004dd7",
          5821 => x"00004ddd",
          5822 => x"00004de3",
          5823 => x"00004de9",
          5824 => x"00004def",
          5825 => x"00004df5",
          5826 => x"25642f25",
          5827 => x"642f2564",
          5828 => x"2025643a",
          5829 => x"25643a25",
          5830 => x"642e2564",
          5831 => x"25640a00",
          5832 => x"536f4320",
          5833 => x"436f6e66",
          5834 => x"69677572",
          5835 => x"6174696f",
          5836 => x"6e000000",
          5837 => x"20286672",
          5838 => x"6f6d2053",
          5839 => x"6f432063",
          5840 => x"6f6e6669",
          5841 => x"67290000",
          5842 => x"3a0a4465",
          5843 => x"76696365",
          5844 => x"7320696d",
          5845 => x"706c656d",
          5846 => x"656e7465",
          5847 => x"643a0a00",
          5848 => x"20202020",
          5849 => x"494e534e",
          5850 => x"20425241",
          5851 => x"4d202853",
          5852 => x"74617274",
          5853 => x"3d253038",
          5854 => x"582c2053",
          5855 => x"697a653d",
          5856 => x"25303858",
          5857 => x"292e0a00",
          5858 => x"20202020",
          5859 => x"4252414d",
          5860 => x"20285374",
          5861 => x"6172743d",
          5862 => x"25303858",
          5863 => x"2c205369",
          5864 => x"7a653d25",
          5865 => x"30385829",
          5866 => x"2e0a0000",
          5867 => x"20202020",
          5868 => x"52414d20",
          5869 => x"28537461",
          5870 => x"72743d25",
          5871 => x"3038582c",
          5872 => x"2053697a",
          5873 => x"653d2530",
          5874 => x"3858292e",
          5875 => x"0a000000",
          5876 => x"20202020",
          5877 => x"494f4354",
          5878 => x"4c0a0000",
          5879 => x"20202020",
          5880 => x"5053320a",
          5881 => x"00000000",
          5882 => x"20202020",
          5883 => x"5350490a",
          5884 => x"00000000",
          5885 => x"20202020",
          5886 => x"53442043",
          5887 => x"61726420",
          5888 => x"28446576",
          5889 => x"69636573",
          5890 => x"3d253032",
          5891 => x"58292e0a",
          5892 => x"00000000",
          5893 => x"20202020",
          5894 => x"494e5445",
          5895 => x"52525550",
          5896 => x"5420434f",
          5897 => x"4e54524f",
          5898 => x"4c4c4552",
          5899 => x"0a000000",
          5900 => x"20202020",
          5901 => x"54494d45",
          5902 => x"52312028",
          5903 => x"54696d65",
          5904 => x"72733d25",
          5905 => x"30315829",
          5906 => x"2e0a0000",
          5907 => x"41646472",
          5908 => x"65737365",
          5909 => x"733a0a00",
          5910 => x"20202020",
          5911 => x"43505520",
          5912 => x"52657365",
          5913 => x"74205665",
          5914 => x"63746f72",
          5915 => x"20416464",
          5916 => x"72657373",
          5917 => x"203d2025",
          5918 => x"3038580a",
          5919 => x"00000000",
          5920 => x"20202020",
          5921 => x"43505520",
          5922 => x"4d656d6f",
          5923 => x"72792053",
          5924 => x"74617274",
          5925 => x"20416464",
          5926 => x"72657373",
          5927 => x"203d2025",
          5928 => x"3038580a",
          5929 => x"00000000",
          5930 => x"20202020",
          5931 => x"53746163",
          5932 => x"6b205374",
          5933 => x"61727420",
          5934 => x"41646472",
          5935 => x"65737320",
          5936 => x"20202020",
          5937 => x"203d2025",
          5938 => x"3038580a",
          5939 => x"00000000",
          5940 => x"20202020",
          5941 => x"5a505520",
          5942 => x"49642020",
          5943 => x"20202020",
          5944 => x"20202020",
          5945 => x"20202020",
          5946 => x"20202020",
          5947 => x"203d2025",
          5948 => x"3038580a",
          5949 => x"00000000",
          5950 => x"20202020",
          5951 => x"53797374",
          5952 => x"656d2043",
          5953 => x"6c6f636b",
          5954 => x"20467265",
          5955 => x"71202020",
          5956 => x"20202020",
          5957 => x"203d2025",
          5958 => x"3038580a",
          5959 => x"00000000",
          5960 => x"536d616c",
          5961 => x"6c000000",
          5962 => x"4d656469",
          5963 => x"756d0000",
          5964 => x"466c6578",
          5965 => x"00000000",
          5966 => x"45564f00",
          5967 => x"45564f6d",
          5968 => x"696e0000",
          5969 => x"556e6b6e",
          5970 => x"6f776e00",
          5971 => x"53440000",
          5972 => x"222a2b2c",
          5973 => x"3a3b3c3d",
          5974 => x"3e3f5b5d",
          5975 => x"7c7f0000",
          5976 => x"46415400",
          5977 => x"46415433",
          5978 => x"32000000",
          5979 => x"ebfe904d",
          5980 => x"53444f53",
          5981 => x"352e3000",
          5982 => x"4e4f204e",
          5983 => x"414d4520",
          5984 => x"20202046",
          5985 => x"41543332",
          5986 => x"20202000",
          5987 => x"4e4f204e",
          5988 => x"414d4520",
          5989 => x"20202046",
          5990 => x"41542020",
          5991 => x"20202000",
          5992 => x"00005d4c",
          5993 => x"00000000",
          5994 => x"00000000",
          5995 => x"00000000",
          5996 => x"809a4541",
          5997 => x"8e418f80",
          5998 => x"45454549",
          5999 => x"49498e8f",
          6000 => x"9092924f",
          6001 => x"994f5555",
          6002 => x"59999a9b",
          6003 => x"9c9d9e9f",
          6004 => x"41494f55",
          6005 => x"a5a5a6a7",
          6006 => x"a8a9aaab",
          6007 => x"acadaeaf",
          6008 => x"b0b1b2b3",
          6009 => x"b4b5b6b7",
          6010 => x"b8b9babb",
          6011 => x"bcbdbebf",
          6012 => x"c0c1c2c3",
          6013 => x"c4c5c6c7",
          6014 => x"c8c9cacb",
          6015 => x"cccdcecf",
          6016 => x"d0d1d2d3",
          6017 => x"d4d5d6d7",
          6018 => x"d8d9dadb",
          6019 => x"dcdddedf",
          6020 => x"e0e1e2e3",
          6021 => x"e4e5e6e7",
          6022 => x"e8e9eaeb",
          6023 => x"ecedeeef",
          6024 => x"f0f1f2f3",
          6025 => x"f4f5f6f7",
          6026 => x"f8f9fafb",
          6027 => x"fcfdfeff",
          6028 => x"2b2e2c3b",
          6029 => x"3d5b5d2f",
          6030 => x"5c222a3a",
          6031 => x"3c3e3f7c",
          6032 => x"7f000000",
          6033 => x"00010004",
          6034 => x"00100040",
          6035 => x"01000200",
          6036 => x"00000000",
          6037 => x"00010002",
          6038 => x"00040008",
          6039 => x"00100020",
          6040 => x"00000000",
          6041 => x"64696e69",
          6042 => x"74000000",
          6043 => x"64696f63",
          6044 => x"746c0000",
          6045 => x"66696e69",
          6046 => x"74000000",
          6047 => x"666c6f61",
          6048 => x"64000000",
          6049 => x"66657865",
          6050 => x"63000000",
          6051 => x"6d636c65",
          6052 => x"61720000",
          6053 => x"6d64756d",
          6054 => x"70000000",
          6055 => x"6d746573",
          6056 => x"74000000",
          6057 => x"6d656200",
          6058 => x"6d656800",
          6059 => x"6d657700",
          6060 => x"68696400",
          6061 => x"68696500",
          6062 => x"68666400",
          6063 => x"68666500",
          6064 => x"63616c6c",
          6065 => x"00000000",
          6066 => x"6a6d7000",
          6067 => x"72657374",
          6068 => x"61727400",
          6069 => x"72657365",
          6070 => x"74000000",
          6071 => x"696e666f",
          6072 => x"00000000",
          6073 => x"74657374",
          6074 => x"00000000",
          6075 => x"4469736b",
          6076 => x"20457272",
          6077 => x"6f720a00",
          6078 => x"496e7465",
          6079 => x"726e616c",
          6080 => x"20657272",
          6081 => x"6f722e0a",
          6082 => x"00000000",
          6083 => x"4469736b",
          6084 => x"206e6f74",
          6085 => x"20726561",
          6086 => x"64792e0a",
          6087 => x"00000000",
          6088 => x"4e6f2066",
          6089 => x"696c6520",
          6090 => x"666f756e",
          6091 => x"642e0a00",
          6092 => x"4e6f2070",
          6093 => x"61746820",
          6094 => x"666f756e",
          6095 => x"642e0a00",
          6096 => x"496e7661",
          6097 => x"6c696420",
          6098 => x"66696c65",
          6099 => x"6e616d65",
          6100 => x"2e0a0000",
          6101 => x"41636365",
          6102 => x"73732064",
          6103 => x"656e6965",
          6104 => x"642e0a00",
          6105 => x"46696c65",
          6106 => x"20616c72",
          6107 => x"65616479",
          6108 => x"20657869",
          6109 => x"7374732e",
          6110 => x"0a000000",
          6111 => x"46696c65",
          6112 => x"2068616e",
          6113 => x"646c6520",
          6114 => x"696e7661",
          6115 => x"6c69642e",
          6116 => x"0a000000",
          6117 => x"53442069",
          6118 => x"73207772",
          6119 => x"69746520",
          6120 => x"70726f74",
          6121 => x"65637465",
          6122 => x"642e0a00",
          6123 => x"44726976",
          6124 => x"65206e75",
          6125 => x"6d626572",
          6126 => x"20697320",
          6127 => x"696e7661",
          6128 => x"6c69642e",
          6129 => x"0a000000",
          6130 => x"4469736b",
          6131 => x"206e6f74",
          6132 => x"20656e61",
          6133 => x"626c6564",
          6134 => x"2e0a0000",
          6135 => x"4e6f2063",
          6136 => x"6f6d7061",
          6137 => x"7469626c",
          6138 => x"65206669",
          6139 => x"6c657379",
          6140 => x"7374656d",
          6141 => x"20666f75",
          6142 => x"6e64206f",
          6143 => x"6e206469",
          6144 => x"736b2e0a",
          6145 => x"00000000",
          6146 => x"466f726d",
          6147 => x"61742061",
          6148 => x"626f7274",
          6149 => x"65642e0a",
          6150 => x"00000000",
          6151 => x"54696d65",
          6152 => x"6f75742c",
          6153 => x"206f7065",
          6154 => x"72617469",
          6155 => x"6f6e2063",
          6156 => x"616e6365",
          6157 => x"6c6c6564",
          6158 => x"2e0a0000",
          6159 => x"46696c65",
          6160 => x"20697320",
          6161 => x"6c6f636b",
          6162 => x"65642e0a",
          6163 => x"00000000",
          6164 => x"496e7375",
          6165 => x"66666963",
          6166 => x"69656e74",
          6167 => x"206d656d",
          6168 => x"6f72792e",
          6169 => x"0a000000",
          6170 => x"546f6f20",
          6171 => x"6d616e79",
          6172 => x"206f7065",
          6173 => x"6e206669",
          6174 => x"6c65732e",
          6175 => x"0a000000",
          6176 => x"50617261",
          6177 => x"6d657465",
          6178 => x"72732069",
          6179 => x"6e636f72",
          6180 => x"72656374",
          6181 => x"2e0a0000",
          6182 => x"53756363",
          6183 => x"6573732e",
          6184 => x"0a000000",
          6185 => x"556e6b6e",
          6186 => x"6f776e20",
          6187 => x"6572726f",
          6188 => x"722e0a00",
          6189 => x"0a256c75",
          6190 => x"20627974",
          6191 => x"65732025",
          6192 => x"73206174",
          6193 => x"20256c75",
          6194 => x"20627974",
          6195 => x"65732f73",
          6196 => x"65632e0a",
          6197 => x"00000000",
          6198 => x"25303858",
          6199 => x"00000000",
          6200 => x"3a202000",
          6201 => x"25303458",
          6202 => x"00000000",
          6203 => x"20202020",
          6204 => x"20202020",
          6205 => x"00000000",
          6206 => x"25303258",
          6207 => x"00000000",
          6208 => x"20200000",
          6209 => x"207c0000",
          6210 => x"7c0d0a00",
          6211 => x"72656164",
          6212 => x"00000000",
          6213 => x"5a505554",
          6214 => x"41000000",
          6215 => x"0a2a2a20",
          6216 => x"25732028",
          6217 => x"00000000",
          6218 => x"31382f30",
          6219 => x"372f3230",
          6220 => x"31390000",
          6221 => x"76312e33",
          6222 => x"00000000",
          6223 => x"205a5055",
          6224 => x"2c207265",
          6225 => x"76202530",
          6226 => x"32782920",
          6227 => x"25732025",
          6228 => x"73202a2a",
          6229 => x"0a0a0000",
          6230 => x"5a505554",
          6231 => x"4120496e",
          6232 => x"74657272",
          6233 => x"75707420",
          6234 => x"48616e64",
          6235 => x"6c65720a",
          6236 => x"00000000",
          6237 => x"54696d65",
          6238 => x"7220696e",
          6239 => x"74657272",
          6240 => x"7570740a",
          6241 => x"00000000",
          6242 => x"50533220",
          6243 => x"696e7465",
          6244 => x"72727570",
          6245 => x"740a0000",
          6246 => x"494f4354",
          6247 => x"4c205244",
          6248 => x"20696e74",
          6249 => x"65727275",
          6250 => x"70740a00",
          6251 => x"494f4354",
          6252 => x"4c205752",
          6253 => x"20696e74",
          6254 => x"65727275",
          6255 => x"70740a00",
          6256 => x"55415254",
          6257 => x"30205258",
          6258 => x"20696e74",
          6259 => x"65727275",
          6260 => x"70740a00",
          6261 => x"55415254",
          6262 => x"30205458",
          6263 => x"20696e74",
          6264 => x"65727275",
          6265 => x"70740a00",
          6266 => x"55415254",
          6267 => x"31205258",
          6268 => x"20696e74",
          6269 => x"65727275",
          6270 => x"70740a00",
          6271 => x"55415254",
          6272 => x"31205458",
          6273 => x"20696e74",
          6274 => x"65727275",
          6275 => x"70740a00",
          6276 => x"53657474",
          6277 => x"696e6720",
          6278 => x"75702074",
          6279 => x"696d6572",
          6280 => x"2e2e2e0a",
          6281 => x"00000000",
          6282 => x"456e6162",
          6283 => x"6c696e67",
          6284 => x"2074696d",
          6285 => x"65722e2e",
          6286 => x"2e0a0000",
          6287 => x"303a0000",
          6288 => x"4661696c",
          6289 => x"65642074",
          6290 => x"6f20696e",
          6291 => x"69746961",
          6292 => x"6c697365",
          6293 => x"20736420",
          6294 => x"63617264",
          6295 => x"20302c20",
          6296 => x"706c6561",
          6297 => x"73652069",
          6298 => x"6e697420",
          6299 => x"6d616e75",
          6300 => x"616c6c79",
          6301 => x"2e0a0000",
          6302 => x"2a200000",
          6303 => x"42616420",
          6304 => x"6469736b",
          6305 => x"20696421",
          6306 => x"0a000000",
          6307 => x"496e6974",
          6308 => x"69616c69",
          6309 => x"7365642e",
          6310 => x"0a000000",
          6311 => x"4661696c",
          6312 => x"65642074",
          6313 => x"6f20696e",
          6314 => x"69746961",
          6315 => x"6c697365",
          6316 => x"2e0a0000",
          6317 => x"72633d25",
          6318 => x"640a0000",
          6319 => x"25753a00",
          6320 => x"436c6561",
          6321 => x"72696e67",
          6322 => x"2e2e2e00",
          6323 => x"44756d70",
          6324 => x"204d656d",
          6325 => x"6f72790a",
          6326 => x"00000000",
          6327 => x"0a436f6d",
          6328 => x"706c6574",
          6329 => x"652e0a00",
          6330 => x"25303858",
          6331 => x"20253032",
          6332 => x"582d0000",
          6333 => x"3f3f3f0a",
          6334 => x"00000000",
          6335 => x"25303858",
          6336 => x"20253034",
          6337 => x"582d0000",
          6338 => x"25303858",
          6339 => x"20253038",
          6340 => x"582d0000",
          6341 => x"44697361",
          6342 => x"626c696e",
          6343 => x"6720696e",
          6344 => x"74657272",
          6345 => x"75707473",
          6346 => x"0a000000",
          6347 => x"456e6162",
          6348 => x"6c696e67",
          6349 => x"20696e74",
          6350 => x"65727275",
          6351 => x"7074730a",
          6352 => x"00000000",
          6353 => x"44697361",
          6354 => x"626c6564",
          6355 => x"20756172",
          6356 => x"74206669",
          6357 => x"666f0a00",
          6358 => x"456e6162",
          6359 => x"6c696e67",
          6360 => x"20756172",
          6361 => x"74206669",
          6362 => x"666f0a00",
          6363 => x"45786563",
          6364 => x"7574696e",
          6365 => x"6720636f",
          6366 => x"64652040",
          6367 => x"20253038",
          6368 => x"78202e2e",
          6369 => x"2e0a0000",
          6370 => x"43616c6c",
          6371 => x"696e6720",
          6372 => x"636f6465",
          6373 => x"20402025",
          6374 => x"30387820",
          6375 => x"2e2e2e0a",
          6376 => x"00000000",
          6377 => x"43616c6c",
          6378 => x"20726574",
          6379 => x"75726e65",
          6380 => x"6420636f",
          6381 => x"64652028",
          6382 => x"2564292e",
          6383 => x"0a000000",
          6384 => x"52657374",
          6385 => x"61727469",
          6386 => x"6e672061",
          6387 => x"70706c69",
          6388 => x"63617469",
          6389 => x"6f6e2e2e",
          6390 => x"2e0a0000",
          6391 => x"436f6c64",
          6392 => x"20726562",
          6393 => x"6f6f7469",
          6394 => x"6e672e2e",
          6395 => x"2e0a0000",
          6396 => x"5a505500",
          6397 => x"62696e00",
          6398 => x"25643a5c",
          6399 => x"25735c25",
          6400 => x"732e2573",
          6401 => x"00000000",
          6402 => x"42616420",
          6403 => x"636f6d6d",
          6404 => x"616e642e",
          6405 => x"0a000000",
          6406 => x"52756e6e",
          6407 => x"696e672e",
          6408 => x"2e2e0a00",
          6409 => x"456e6162",
          6410 => x"6c696e67",
          6411 => x"20696e74",
          6412 => x"65727275",
          6413 => x"7074732e",
          6414 => x"2e2e0a00",
          6415 => x"00000000",
          6416 => x"00000000",
          6417 => x"00007fff",
          6418 => x"00000000",
          6419 => x"00007fff",
          6420 => x"00010000",
          6421 => x"00007fff",
          6422 => x"00000000",
          6423 => x"00000000",
          6424 => x"00007800",
          6425 => x"00000000",
          6426 => x"05f5e100",
          6427 => x"00010101",
          6428 => x"01010101",
          6429 => x"80010101",
          6430 => x"01000000",
          6431 => x"00000000",
          6432 => x"01000000",
          6433 => x"00005e64",
          6434 => x"01020100",
          6435 => x"00000000",
          6436 => x"00000000",
          6437 => x"00005e6c",
          6438 => x"01040100",
          6439 => x"00000000",
          6440 => x"00000000",
          6441 => x"00005e74",
          6442 => x"01140300",
          6443 => x"00000000",
          6444 => x"00000000",
          6445 => x"00005e7c",
          6446 => x"012b0300",
          6447 => x"00000000",
          6448 => x"00000000",
          6449 => x"00005e84",
          6450 => x"01300300",
          6451 => x"00000000",
          6452 => x"00000000",
          6453 => x"00005e8c",
          6454 => x"013c0400",
          6455 => x"00000000",
          6456 => x"00000000",
          6457 => x"00005e94",
          6458 => x"01400400",
          6459 => x"00000000",
          6460 => x"00000000",
          6461 => x"00005e9c",
          6462 => x"01440400",
          6463 => x"00000000",
          6464 => x"00000000",
          6465 => x"00005ea4",
          6466 => x"01410400",
          6467 => x"00000000",
          6468 => x"00000000",
          6469 => x"00005ea8",
          6470 => x"01420400",
          6471 => x"00000000",
          6472 => x"00000000",
          6473 => x"00005eac",
          6474 => x"01430400",
          6475 => x"00000000",
          6476 => x"00000000",
          6477 => x"00005eb0",
          6478 => x"01500500",
          6479 => x"00000000",
          6480 => x"00000000",
          6481 => x"00005eb4",
          6482 => x"01510500",
          6483 => x"00000000",
          6484 => x"00000000",
          6485 => x"00005eb8",
          6486 => x"01540500",
          6487 => x"00000000",
          6488 => x"00000000",
          6489 => x"00005ebc",
          6490 => x"01550500",
          6491 => x"00000000",
          6492 => x"00000000",
          6493 => x"00005ec0",
          6494 => x"01790700",
          6495 => x"00000000",
          6496 => x"00000000",
          6497 => x"00005ec8",
          6498 => x"01780700",
          6499 => x"00000000",
          6500 => x"00000000",
          6501 => x"00005ecc",
          6502 => x"01820800",
          6503 => x"00000000",
          6504 => x"00000000",
          6505 => x"00005ed4",
          6506 => x"01830800",
          6507 => x"00000000",
          6508 => x"00000000",
          6509 => x"00005edc",
          6510 => x"01850800",
          6511 => x"00000000",
          6512 => x"00000000",
          6513 => x"00005ee4",
          6514 => x"01870800",
          6515 => x"00000000",
          6516 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;


end arch;

