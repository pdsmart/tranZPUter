-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"88",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"0b",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"88",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"a7",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"9f",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"89",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"8b",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"00",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"53",
           266 => x"00",
           267 => x"06",
           268 => x"09",
           269 => x"05",
           270 => x"2b",
           271 => x"06",
           272 => x"04",
           273 => x"72",
           274 => x"05",
           275 => x"05",
           276 => x"72",
           277 => x"53",
           278 => x"51",
           279 => x"04",
           280 => x"a0",
           281 => x"38",
           282 => x"84",
           283 => x"0b",
           284 => x"e2",
           285 => x"51",
           286 => x"00",
           287 => x"88",
           288 => x"00",
           289 => x"02",
           290 => x"3d",
           291 => x"94",
           292 => x"08",
           293 => x"88",
           294 => x"82",
           295 => x"08",
           296 => x"54",
           297 => x"94",
           298 => x"08",
           299 => x"fd",
           300 => x"53",
           301 => x"05",
           302 => x"08",
           303 => x"51",
           304 => x"88",
           305 => x"0c",
           306 => x"0d",
           307 => x"94",
           308 => x"0c",
           309 => x"80",
           310 => x"fc",
           311 => x"08",
           312 => x"80",
           313 => x"94",
           314 => x"08",
           315 => x"88",
           316 => x"0b",
           317 => x"05",
           318 => x"fc",
           319 => x"38",
           320 => x"08",
           321 => x"94",
           322 => x"08",
           323 => x"05",
           324 => x"8c",
           325 => x"25",
           326 => x"08",
           327 => x"30",
           328 => x"05",
           329 => x"94",
           330 => x"0c",
           331 => x"05",
           332 => x"81",
           333 => x"f0",
           334 => x"08",
           335 => x"94",
           336 => x"0c",
           337 => x"08",
           338 => x"52",
           339 => x"05",
           340 => x"a7",
           341 => x"70",
           342 => x"05",
           343 => x"08",
           344 => x"80",
           345 => x"94",
           346 => x"08",
           347 => x"f8",
           348 => x"08",
           349 => x"70",
           350 => x"89",
           351 => x"0c",
           352 => x"02",
           353 => x"3d",
           354 => x"94",
           355 => x"0c",
           356 => x"05",
           357 => x"93",
           358 => x"88",
           359 => x"94",
           360 => x"0c",
           361 => x"08",
           362 => x"94",
           363 => x"08",
           364 => x"38",
           365 => x"05",
           366 => x"08",
           367 => x"81",
           368 => x"8c",
           369 => x"94",
           370 => x"08",
           371 => x"88",
           372 => x"08",
           373 => x"54",
           374 => x"05",
           375 => x"8c",
           376 => x"f8",
           377 => x"94",
           378 => x"0c",
           379 => x"05",
           380 => x"0c",
           381 => x"0d",
           382 => x"94",
           383 => x"0c",
           384 => x"81",
           385 => x"fc",
           386 => x"0b",
           387 => x"05",
           388 => x"8c",
           389 => x"08",
           390 => x"27",
           391 => x"08",
           392 => x"80",
           393 => x"80",
           394 => x"8c",
           395 => x"99",
           396 => x"8c",
           397 => x"94",
           398 => x"0c",
           399 => x"05",
           400 => x"08",
           401 => x"c9",
           402 => x"fc",
           403 => x"2e",
           404 => x"94",
           405 => x"08",
           406 => x"05",
           407 => x"38",
           408 => x"05",
           409 => x"8c",
           410 => x"94",
           411 => x"0c",
           412 => x"05",
           413 => x"fc",
           414 => x"94",
           415 => x"0c",
           416 => x"05",
           417 => x"94",
           418 => x"0c",
           419 => x"05",
           420 => x"94",
           421 => x"0c",
           422 => x"94",
           423 => x"08",
           424 => x"38",
           425 => x"05",
           426 => x"08",
           427 => x"51",
           428 => x"08",
           429 => x"70",
           430 => x"05",
           431 => x"08",
           432 => x"88",
           433 => x"0d",
           434 => x"ff",
           435 => x"88",
           436 => x"92",
           437 => x"0b",
           438 => x"8c",
           439 => x"87",
           440 => x"0c",
           441 => x"8c",
           442 => x"06",
           443 => x"80",
           444 => x"87",
           445 => x"08",
           446 => x"38",
           447 => x"8c",
           448 => x"80",
           449 => x"93",
           450 => x"98",
           451 => x"70",
           452 => x"38",
           453 => x"0b",
           454 => x"0b",
           455 => x"f0",
           456 => x"83",
           457 => x"fa",
           458 => x"7b",
           459 => x"56",
           460 => x"0b",
           461 => x"33",
           462 => x"55",
           463 => x"75",
           464 => x"06",
           465 => x"85",
           466 => x"98",
           467 => x"87",
           468 => x"0c",
           469 => x"c0",
           470 => x"87",
           471 => x"08",
           472 => x"70",
           473 => x"52",
           474 => x"2e",
           475 => x"c0",
           476 => x"70",
           477 => x"76",
           478 => x"53",
           479 => x"2e",
           480 => x"80",
           481 => x"71",
           482 => x"05",
           483 => x"14",
           484 => x"55",
           485 => x"51",
           486 => x"8b",
           487 => x"98",
           488 => x"70",
           489 => x"87",
           490 => x"08",
           491 => x"38",
           492 => x"c0",
           493 => x"87",
           494 => x"08",
           495 => x"51",
           496 => x"38",
           497 => x"80",
           498 => x"52",
           499 => x"09",
           500 => x"38",
           501 => x"8c",
           502 => x"72",
           503 => x"06",
           504 => x"52",
           505 => x"88",
           506 => x"fe",
           507 => x"81",
           508 => x"33",
           509 => x"07",
           510 => x"51",
           511 => x"04",
           512 => x"75",
           513 => x"82",
           514 => x"90",
           515 => x"2b",
           516 => x"33",
           517 => x"88",
           518 => x"71",
           519 => x"52",
           520 => x"54",
           521 => x"0d",
           522 => x"0d",
           523 => x"0b",
           524 => x"57",
           525 => x"27",
           526 => x"76",
           527 => x"27",
           528 => x"75",
           529 => x"82",
           530 => x"74",
           531 => x"38",
           532 => x"74",
           533 => x"83",
           534 => x"76",
           535 => x"17",
           536 => x"88",
           537 => x"55",
           538 => x"88",
           539 => x"74",
           540 => x"3f",
           541 => x"ff",
           542 => x"ad",
           543 => x"76",
           544 => x"fc",
           545 => x"87",
           546 => x"08",
           547 => x"3d",
           548 => x"fd",
           549 => x"08",
           550 => x"51",
           551 => x"88",
           552 => x"06",
           553 => x"81",
           554 => x"0c",
           555 => x"04",
           556 => x"0b",
           557 => x"f4",
           558 => x"88",
           559 => x"05",
           560 => x"80",
           561 => x"27",
           562 => x"14",
           563 => x"29",
           564 => x"05",
           565 => x"88",
           566 => x"0d",
           567 => x"0d",
           568 => x"0b",
           569 => x"9f",
           570 => x"33",
           571 => x"71",
           572 => x"81",
           573 => x"94",
           574 => x"ef",
           575 => x"90",
           576 => x"14",
           577 => x"3f",
           578 => x"ff",
           579 => x"07",
           580 => x"3d",
           581 => x"3d",
           582 => x"0b",
           583 => x"08",
           584 => x"75",
           585 => x"08",
           586 => x"2e",
           587 => x"14",
           588 => x"85",
           589 => x"b0",
           590 => x"38",
           591 => x"71",
           592 => x"81",
           593 => x"90",
           594 => x"72",
           595 => x"72",
           596 => x"38",
           597 => x"d8",
           598 => x"52",
           599 => x"14",
           600 => x"90",
           601 => x"52",
           602 => x"86",
           603 => x"fa",
           604 => x"0b",
           605 => x"f4",
           606 => x"81",
           607 => x"ff",
           608 => x"54",
           609 => x"80",
           610 => x"90",
           611 => x"72",
           612 => x"52",
           613 => x"73",
           614 => x"71",
           615 => x"81",
           616 => x"0c",
           617 => x"53",
           618 => x"83",
           619 => x"22",
           620 => x"76",
           621 => x"b5",
           622 => x"33",
           623 => x"84",
           624 => x"71",
           625 => x"51",
           626 => x"81",
           627 => x"08",
           628 => x"83",
           629 => x"88",
           630 => x"96",
           631 => x"8c",
           632 => x"08",
           633 => x"3f",
           634 => x"16",
           635 => x"23",
           636 => x"88",
           637 => x"0d",
           638 => x"0d",
           639 => x"58",
           640 => x"33",
           641 => x"2e",
           642 => x"88",
           643 => x"70",
           644 => x"39",
           645 => x"56",
           646 => x"2e",
           647 => x"84",
           648 => x"43",
           649 => x"1d",
           650 => x"33",
           651 => x"9f",
           652 => x"7b",
           653 => x"3f",
           654 => x"80",
           655 => x"d3",
           656 => x"84",
           657 => x"58",
           658 => x"55",
           659 => x"81",
           660 => x"ff",
           661 => x"ff",
           662 => x"06",
           663 => x"70",
           664 => x"7f",
           665 => x"7a",
           666 => x"81",
           667 => x"13",
           668 => x"af",
           669 => x"a0",
           670 => x"80",
           671 => x"51",
           672 => x"5d",
           673 => x"80",
           674 => x"ae",
           675 => x"06",
           676 => x"55",
           677 => x"75",
           678 => x"80",
           679 => x"79",
           680 => x"30",
           681 => x"70",
           682 => x"07",
           683 => x"51",
           684 => x"75",
           685 => x"58",
           686 => x"ab",
           687 => x"19",
           688 => x"06",
           689 => x"5a",
           690 => x"75",
           691 => x"39",
           692 => x"0c",
           693 => x"a0",
           694 => x"81",
           695 => x"1a",
           696 => x"fc",
           697 => x"08",
           698 => x"a0",
           699 => x"70",
           700 => x"e0",
           701 => x"90",
           702 => x"7c",
           703 => x"3f",
           704 => x"88",
           705 => x"38",
           706 => x"74",
           707 => x"ee",
           708 => x"33",
           709 => x"70",
           710 => x"56",
           711 => x"38",
           712 => x"1e",
           713 => x"59",
           714 => x"ff",
           715 => x"ff",
           716 => x"79",
           717 => x"5b",
           718 => x"81",
           719 => x"71",
           720 => x"56",
           721 => x"2e",
           722 => x"39",
           723 => x"92",
           724 => x"fc",
           725 => x"8e",
           726 => x"56",
           727 => x"38",
           728 => x"56",
           729 => x"8b",
           730 => x"55",
           731 => x"8b",
           732 => x"84",
           733 => x"06",
           734 => x"74",
           735 => x"56",
           736 => x"56",
           737 => x"51",
           738 => x"88",
           739 => x"0c",
           740 => x"75",
           741 => x"3d",
           742 => x"3d",
           743 => x"59",
           744 => x"83",
           745 => x"52",
           746 => x"fb",
           747 => x"88",
           748 => x"38",
           749 => x"b3",
           750 => x"83",
           751 => x"55",
           752 => x"82",
           753 => x"09",
           754 => x"ce",
           755 => x"b6",
           756 => x"76",
           757 => x"3f",
           758 => x"88",
           759 => x"76",
           760 => x"3f",
           761 => x"ff",
           762 => x"74",
           763 => x"2e",
           764 => x"54",
           765 => x"77",
           766 => x"f6",
           767 => x"08",
           768 => x"94",
           769 => x"f7",
           770 => x"08",
           771 => x"06",
           772 => x"82",
           773 => x"38",
           774 => x"88",
           775 => x"0d",
           776 => x"0d",
           777 => x"0b",
           778 => x"9f",
           779 => x"9b",
           780 => x"81",
           781 => x"56",
           782 => x"38",
           783 => x"8d",
           784 => x"57",
           785 => x"3f",
           786 => x"ff",
           787 => x"81",
           788 => x"06",
           789 => x"54",
           790 => x"74",
           791 => x"f5",
           792 => x"08",
           793 => x"3d",
           794 => x"80",
           795 => x"95",
           796 => x"51",
           797 => x"88",
           798 => x"53",
           799 => x"fe",
           800 => x"08",
           801 => x"57",
           802 => x"09",
           803 => x"38",
           804 => x"99",
           805 => x"2e",
           806 => x"56",
           807 => x"a4",
           808 => x"79",
           809 => x"f4",
           810 => x"56",
           811 => x"fd",
           812 => x"e5",
           813 => x"b3",
           814 => x"83",
           815 => x"58",
           816 => x"95",
           817 => x"51",
           818 => x"88",
           819 => x"af",
           820 => x"71",
           821 => x"05",
           822 => x"54",
           823 => x"f6",
           824 => x"08",
           825 => x"06",
           826 => x"1a",
           827 => x"33",
           828 => x"95",
           829 => x"51",
           830 => x"88",
           831 => x"23",
           832 => x"05",
           833 => x"3f",
           834 => x"ff",
           835 => x"75",
           836 => x"3d",
           837 => x"f5",
           838 => x"08",
           839 => x"f5",
           840 => x"08",
           841 => x"06",
           842 => x"79",
           843 => x"22",
           844 => x"82",
           845 => x"72",
           846 => x"59",
           847 => x"ee",
           848 => x"08",
           849 => x"88",
           850 => x"08",
           851 => x"56",
           852 => x"df",
           853 => x"38",
           854 => x"ff",
           855 => x"85",
           856 => x"89",
           857 => x"76",
           858 => x"c1",
           859 => x"34",
           860 => x"09",
           861 => x"38",
           862 => x"05",
           863 => x"3f",
           864 => x"1a",
           865 => x"8c",
           866 => x"90",
           867 => x"83",
           868 => x"8c",
           869 => x"71",
           870 => x"94",
           871 => x"80",
           872 => x"34",
           873 => x"0b",
           874 => x"80",
           875 => x"0c",
           876 => x"04",
           877 => x"0b",
           878 => x"f4",
           879 => x"54",
           880 => x"80",
           881 => x"0b",
           882 => x"98",
           883 => x"45",
           884 => x"3d",
           885 => x"ec",
           886 => x"9d",
           887 => x"54",
           888 => x"c0",
           889 => x"33",
           890 => x"2e",
           891 => x"a7",
           892 => x"84",
           893 => x"06",
           894 => x"73",
           895 => x"38",
           896 => x"39",
           897 => x"d5",
           898 => x"a0",
           899 => x"3d",
           900 => x"f3",
           901 => x"08",
           902 => x"73",
           903 => x"81",
           904 => x"34",
           905 => x"98",
           906 => x"f6",
           907 => x"7f",
           908 => x"0b",
           909 => x"59",
           910 => x"80",
           911 => x"57",
           912 => x"81",
           913 => x"16",
           914 => x"55",
           915 => x"80",
           916 => x"38",
           917 => x"81",
           918 => x"39",
           919 => x"17",
           920 => x"81",
           921 => x"16",
           922 => x"08",
           923 => x"78",
           924 => x"74",
           925 => x"2e",
           926 => x"98",
           927 => x"83",
           928 => x"57",
           929 => x"38",
           930 => x"ff",
           931 => x"2a",
           932 => x"ff",
           933 => x"79",
           934 => x"87",
           935 => x"08",
           936 => x"a4",
           937 => x"f3",
           938 => x"08",
           939 => x"27",
           940 => x"74",
           941 => x"a4",
           942 => x"f3",
           943 => x"08",
           944 => x"80",
           945 => x"38",
           946 => x"a8",
           947 => x"16",
           948 => x"06",
           949 => x"31",
           950 => x"75",
           951 => x"77",
           952 => x"98",
           953 => x"ff",
           954 => x"16",
           955 => x"51",
           956 => x"88",
           957 => x"38",
           958 => x"15",
           959 => x"77",
           960 => x"08",
           961 => x"58",
           962 => x"fe",
           963 => x"19",
           964 => x"39",
           965 => x"88",
           966 => x"0d",
           967 => x"0d",
           968 => x"8c",
           969 => x"84",
           970 => x"51",
           971 => x"88",
           972 => x"87",
           973 => x"08",
           974 => x"84",
           975 => x"51",
           976 => x"73",
           977 => x"87",
           978 => x"0c",
           979 => x"9c",
           980 => x"84",
           981 => x"51",
           982 => x"88",
           983 => x"87",
           984 => x"08",
           985 => x"84",
           986 => x"51",
           987 => x"73",
           988 => x"87",
           989 => x"0c",
           990 => x"0b",
           991 => x"84",
           992 => x"83",
           993 => x"94",
           994 => x"f8",
           995 => x"3f",
           996 => x"38",
           997 => x"fc",
           998 => x"08",
           999 => x"80",
          1000 => x"87",
          1001 => x"0c",
          1002 => x"fc",
          1003 => x"80",
          1004 => x"fc",
          1005 => x"08",
          1006 => x"54",
          1007 => x"86",
          1008 => x"55",
          1009 => x"80",
          1010 => x"80",
          1011 => x"00",
          1012 => x"ff",
          1013 => x"ff",
          1014 => x"ff",
          1015 => x"00",
          1016 => x"54",
          1017 => x"59",
          1018 => x"4d",
          1019 => x"00",
          1020 => x"00",
          2048 => x"c4",
          2049 => x"0b",
          2050 => x"04",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"c4",
          2057 => x"0b",
          2058 => x"04",
          2059 => x"c4",
          2060 => x"0b",
          2061 => x"04",
          2062 => x"c4",
          2063 => x"0b",
          2064 => x"04",
          2065 => x"c4",
          2066 => x"0b",
          2067 => x"04",
          2068 => x"c4",
          2069 => x"0b",
          2070 => x"04",
          2071 => x"c5",
          2072 => x"0b",
          2073 => x"04",
          2074 => x"c5",
          2075 => x"0b",
          2076 => x"04",
          2077 => x"c5",
          2078 => x"0b",
          2079 => x"04",
          2080 => x"c5",
          2081 => x"0b",
          2082 => x"04",
          2083 => x"c6",
          2084 => x"0b",
          2085 => x"04",
          2086 => x"c6",
          2087 => x"0b",
          2088 => x"04",
          2089 => x"c6",
          2090 => x"0b",
          2091 => x"04",
          2092 => x"c6",
          2093 => x"0b",
          2094 => x"04",
          2095 => x"c7",
          2096 => x"0b",
          2097 => x"04",
          2098 => x"c7",
          2099 => x"0b",
          2100 => x"04",
          2101 => x"c7",
          2102 => x"0b",
          2103 => x"04",
          2104 => x"c7",
          2105 => x"0b",
          2106 => x"04",
          2107 => x"c8",
          2108 => x"0b",
          2109 => x"04",
          2110 => x"c8",
          2111 => x"0b",
          2112 => x"04",
          2113 => x"c8",
          2114 => x"0b",
          2115 => x"04",
          2116 => x"c8",
          2117 => x"0b",
          2118 => x"04",
          2119 => x"c9",
          2120 => x"0b",
          2121 => x"04",
          2122 => x"c9",
          2123 => x"0b",
          2124 => x"04",
          2125 => x"c9",
          2126 => x"0b",
          2127 => x"04",
          2128 => x"c9",
          2129 => x"0b",
          2130 => x"04",
          2131 => x"00",
          2132 => x"00",
          2133 => x"00",
          2134 => x"00",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"80",
          2177 => x"f8",
          2178 => x"de",
          2179 => x"f8",
          2180 => x"90",
          2181 => x"f8",
          2182 => x"d3",
          2183 => x"f8",
          2184 => x"90",
          2185 => x"f8",
          2186 => x"92",
          2187 => x"f8",
          2188 => x"90",
          2189 => x"f8",
          2190 => x"b0",
          2191 => x"f8",
          2192 => x"90",
          2193 => x"f8",
          2194 => x"ee",
          2195 => x"f8",
          2196 => x"90",
          2197 => x"f8",
          2198 => x"ec",
          2199 => x"f8",
          2200 => x"90",
          2201 => x"f8",
          2202 => x"d3",
          2203 => x"f8",
          2204 => x"90",
          2205 => x"f8",
          2206 => x"89",
          2207 => x"f8",
          2208 => x"90",
          2209 => x"f8",
          2210 => x"fb",
          2211 => x"f8",
          2212 => x"90",
          2213 => x"f8",
          2214 => x"94",
          2215 => x"f8",
          2216 => x"90",
          2217 => x"f8",
          2218 => x"aa",
          2219 => x"f8",
          2220 => x"90",
          2221 => x"f8",
          2222 => x"ce",
          2223 => x"f8",
          2224 => x"90",
          2225 => x"f8",
          2226 => x"eb",
          2227 => x"f8",
          2228 => x"90",
          2229 => x"f8",
          2230 => x"bc",
          2231 => x"f8",
          2232 => x"90",
          2233 => x"f8",
          2234 => x"d8",
          2235 => x"f8",
          2236 => x"90",
          2237 => x"f8",
          2238 => x"8d",
          2239 => x"f8",
          2240 => x"90",
          2241 => x"f8",
          2242 => x"c0",
          2243 => x"f8",
          2244 => x"90",
          2245 => x"f8",
          2246 => x"b0",
          2247 => x"f8",
          2248 => x"90",
          2249 => x"f8",
          2250 => x"a1",
          2251 => x"f8",
          2252 => x"90",
          2253 => x"f8",
          2254 => x"95",
          2255 => x"f8",
          2256 => x"90",
          2257 => x"f8",
          2258 => x"92",
          2259 => x"f8",
          2260 => x"90",
          2261 => x"f8",
          2262 => x"b0",
          2263 => x"f8",
          2264 => x"90",
          2265 => x"f8",
          2266 => x"90",
          2267 => x"f8",
          2268 => x"90",
          2269 => x"f8",
          2270 => x"83",
          2271 => x"f8",
          2272 => x"90",
          2273 => x"f8",
          2274 => x"cf",
          2275 => x"f8",
          2276 => x"90",
          2277 => x"f8",
          2278 => x"ee",
          2279 => x"f8",
          2280 => x"90",
          2281 => x"f8",
          2282 => x"8d",
          2283 => x"f8",
          2284 => x"90",
          2285 => x"f8",
          2286 => x"f7",
          2287 => x"f8",
          2288 => x"90",
          2289 => x"f8",
          2290 => x"dd",
          2291 => x"f8",
          2292 => x"90",
          2293 => x"f8",
          2294 => x"cb",
          2295 => x"f8",
          2296 => x"90",
          2297 => x"f8",
          2298 => x"91",
          2299 => x"f8",
          2300 => x"90",
          2301 => x"f8",
          2302 => x"cb",
          2303 => x"f8",
          2304 => x"90",
          2305 => x"f8",
          2306 => x"cc",
          2307 => x"f8",
          2308 => x"90",
          2309 => x"f8",
          2310 => x"81",
          2311 => x"f8",
          2312 => x"90",
          2313 => x"f8",
          2314 => x"da",
          2315 => x"f8",
          2316 => x"90",
          2317 => x"f8",
          2318 => x"85",
          2319 => x"f8",
          2320 => x"90",
          2321 => x"f8",
          2322 => x"e8",
          2323 => x"f8",
          2324 => x"90",
          2325 => x"f8",
          2326 => x"bd",
          2327 => x"f8",
          2328 => x"90",
          2329 => x"f8",
          2330 => x"c7",
          2331 => x"f8",
          2332 => x"90",
          2333 => x"f8",
          2334 => x"89",
          2335 => x"f8",
          2336 => x"90",
          2337 => x"f8",
          2338 => x"cf",
          2339 => x"f8",
          2340 => x"90",
          2341 => x"f8",
          2342 => x"f5",
          2343 => x"f8",
          2344 => x"90",
          2345 => x"f8",
          2346 => x"8a",
          2347 => x"f8",
          2348 => x"90",
          2349 => x"f8",
          2350 => x"f4",
          2351 => x"f8",
          2352 => x"90",
          2353 => x"f8",
          2354 => x"d8",
          2355 => x"f8",
          2356 => x"90",
          2357 => x"f8",
          2358 => x"81",
          2359 => x"f8",
          2360 => x"90",
          2361 => x"f8",
          2362 => x"e3",
          2363 => x"f8",
          2364 => x"90",
          2365 => x"f8",
          2366 => x"d0",
          2367 => x"f8",
          2368 => x"90",
          2369 => x"f8",
          2370 => x"f2",
          2371 => x"f8",
          2372 => x"90",
          2373 => x"ec",
          2374 => x"98",
          2375 => x"80",
          2376 => x"05",
          2377 => x"0b",
          2378 => x"04",
          2379 => x"51",
          2380 => x"04",
          2381 => x"8c",
          2382 => x"82",
          2383 => x"fd",
          2384 => x"53",
          2385 => x"08",
          2386 => x"52",
          2387 => x"08",
          2388 => x"51",
          2389 => x"82",
          2390 => x"70",
          2391 => x"0c",
          2392 => x"0d",
          2393 => x"0c",
          2394 => x"f8",
          2395 => x"8c",
          2396 => x"3d",
          2397 => x"82",
          2398 => x"8c",
          2399 => x"82",
          2400 => x"88",
          2401 => x"93",
          2402 => x"ec",
          2403 => x"8c",
          2404 => x"85",
          2405 => x"8c",
          2406 => x"82",
          2407 => x"02",
          2408 => x"0c",
          2409 => x"81",
          2410 => x"f8",
          2411 => x"0c",
          2412 => x"8c",
          2413 => x"05",
          2414 => x"f8",
          2415 => x"08",
          2416 => x"08",
          2417 => x"27",
          2418 => x"8c",
          2419 => x"05",
          2420 => x"ae",
          2421 => x"82",
          2422 => x"8c",
          2423 => x"a2",
          2424 => x"f8",
          2425 => x"08",
          2426 => x"f8",
          2427 => x"0c",
          2428 => x"08",
          2429 => x"10",
          2430 => x"08",
          2431 => x"ff",
          2432 => x"8c",
          2433 => x"05",
          2434 => x"80",
          2435 => x"8c",
          2436 => x"05",
          2437 => x"f8",
          2438 => x"08",
          2439 => x"82",
          2440 => x"88",
          2441 => x"8c",
          2442 => x"05",
          2443 => x"8c",
          2444 => x"05",
          2445 => x"f8",
          2446 => x"08",
          2447 => x"08",
          2448 => x"07",
          2449 => x"08",
          2450 => x"82",
          2451 => x"fc",
          2452 => x"2a",
          2453 => x"08",
          2454 => x"82",
          2455 => x"8c",
          2456 => x"2a",
          2457 => x"08",
          2458 => x"ff",
          2459 => x"8c",
          2460 => x"05",
          2461 => x"93",
          2462 => x"f8",
          2463 => x"08",
          2464 => x"f8",
          2465 => x"0c",
          2466 => x"82",
          2467 => x"f8",
          2468 => x"82",
          2469 => x"f4",
          2470 => x"82",
          2471 => x"f4",
          2472 => x"8c",
          2473 => x"3d",
          2474 => x"f8",
          2475 => x"3d",
          2476 => x"71",
          2477 => x"9f",
          2478 => x"55",
          2479 => x"72",
          2480 => x"74",
          2481 => x"70",
          2482 => x"38",
          2483 => x"71",
          2484 => x"38",
          2485 => x"81",
          2486 => x"ff",
          2487 => x"ff",
          2488 => x"06",
          2489 => x"82",
          2490 => x"86",
          2491 => x"74",
          2492 => x"75",
          2493 => x"90",
          2494 => x"54",
          2495 => x"27",
          2496 => x"71",
          2497 => x"53",
          2498 => x"70",
          2499 => x"0c",
          2500 => x"84",
          2501 => x"72",
          2502 => x"05",
          2503 => x"12",
          2504 => x"26",
          2505 => x"72",
          2506 => x"72",
          2507 => x"05",
          2508 => x"12",
          2509 => x"26",
          2510 => x"53",
          2511 => x"fb",
          2512 => x"79",
          2513 => x"83",
          2514 => x"52",
          2515 => x"71",
          2516 => x"54",
          2517 => x"73",
          2518 => x"c6",
          2519 => x"54",
          2520 => x"70",
          2521 => x"52",
          2522 => x"2e",
          2523 => x"33",
          2524 => x"2e",
          2525 => x"95",
          2526 => x"81",
          2527 => x"70",
          2528 => x"54",
          2529 => x"70",
          2530 => x"33",
          2531 => x"ff",
          2532 => x"ff",
          2533 => x"31",
          2534 => x"0c",
          2535 => x"3d",
          2536 => x"09",
          2537 => x"fd",
          2538 => x"70",
          2539 => x"81",
          2540 => x"51",
          2541 => x"38",
          2542 => x"16",
          2543 => x"56",
          2544 => x"08",
          2545 => x"73",
          2546 => x"ff",
          2547 => x"0b",
          2548 => x"0c",
          2549 => x"04",
          2550 => x"80",
          2551 => x"71",
          2552 => x"87",
          2553 => x"8c",
          2554 => x"ff",
          2555 => x"ff",
          2556 => x"72",
          2557 => x"38",
          2558 => x"ec",
          2559 => x"0d",
          2560 => x"0d",
          2561 => x"70",
          2562 => x"71",
          2563 => x"ca",
          2564 => x"51",
          2565 => x"09",
          2566 => x"38",
          2567 => x"f1",
          2568 => x"84",
          2569 => x"53",
          2570 => x"70",
          2571 => x"53",
          2572 => x"a0",
          2573 => x"81",
          2574 => x"2e",
          2575 => x"e5",
          2576 => x"ff",
          2577 => x"a0",
          2578 => x"06",
          2579 => x"73",
          2580 => x"55",
          2581 => x"0c",
          2582 => x"82",
          2583 => x"87",
          2584 => x"fc",
          2585 => x"53",
          2586 => x"2e",
          2587 => x"3d",
          2588 => x"72",
          2589 => x"3f",
          2590 => x"08",
          2591 => x"53",
          2592 => x"53",
          2593 => x"ec",
          2594 => x"0d",
          2595 => x"0d",
          2596 => x"33",
          2597 => x"53",
          2598 => x"8b",
          2599 => x"38",
          2600 => x"ff",
          2601 => x"52",
          2602 => x"81",
          2603 => x"13",
          2604 => x"52",
          2605 => x"80",
          2606 => x"13",
          2607 => x"52",
          2608 => x"80",
          2609 => x"13",
          2610 => x"52",
          2611 => x"80",
          2612 => x"13",
          2613 => x"52",
          2614 => x"26",
          2615 => x"8a",
          2616 => x"87",
          2617 => x"e7",
          2618 => x"38",
          2619 => x"c0",
          2620 => x"72",
          2621 => x"98",
          2622 => x"13",
          2623 => x"98",
          2624 => x"13",
          2625 => x"98",
          2626 => x"13",
          2627 => x"98",
          2628 => x"13",
          2629 => x"98",
          2630 => x"13",
          2631 => x"98",
          2632 => x"87",
          2633 => x"0c",
          2634 => x"98",
          2635 => x"0b",
          2636 => x"9c",
          2637 => x"71",
          2638 => x"0c",
          2639 => x"04",
          2640 => x"7f",
          2641 => x"98",
          2642 => x"7d",
          2643 => x"98",
          2644 => x"7d",
          2645 => x"c0",
          2646 => x"5a",
          2647 => x"34",
          2648 => x"b4",
          2649 => x"83",
          2650 => x"c0",
          2651 => x"5a",
          2652 => x"34",
          2653 => x"ac",
          2654 => x"85",
          2655 => x"c0",
          2656 => x"5a",
          2657 => x"34",
          2658 => x"a4",
          2659 => x"88",
          2660 => x"c0",
          2661 => x"5a",
          2662 => x"23",
          2663 => x"79",
          2664 => x"06",
          2665 => x"ff",
          2666 => x"86",
          2667 => x"85",
          2668 => x"84",
          2669 => x"83",
          2670 => x"82",
          2671 => x"7d",
          2672 => x"06",
          2673 => x"ec",
          2674 => x"3f",
          2675 => x"04",
          2676 => x"02",
          2677 => x"70",
          2678 => x"2a",
          2679 => x"70",
          2680 => x"89",
          2681 => x"3d",
          2682 => x"3d",
          2683 => x"0b",
          2684 => x"33",
          2685 => x"06",
          2686 => x"87",
          2687 => x"51",
          2688 => x"86",
          2689 => x"94",
          2690 => x"08",
          2691 => x"70",
          2692 => x"54",
          2693 => x"2e",
          2694 => x"91",
          2695 => x"06",
          2696 => x"d7",
          2697 => x"32",
          2698 => x"51",
          2699 => x"2e",
          2700 => x"93",
          2701 => x"06",
          2702 => x"ff",
          2703 => x"81",
          2704 => x"87",
          2705 => x"52",
          2706 => x"86",
          2707 => x"94",
          2708 => x"72",
          2709 => x"8c",
          2710 => x"3d",
          2711 => x"3d",
          2712 => x"05",
          2713 => x"82",
          2714 => x"70",
          2715 => x"57",
          2716 => x"c0",
          2717 => x"74",
          2718 => x"38",
          2719 => x"94",
          2720 => x"70",
          2721 => x"81",
          2722 => x"52",
          2723 => x"8c",
          2724 => x"2a",
          2725 => x"51",
          2726 => x"38",
          2727 => x"70",
          2728 => x"51",
          2729 => x"8d",
          2730 => x"2a",
          2731 => x"51",
          2732 => x"be",
          2733 => x"ff",
          2734 => x"c0",
          2735 => x"70",
          2736 => x"38",
          2737 => x"90",
          2738 => x"0c",
          2739 => x"04",
          2740 => x"79",
          2741 => x"33",
          2742 => x"06",
          2743 => x"70",
          2744 => x"fe",
          2745 => x"ff",
          2746 => x"0b",
          2747 => x"94",
          2748 => x"ff",
          2749 => x"55",
          2750 => x"94",
          2751 => x"80",
          2752 => x"87",
          2753 => x"51",
          2754 => x"96",
          2755 => x"06",
          2756 => x"70",
          2757 => x"38",
          2758 => x"70",
          2759 => x"51",
          2760 => x"72",
          2761 => x"81",
          2762 => x"70",
          2763 => x"38",
          2764 => x"70",
          2765 => x"51",
          2766 => x"38",
          2767 => x"06",
          2768 => x"94",
          2769 => x"80",
          2770 => x"87",
          2771 => x"52",
          2772 => x"81",
          2773 => x"70",
          2774 => x"53",
          2775 => x"ff",
          2776 => x"82",
          2777 => x"89",
          2778 => x"fe",
          2779 => x"0b",
          2780 => x"33",
          2781 => x"06",
          2782 => x"c0",
          2783 => x"72",
          2784 => x"38",
          2785 => x"94",
          2786 => x"70",
          2787 => x"81",
          2788 => x"51",
          2789 => x"e2",
          2790 => x"ff",
          2791 => x"c0",
          2792 => x"70",
          2793 => x"38",
          2794 => x"90",
          2795 => x"70",
          2796 => x"82",
          2797 => x"51",
          2798 => x"04",
          2799 => x"0b",
          2800 => x"94",
          2801 => x"ff",
          2802 => x"87",
          2803 => x"52",
          2804 => x"86",
          2805 => x"94",
          2806 => x"08",
          2807 => x"70",
          2808 => x"51",
          2809 => x"70",
          2810 => x"38",
          2811 => x"06",
          2812 => x"94",
          2813 => x"80",
          2814 => x"87",
          2815 => x"52",
          2816 => x"98",
          2817 => x"2c",
          2818 => x"71",
          2819 => x"0c",
          2820 => x"04",
          2821 => x"87",
          2822 => x"08",
          2823 => x"8a",
          2824 => x"70",
          2825 => x"b4",
          2826 => x"9e",
          2827 => x"89",
          2828 => x"c0",
          2829 => x"82",
          2830 => x"87",
          2831 => x"08",
          2832 => x"0c",
          2833 => x"98",
          2834 => x"a4",
          2835 => x"9e",
          2836 => x"89",
          2837 => x"c0",
          2838 => x"82",
          2839 => x"87",
          2840 => x"08",
          2841 => x"0c",
          2842 => x"b0",
          2843 => x"b4",
          2844 => x"9e",
          2845 => x"89",
          2846 => x"c0",
          2847 => x"82",
          2848 => x"87",
          2849 => x"08",
          2850 => x"0c",
          2851 => x"c0",
          2852 => x"c4",
          2853 => x"9e",
          2854 => x"89",
          2855 => x"c0",
          2856 => x"51",
          2857 => x"cc",
          2858 => x"9e",
          2859 => x"89",
          2860 => x"c0",
          2861 => x"82",
          2862 => x"87",
          2863 => x"08",
          2864 => x"0c",
          2865 => x"89",
          2866 => x"0b",
          2867 => x"90",
          2868 => x"80",
          2869 => x"52",
          2870 => x"2e",
          2871 => x"52",
          2872 => x"dd",
          2873 => x"87",
          2874 => x"08",
          2875 => x"0a",
          2876 => x"52",
          2877 => x"83",
          2878 => x"71",
          2879 => x"34",
          2880 => x"c0",
          2881 => x"70",
          2882 => x"06",
          2883 => x"70",
          2884 => x"38",
          2885 => x"82",
          2886 => x"80",
          2887 => x"9e",
          2888 => x"88",
          2889 => x"51",
          2890 => x"80",
          2891 => x"81",
          2892 => x"89",
          2893 => x"0b",
          2894 => x"90",
          2895 => x"80",
          2896 => x"52",
          2897 => x"2e",
          2898 => x"52",
          2899 => x"e1",
          2900 => x"87",
          2901 => x"08",
          2902 => x"80",
          2903 => x"52",
          2904 => x"83",
          2905 => x"71",
          2906 => x"34",
          2907 => x"c0",
          2908 => x"70",
          2909 => x"06",
          2910 => x"70",
          2911 => x"38",
          2912 => x"82",
          2913 => x"80",
          2914 => x"9e",
          2915 => x"82",
          2916 => x"51",
          2917 => x"80",
          2918 => x"81",
          2919 => x"89",
          2920 => x"0b",
          2921 => x"90",
          2922 => x"80",
          2923 => x"52",
          2924 => x"2e",
          2925 => x"52",
          2926 => x"e5",
          2927 => x"87",
          2928 => x"08",
          2929 => x"80",
          2930 => x"52",
          2931 => x"83",
          2932 => x"71",
          2933 => x"34",
          2934 => x"c0",
          2935 => x"70",
          2936 => x"51",
          2937 => x"80",
          2938 => x"81",
          2939 => x"89",
          2940 => x"c0",
          2941 => x"70",
          2942 => x"70",
          2943 => x"51",
          2944 => x"89",
          2945 => x"0b",
          2946 => x"90",
          2947 => x"80",
          2948 => x"52",
          2949 => x"83",
          2950 => x"71",
          2951 => x"34",
          2952 => x"90",
          2953 => x"f0",
          2954 => x"2a",
          2955 => x"70",
          2956 => x"34",
          2957 => x"c0",
          2958 => x"70",
          2959 => x"52",
          2960 => x"2e",
          2961 => x"52",
          2962 => x"eb",
          2963 => x"9e",
          2964 => x"87",
          2965 => x"70",
          2966 => x"34",
          2967 => x"04",
          2968 => x"81",
          2969 => x"85",
          2970 => x"89",
          2971 => x"73",
          2972 => x"38",
          2973 => x"51",
          2974 => x"81",
          2975 => x"85",
          2976 => x"89",
          2977 => x"73",
          2978 => x"38",
          2979 => x"08",
          2980 => x"08",
          2981 => x"81",
          2982 => x"8a",
          2983 => x"89",
          2984 => x"73",
          2985 => x"38",
          2986 => x"08",
          2987 => x"08",
          2988 => x"81",
          2989 => x"8a",
          2990 => x"89",
          2991 => x"73",
          2992 => x"38",
          2993 => x"08",
          2994 => x"08",
          2995 => x"81",
          2996 => x"8a",
          2997 => x"89",
          2998 => x"73",
          2999 => x"38",
          3000 => x"08",
          3001 => x"08",
          3002 => x"81",
          3003 => x"8a",
          3004 => x"89",
          3005 => x"73",
          3006 => x"38",
          3007 => x"08",
          3008 => x"08",
          3009 => x"81",
          3010 => x"8a",
          3011 => x"89",
          3012 => x"73",
          3013 => x"38",
          3014 => x"33",
          3015 => x"d0",
          3016 => x"3f",
          3017 => x"33",
          3018 => x"2e",
          3019 => x"89",
          3020 => x"81",
          3021 => x"89",
          3022 => x"89",
          3023 => x"73",
          3024 => x"38",
          3025 => x"33",
          3026 => x"90",
          3027 => x"3f",
          3028 => x"33",
          3029 => x"2e",
          3030 => x"f8",
          3031 => x"d0",
          3032 => x"df",
          3033 => x"80",
          3034 => x"81",
          3035 => x"83",
          3036 => x"89",
          3037 => x"73",
          3038 => x"38",
          3039 => x"51",
          3040 => x"82",
          3041 => x"54",
          3042 => x"88",
          3043 => x"dc",
          3044 => x"3f",
          3045 => x"33",
          3046 => x"2e",
          3047 => x"f8",
          3048 => x"8c",
          3049 => x"f4",
          3050 => x"3f",
          3051 => x"08",
          3052 => x"80",
          3053 => x"3f",
          3054 => x"08",
          3055 => x"a8",
          3056 => x"3f",
          3057 => x"08",
          3058 => x"d0",
          3059 => x"3f",
          3060 => x"51",
          3061 => x"82",
          3062 => x"52",
          3063 => x"51",
          3064 => x"82",
          3065 => x"56",
          3066 => x"52",
          3067 => x"c6",
          3068 => x"ec",
          3069 => x"c0",
          3070 => x"31",
          3071 => x"8c",
          3072 => x"81",
          3073 => x"88",
          3074 => x"89",
          3075 => x"73",
          3076 => x"38",
          3077 => x"08",
          3078 => x"c0",
          3079 => x"ea",
          3080 => x"8c",
          3081 => x"84",
          3082 => x"71",
          3083 => x"82",
          3084 => x"52",
          3085 => x"51",
          3086 => x"82",
          3087 => x"54",
          3088 => x"a8",
          3089 => x"d8",
          3090 => x"84",
          3091 => x"51",
          3092 => x"82",
          3093 => x"bd",
          3094 => x"76",
          3095 => x"54",
          3096 => x"08",
          3097 => x"80",
          3098 => x"3f",
          3099 => x"51",
          3100 => x"87",
          3101 => x"fe",
          3102 => x"92",
          3103 => x"05",
          3104 => x"26",
          3105 => x"84",
          3106 => x"81",
          3107 => x"52",
          3108 => x"81",
          3109 => x"9d",
          3110 => x"b4",
          3111 => x"81",
          3112 => x"91",
          3113 => x"c4",
          3114 => x"81",
          3115 => x"85",
          3116 => x"d0",
          3117 => x"3f",
          3118 => x"04",
          3119 => x"0c",
          3120 => x"87",
          3121 => x"0c",
          3122 => x"f0",
          3123 => x"96",
          3124 => x"fe",
          3125 => x"93",
          3126 => x"72",
          3127 => x"81",
          3128 => x"8d",
          3129 => x"82",
          3130 => x"52",
          3131 => x"90",
          3132 => x"34",
          3133 => x"08",
          3134 => x"8d",
          3135 => x"39",
          3136 => x"08",
          3137 => x"2e",
          3138 => x"51",
          3139 => x"3d",
          3140 => x"3d",
          3141 => x"05",
          3142 => x"fc",
          3143 => x"8c",
          3144 => x"51",
          3145 => x"72",
          3146 => x"0c",
          3147 => x"04",
          3148 => x"75",
          3149 => x"70",
          3150 => x"53",
          3151 => x"2e",
          3152 => x"81",
          3153 => x"81",
          3154 => x"87",
          3155 => x"85",
          3156 => x"fc",
          3157 => x"82",
          3158 => x"78",
          3159 => x"0c",
          3160 => x"33",
          3161 => x"06",
          3162 => x"80",
          3163 => x"72",
          3164 => x"51",
          3165 => x"fe",
          3166 => x"39",
          3167 => x"fc",
          3168 => x"0d",
          3169 => x"0d",
          3170 => x"59",
          3171 => x"05",
          3172 => x"75",
          3173 => x"f8",
          3174 => x"2e",
          3175 => x"82",
          3176 => x"70",
          3177 => x"05",
          3178 => x"5b",
          3179 => x"2e",
          3180 => x"85",
          3181 => x"8b",
          3182 => x"2e",
          3183 => x"8a",
          3184 => x"78",
          3185 => x"5a",
          3186 => x"aa",
          3187 => x"06",
          3188 => x"84",
          3189 => x"7b",
          3190 => x"5d",
          3191 => x"59",
          3192 => x"d0",
          3193 => x"89",
          3194 => x"7a",
          3195 => x"10",
          3196 => x"d0",
          3197 => x"81",
          3198 => x"57",
          3199 => x"75",
          3200 => x"70",
          3201 => x"07",
          3202 => x"80",
          3203 => x"30",
          3204 => x"80",
          3205 => x"53",
          3206 => x"55",
          3207 => x"2e",
          3208 => x"84",
          3209 => x"81",
          3210 => x"57",
          3211 => x"2e",
          3212 => x"75",
          3213 => x"76",
          3214 => x"e0",
          3215 => x"ff",
          3216 => x"73",
          3217 => x"81",
          3218 => x"80",
          3219 => x"38",
          3220 => x"2e",
          3221 => x"73",
          3222 => x"8b",
          3223 => x"c2",
          3224 => x"38",
          3225 => x"73",
          3226 => x"81",
          3227 => x"8f",
          3228 => x"d5",
          3229 => x"38",
          3230 => x"24",
          3231 => x"80",
          3232 => x"38",
          3233 => x"73",
          3234 => x"80",
          3235 => x"ef",
          3236 => x"19",
          3237 => x"59",
          3238 => x"33",
          3239 => x"75",
          3240 => x"81",
          3241 => x"70",
          3242 => x"55",
          3243 => x"79",
          3244 => x"90",
          3245 => x"16",
          3246 => x"7b",
          3247 => x"a0",
          3248 => x"3f",
          3249 => x"53",
          3250 => x"e9",
          3251 => x"fc",
          3252 => x"81",
          3253 => x"72",
          3254 => x"b0",
          3255 => x"fb",
          3256 => x"39",
          3257 => x"83",
          3258 => x"59",
          3259 => x"82",
          3260 => x"88",
          3261 => x"8a",
          3262 => x"90",
          3263 => x"75",
          3264 => x"3f",
          3265 => x"79",
          3266 => x"81",
          3267 => x"72",
          3268 => x"38",
          3269 => x"59",
          3270 => x"84",
          3271 => x"58",
          3272 => x"80",
          3273 => x"30",
          3274 => x"80",
          3275 => x"55",
          3276 => x"25",
          3277 => x"80",
          3278 => x"74",
          3279 => x"07",
          3280 => x"0b",
          3281 => x"57",
          3282 => x"51",
          3283 => x"82",
          3284 => x"81",
          3285 => x"53",
          3286 => x"e3",
          3287 => x"8c",
          3288 => x"89",
          3289 => x"38",
          3290 => x"75",
          3291 => x"84",
          3292 => x"53",
          3293 => x"06",
          3294 => x"53",
          3295 => x"81",
          3296 => x"81",
          3297 => x"70",
          3298 => x"2a",
          3299 => x"76",
          3300 => x"38",
          3301 => x"38",
          3302 => x"70",
          3303 => x"53",
          3304 => x"8e",
          3305 => x"77",
          3306 => x"53",
          3307 => x"81",
          3308 => x"7a",
          3309 => x"55",
          3310 => x"83",
          3311 => x"79",
          3312 => x"81",
          3313 => x"72",
          3314 => x"17",
          3315 => x"27",
          3316 => x"51",
          3317 => x"75",
          3318 => x"72",
          3319 => x"81",
          3320 => x"7a",
          3321 => x"38",
          3322 => x"05",
          3323 => x"ff",
          3324 => x"70",
          3325 => x"57",
          3326 => x"76",
          3327 => x"81",
          3328 => x"72",
          3329 => x"84",
          3330 => x"f9",
          3331 => x"39",
          3332 => x"04",
          3333 => x"86",
          3334 => x"84",
          3335 => x"55",
          3336 => x"fa",
          3337 => x"3d",
          3338 => x"3d",
          3339 => x"8d",
          3340 => x"3d",
          3341 => x"75",
          3342 => x"3f",
          3343 => x"08",
          3344 => x"34",
          3345 => x"8d",
          3346 => x"3d",
          3347 => x"3d",
          3348 => x"fc",
          3349 => x"8c",
          3350 => x"3d",
          3351 => x"77",
          3352 => x"a1",
          3353 => x"8c",
          3354 => x"3d",
          3355 => x"3d",
          3356 => x"82",
          3357 => x"70",
          3358 => x"55",
          3359 => x"80",
          3360 => x"38",
          3361 => x"08",
          3362 => x"82",
          3363 => x"81",
          3364 => x"72",
          3365 => x"cb",
          3366 => x"2e",
          3367 => x"88",
          3368 => x"70",
          3369 => x"51",
          3370 => x"2e",
          3371 => x"80",
          3372 => x"ff",
          3373 => x"39",
          3374 => x"c8",
          3375 => x"52",
          3376 => x"c0",
          3377 => x"52",
          3378 => x"81",
          3379 => x"51",
          3380 => x"ff",
          3381 => x"15",
          3382 => x"34",
          3383 => x"f3",
          3384 => x"72",
          3385 => x"0c",
          3386 => x"04",
          3387 => x"82",
          3388 => x"75",
          3389 => x"0c",
          3390 => x"52",
          3391 => x"3f",
          3392 => x"80",
          3393 => x"0d",
          3394 => x"0d",
          3395 => x"56",
          3396 => x"0c",
          3397 => x"70",
          3398 => x"73",
          3399 => x"81",
          3400 => x"81",
          3401 => x"ed",
          3402 => x"2e",
          3403 => x"8e",
          3404 => x"08",
          3405 => x"76",
          3406 => x"56",
          3407 => x"b0",
          3408 => x"06",
          3409 => x"75",
          3410 => x"76",
          3411 => x"70",
          3412 => x"73",
          3413 => x"8b",
          3414 => x"73",
          3415 => x"85",
          3416 => x"82",
          3417 => x"76",
          3418 => x"70",
          3419 => x"ac",
          3420 => x"a0",
          3421 => x"fa",
          3422 => x"53",
          3423 => x"57",
          3424 => x"98",
          3425 => x"39",
          3426 => x"80",
          3427 => x"26",
          3428 => x"86",
          3429 => x"80",
          3430 => x"57",
          3431 => x"74",
          3432 => x"38",
          3433 => x"27",
          3434 => x"14",
          3435 => x"06",
          3436 => x"14",
          3437 => x"06",
          3438 => x"74",
          3439 => x"f9",
          3440 => x"ff",
          3441 => x"89",
          3442 => x"38",
          3443 => x"c5",
          3444 => x"29",
          3445 => x"81",
          3446 => x"76",
          3447 => x"56",
          3448 => x"ba",
          3449 => x"2e",
          3450 => x"30",
          3451 => x"0c",
          3452 => x"82",
          3453 => x"8a",
          3454 => x"f8",
          3455 => x"7c",
          3456 => x"70",
          3457 => x"75",
          3458 => x"55",
          3459 => x"2e",
          3460 => x"87",
          3461 => x"76",
          3462 => x"73",
          3463 => x"81",
          3464 => x"81",
          3465 => x"77",
          3466 => x"70",
          3467 => x"58",
          3468 => x"09",
          3469 => x"c2",
          3470 => x"81",
          3471 => x"75",
          3472 => x"55",
          3473 => x"e2",
          3474 => x"90",
          3475 => x"f8",
          3476 => x"8f",
          3477 => x"81",
          3478 => x"75",
          3479 => x"55",
          3480 => x"81",
          3481 => x"27",
          3482 => x"d0",
          3483 => x"55",
          3484 => x"73",
          3485 => x"80",
          3486 => x"14",
          3487 => x"72",
          3488 => x"e0",
          3489 => x"80",
          3490 => x"39",
          3491 => x"55",
          3492 => x"80",
          3493 => x"e0",
          3494 => x"38",
          3495 => x"81",
          3496 => x"53",
          3497 => x"81",
          3498 => x"53",
          3499 => x"8e",
          3500 => x"70",
          3501 => x"55",
          3502 => x"27",
          3503 => x"77",
          3504 => x"74",
          3505 => x"76",
          3506 => x"77",
          3507 => x"70",
          3508 => x"55",
          3509 => x"77",
          3510 => x"38",
          3511 => x"74",
          3512 => x"55",
          3513 => x"ec",
          3514 => x"0d",
          3515 => x"0d",
          3516 => x"33",
          3517 => x"70",
          3518 => x"38",
          3519 => x"11",
          3520 => x"82",
          3521 => x"83",
          3522 => x"fc",
          3523 => x"9b",
          3524 => x"84",
          3525 => x"33",
          3526 => x"51",
          3527 => x"80",
          3528 => x"84",
          3529 => x"92",
          3530 => x"51",
          3531 => x"80",
          3532 => x"81",
          3533 => x"72",
          3534 => x"92",
          3535 => x"81",
          3536 => x"0b",
          3537 => x"8c",
          3538 => x"71",
          3539 => x"06",
          3540 => x"80",
          3541 => x"87",
          3542 => x"08",
          3543 => x"38",
          3544 => x"80",
          3545 => x"71",
          3546 => x"c0",
          3547 => x"51",
          3548 => x"87",
          3549 => x"89",
          3550 => x"82",
          3551 => x"33",
          3552 => x"8c",
          3553 => x"3d",
          3554 => x"3d",
          3555 => x"64",
          3556 => x"bf",
          3557 => x"40",
          3558 => x"74",
          3559 => x"cd",
          3560 => x"ec",
          3561 => x"7a",
          3562 => x"81",
          3563 => x"72",
          3564 => x"87",
          3565 => x"11",
          3566 => x"8c",
          3567 => x"92",
          3568 => x"5a",
          3569 => x"58",
          3570 => x"c0",
          3571 => x"76",
          3572 => x"76",
          3573 => x"70",
          3574 => x"81",
          3575 => x"54",
          3576 => x"8e",
          3577 => x"52",
          3578 => x"81",
          3579 => x"81",
          3580 => x"74",
          3581 => x"53",
          3582 => x"83",
          3583 => x"78",
          3584 => x"8f",
          3585 => x"2e",
          3586 => x"c0",
          3587 => x"52",
          3588 => x"87",
          3589 => x"08",
          3590 => x"2e",
          3591 => x"84",
          3592 => x"38",
          3593 => x"87",
          3594 => x"15",
          3595 => x"70",
          3596 => x"52",
          3597 => x"ff",
          3598 => x"39",
          3599 => x"81",
          3600 => x"ff",
          3601 => x"57",
          3602 => x"90",
          3603 => x"80",
          3604 => x"71",
          3605 => x"78",
          3606 => x"38",
          3607 => x"80",
          3608 => x"80",
          3609 => x"81",
          3610 => x"72",
          3611 => x"0c",
          3612 => x"04",
          3613 => x"60",
          3614 => x"8c",
          3615 => x"33",
          3616 => x"5b",
          3617 => x"74",
          3618 => x"e1",
          3619 => x"ec",
          3620 => x"79",
          3621 => x"78",
          3622 => x"06",
          3623 => x"77",
          3624 => x"87",
          3625 => x"11",
          3626 => x"8c",
          3627 => x"92",
          3628 => x"59",
          3629 => x"85",
          3630 => x"98",
          3631 => x"7d",
          3632 => x"0c",
          3633 => x"08",
          3634 => x"70",
          3635 => x"53",
          3636 => x"2e",
          3637 => x"70",
          3638 => x"33",
          3639 => x"18",
          3640 => x"2a",
          3641 => x"51",
          3642 => x"2e",
          3643 => x"c0",
          3644 => x"52",
          3645 => x"87",
          3646 => x"08",
          3647 => x"2e",
          3648 => x"84",
          3649 => x"38",
          3650 => x"87",
          3651 => x"15",
          3652 => x"70",
          3653 => x"52",
          3654 => x"ff",
          3655 => x"39",
          3656 => x"81",
          3657 => x"80",
          3658 => x"52",
          3659 => x"90",
          3660 => x"80",
          3661 => x"71",
          3662 => x"7a",
          3663 => x"38",
          3664 => x"80",
          3665 => x"80",
          3666 => x"81",
          3667 => x"72",
          3668 => x"0c",
          3669 => x"04",
          3670 => x"7a",
          3671 => x"a3",
          3672 => x"88",
          3673 => x"33",
          3674 => x"56",
          3675 => x"3f",
          3676 => x"08",
          3677 => x"83",
          3678 => x"fe",
          3679 => x"87",
          3680 => x"0c",
          3681 => x"76",
          3682 => x"38",
          3683 => x"93",
          3684 => x"2b",
          3685 => x"8c",
          3686 => x"71",
          3687 => x"38",
          3688 => x"71",
          3689 => x"c6",
          3690 => x"39",
          3691 => x"81",
          3692 => x"06",
          3693 => x"71",
          3694 => x"38",
          3695 => x"8c",
          3696 => x"e8",
          3697 => x"98",
          3698 => x"71",
          3699 => x"73",
          3700 => x"92",
          3701 => x"72",
          3702 => x"06",
          3703 => x"f7",
          3704 => x"80",
          3705 => x"88",
          3706 => x"0c",
          3707 => x"80",
          3708 => x"56",
          3709 => x"56",
          3710 => x"82",
          3711 => x"88",
          3712 => x"fe",
          3713 => x"81",
          3714 => x"33",
          3715 => x"07",
          3716 => x"0c",
          3717 => x"3d",
          3718 => x"3d",
          3719 => x"11",
          3720 => x"33",
          3721 => x"71",
          3722 => x"81",
          3723 => x"72",
          3724 => x"75",
          3725 => x"82",
          3726 => x"52",
          3727 => x"54",
          3728 => x"0d",
          3729 => x"0d",
          3730 => x"05",
          3731 => x"52",
          3732 => x"70",
          3733 => x"34",
          3734 => x"51",
          3735 => x"83",
          3736 => x"ff",
          3737 => x"75",
          3738 => x"72",
          3739 => x"54",
          3740 => x"2a",
          3741 => x"70",
          3742 => x"34",
          3743 => x"51",
          3744 => x"81",
          3745 => x"70",
          3746 => x"70",
          3747 => x"3d",
          3748 => x"3d",
          3749 => x"77",
          3750 => x"70",
          3751 => x"38",
          3752 => x"05",
          3753 => x"70",
          3754 => x"34",
          3755 => x"eb",
          3756 => x"0d",
          3757 => x"0d",
          3758 => x"54",
          3759 => x"72",
          3760 => x"54",
          3761 => x"51",
          3762 => x"84",
          3763 => x"fc",
          3764 => x"77",
          3765 => x"53",
          3766 => x"05",
          3767 => x"70",
          3768 => x"33",
          3769 => x"ff",
          3770 => x"52",
          3771 => x"2e",
          3772 => x"80",
          3773 => x"71",
          3774 => x"0c",
          3775 => x"04",
          3776 => x"74",
          3777 => x"89",
          3778 => x"2e",
          3779 => x"11",
          3780 => x"52",
          3781 => x"70",
          3782 => x"ec",
          3783 => x"0d",
          3784 => x"82",
          3785 => x"04",
          3786 => x"8c",
          3787 => x"f7",
          3788 => x"56",
          3789 => x"17",
          3790 => x"74",
          3791 => x"d6",
          3792 => x"b0",
          3793 => x"b4",
          3794 => x"81",
          3795 => x"59",
          3796 => x"82",
          3797 => x"7a",
          3798 => x"06",
          3799 => x"8c",
          3800 => x"17",
          3801 => x"08",
          3802 => x"08",
          3803 => x"08",
          3804 => x"74",
          3805 => x"38",
          3806 => x"55",
          3807 => x"09",
          3808 => x"38",
          3809 => x"18",
          3810 => x"81",
          3811 => x"f9",
          3812 => x"39",
          3813 => x"82",
          3814 => x"8b",
          3815 => x"fa",
          3816 => x"7a",
          3817 => x"57",
          3818 => x"08",
          3819 => x"75",
          3820 => x"3f",
          3821 => x"08",
          3822 => x"ec",
          3823 => x"81",
          3824 => x"b4",
          3825 => x"16",
          3826 => x"be",
          3827 => x"ec",
          3828 => x"85",
          3829 => x"81",
          3830 => x"17",
          3831 => x"8c",
          3832 => x"3d",
          3833 => x"3d",
          3834 => x"52",
          3835 => x"3f",
          3836 => x"08",
          3837 => x"ec",
          3838 => x"38",
          3839 => x"74",
          3840 => x"81",
          3841 => x"38",
          3842 => x"59",
          3843 => x"09",
          3844 => x"e3",
          3845 => x"53",
          3846 => x"08",
          3847 => x"70",
          3848 => x"91",
          3849 => x"d5",
          3850 => x"17",
          3851 => x"3f",
          3852 => x"a4",
          3853 => x"51",
          3854 => x"86",
          3855 => x"f2",
          3856 => x"17",
          3857 => x"3f",
          3858 => x"52",
          3859 => x"51",
          3860 => x"8c",
          3861 => x"84",
          3862 => x"fc",
          3863 => x"17",
          3864 => x"70",
          3865 => x"79",
          3866 => x"52",
          3867 => x"51",
          3868 => x"77",
          3869 => x"80",
          3870 => x"81",
          3871 => x"f9",
          3872 => x"8c",
          3873 => x"2e",
          3874 => x"58",
          3875 => x"ec",
          3876 => x"0d",
          3877 => x"0d",
          3878 => x"98",
          3879 => x"05",
          3880 => x"80",
          3881 => x"27",
          3882 => x"14",
          3883 => x"29",
          3884 => x"05",
          3885 => x"82",
          3886 => x"87",
          3887 => x"f9",
          3888 => x"7a",
          3889 => x"54",
          3890 => x"27",
          3891 => x"76",
          3892 => x"27",
          3893 => x"ff",
          3894 => x"58",
          3895 => x"80",
          3896 => x"82",
          3897 => x"72",
          3898 => x"38",
          3899 => x"72",
          3900 => x"8e",
          3901 => x"39",
          3902 => x"17",
          3903 => x"a4",
          3904 => x"53",
          3905 => x"fd",
          3906 => x"8c",
          3907 => x"9f",
          3908 => x"ff",
          3909 => x"11",
          3910 => x"70",
          3911 => x"18",
          3912 => x"76",
          3913 => x"53",
          3914 => x"82",
          3915 => x"80",
          3916 => x"83",
          3917 => x"b4",
          3918 => x"88",
          3919 => x"79",
          3920 => x"84",
          3921 => x"58",
          3922 => x"80",
          3923 => x"9f",
          3924 => x"80",
          3925 => x"88",
          3926 => x"08",
          3927 => x"51",
          3928 => x"82",
          3929 => x"80",
          3930 => x"10",
          3931 => x"74",
          3932 => x"51",
          3933 => x"82",
          3934 => x"83",
          3935 => x"58",
          3936 => x"87",
          3937 => x"08",
          3938 => x"51",
          3939 => x"82",
          3940 => x"9b",
          3941 => x"2b",
          3942 => x"74",
          3943 => x"51",
          3944 => x"82",
          3945 => x"f0",
          3946 => x"83",
          3947 => x"77",
          3948 => x"0c",
          3949 => x"04",
          3950 => x"7a",
          3951 => x"58",
          3952 => x"81",
          3953 => x"9e",
          3954 => x"17",
          3955 => x"96",
          3956 => x"53",
          3957 => x"81",
          3958 => x"79",
          3959 => x"72",
          3960 => x"38",
          3961 => x"72",
          3962 => x"b8",
          3963 => x"39",
          3964 => x"17",
          3965 => x"a4",
          3966 => x"53",
          3967 => x"fb",
          3968 => x"8c",
          3969 => x"82",
          3970 => x"81",
          3971 => x"83",
          3972 => x"b4",
          3973 => x"78",
          3974 => x"56",
          3975 => x"76",
          3976 => x"38",
          3977 => x"9f",
          3978 => x"33",
          3979 => x"07",
          3980 => x"74",
          3981 => x"83",
          3982 => x"89",
          3983 => x"08",
          3984 => x"51",
          3985 => x"82",
          3986 => x"59",
          3987 => x"08",
          3988 => x"74",
          3989 => x"16",
          3990 => x"84",
          3991 => x"76",
          3992 => x"88",
          3993 => x"81",
          3994 => x"8f",
          3995 => x"53",
          3996 => x"80",
          3997 => x"88",
          3998 => x"08",
          3999 => x"51",
          4000 => x"82",
          4001 => x"59",
          4002 => x"08",
          4003 => x"77",
          4004 => x"06",
          4005 => x"83",
          4006 => x"05",
          4007 => x"f7",
          4008 => x"39",
          4009 => x"a4",
          4010 => x"52",
          4011 => x"ef",
          4012 => x"ec",
          4013 => x"8c",
          4014 => x"38",
          4015 => x"06",
          4016 => x"83",
          4017 => x"18",
          4018 => x"54",
          4019 => x"f6",
          4020 => x"8c",
          4021 => x"0a",
          4022 => x"52",
          4023 => x"83",
          4024 => x"83",
          4025 => x"82",
          4026 => x"8a",
          4027 => x"f8",
          4028 => x"7c",
          4029 => x"59",
          4030 => x"81",
          4031 => x"38",
          4032 => x"08",
          4033 => x"73",
          4034 => x"38",
          4035 => x"52",
          4036 => x"a4",
          4037 => x"ec",
          4038 => x"8c",
          4039 => x"f2",
          4040 => x"82",
          4041 => x"39",
          4042 => x"e6",
          4043 => x"ec",
          4044 => x"de",
          4045 => x"78",
          4046 => x"3f",
          4047 => x"08",
          4048 => x"ec",
          4049 => x"80",
          4050 => x"8c",
          4051 => x"2e",
          4052 => x"8c",
          4053 => x"2e",
          4054 => x"53",
          4055 => x"51",
          4056 => x"82",
          4057 => x"c5",
          4058 => x"08",
          4059 => x"18",
          4060 => x"57",
          4061 => x"90",
          4062 => x"90",
          4063 => x"16",
          4064 => x"54",
          4065 => x"34",
          4066 => x"78",
          4067 => x"38",
          4068 => x"82",
          4069 => x"8a",
          4070 => x"f6",
          4071 => x"7e",
          4072 => x"5b",
          4073 => x"38",
          4074 => x"58",
          4075 => x"88",
          4076 => x"08",
          4077 => x"38",
          4078 => x"39",
          4079 => x"51",
          4080 => x"81",
          4081 => x"8c",
          4082 => x"82",
          4083 => x"8c",
          4084 => x"82",
          4085 => x"ff",
          4086 => x"38",
          4087 => x"82",
          4088 => x"26",
          4089 => x"79",
          4090 => x"08",
          4091 => x"73",
          4092 => x"b9",
          4093 => x"2e",
          4094 => x"80",
          4095 => x"1a",
          4096 => x"08",
          4097 => x"38",
          4098 => x"52",
          4099 => x"af",
          4100 => x"82",
          4101 => x"81",
          4102 => x"06",
          4103 => x"8c",
          4104 => x"82",
          4105 => x"09",
          4106 => x"72",
          4107 => x"70",
          4108 => x"8c",
          4109 => x"51",
          4110 => x"73",
          4111 => x"82",
          4112 => x"80",
          4113 => x"8c",
          4114 => x"81",
          4115 => x"38",
          4116 => x"08",
          4117 => x"73",
          4118 => x"75",
          4119 => x"77",
          4120 => x"56",
          4121 => x"76",
          4122 => x"82",
          4123 => x"26",
          4124 => x"75",
          4125 => x"f8",
          4126 => x"8c",
          4127 => x"2e",
          4128 => x"59",
          4129 => x"08",
          4130 => x"81",
          4131 => x"82",
          4132 => x"59",
          4133 => x"08",
          4134 => x"70",
          4135 => x"25",
          4136 => x"51",
          4137 => x"73",
          4138 => x"75",
          4139 => x"81",
          4140 => x"38",
          4141 => x"f5",
          4142 => x"75",
          4143 => x"f9",
          4144 => x"8c",
          4145 => x"8c",
          4146 => x"70",
          4147 => x"08",
          4148 => x"51",
          4149 => x"80",
          4150 => x"73",
          4151 => x"38",
          4152 => x"52",
          4153 => x"d0",
          4154 => x"ec",
          4155 => x"a5",
          4156 => x"18",
          4157 => x"08",
          4158 => x"18",
          4159 => x"74",
          4160 => x"38",
          4161 => x"18",
          4162 => x"33",
          4163 => x"73",
          4164 => x"97",
          4165 => x"74",
          4166 => x"38",
          4167 => x"55",
          4168 => x"8c",
          4169 => x"85",
          4170 => x"75",
          4171 => x"8c",
          4172 => x"3d",
          4173 => x"3d",
          4174 => x"52",
          4175 => x"3f",
          4176 => x"08",
          4177 => x"82",
          4178 => x"80",
          4179 => x"52",
          4180 => x"c1",
          4181 => x"ec",
          4182 => x"ec",
          4183 => x"0c",
          4184 => x"53",
          4185 => x"15",
          4186 => x"f2",
          4187 => x"56",
          4188 => x"16",
          4189 => x"22",
          4190 => x"27",
          4191 => x"54",
          4192 => x"76",
          4193 => x"33",
          4194 => x"3f",
          4195 => x"08",
          4196 => x"38",
          4197 => x"76",
          4198 => x"70",
          4199 => x"9f",
          4200 => x"56",
          4201 => x"8c",
          4202 => x"3d",
          4203 => x"3d",
          4204 => x"71",
          4205 => x"57",
          4206 => x"0a",
          4207 => x"38",
          4208 => x"53",
          4209 => x"38",
          4210 => x"0c",
          4211 => x"54",
          4212 => x"75",
          4213 => x"73",
          4214 => x"a8",
          4215 => x"73",
          4216 => x"85",
          4217 => x"0b",
          4218 => x"5a",
          4219 => x"27",
          4220 => x"a8",
          4221 => x"18",
          4222 => x"39",
          4223 => x"70",
          4224 => x"58",
          4225 => x"b2",
          4226 => x"76",
          4227 => x"3f",
          4228 => x"08",
          4229 => x"ec",
          4230 => x"bd",
          4231 => x"82",
          4232 => x"27",
          4233 => x"16",
          4234 => x"ec",
          4235 => x"38",
          4236 => x"39",
          4237 => x"55",
          4238 => x"52",
          4239 => x"d5",
          4240 => x"ec",
          4241 => x"0c",
          4242 => x"0c",
          4243 => x"53",
          4244 => x"80",
          4245 => x"85",
          4246 => x"94",
          4247 => x"2a",
          4248 => x"0c",
          4249 => x"06",
          4250 => x"9c",
          4251 => x"58",
          4252 => x"ec",
          4253 => x"0d",
          4254 => x"0d",
          4255 => x"90",
          4256 => x"05",
          4257 => x"f0",
          4258 => x"27",
          4259 => x"0b",
          4260 => x"98",
          4261 => x"84",
          4262 => x"2e",
          4263 => x"76",
          4264 => x"58",
          4265 => x"38",
          4266 => x"15",
          4267 => x"08",
          4268 => x"38",
          4269 => x"88",
          4270 => x"53",
          4271 => x"81",
          4272 => x"c0",
          4273 => x"22",
          4274 => x"89",
          4275 => x"72",
          4276 => x"74",
          4277 => x"f3",
          4278 => x"8c",
          4279 => x"82",
          4280 => x"82",
          4281 => x"27",
          4282 => x"81",
          4283 => x"ec",
          4284 => x"80",
          4285 => x"16",
          4286 => x"ec",
          4287 => x"ca",
          4288 => x"38",
          4289 => x"0c",
          4290 => x"dd",
          4291 => x"08",
          4292 => x"f9",
          4293 => x"8c",
          4294 => x"87",
          4295 => x"ec",
          4296 => x"80",
          4297 => x"55",
          4298 => x"08",
          4299 => x"38",
          4300 => x"8c",
          4301 => x"2e",
          4302 => x"8c",
          4303 => x"75",
          4304 => x"3f",
          4305 => x"08",
          4306 => x"94",
          4307 => x"52",
          4308 => x"c1",
          4309 => x"ec",
          4310 => x"0c",
          4311 => x"0c",
          4312 => x"05",
          4313 => x"80",
          4314 => x"8c",
          4315 => x"3d",
          4316 => x"3d",
          4317 => x"71",
          4318 => x"57",
          4319 => x"51",
          4320 => x"82",
          4321 => x"54",
          4322 => x"08",
          4323 => x"82",
          4324 => x"56",
          4325 => x"52",
          4326 => x"83",
          4327 => x"ec",
          4328 => x"8c",
          4329 => x"d2",
          4330 => x"ec",
          4331 => x"08",
          4332 => x"54",
          4333 => x"e5",
          4334 => x"06",
          4335 => x"58",
          4336 => x"08",
          4337 => x"38",
          4338 => x"75",
          4339 => x"80",
          4340 => x"81",
          4341 => x"7a",
          4342 => x"06",
          4343 => x"39",
          4344 => x"08",
          4345 => x"76",
          4346 => x"3f",
          4347 => x"08",
          4348 => x"ec",
          4349 => x"ff",
          4350 => x"84",
          4351 => x"06",
          4352 => x"54",
          4353 => x"ec",
          4354 => x"0d",
          4355 => x"0d",
          4356 => x"52",
          4357 => x"3f",
          4358 => x"08",
          4359 => x"06",
          4360 => x"51",
          4361 => x"83",
          4362 => x"06",
          4363 => x"14",
          4364 => x"3f",
          4365 => x"08",
          4366 => x"07",
          4367 => x"8c",
          4368 => x"3d",
          4369 => x"3d",
          4370 => x"70",
          4371 => x"06",
          4372 => x"53",
          4373 => x"ed",
          4374 => x"33",
          4375 => x"83",
          4376 => x"06",
          4377 => x"90",
          4378 => x"15",
          4379 => x"3f",
          4380 => x"04",
          4381 => x"7b",
          4382 => x"84",
          4383 => x"58",
          4384 => x"80",
          4385 => x"38",
          4386 => x"52",
          4387 => x"8f",
          4388 => x"ec",
          4389 => x"8c",
          4390 => x"f5",
          4391 => x"08",
          4392 => x"53",
          4393 => x"84",
          4394 => x"39",
          4395 => x"70",
          4396 => x"81",
          4397 => x"51",
          4398 => x"16",
          4399 => x"ec",
          4400 => x"81",
          4401 => x"38",
          4402 => x"ae",
          4403 => x"81",
          4404 => x"54",
          4405 => x"2e",
          4406 => x"8f",
          4407 => x"82",
          4408 => x"76",
          4409 => x"54",
          4410 => x"09",
          4411 => x"38",
          4412 => x"7a",
          4413 => x"80",
          4414 => x"fa",
          4415 => x"8c",
          4416 => x"82",
          4417 => x"89",
          4418 => x"08",
          4419 => x"86",
          4420 => x"98",
          4421 => x"82",
          4422 => x"8b",
          4423 => x"fb",
          4424 => x"70",
          4425 => x"81",
          4426 => x"fc",
          4427 => x"8c",
          4428 => x"82",
          4429 => x"b4",
          4430 => x"08",
          4431 => x"ec",
          4432 => x"8c",
          4433 => x"82",
          4434 => x"a0",
          4435 => x"82",
          4436 => x"52",
          4437 => x"51",
          4438 => x"8b",
          4439 => x"52",
          4440 => x"51",
          4441 => x"81",
          4442 => x"34",
          4443 => x"ec",
          4444 => x"0d",
          4445 => x"0d",
          4446 => x"98",
          4447 => x"70",
          4448 => x"ec",
          4449 => x"8c",
          4450 => x"38",
          4451 => x"53",
          4452 => x"81",
          4453 => x"34",
          4454 => x"04",
          4455 => x"78",
          4456 => x"80",
          4457 => x"34",
          4458 => x"80",
          4459 => x"38",
          4460 => x"18",
          4461 => x"9c",
          4462 => x"70",
          4463 => x"56",
          4464 => x"a0",
          4465 => x"71",
          4466 => x"81",
          4467 => x"81",
          4468 => x"89",
          4469 => x"06",
          4470 => x"73",
          4471 => x"55",
          4472 => x"55",
          4473 => x"81",
          4474 => x"81",
          4475 => x"74",
          4476 => x"75",
          4477 => x"52",
          4478 => x"13",
          4479 => x"08",
          4480 => x"33",
          4481 => x"9c",
          4482 => x"11",
          4483 => x"8a",
          4484 => x"ec",
          4485 => x"96",
          4486 => x"e7",
          4487 => x"ec",
          4488 => x"23",
          4489 => x"e7",
          4490 => x"8c",
          4491 => x"17",
          4492 => x"0d",
          4493 => x"0d",
          4494 => x"5e",
          4495 => x"70",
          4496 => x"55",
          4497 => x"83",
          4498 => x"73",
          4499 => x"91",
          4500 => x"2e",
          4501 => x"1d",
          4502 => x"0c",
          4503 => x"15",
          4504 => x"70",
          4505 => x"56",
          4506 => x"09",
          4507 => x"38",
          4508 => x"80",
          4509 => x"30",
          4510 => x"78",
          4511 => x"54",
          4512 => x"73",
          4513 => x"60",
          4514 => x"54",
          4515 => x"96",
          4516 => x"0b",
          4517 => x"80",
          4518 => x"f6",
          4519 => x"8c",
          4520 => x"85",
          4521 => x"3d",
          4522 => x"5c",
          4523 => x"53",
          4524 => x"51",
          4525 => x"80",
          4526 => x"88",
          4527 => x"5c",
          4528 => x"09",
          4529 => x"d4",
          4530 => x"70",
          4531 => x"71",
          4532 => x"30",
          4533 => x"73",
          4534 => x"51",
          4535 => x"57",
          4536 => x"38",
          4537 => x"75",
          4538 => x"17",
          4539 => x"75",
          4540 => x"30",
          4541 => x"51",
          4542 => x"80",
          4543 => x"38",
          4544 => x"87",
          4545 => x"26",
          4546 => x"77",
          4547 => x"a4",
          4548 => x"27",
          4549 => x"a0",
          4550 => x"39",
          4551 => x"33",
          4552 => x"57",
          4553 => x"27",
          4554 => x"75",
          4555 => x"30",
          4556 => x"32",
          4557 => x"80",
          4558 => x"25",
          4559 => x"56",
          4560 => x"80",
          4561 => x"84",
          4562 => x"58",
          4563 => x"70",
          4564 => x"55",
          4565 => x"09",
          4566 => x"38",
          4567 => x"80",
          4568 => x"30",
          4569 => x"77",
          4570 => x"54",
          4571 => x"81",
          4572 => x"ae",
          4573 => x"06",
          4574 => x"54",
          4575 => x"74",
          4576 => x"80",
          4577 => x"7b",
          4578 => x"30",
          4579 => x"70",
          4580 => x"25",
          4581 => x"07",
          4582 => x"51",
          4583 => x"a7",
          4584 => x"8b",
          4585 => x"39",
          4586 => x"54",
          4587 => x"8c",
          4588 => x"ff",
          4589 => x"bc",
          4590 => x"54",
          4591 => x"e1",
          4592 => x"ec",
          4593 => x"b2",
          4594 => x"70",
          4595 => x"71",
          4596 => x"54",
          4597 => x"82",
          4598 => x"80",
          4599 => x"38",
          4600 => x"76",
          4601 => x"df",
          4602 => x"54",
          4603 => x"81",
          4604 => x"55",
          4605 => x"34",
          4606 => x"52",
          4607 => x"51",
          4608 => x"82",
          4609 => x"bf",
          4610 => x"16",
          4611 => x"26",
          4612 => x"16",
          4613 => x"06",
          4614 => x"17",
          4615 => x"34",
          4616 => x"fd",
          4617 => x"19",
          4618 => x"80",
          4619 => x"79",
          4620 => x"81",
          4621 => x"81",
          4622 => x"85",
          4623 => x"54",
          4624 => x"8f",
          4625 => x"86",
          4626 => x"39",
          4627 => x"f3",
          4628 => x"73",
          4629 => x"80",
          4630 => x"52",
          4631 => x"ce",
          4632 => x"ec",
          4633 => x"8c",
          4634 => x"d7",
          4635 => x"08",
          4636 => x"e6",
          4637 => x"8c",
          4638 => x"82",
          4639 => x"80",
          4640 => x"1b",
          4641 => x"55",
          4642 => x"2e",
          4643 => x"8b",
          4644 => x"06",
          4645 => x"1c",
          4646 => x"33",
          4647 => x"70",
          4648 => x"55",
          4649 => x"38",
          4650 => x"52",
          4651 => x"9f",
          4652 => x"ec",
          4653 => x"8b",
          4654 => x"7a",
          4655 => x"3f",
          4656 => x"75",
          4657 => x"57",
          4658 => x"2e",
          4659 => x"84",
          4660 => x"06",
          4661 => x"75",
          4662 => x"81",
          4663 => x"2a",
          4664 => x"73",
          4665 => x"38",
          4666 => x"54",
          4667 => x"fb",
          4668 => x"80",
          4669 => x"34",
          4670 => x"c1",
          4671 => x"06",
          4672 => x"38",
          4673 => x"39",
          4674 => x"70",
          4675 => x"54",
          4676 => x"86",
          4677 => x"84",
          4678 => x"06",
          4679 => x"73",
          4680 => x"38",
          4681 => x"83",
          4682 => x"b4",
          4683 => x"51",
          4684 => x"82",
          4685 => x"88",
          4686 => x"ea",
          4687 => x"8c",
          4688 => x"3d",
          4689 => x"3d",
          4690 => x"ff",
          4691 => x"71",
          4692 => x"5c",
          4693 => x"80",
          4694 => x"38",
          4695 => x"05",
          4696 => x"a0",
          4697 => x"71",
          4698 => x"38",
          4699 => x"71",
          4700 => x"81",
          4701 => x"38",
          4702 => x"11",
          4703 => x"06",
          4704 => x"70",
          4705 => x"38",
          4706 => x"81",
          4707 => x"05",
          4708 => x"76",
          4709 => x"38",
          4710 => x"fc",
          4711 => x"77",
          4712 => x"57",
          4713 => x"05",
          4714 => x"70",
          4715 => x"33",
          4716 => x"53",
          4717 => x"99",
          4718 => x"e0",
          4719 => x"ff",
          4720 => x"ff",
          4721 => x"70",
          4722 => x"38",
          4723 => x"81",
          4724 => x"51",
          4725 => x"9f",
          4726 => x"72",
          4727 => x"81",
          4728 => x"70",
          4729 => x"72",
          4730 => x"32",
          4731 => x"72",
          4732 => x"73",
          4733 => x"53",
          4734 => x"70",
          4735 => x"38",
          4736 => x"19",
          4737 => x"75",
          4738 => x"38",
          4739 => x"83",
          4740 => x"74",
          4741 => x"59",
          4742 => x"39",
          4743 => x"33",
          4744 => x"8c",
          4745 => x"3d",
          4746 => x"3d",
          4747 => x"80",
          4748 => x"34",
          4749 => x"17",
          4750 => x"75",
          4751 => x"3f",
          4752 => x"8c",
          4753 => x"80",
          4754 => x"16",
          4755 => x"3f",
          4756 => x"08",
          4757 => x"06",
          4758 => x"73",
          4759 => x"2e",
          4760 => x"80",
          4761 => x"0b",
          4762 => x"56",
          4763 => x"e9",
          4764 => x"06",
          4765 => x"57",
          4766 => x"32",
          4767 => x"80",
          4768 => x"51",
          4769 => x"8a",
          4770 => x"e8",
          4771 => x"06",
          4772 => x"53",
          4773 => x"52",
          4774 => x"51",
          4775 => x"82",
          4776 => x"55",
          4777 => x"08",
          4778 => x"38",
          4779 => x"fb",
          4780 => x"86",
          4781 => x"97",
          4782 => x"ec",
          4783 => x"8c",
          4784 => x"2e",
          4785 => x"55",
          4786 => x"ec",
          4787 => x"0d",
          4788 => x"0d",
          4789 => x"05",
          4790 => x"33",
          4791 => x"75",
          4792 => x"fc",
          4793 => x"8c",
          4794 => x"8b",
          4795 => x"82",
          4796 => x"24",
          4797 => x"82",
          4798 => x"84",
          4799 => x"88",
          4800 => x"55",
          4801 => x"73",
          4802 => x"e6",
          4803 => x"0c",
          4804 => x"06",
          4805 => x"57",
          4806 => x"ae",
          4807 => x"33",
          4808 => x"3f",
          4809 => x"08",
          4810 => x"70",
          4811 => x"55",
          4812 => x"76",
          4813 => x"b8",
          4814 => x"2a",
          4815 => x"51",
          4816 => x"72",
          4817 => x"86",
          4818 => x"74",
          4819 => x"15",
          4820 => x"81",
          4821 => x"d7",
          4822 => x"8c",
          4823 => x"ff",
          4824 => x"06",
          4825 => x"56",
          4826 => x"38",
          4827 => x"8f",
          4828 => x"2a",
          4829 => x"51",
          4830 => x"72",
          4831 => x"80",
          4832 => x"52",
          4833 => x"3f",
          4834 => x"08",
          4835 => x"57",
          4836 => x"09",
          4837 => x"e2",
          4838 => x"74",
          4839 => x"56",
          4840 => x"33",
          4841 => x"72",
          4842 => x"38",
          4843 => x"51",
          4844 => x"82",
          4845 => x"57",
          4846 => x"84",
          4847 => x"ff",
          4848 => x"56",
          4849 => x"25",
          4850 => x"0b",
          4851 => x"56",
          4852 => x"05",
          4853 => x"83",
          4854 => x"2e",
          4855 => x"52",
          4856 => x"c6",
          4857 => x"ec",
          4858 => x"06",
          4859 => x"27",
          4860 => x"16",
          4861 => x"27",
          4862 => x"56",
          4863 => x"84",
          4864 => x"56",
          4865 => x"84",
          4866 => x"14",
          4867 => x"3f",
          4868 => x"08",
          4869 => x"06",
          4870 => x"80",
          4871 => x"06",
          4872 => x"80",
          4873 => x"db",
          4874 => x"8c",
          4875 => x"ff",
          4876 => x"77",
          4877 => x"d8",
          4878 => x"de",
          4879 => x"ec",
          4880 => x"9c",
          4881 => x"c4",
          4882 => x"15",
          4883 => x"14",
          4884 => x"70",
          4885 => x"51",
          4886 => x"56",
          4887 => x"84",
          4888 => x"81",
          4889 => x"71",
          4890 => x"16",
          4891 => x"53",
          4892 => x"23",
          4893 => x"8b",
          4894 => x"73",
          4895 => x"80",
          4896 => x"8d",
          4897 => x"39",
          4898 => x"51",
          4899 => x"82",
          4900 => x"53",
          4901 => x"08",
          4902 => x"72",
          4903 => x"8d",
          4904 => x"ce",
          4905 => x"14",
          4906 => x"3f",
          4907 => x"08",
          4908 => x"06",
          4909 => x"38",
          4910 => x"51",
          4911 => x"82",
          4912 => x"55",
          4913 => x"51",
          4914 => x"82",
          4915 => x"83",
          4916 => x"53",
          4917 => x"80",
          4918 => x"38",
          4919 => x"78",
          4920 => x"2a",
          4921 => x"78",
          4922 => x"86",
          4923 => x"22",
          4924 => x"31",
          4925 => x"be",
          4926 => x"ec",
          4927 => x"8c",
          4928 => x"2e",
          4929 => x"82",
          4930 => x"80",
          4931 => x"f5",
          4932 => x"83",
          4933 => x"ff",
          4934 => x"38",
          4935 => x"9f",
          4936 => x"38",
          4937 => x"39",
          4938 => x"80",
          4939 => x"38",
          4940 => x"98",
          4941 => x"a0",
          4942 => x"1c",
          4943 => x"0c",
          4944 => x"17",
          4945 => x"76",
          4946 => x"81",
          4947 => x"80",
          4948 => x"d9",
          4949 => x"8c",
          4950 => x"ff",
          4951 => x"8d",
          4952 => x"8e",
          4953 => x"8a",
          4954 => x"14",
          4955 => x"3f",
          4956 => x"08",
          4957 => x"74",
          4958 => x"a2",
          4959 => x"79",
          4960 => x"ee",
          4961 => x"a8",
          4962 => x"15",
          4963 => x"2e",
          4964 => x"10",
          4965 => x"2a",
          4966 => x"05",
          4967 => x"ff",
          4968 => x"53",
          4969 => x"9c",
          4970 => x"81",
          4971 => x"0b",
          4972 => x"ff",
          4973 => x"0c",
          4974 => x"84",
          4975 => x"83",
          4976 => x"06",
          4977 => x"80",
          4978 => x"d8",
          4979 => x"8c",
          4980 => x"ff",
          4981 => x"72",
          4982 => x"81",
          4983 => x"38",
          4984 => x"73",
          4985 => x"3f",
          4986 => x"08",
          4987 => x"82",
          4988 => x"84",
          4989 => x"b2",
          4990 => x"87",
          4991 => x"ec",
          4992 => x"ff",
          4993 => x"82",
          4994 => x"09",
          4995 => x"c8",
          4996 => x"51",
          4997 => x"82",
          4998 => x"84",
          4999 => x"d2",
          5000 => x"06",
          5001 => x"98",
          5002 => x"ee",
          5003 => x"ec",
          5004 => x"85",
          5005 => x"09",
          5006 => x"38",
          5007 => x"51",
          5008 => x"82",
          5009 => x"90",
          5010 => x"a0",
          5011 => x"ca",
          5012 => x"ec",
          5013 => x"0c",
          5014 => x"82",
          5015 => x"81",
          5016 => x"82",
          5017 => x"72",
          5018 => x"80",
          5019 => x"0c",
          5020 => x"82",
          5021 => x"90",
          5022 => x"fb",
          5023 => x"54",
          5024 => x"80",
          5025 => x"73",
          5026 => x"80",
          5027 => x"72",
          5028 => x"80",
          5029 => x"86",
          5030 => x"15",
          5031 => x"71",
          5032 => x"81",
          5033 => x"81",
          5034 => x"d0",
          5035 => x"8c",
          5036 => x"06",
          5037 => x"38",
          5038 => x"54",
          5039 => x"80",
          5040 => x"71",
          5041 => x"82",
          5042 => x"87",
          5043 => x"fa",
          5044 => x"ab",
          5045 => x"58",
          5046 => x"05",
          5047 => x"e6",
          5048 => x"80",
          5049 => x"ec",
          5050 => x"38",
          5051 => x"08",
          5052 => x"8d",
          5053 => x"08",
          5054 => x"80",
          5055 => x"80",
          5056 => x"54",
          5057 => x"84",
          5058 => x"34",
          5059 => x"75",
          5060 => x"2e",
          5061 => x"53",
          5062 => x"53",
          5063 => x"f7",
          5064 => x"8c",
          5065 => x"73",
          5066 => x"0c",
          5067 => x"04",
          5068 => x"67",
          5069 => x"80",
          5070 => x"59",
          5071 => x"78",
          5072 => x"c8",
          5073 => x"06",
          5074 => x"3d",
          5075 => x"99",
          5076 => x"52",
          5077 => x"3f",
          5078 => x"08",
          5079 => x"ec",
          5080 => x"38",
          5081 => x"52",
          5082 => x"52",
          5083 => x"3f",
          5084 => x"08",
          5085 => x"ec",
          5086 => x"02",
          5087 => x"33",
          5088 => x"55",
          5089 => x"25",
          5090 => x"55",
          5091 => x"54",
          5092 => x"81",
          5093 => x"80",
          5094 => x"74",
          5095 => x"81",
          5096 => x"75",
          5097 => x"3f",
          5098 => x"08",
          5099 => x"02",
          5100 => x"91",
          5101 => x"81",
          5102 => x"82",
          5103 => x"06",
          5104 => x"80",
          5105 => x"88",
          5106 => x"39",
          5107 => x"58",
          5108 => x"38",
          5109 => x"70",
          5110 => x"54",
          5111 => x"81",
          5112 => x"52",
          5113 => x"a5",
          5114 => x"ec",
          5115 => x"88",
          5116 => x"62",
          5117 => x"d4",
          5118 => x"54",
          5119 => x"15",
          5120 => x"62",
          5121 => x"e8",
          5122 => x"52",
          5123 => x"51",
          5124 => x"7a",
          5125 => x"83",
          5126 => x"80",
          5127 => x"38",
          5128 => x"08",
          5129 => x"53",
          5130 => x"3d",
          5131 => x"dd",
          5132 => x"8c",
          5133 => x"82",
          5134 => x"82",
          5135 => x"39",
          5136 => x"38",
          5137 => x"33",
          5138 => x"70",
          5139 => x"55",
          5140 => x"2e",
          5141 => x"55",
          5142 => x"77",
          5143 => x"81",
          5144 => x"73",
          5145 => x"38",
          5146 => x"54",
          5147 => x"a0",
          5148 => x"82",
          5149 => x"52",
          5150 => x"a3",
          5151 => x"ec",
          5152 => x"18",
          5153 => x"55",
          5154 => x"ec",
          5155 => x"38",
          5156 => x"70",
          5157 => x"54",
          5158 => x"86",
          5159 => x"c0",
          5160 => x"b0",
          5161 => x"1b",
          5162 => x"1b",
          5163 => x"70",
          5164 => x"d9",
          5165 => x"ec",
          5166 => x"ec",
          5167 => x"0c",
          5168 => x"52",
          5169 => x"3f",
          5170 => x"08",
          5171 => x"08",
          5172 => x"77",
          5173 => x"86",
          5174 => x"1a",
          5175 => x"1a",
          5176 => x"91",
          5177 => x"0b",
          5178 => x"80",
          5179 => x"0c",
          5180 => x"70",
          5181 => x"54",
          5182 => x"81",
          5183 => x"8c",
          5184 => x"2e",
          5185 => x"82",
          5186 => x"94",
          5187 => x"17",
          5188 => x"2b",
          5189 => x"57",
          5190 => x"52",
          5191 => x"9f",
          5192 => x"ec",
          5193 => x"8c",
          5194 => x"26",
          5195 => x"55",
          5196 => x"08",
          5197 => x"81",
          5198 => x"79",
          5199 => x"31",
          5200 => x"70",
          5201 => x"25",
          5202 => x"76",
          5203 => x"81",
          5204 => x"55",
          5205 => x"38",
          5206 => x"0c",
          5207 => x"75",
          5208 => x"54",
          5209 => x"a2",
          5210 => x"7a",
          5211 => x"3f",
          5212 => x"08",
          5213 => x"55",
          5214 => x"89",
          5215 => x"ec",
          5216 => x"1a",
          5217 => x"80",
          5218 => x"54",
          5219 => x"ec",
          5220 => x"0d",
          5221 => x"0d",
          5222 => x"64",
          5223 => x"59",
          5224 => x"90",
          5225 => x"52",
          5226 => x"cf",
          5227 => x"ec",
          5228 => x"8c",
          5229 => x"38",
          5230 => x"55",
          5231 => x"86",
          5232 => x"82",
          5233 => x"19",
          5234 => x"55",
          5235 => x"80",
          5236 => x"38",
          5237 => x"0b",
          5238 => x"82",
          5239 => x"39",
          5240 => x"1a",
          5241 => x"82",
          5242 => x"19",
          5243 => x"08",
          5244 => x"7c",
          5245 => x"74",
          5246 => x"2e",
          5247 => x"94",
          5248 => x"83",
          5249 => x"56",
          5250 => x"38",
          5251 => x"22",
          5252 => x"89",
          5253 => x"55",
          5254 => x"75",
          5255 => x"19",
          5256 => x"39",
          5257 => x"52",
          5258 => x"93",
          5259 => x"ec",
          5260 => x"75",
          5261 => x"38",
          5262 => x"ff",
          5263 => x"98",
          5264 => x"19",
          5265 => x"51",
          5266 => x"82",
          5267 => x"80",
          5268 => x"38",
          5269 => x"08",
          5270 => x"2a",
          5271 => x"80",
          5272 => x"38",
          5273 => x"8a",
          5274 => x"5c",
          5275 => x"27",
          5276 => x"7a",
          5277 => x"54",
          5278 => x"52",
          5279 => x"51",
          5280 => x"82",
          5281 => x"fe",
          5282 => x"83",
          5283 => x"56",
          5284 => x"9f",
          5285 => x"08",
          5286 => x"74",
          5287 => x"38",
          5288 => x"b4",
          5289 => x"16",
          5290 => x"89",
          5291 => x"51",
          5292 => x"77",
          5293 => x"b9",
          5294 => x"1a",
          5295 => x"08",
          5296 => x"84",
          5297 => x"57",
          5298 => x"27",
          5299 => x"56",
          5300 => x"52",
          5301 => x"c7",
          5302 => x"ec",
          5303 => x"38",
          5304 => x"19",
          5305 => x"06",
          5306 => x"52",
          5307 => x"a2",
          5308 => x"31",
          5309 => x"7f",
          5310 => x"94",
          5311 => x"94",
          5312 => x"5c",
          5313 => x"80",
          5314 => x"8c",
          5315 => x"3d",
          5316 => x"3d",
          5317 => x"65",
          5318 => x"5d",
          5319 => x"0c",
          5320 => x"05",
          5321 => x"f6",
          5322 => x"8c",
          5323 => x"82",
          5324 => x"8a",
          5325 => x"33",
          5326 => x"2e",
          5327 => x"56",
          5328 => x"90",
          5329 => x"81",
          5330 => x"06",
          5331 => x"87",
          5332 => x"2e",
          5333 => x"95",
          5334 => x"91",
          5335 => x"56",
          5336 => x"81",
          5337 => x"34",
          5338 => x"8e",
          5339 => x"08",
          5340 => x"56",
          5341 => x"84",
          5342 => x"5c",
          5343 => x"82",
          5344 => x"18",
          5345 => x"ff",
          5346 => x"74",
          5347 => x"7e",
          5348 => x"ff",
          5349 => x"2a",
          5350 => x"7a",
          5351 => x"8c",
          5352 => x"08",
          5353 => x"38",
          5354 => x"39",
          5355 => x"52",
          5356 => x"e7",
          5357 => x"ec",
          5358 => x"8c",
          5359 => x"2e",
          5360 => x"74",
          5361 => x"91",
          5362 => x"2e",
          5363 => x"74",
          5364 => x"88",
          5365 => x"38",
          5366 => x"0c",
          5367 => x"15",
          5368 => x"08",
          5369 => x"06",
          5370 => x"51",
          5371 => x"82",
          5372 => x"fe",
          5373 => x"18",
          5374 => x"51",
          5375 => x"82",
          5376 => x"80",
          5377 => x"38",
          5378 => x"08",
          5379 => x"2a",
          5380 => x"80",
          5381 => x"38",
          5382 => x"8a",
          5383 => x"5b",
          5384 => x"27",
          5385 => x"7b",
          5386 => x"54",
          5387 => x"52",
          5388 => x"51",
          5389 => x"82",
          5390 => x"fe",
          5391 => x"b0",
          5392 => x"31",
          5393 => x"79",
          5394 => x"84",
          5395 => x"16",
          5396 => x"89",
          5397 => x"52",
          5398 => x"cc",
          5399 => x"55",
          5400 => x"16",
          5401 => x"2b",
          5402 => x"39",
          5403 => x"94",
          5404 => x"93",
          5405 => x"cd",
          5406 => x"8c",
          5407 => x"e3",
          5408 => x"b0",
          5409 => x"76",
          5410 => x"94",
          5411 => x"ff",
          5412 => x"71",
          5413 => x"7b",
          5414 => x"38",
          5415 => x"18",
          5416 => x"51",
          5417 => x"82",
          5418 => x"fd",
          5419 => x"53",
          5420 => x"18",
          5421 => x"06",
          5422 => x"51",
          5423 => x"7e",
          5424 => x"83",
          5425 => x"76",
          5426 => x"17",
          5427 => x"1e",
          5428 => x"18",
          5429 => x"0c",
          5430 => x"58",
          5431 => x"74",
          5432 => x"38",
          5433 => x"8c",
          5434 => x"90",
          5435 => x"33",
          5436 => x"55",
          5437 => x"34",
          5438 => x"82",
          5439 => x"90",
          5440 => x"f8",
          5441 => x"8b",
          5442 => x"53",
          5443 => x"f2",
          5444 => x"8c",
          5445 => x"82",
          5446 => x"80",
          5447 => x"16",
          5448 => x"2a",
          5449 => x"51",
          5450 => x"80",
          5451 => x"38",
          5452 => x"52",
          5453 => x"e7",
          5454 => x"ec",
          5455 => x"8c",
          5456 => x"d4",
          5457 => x"08",
          5458 => x"a0",
          5459 => x"73",
          5460 => x"88",
          5461 => x"74",
          5462 => x"51",
          5463 => x"8c",
          5464 => x"9c",
          5465 => x"fb",
          5466 => x"b2",
          5467 => x"15",
          5468 => x"3f",
          5469 => x"15",
          5470 => x"3f",
          5471 => x"0b",
          5472 => x"78",
          5473 => x"3f",
          5474 => x"08",
          5475 => x"81",
          5476 => x"57",
          5477 => x"34",
          5478 => x"ec",
          5479 => x"0d",
          5480 => x"0d",
          5481 => x"54",
          5482 => x"82",
          5483 => x"53",
          5484 => x"08",
          5485 => x"3d",
          5486 => x"73",
          5487 => x"3f",
          5488 => x"08",
          5489 => x"ec",
          5490 => x"82",
          5491 => x"74",
          5492 => x"8c",
          5493 => x"3d",
          5494 => x"3d",
          5495 => x"51",
          5496 => x"8b",
          5497 => x"82",
          5498 => x"24",
          5499 => x"8c",
          5500 => x"8d",
          5501 => x"52",
          5502 => x"ec",
          5503 => x"0d",
          5504 => x"0d",
          5505 => x"3d",
          5506 => x"94",
          5507 => x"c1",
          5508 => x"ec",
          5509 => x"8c",
          5510 => x"e0",
          5511 => x"63",
          5512 => x"d4",
          5513 => x"8d",
          5514 => x"ec",
          5515 => x"8c",
          5516 => x"38",
          5517 => x"05",
          5518 => x"2b",
          5519 => x"80",
          5520 => x"76",
          5521 => x"0c",
          5522 => x"02",
          5523 => x"70",
          5524 => x"81",
          5525 => x"56",
          5526 => x"9e",
          5527 => x"53",
          5528 => x"db",
          5529 => x"8c",
          5530 => x"15",
          5531 => x"82",
          5532 => x"84",
          5533 => x"06",
          5534 => x"55",
          5535 => x"ec",
          5536 => x"0d",
          5537 => x"0d",
          5538 => x"5b",
          5539 => x"80",
          5540 => x"ff",
          5541 => x"9f",
          5542 => x"b5",
          5543 => x"ec",
          5544 => x"8c",
          5545 => x"fc",
          5546 => x"7a",
          5547 => x"08",
          5548 => x"64",
          5549 => x"2e",
          5550 => x"a0",
          5551 => x"70",
          5552 => x"ea",
          5553 => x"ec",
          5554 => x"8c",
          5555 => x"d4",
          5556 => x"7b",
          5557 => x"3f",
          5558 => x"08",
          5559 => x"ec",
          5560 => x"38",
          5561 => x"51",
          5562 => x"82",
          5563 => x"45",
          5564 => x"51",
          5565 => x"82",
          5566 => x"57",
          5567 => x"08",
          5568 => x"80",
          5569 => x"da",
          5570 => x"8c",
          5571 => x"82",
          5572 => x"a4",
          5573 => x"7b",
          5574 => x"3f",
          5575 => x"ec",
          5576 => x"38",
          5577 => x"51",
          5578 => x"82",
          5579 => x"57",
          5580 => x"08",
          5581 => x"38",
          5582 => x"09",
          5583 => x"38",
          5584 => x"e0",
          5585 => x"dc",
          5586 => x"ff",
          5587 => x"74",
          5588 => x"3f",
          5589 => x"78",
          5590 => x"33",
          5591 => x"56",
          5592 => x"91",
          5593 => x"05",
          5594 => x"81",
          5595 => x"56",
          5596 => x"f5",
          5597 => x"54",
          5598 => x"81",
          5599 => x"80",
          5600 => x"78",
          5601 => x"55",
          5602 => x"11",
          5603 => x"18",
          5604 => x"58",
          5605 => x"34",
          5606 => x"ff",
          5607 => x"55",
          5608 => x"34",
          5609 => x"77",
          5610 => x"81",
          5611 => x"ff",
          5612 => x"55",
          5613 => x"34",
          5614 => x"8d",
          5615 => x"84",
          5616 => x"ac",
          5617 => x"70",
          5618 => x"56",
          5619 => x"76",
          5620 => x"81",
          5621 => x"70",
          5622 => x"56",
          5623 => x"82",
          5624 => x"78",
          5625 => x"80",
          5626 => x"27",
          5627 => x"19",
          5628 => x"7a",
          5629 => x"5c",
          5630 => x"55",
          5631 => x"7a",
          5632 => x"5c",
          5633 => x"2e",
          5634 => x"85",
          5635 => x"94",
          5636 => x"81",
          5637 => x"73",
          5638 => x"81",
          5639 => x"7a",
          5640 => x"38",
          5641 => x"76",
          5642 => x"0c",
          5643 => x"04",
          5644 => x"7b",
          5645 => x"fc",
          5646 => x"53",
          5647 => x"bb",
          5648 => x"ec",
          5649 => x"8c",
          5650 => x"fa",
          5651 => x"33",
          5652 => x"f2",
          5653 => x"08",
          5654 => x"27",
          5655 => x"15",
          5656 => x"2a",
          5657 => x"51",
          5658 => x"83",
          5659 => x"94",
          5660 => x"80",
          5661 => x"0c",
          5662 => x"2e",
          5663 => x"79",
          5664 => x"70",
          5665 => x"51",
          5666 => x"2e",
          5667 => x"52",
          5668 => x"ff",
          5669 => x"82",
          5670 => x"ff",
          5671 => x"70",
          5672 => x"ff",
          5673 => x"82",
          5674 => x"73",
          5675 => x"76",
          5676 => x"06",
          5677 => x"0c",
          5678 => x"98",
          5679 => x"58",
          5680 => x"39",
          5681 => x"54",
          5682 => x"73",
          5683 => x"cd",
          5684 => x"8c",
          5685 => x"82",
          5686 => x"81",
          5687 => x"38",
          5688 => x"08",
          5689 => x"9b",
          5690 => x"ec",
          5691 => x"0c",
          5692 => x"0c",
          5693 => x"81",
          5694 => x"76",
          5695 => x"38",
          5696 => x"94",
          5697 => x"94",
          5698 => x"16",
          5699 => x"2a",
          5700 => x"51",
          5701 => x"72",
          5702 => x"38",
          5703 => x"51",
          5704 => x"82",
          5705 => x"54",
          5706 => x"08",
          5707 => x"8c",
          5708 => x"a7",
          5709 => x"74",
          5710 => x"3f",
          5711 => x"08",
          5712 => x"2e",
          5713 => x"74",
          5714 => x"79",
          5715 => x"14",
          5716 => x"38",
          5717 => x"0c",
          5718 => x"94",
          5719 => x"94",
          5720 => x"83",
          5721 => x"72",
          5722 => x"38",
          5723 => x"51",
          5724 => x"82",
          5725 => x"94",
          5726 => x"91",
          5727 => x"53",
          5728 => x"81",
          5729 => x"34",
          5730 => x"39",
          5731 => x"82",
          5732 => x"05",
          5733 => x"08",
          5734 => x"08",
          5735 => x"38",
          5736 => x"0c",
          5737 => x"80",
          5738 => x"72",
          5739 => x"73",
          5740 => x"53",
          5741 => x"8c",
          5742 => x"16",
          5743 => x"38",
          5744 => x"0c",
          5745 => x"82",
          5746 => x"8b",
          5747 => x"f9",
          5748 => x"56",
          5749 => x"80",
          5750 => x"38",
          5751 => x"3d",
          5752 => x"8a",
          5753 => x"51",
          5754 => x"82",
          5755 => x"55",
          5756 => x"08",
          5757 => x"77",
          5758 => x"52",
          5759 => x"b5",
          5760 => x"ec",
          5761 => x"8c",
          5762 => x"c3",
          5763 => x"33",
          5764 => x"55",
          5765 => x"24",
          5766 => x"16",
          5767 => x"2a",
          5768 => x"51",
          5769 => x"80",
          5770 => x"9c",
          5771 => x"77",
          5772 => x"3f",
          5773 => x"08",
          5774 => x"77",
          5775 => x"22",
          5776 => x"74",
          5777 => x"ce",
          5778 => x"8c",
          5779 => x"74",
          5780 => x"81",
          5781 => x"85",
          5782 => x"74",
          5783 => x"38",
          5784 => x"74",
          5785 => x"8c",
          5786 => x"3d",
          5787 => x"3d",
          5788 => x"3d",
          5789 => x"70",
          5790 => x"ff",
          5791 => x"ec",
          5792 => x"82",
          5793 => x"73",
          5794 => x"0d",
          5795 => x"0d",
          5796 => x"3d",
          5797 => x"71",
          5798 => x"e7",
          5799 => x"8c",
          5800 => x"82",
          5801 => x"80",
          5802 => x"93",
          5803 => x"ec",
          5804 => x"51",
          5805 => x"82",
          5806 => x"53",
          5807 => x"82",
          5808 => x"52",
          5809 => x"ac",
          5810 => x"ec",
          5811 => x"8c",
          5812 => x"2e",
          5813 => x"85",
          5814 => x"87",
          5815 => x"ec",
          5816 => x"74",
          5817 => x"d5",
          5818 => x"52",
          5819 => x"89",
          5820 => x"ec",
          5821 => x"70",
          5822 => x"07",
          5823 => x"82",
          5824 => x"06",
          5825 => x"54",
          5826 => x"ec",
          5827 => x"0d",
          5828 => x"0d",
          5829 => x"53",
          5830 => x"53",
          5831 => x"56",
          5832 => x"82",
          5833 => x"55",
          5834 => x"08",
          5835 => x"52",
          5836 => x"81",
          5837 => x"ec",
          5838 => x"8c",
          5839 => x"38",
          5840 => x"05",
          5841 => x"2b",
          5842 => x"80",
          5843 => x"86",
          5844 => x"76",
          5845 => x"38",
          5846 => x"51",
          5847 => x"74",
          5848 => x"0c",
          5849 => x"04",
          5850 => x"63",
          5851 => x"80",
          5852 => x"ec",
          5853 => x"3d",
          5854 => x"3f",
          5855 => x"08",
          5856 => x"ec",
          5857 => x"38",
          5858 => x"73",
          5859 => x"08",
          5860 => x"13",
          5861 => x"58",
          5862 => x"26",
          5863 => x"7c",
          5864 => x"39",
          5865 => x"cc",
          5866 => x"81",
          5867 => x"8c",
          5868 => x"33",
          5869 => x"81",
          5870 => x"06",
          5871 => x"75",
          5872 => x"52",
          5873 => x"05",
          5874 => x"3f",
          5875 => x"08",
          5876 => x"38",
          5877 => x"08",
          5878 => x"38",
          5879 => x"08",
          5880 => x"8c",
          5881 => x"80",
          5882 => x"81",
          5883 => x"59",
          5884 => x"14",
          5885 => x"ca",
          5886 => x"39",
          5887 => x"82",
          5888 => x"57",
          5889 => x"38",
          5890 => x"18",
          5891 => x"ff",
          5892 => x"82",
          5893 => x"5b",
          5894 => x"08",
          5895 => x"7c",
          5896 => x"12",
          5897 => x"52",
          5898 => x"82",
          5899 => x"06",
          5900 => x"14",
          5901 => x"cb",
          5902 => x"ec",
          5903 => x"ff",
          5904 => x"70",
          5905 => x"82",
          5906 => x"51",
          5907 => x"b4",
          5908 => x"bb",
          5909 => x"8c",
          5910 => x"0a",
          5911 => x"70",
          5912 => x"84",
          5913 => x"51",
          5914 => x"ff",
          5915 => x"56",
          5916 => x"38",
          5917 => x"7c",
          5918 => x"0c",
          5919 => x"81",
          5920 => x"74",
          5921 => x"7a",
          5922 => x"0c",
          5923 => x"04",
          5924 => x"79",
          5925 => x"05",
          5926 => x"57",
          5927 => x"82",
          5928 => x"56",
          5929 => x"08",
          5930 => x"91",
          5931 => x"75",
          5932 => x"90",
          5933 => x"81",
          5934 => x"06",
          5935 => x"87",
          5936 => x"2e",
          5937 => x"94",
          5938 => x"73",
          5939 => x"27",
          5940 => x"73",
          5941 => x"8c",
          5942 => x"88",
          5943 => x"76",
          5944 => x"3f",
          5945 => x"08",
          5946 => x"0c",
          5947 => x"39",
          5948 => x"52",
          5949 => x"bf",
          5950 => x"8c",
          5951 => x"2e",
          5952 => x"83",
          5953 => x"82",
          5954 => x"81",
          5955 => x"06",
          5956 => x"56",
          5957 => x"a0",
          5958 => x"82",
          5959 => x"98",
          5960 => x"94",
          5961 => x"08",
          5962 => x"ec",
          5963 => x"51",
          5964 => x"82",
          5965 => x"56",
          5966 => x"8c",
          5967 => x"17",
          5968 => x"07",
          5969 => x"18",
          5970 => x"2e",
          5971 => x"91",
          5972 => x"55",
          5973 => x"ec",
          5974 => x"0d",
          5975 => x"0d",
          5976 => x"3d",
          5977 => x"52",
          5978 => x"da",
          5979 => x"8c",
          5980 => x"82",
          5981 => x"81",
          5982 => x"45",
          5983 => x"52",
          5984 => x"52",
          5985 => x"3f",
          5986 => x"08",
          5987 => x"ec",
          5988 => x"38",
          5989 => x"05",
          5990 => x"2a",
          5991 => x"51",
          5992 => x"55",
          5993 => x"38",
          5994 => x"54",
          5995 => x"81",
          5996 => x"80",
          5997 => x"70",
          5998 => x"54",
          5999 => x"81",
          6000 => x"52",
          6001 => x"c5",
          6002 => x"ec",
          6003 => x"2a",
          6004 => x"51",
          6005 => x"80",
          6006 => x"38",
          6007 => x"8c",
          6008 => x"15",
          6009 => x"86",
          6010 => x"82",
          6011 => x"5c",
          6012 => x"3d",
          6013 => x"c7",
          6014 => x"8c",
          6015 => x"82",
          6016 => x"80",
          6017 => x"8c",
          6018 => x"73",
          6019 => x"3f",
          6020 => x"08",
          6021 => x"ec",
          6022 => x"87",
          6023 => x"39",
          6024 => x"08",
          6025 => x"38",
          6026 => x"08",
          6027 => x"77",
          6028 => x"3f",
          6029 => x"08",
          6030 => x"08",
          6031 => x"8c",
          6032 => x"80",
          6033 => x"55",
          6034 => x"94",
          6035 => x"2e",
          6036 => x"53",
          6037 => x"51",
          6038 => x"82",
          6039 => x"55",
          6040 => x"78",
          6041 => x"fe",
          6042 => x"ec",
          6043 => x"82",
          6044 => x"a0",
          6045 => x"e9",
          6046 => x"53",
          6047 => x"05",
          6048 => x"51",
          6049 => x"82",
          6050 => x"54",
          6051 => x"08",
          6052 => x"78",
          6053 => x"8e",
          6054 => x"58",
          6055 => x"82",
          6056 => x"54",
          6057 => x"08",
          6058 => x"54",
          6059 => x"82",
          6060 => x"84",
          6061 => x"06",
          6062 => x"02",
          6063 => x"33",
          6064 => x"81",
          6065 => x"86",
          6066 => x"f6",
          6067 => x"74",
          6068 => x"70",
          6069 => x"c3",
          6070 => x"ec",
          6071 => x"56",
          6072 => x"08",
          6073 => x"54",
          6074 => x"08",
          6075 => x"81",
          6076 => x"82",
          6077 => x"ec",
          6078 => x"09",
          6079 => x"38",
          6080 => x"b4",
          6081 => x"b0",
          6082 => x"ec",
          6083 => x"51",
          6084 => x"82",
          6085 => x"54",
          6086 => x"08",
          6087 => x"8b",
          6088 => x"b4",
          6089 => x"b7",
          6090 => x"54",
          6091 => x"15",
          6092 => x"90",
          6093 => x"34",
          6094 => x"0a",
          6095 => x"19",
          6096 => x"9f",
          6097 => x"78",
          6098 => x"51",
          6099 => x"a0",
          6100 => x"11",
          6101 => x"05",
          6102 => x"b6",
          6103 => x"ae",
          6104 => x"15",
          6105 => x"78",
          6106 => x"53",
          6107 => x"3f",
          6108 => x"0b",
          6109 => x"77",
          6110 => x"3f",
          6111 => x"08",
          6112 => x"ec",
          6113 => x"82",
          6114 => x"52",
          6115 => x"51",
          6116 => x"3f",
          6117 => x"52",
          6118 => x"aa",
          6119 => x"90",
          6120 => x"34",
          6121 => x"0b",
          6122 => x"78",
          6123 => x"b6",
          6124 => x"ec",
          6125 => x"39",
          6126 => x"52",
          6127 => x"be",
          6128 => x"82",
          6129 => x"99",
          6130 => x"da",
          6131 => x"3d",
          6132 => x"d2",
          6133 => x"53",
          6134 => x"84",
          6135 => x"3d",
          6136 => x"3f",
          6137 => x"08",
          6138 => x"ec",
          6139 => x"38",
          6140 => x"3d",
          6141 => x"3d",
          6142 => x"cc",
          6143 => x"8c",
          6144 => x"82",
          6145 => x"82",
          6146 => x"81",
          6147 => x"81",
          6148 => x"86",
          6149 => x"aa",
          6150 => x"a4",
          6151 => x"a8",
          6152 => x"05",
          6153 => x"ea",
          6154 => x"77",
          6155 => x"70",
          6156 => x"b4",
          6157 => x"3d",
          6158 => x"51",
          6159 => x"82",
          6160 => x"55",
          6161 => x"08",
          6162 => x"6f",
          6163 => x"06",
          6164 => x"a2",
          6165 => x"92",
          6166 => x"81",
          6167 => x"8c",
          6168 => x"2e",
          6169 => x"81",
          6170 => x"51",
          6171 => x"82",
          6172 => x"55",
          6173 => x"08",
          6174 => x"68",
          6175 => x"a8",
          6176 => x"05",
          6177 => x"51",
          6178 => x"3f",
          6179 => x"33",
          6180 => x"8b",
          6181 => x"84",
          6182 => x"06",
          6183 => x"73",
          6184 => x"a0",
          6185 => x"8b",
          6186 => x"54",
          6187 => x"15",
          6188 => x"33",
          6189 => x"70",
          6190 => x"55",
          6191 => x"2e",
          6192 => x"6e",
          6193 => x"df",
          6194 => x"78",
          6195 => x"3f",
          6196 => x"08",
          6197 => x"ff",
          6198 => x"82",
          6199 => x"ec",
          6200 => x"80",
          6201 => x"8c",
          6202 => x"78",
          6203 => x"af",
          6204 => x"ec",
          6205 => x"d4",
          6206 => x"55",
          6207 => x"08",
          6208 => x"81",
          6209 => x"73",
          6210 => x"81",
          6211 => x"63",
          6212 => x"76",
          6213 => x"3f",
          6214 => x"0b",
          6215 => x"87",
          6216 => x"ec",
          6217 => x"77",
          6218 => x"3f",
          6219 => x"08",
          6220 => x"ec",
          6221 => x"78",
          6222 => x"aa",
          6223 => x"ec",
          6224 => x"82",
          6225 => x"a8",
          6226 => x"ed",
          6227 => x"80",
          6228 => x"02",
          6229 => x"df",
          6230 => x"57",
          6231 => x"3d",
          6232 => x"96",
          6233 => x"e9",
          6234 => x"ec",
          6235 => x"8c",
          6236 => x"cf",
          6237 => x"65",
          6238 => x"d4",
          6239 => x"b5",
          6240 => x"ec",
          6241 => x"8c",
          6242 => x"38",
          6243 => x"05",
          6244 => x"06",
          6245 => x"73",
          6246 => x"a7",
          6247 => x"09",
          6248 => x"71",
          6249 => x"06",
          6250 => x"55",
          6251 => x"15",
          6252 => x"81",
          6253 => x"34",
          6254 => x"b4",
          6255 => x"8c",
          6256 => x"74",
          6257 => x"0c",
          6258 => x"04",
          6259 => x"64",
          6260 => x"93",
          6261 => x"52",
          6262 => x"d1",
          6263 => x"8c",
          6264 => x"82",
          6265 => x"80",
          6266 => x"58",
          6267 => x"3d",
          6268 => x"c8",
          6269 => x"8c",
          6270 => x"82",
          6271 => x"b4",
          6272 => x"c7",
          6273 => x"a0",
          6274 => x"55",
          6275 => x"84",
          6276 => x"17",
          6277 => x"2b",
          6278 => x"96",
          6279 => x"b0",
          6280 => x"54",
          6281 => x"15",
          6282 => x"ff",
          6283 => x"82",
          6284 => x"55",
          6285 => x"ec",
          6286 => x"0d",
          6287 => x"0d",
          6288 => x"5a",
          6289 => x"3d",
          6290 => x"99",
          6291 => x"81",
          6292 => x"ec",
          6293 => x"ec",
          6294 => x"82",
          6295 => x"07",
          6296 => x"55",
          6297 => x"2e",
          6298 => x"81",
          6299 => x"55",
          6300 => x"2e",
          6301 => x"7b",
          6302 => x"80",
          6303 => x"70",
          6304 => x"be",
          6305 => x"8c",
          6306 => x"82",
          6307 => x"80",
          6308 => x"52",
          6309 => x"dc",
          6310 => x"ec",
          6311 => x"8c",
          6312 => x"38",
          6313 => x"08",
          6314 => x"08",
          6315 => x"56",
          6316 => x"19",
          6317 => x"59",
          6318 => x"74",
          6319 => x"56",
          6320 => x"ec",
          6321 => x"75",
          6322 => x"74",
          6323 => x"2e",
          6324 => x"16",
          6325 => x"33",
          6326 => x"73",
          6327 => x"38",
          6328 => x"84",
          6329 => x"06",
          6330 => x"7a",
          6331 => x"76",
          6332 => x"07",
          6333 => x"54",
          6334 => x"80",
          6335 => x"80",
          6336 => x"7b",
          6337 => x"53",
          6338 => x"93",
          6339 => x"ec",
          6340 => x"8c",
          6341 => x"38",
          6342 => x"55",
          6343 => x"56",
          6344 => x"8b",
          6345 => x"56",
          6346 => x"83",
          6347 => x"75",
          6348 => x"51",
          6349 => x"3f",
          6350 => x"08",
          6351 => x"82",
          6352 => x"98",
          6353 => x"e6",
          6354 => x"53",
          6355 => x"b8",
          6356 => x"3d",
          6357 => x"3f",
          6358 => x"08",
          6359 => x"08",
          6360 => x"8c",
          6361 => x"98",
          6362 => x"a0",
          6363 => x"70",
          6364 => x"ae",
          6365 => x"6d",
          6366 => x"81",
          6367 => x"57",
          6368 => x"74",
          6369 => x"38",
          6370 => x"81",
          6371 => x"81",
          6372 => x"52",
          6373 => x"89",
          6374 => x"ec",
          6375 => x"a5",
          6376 => x"33",
          6377 => x"54",
          6378 => x"3f",
          6379 => x"08",
          6380 => x"38",
          6381 => x"76",
          6382 => x"05",
          6383 => x"39",
          6384 => x"08",
          6385 => x"15",
          6386 => x"ff",
          6387 => x"73",
          6388 => x"38",
          6389 => x"83",
          6390 => x"56",
          6391 => x"75",
          6392 => x"81",
          6393 => x"33",
          6394 => x"2e",
          6395 => x"52",
          6396 => x"51",
          6397 => x"3f",
          6398 => x"08",
          6399 => x"ff",
          6400 => x"38",
          6401 => x"88",
          6402 => x"8a",
          6403 => x"38",
          6404 => x"ec",
          6405 => x"75",
          6406 => x"74",
          6407 => x"73",
          6408 => x"05",
          6409 => x"17",
          6410 => x"70",
          6411 => x"34",
          6412 => x"70",
          6413 => x"ff",
          6414 => x"55",
          6415 => x"26",
          6416 => x"8b",
          6417 => x"86",
          6418 => x"e5",
          6419 => x"38",
          6420 => x"99",
          6421 => x"05",
          6422 => x"70",
          6423 => x"73",
          6424 => x"81",
          6425 => x"ff",
          6426 => x"ed",
          6427 => x"80",
          6428 => x"91",
          6429 => x"55",
          6430 => x"3f",
          6431 => x"08",
          6432 => x"ec",
          6433 => x"38",
          6434 => x"51",
          6435 => x"3f",
          6436 => x"08",
          6437 => x"ec",
          6438 => x"76",
          6439 => x"67",
          6440 => x"34",
          6441 => x"82",
          6442 => x"84",
          6443 => x"06",
          6444 => x"80",
          6445 => x"2e",
          6446 => x"81",
          6447 => x"ff",
          6448 => x"82",
          6449 => x"54",
          6450 => x"08",
          6451 => x"53",
          6452 => x"08",
          6453 => x"ff",
          6454 => x"67",
          6455 => x"8b",
          6456 => x"53",
          6457 => x"51",
          6458 => x"3f",
          6459 => x"0b",
          6460 => x"79",
          6461 => x"ee",
          6462 => x"ec",
          6463 => x"55",
          6464 => x"ec",
          6465 => x"0d",
          6466 => x"0d",
          6467 => x"88",
          6468 => x"05",
          6469 => x"fc",
          6470 => x"54",
          6471 => x"d2",
          6472 => x"8c",
          6473 => x"82",
          6474 => x"82",
          6475 => x"1a",
          6476 => x"82",
          6477 => x"80",
          6478 => x"8c",
          6479 => x"78",
          6480 => x"1a",
          6481 => x"2a",
          6482 => x"51",
          6483 => x"90",
          6484 => x"82",
          6485 => x"58",
          6486 => x"81",
          6487 => x"39",
          6488 => x"22",
          6489 => x"70",
          6490 => x"56",
          6491 => x"ff",
          6492 => x"14",
          6493 => x"30",
          6494 => x"9f",
          6495 => x"ec",
          6496 => x"19",
          6497 => x"5a",
          6498 => x"81",
          6499 => x"38",
          6500 => x"77",
          6501 => x"82",
          6502 => x"56",
          6503 => x"74",
          6504 => x"ff",
          6505 => x"81",
          6506 => x"55",
          6507 => x"75",
          6508 => x"82",
          6509 => x"ec",
          6510 => x"ff",
          6511 => x"8c",
          6512 => x"2e",
          6513 => x"82",
          6514 => x"8e",
          6515 => x"56",
          6516 => x"09",
          6517 => x"38",
          6518 => x"59",
          6519 => x"77",
          6520 => x"06",
          6521 => x"87",
          6522 => x"39",
          6523 => x"ba",
          6524 => x"55",
          6525 => x"2e",
          6526 => x"15",
          6527 => x"2e",
          6528 => x"83",
          6529 => x"75",
          6530 => x"7e",
          6531 => x"a8",
          6532 => x"ec",
          6533 => x"8c",
          6534 => x"ce",
          6535 => x"16",
          6536 => x"56",
          6537 => x"38",
          6538 => x"19",
          6539 => x"8c",
          6540 => x"7d",
          6541 => x"38",
          6542 => x"0c",
          6543 => x"0c",
          6544 => x"80",
          6545 => x"73",
          6546 => x"98",
          6547 => x"05",
          6548 => x"57",
          6549 => x"26",
          6550 => x"7b",
          6551 => x"0c",
          6552 => x"81",
          6553 => x"84",
          6554 => x"54",
          6555 => x"ec",
          6556 => x"0d",
          6557 => x"0d",
          6558 => x"88",
          6559 => x"05",
          6560 => x"54",
          6561 => x"c5",
          6562 => x"56",
          6563 => x"8c",
          6564 => x"8b",
          6565 => x"8c",
          6566 => x"29",
          6567 => x"05",
          6568 => x"55",
          6569 => x"84",
          6570 => x"34",
          6571 => x"08",
          6572 => x"5f",
          6573 => x"51",
          6574 => x"3f",
          6575 => x"08",
          6576 => x"70",
          6577 => x"57",
          6578 => x"8b",
          6579 => x"82",
          6580 => x"06",
          6581 => x"56",
          6582 => x"38",
          6583 => x"05",
          6584 => x"7e",
          6585 => x"f0",
          6586 => x"ec",
          6587 => x"67",
          6588 => x"2e",
          6589 => x"82",
          6590 => x"8b",
          6591 => x"75",
          6592 => x"80",
          6593 => x"81",
          6594 => x"2e",
          6595 => x"80",
          6596 => x"38",
          6597 => x"0a",
          6598 => x"ff",
          6599 => x"55",
          6600 => x"86",
          6601 => x"8a",
          6602 => x"89",
          6603 => x"2a",
          6604 => x"77",
          6605 => x"59",
          6606 => x"81",
          6607 => x"70",
          6608 => x"07",
          6609 => x"56",
          6610 => x"38",
          6611 => x"05",
          6612 => x"7e",
          6613 => x"80",
          6614 => x"82",
          6615 => x"8a",
          6616 => x"83",
          6617 => x"06",
          6618 => x"08",
          6619 => x"74",
          6620 => x"41",
          6621 => x"56",
          6622 => x"8a",
          6623 => x"61",
          6624 => x"55",
          6625 => x"27",
          6626 => x"93",
          6627 => x"80",
          6628 => x"38",
          6629 => x"70",
          6630 => x"43",
          6631 => x"95",
          6632 => x"06",
          6633 => x"2e",
          6634 => x"77",
          6635 => x"74",
          6636 => x"83",
          6637 => x"06",
          6638 => x"82",
          6639 => x"2e",
          6640 => x"78",
          6641 => x"2e",
          6642 => x"80",
          6643 => x"ae",
          6644 => x"2a",
          6645 => x"81",
          6646 => x"56",
          6647 => x"2e",
          6648 => x"77",
          6649 => x"81",
          6650 => x"79",
          6651 => x"70",
          6652 => x"5a",
          6653 => x"86",
          6654 => x"27",
          6655 => x"52",
          6656 => x"fa",
          6657 => x"8c",
          6658 => x"29",
          6659 => x"70",
          6660 => x"55",
          6661 => x"0b",
          6662 => x"08",
          6663 => x"05",
          6664 => x"ff",
          6665 => x"27",
          6666 => x"88",
          6667 => x"ae",
          6668 => x"2a",
          6669 => x"81",
          6670 => x"56",
          6671 => x"2e",
          6672 => x"77",
          6673 => x"81",
          6674 => x"79",
          6675 => x"70",
          6676 => x"5a",
          6677 => x"86",
          6678 => x"27",
          6679 => x"52",
          6680 => x"f9",
          6681 => x"8c",
          6682 => x"84",
          6683 => x"8c",
          6684 => x"f5",
          6685 => x"81",
          6686 => x"ec",
          6687 => x"8c",
          6688 => x"71",
          6689 => x"83",
          6690 => x"5e",
          6691 => x"89",
          6692 => x"5c",
          6693 => x"1c",
          6694 => x"05",
          6695 => x"ff",
          6696 => x"70",
          6697 => x"31",
          6698 => x"57",
          6699 => x"83",
          6700 => x"06",
          6701 => x"1c",
          6702 => x"5c",
          6703 => x"1d",
          6704 => x"29",
          6705 => x"31",
          6706 => x"55",
          6707 => x"87",
          6708 => x"7c",
          6709 => x"7a",
          6710 => x"31",
          6711 => x"f8",
          6712 => x"8c",
          6713 => x"7d",
          6714 => x"81",
          6715 => x"82",
          6716 => x"83",
          6717 => x"80",
          6718 => x"87",
          6719 => x"81",
          6720 => x"fd",
          6721 => x"f8",
          6722 => x"2e",
          6723 => x"80",
          6724 => x"ff",
          6725 => x"8c",
          6726 => x"a0",
          6727 => x"38",
          6728 => x"74",
          6729 => x"86",
          6730 => x"fd",
          6731 => x"81",
          6732 => x"80",
          6733 => x"83",
          6734 => x"39",
          6735 => x"08",
          6736 => x"92",
          6737 => x"b8",
          6738 => x"59",
          6739 => x"27",
          6740 => x"86",
          6741 => x"55",
          6742 => x"09",
          6743 => x"38",
          6744 => x"f5",
          6745 => x"38",
          6746 => x"55",
          6747 => x"86",
          6748 => x"80",
          6749 => x"7a",
          6750 => x"b9",
          6751 => x"81",
          6752 => x"7a",
          6753 => x"8a",
          6754 => x"52",
          6755 => x"ff",
          6756 => x"79",
          6757 => x"7b",
          6758 => x"06",
          6759 => x"51",
          6760 => x"3f",
          6761 => x"1c",
          6762 => x"32",
          6763 => x"96",
          6764 => x"06",
          6765 => x"91",
          6766 => x"a1",
          6767 => x"55",
          6768 => x"ff",
          6769 => x"74",
          6770 => x"06",
          6771 => x"51",
          6772 => x"3f",
          6773 => x"52",
          6774 => x"ff",
          6775 => x"f8",
          6776 => x"34",
          6777 => x"1b",
          6778 => x"d9",
          6779 => x"52",
          6780 => x"ff",
          6781 => x"60",
          6782 => x"51",
          6783 => x"3f",
          6784 => x"09",
          6785 => x"cb",
          6786 => x"b2",
          6787 => x"c3",
          6788 => x"a0",
          6789 => x"52",
          6790 => x"ff",
          6791 => x"82",
          6792 => x"51",
          6793 => x"3f",
          6794 => x"1b",
          6795 => x"95",
          6796 => x"b2",
          6797 => x"a0",
          6798 => x"80",
          6799 => x"1c",
          6800 => x"80",
          6801 => x"93",
          6802 => x"84",
          6803 => x"1b",
          6804 => x"82",
          6805 => x"52",
          6806 => x"ff",
          6807 => x"7c",
          6808 => x"06",
          6809 => x"51",
          6810 => x"3f",
          6811 => x"a4",
          6812 => x"0b",
          6813 => x"93",
          6814 => x"98",
          6815 => x"51",
          6816 => x"3f",
          6817 => x"52",
          6818 => x"70",
          6819 => x"9f",
          6820 => x"54",
          6821 => x"52",
          6822 => x"9b",
          6823 => x"56",
          6824 => x"08",
          6825 => x"7d",
          6826 => x"81",
          6827 => x"38",
          6828 => x"86",
          6829 => x"52",
          6830 => x"9b",
          6831 => x"80",
          6832 => x"7a",
          6833 => x"ed",
          6834 => x"85",
          6835 => x"7a",
          6836 => x"8f",
          6837 => x"85",
          6838 => x"83",
          6839 => x"ff",
          6840 => x"ff",
          6841 => x"e8",
          6842 => x"9e",
          6843 => x"52",
          6844 => x"51",
          6845 => x"3f",
          6846 => x"52",
          6847 => x"9e",
          6848 => x"54",
          6849 => x"53",
          6850 => x"51",
          6851 => x"3f",
          6852 => x"16",
          6853 => x"7e",
          6854 => x"d8",
          6855 => x"80",
          6856 => x"ff",
          6857 => x"7f",
          6858 => x"7d",
          6859 => x"81",
          6860 => x"f8",
          6861 => x"ff",
          6862 => x"ff",
          6863 => x"51",
          6864 => x"3f",
          6865 => x"88",
          6866 => x"39",
          6867 => x"f8",
          6868 => x"2e",
          6869 => x"55",
          6870 => x"51",
          6871 => x"3f",
          6872 => x"57",
          6873 => x"83",
          6874 => x"76",
          6875 => x"7a",
          6876 => x"ff",
          6877 => x"82",
          6878 => x"82",
          6879 => x"80",
          6880 => x"ec",
          6881 => x"51",
          6882 => x"3f",
          6883 => x"78",
          6884 => x"74",
          6885 => x"18",
          6886 => x"2e",
          6887 => x"79",
          6888 => x"2e",
          6889 => x"55",
          6890 => x"62",
          6891 => x"74",
          6892 => x"75",
          6893 => x"7e",
          6894 => x"b8",
          6895 => x"ec",
          6896 => x"38",
          6897 => x"78",
          6898 => x"74",
          6899 => x"56",
          6900 => x"93",
          6901 => x"66",
          6902 => x"26",
          6903 => x"56",
          6904 => x"83",
          6905 => x"64",
          6906 => x"77",
          6907 => x"84",
          6908 => x"52",
          6909 => x"9d",
          6910 => x"d4",
          6911 => x"51",
          6912 => x"3f",
          6913 => x"55",
          6914 => x"81",
          6915 => x"34",
          6916 => x"16",
          6917 => x"16",
          6918 => x"16",
          6919 => x"05",
          6920 => x"c1",
          6921 => x"fe",
          6922 => x"fe",
          6923 => x"34",
          6924 => x"08",
          6925 => x"07",
          6926 => x"16",
          6927 => x"ec",
          6928 => x"34",
          6929 => x"c6",
          6930 => x"9c",
          6931 => x"52",
          6932 => x"51",
          6933 => x"3f",
          6934 => x"53",
          6935 => x"51",
          6936 => x"3f",
          6937 => x"8c",
          6938 => x"38",
          6939 => x"52",
          6940 => x"99",
          6941 => x"56",
          6942 => x"08",
          6943 => x"39",
          6944 => x"39",
          6945 => x"39",
          6946 => x"08",
          6947 => x"8c",
          6948 => x"3d",
          6949 => x"3d",
          6950 => x"5b",
          6951 => x"60",
          6952 => x"57",
          6953 => x"25",
          6954 => x"3d",
          6955 => x"55",
          6956 => x"15",
          6957 => x"c9",
          6958 => x"81",
          6959 => x"06",
          6960 => x"3d",
          6961 => x"8d",
          6962 => x"74",
          6963 => x"05",
          6964 => x"17",
          6965 => x"2e",
          6966 => x"c9",
          6967 => x"34",
          6968 => x"83",
          6969 => x"74",
          6970 => x"0c",
          6971 => x"04",
          6972 => x"78",
          6973 => x"55",
          6974 => x"80",
          6975 => x"38",
          6976 => x"77",
          6977 => x"33",
          6978 => x"39",
          6979 => x"80",
          6980 => x"56",
          6981 => x"83",
          6982 => x"73",
          6983 => x"2a",
          6984 => x"53",
          6985 => x"73",
          6986 => x"81",
          6987 => x"72",
          6988 => x"05",
          6989 => x"56",
          6990 => x"82",
          6991 => x"77",
          6992 => x"08",
          6993 => x"f3",
          6994 => x"8c",
          6995 => x"38",
          6996 => x"53",
          6997 => x"ff",
          6998 => x"16",
          6999 => x"06",
          7000 => x"76",
          7001 => x"ff",
          7002 => x"8c",
          7003 => x"3d",
          7004 => x"3d",
          7005 => x"71",
          7006 => x"8e",
          7007 => x"29",
          7008 => x"05",
          7009 => x"04",
          7010 => x"51",
          7011 => x"81",
          7012 => x"80",
          7013 => x"ff",
          7014 => x"f2",
          7015 => x"bc",
          7016 => x"39",
          7017 => x"51",
          7018 => x"81",
          7019 => x"80",
          7020 => x"ff",
          7021 => x"d6",
          7022 => x"80",
          7023 => x"39",
          7024 => x"51",
          7025 => x"82",
          7026 => x"80",
          7027 => x"80",
          7028 => x"39",
          7029 => x"51",
          7030 => x"80",
          7031 => x"39",
          7032 => x"51",
          7033 => x"81",
          7034 => x"39",
          7035 => x"51",
          7036 => x"81",
          7037 => x"39",
          7038 => x"51",
          7039 => x"82",
          7040 => x"39",
          7041 => x"51",
          7042 => x"82",
          7043 => x"86",
          7044 => x"3d",
          7045 => x"3d",
          7046 => x"56",
          7047 => x"e7",
          7048 => x"74",
          7049 => x"e8",
          7050 => x"39",
          7051 => x"74",
          7052 => x"82",
          7053 => x"ec",
          7054 => x"51",
          7055 => x"3f",
          7056 => x"08",
          7057 => x"75",
          7058 => x"d0",
          7059 => x"c4",
          7060 => x"0d",
          7061 => x"0d",
          7062 => x"05",
          7063 => x"33",
          7064 => x"68",
          7065 => x"7a",
          7066 => x"51",
          7067 => x"78",
          7068 => x"ff",
          7069 => x"81",
          7070 => x"07",
          7071 => x"06",
          7072 => x"56",
          7073 => x"38",
          7074 => x"52",
          7075 => x"52",
          7076 => x"3f",
          7077 => x"08",
          7078 => x"ec",
          7079 => x"82",
          7080 => x"87",
          7081 => x"0c",
          7082 => x"08",
          7083 => x"d4",
          7084 => x"80",
          7085 => x"75",
          7086 => x"3f",
          7087 => x"08",
          7088 => x"ec",
          7089 => x"7a",
          7090 => x"2e",
          7091 => x"19",
          7092 => x"59",
          7093 => x"3d",
          7094 => x"cd",
          7095 => x"30",
          7096 => x"80",
          7097 => x"70",
          7098 => x"06",
          7099 => x"56",
          7100 => x"90",
          7101 => x"f4",
          7102 => x"98",
          7103 => x"78",
          7104 => x"3f",
          7105 => x"82",
          7106 => x"96",
          7107 => x"f9",
          7108 => x"02",
          7109 => x"05",
          7110 => x"ff",
          7111 => x"7a",
          7112 => x"fe",
          7113 => x"8c",
          7114 => x"38",
          7115 => x"88",
          7116 => x"2e",
          7117 => x"39",
          7118 => x"54",
          7119 => x"53",
          7120 => x"51",
          7121 => x"8c",
          7122 => x"83",
          7123 => x"76",
          7124 => x"0c",
          7125 => x"04",
          7126 => x"7f",
          7127 => x"8c",
          7128 => x"05",
          7129 => x"15",
          7130 => x"5c",
          7131 => x"5e",
          7132 => x"82",
          7133 => x"89",
          7134 => x"83",
          7135 => x"83",
          7136 => x"55",
          7137 => x"80",
          7138 => x"90",
          7139 => x"7b",
          7140 => x"38",
          7141 => x"74",
          7142 => x"7a",
          7143 => x"72",
          7144 => x"83",
          7145 => x"88",
          7146 => x"39",
          7147 => x"51",
          7148 => x"3f",
          7149 => x"80",
          7150 => x"18",
          7151 => x"27",
          7152 => x"08",
          7153 => x"fc",
          7154 => x"c8",
          7155 => x"82",
          7156 => x"ff",
          7157 => x"84",
          7158 => x"39",
          7159 => x"72",
          7160 => x"38",
          7161 => x"82",
          7162 => x"ff",
          7163 => x"89",
          7164 => x"a4",
          7165 => x"b8",
          7166 => x"55",
          7167 => x"81",
          7168 => x"80",
          7169 => x"a8",
          7170 => x"a4",
          7171 => x"74",
          7172 => x"38",
          7173 => x"33",
          7174 => x"56",
          7175 => x"83",
          7176 => x"80",
          7177 => x"27",
          7178 => x"53",
          7179 => x"70",
          7180 => x"51",
          7181 => x"2e",
          7182 => x"80",
          7183 => x"38",
          7184 => x"39",
          7185 => x"81",
          7186 => x"15",
          7187 => x"82",
          7188 => x"ff",
          7189 => x"78",
          7190 => x"5c",
          7191 => x"dc",
          7192 => x"ec",
          7193 => x"70",
          7194 => x"57",
          7195 => x"09",
          7196 => x"38",
          7197 => x"3f",
          7198 => x"08",
          7199 => x"98",
          7200 => x"32",
          7201 => x"9b",
          7202 => x"70",
          7203 => x"75",
          7204 => x"58",
          7205 => x"51",
          7206 => x"24",
          7207 => x"9b",
          7208 => x"06",
          7209 => x"53",
          7210 => x"1e",
          7211 => x"26",
          7212 => x"ff",
          7213 => x"8c",
          7214 => x"3d",
          7215 => x"3d",
          7216 => x"05",
          7217 => x"b0",
          7218 => x"b4",
          7219 => x"86",
          7220 => x"89",
          7221 => x"fe",
          7222 => x"82",
          7223 => x"82",
          7224 => x"82",
          7225 => x"52",
          7226 => x"51",
          7227 => x"3f",
          7228 => x"85",
          7229 => x"e8",
          7230 => x"0d",
          7231 => x"0d",
          7232 => x"80",
          7233 => x"ff",
          7234 => x"51",
          7235 => x"3f",
          7236 => x"51",
          7237 => x"3f",
          7238 => x"f1",
          7239 => x"81",
          7240 => x"06",
          7241 => x"80",
          7242 => x"81",
          7243 => x"a0",
          7244 => x"88",
          7245 => x"98",
          7246 => x"fe",
          7247 => x"72",
          7248 => x"81",
          7249 => x"71",
          7250 => x"38",
          7251 => x"f0",
          7252 => x"84",
          7253 => x"f2",
          7254 => x"51",
          7255 => x"3f",
          7256 => x"70",
          7257 => x"52",
          7258 => x"95",
          7259 => x"fe",
          7260 => x"82",
          7261 => x"fe",
          7262 => x"80",
          7263 => x"d0",
          7264 => x"2a",
          7265 => x"51",
          7266 => x"2e",
          7267 => x"51",
          7268 => x"3f",
          7269 => x"51",
          7270 => x"3f",
          7271 => x"f0",
          7272 => x"85",
          7273 => x"06",
          7274 => x"80",
          7275 => x"81",
          7276 => x"9c",
          7277 => x"d4",
          7278 => x"94",
          7279 => x"fe",
          7280 => x"72",
          7281 => x"81",
          7282 => x"71",
          7283 => x"38",
          7284 => x"ef",
          7285 => x"84",
          7286 => x"f1",
          7287 => x"51",
          7288 => x"3f",
          7289 => x"70",
          7290 => x"52",
          7291 => x"95",
          7292 => x"fe",
          7293 => x"82",
          7294 => x"fe",
          7295 => x"80",
          7296 => x"cc",
          7297 => x"2a",
          7298 => x"51",
          7299 => x"2e",
          7300 => x"51",
          7301 => x"3f",
          7302 => x"51",
          7303 => x"3f",
          7304 => x"ef",
          7305 => x"fd",
          7306 => x"3d",
          7307 => x"3d",
          7308 => x"70",
          7309 => x"80",
          7310 => x"fe",
          7311 => x"82",
          7312 => x"54",
          7313 => x"81",
          7314 => x"d0",
          7315 => x"f0",
          7316 => x"dc",
          7317 => x"ec",
          7318 => x"82",
          7319 => x"07",
          7320 => x"71",
          7321 => x"54",
          7322 => x"f8",
          7323 => x"f8",
          7324 => x"81",
          7325 => x"06",
          7326 => x"a3",
          7327 => x"52",
          7328 => x"92",
          7329 => x"ec",
          7330 => x"8c",
          7331 => x"ec",
          7332 => x"fd",
          7333 => x"39",
          7334 => x"51",
          7335 => x"82",
          7336 => x"f8",
          7337 => x"f8",
          7338 => x"82",
          7339 => x"06",
          7340 => x"52",
          7341 => x"83",
          7342 => x"0b",
          7343 => x"0c",
          7344 => x"04",
          7345 => x"80",
          7346 => x"a3",
          7347 => x"5d",
          7348 => x"51",
          7349 => x"3f",
          7350 => x"08",
          7351 => x"59",
          7352 => x"09",
          7353 => x"38",
          7354 => x"52",
          7355 => x"52",
          7356 => x"b6",
          7357 => x"78",
          7358 => x"9c",
          7359 => x"cf",
          7360 => x"ec",
          7361 => x"88",
          7362 => x"e4",
          7363 => x"39",
          7364 => x"5d",
          7365 => x"51",
          7366 => x"3f",
          7367 => x"46",
          7368 => x"52",
          7369 => x"86",
          7370 => x"ff",
          7371 => x"f3",
          7372 => x"8c",
          7373 => x"2b",
          7374 => x"51",
          7375 => x"c2",
          7376 => x"38",
          7377 => x"24",
          7378 => x"bd",
          7379 => x"38",
          7380 => x"90",
          7381 => x"2e",
          7382 => x"78",
          7383 => x"da",
          7384 => x"39",
          7385 => x"2e",
          7386 => x"78",
          7387 => x"85",
          7388 => x"bf",
          7389 => x"38",
          7390 => x"78",
          7391 => x"89",
          7392 => x"80",
          7393 => x"38",
          7394 => x"2e",
          7395 => x"78",
          7396 => x"89",
          7397 => x"b4",
          7398 => x"83",
          7399 => x"38",
          7400 => x"24",
          7401 => x"81",
          7402 => x"fd",
          7403 => x"39",
          7404 => x"2e",
          7405 => x"8a",
          7406 => x"3d",
          7407 => x"53",
          7408 => x"51",
          7409 => x"3f",
          7410 => x"08",
          7411 => x"c4",
          7412 => x"fe",
          7413 => x"ff",
          7414 => x"ff",
          7415 => x"82",
          7416 => x"80",
          7417 => x"38",
          7418 => x"f8",
          7419 => x"84",
          7420 => x"82",
          7421 => x"8c",
          7422 => x"38",
          7423 => x"08",
          7424 => x"a0",
          7425 => x"a8",
          7426 => x"5c",
          7427 => x"27",
          7428 => x"61",
          7429 => x"70",
          7430 => x"0c",
          7431 => x"f5",
          7432 => x"39",
          7433 => x"80",
          7434 => x"84",
          7435 => x"81",
          7436 => x"8c",
          7437 => x"2e",
          7438 => x"b4",
          7439 => x"11",
          7440 => x"05",
          7441 => x"c1",
          7442 => x"ec",
          7443 => x"fd",
          7444 => x"3d",
          7445 => x"53",
          7446 => x"51",
          7447 => x"3f",
          7448 => x"08",
          7449 => x"ac",
          7450 => x"b0",
          7451 => x"c0",
          7452 => x"79",
          7453 => x"8c",
          7454 => x"79",
          7455 => x"5b",
          7456 => x"61",
          7457 => x"eb",
          7458 => x"ff",
          7459 => x"ff",
          7460 => x"ff",
          7461 => x"82",
          7462 => x"80",
          7463 => x"38",
          7464 => x"fc",
          7465 => x"84",
          7466 => x"80",
          7467 => x"8c",
          7468 => x"2e",
          7469 => x"b4",
          7470 => x"11",
          7471 => x"05",
          7472 => x"c5",
          7473 => x"ec",
          7474 => x"fc",
          7475 => x"86",
          7476 => x"f8",
          7477 => x"5a",
          7478 => x"a8",
          7479 => x"33",
          7480 => x"5a",
          7481 => x"2e",
          7482 => x"55",
          7483 => x"33",
          7484 => x"82",
          7485 => x"fe",
          7486 => x"81",
          7487 => x"05",
          7488 => x"39",
          7489 => x"51",
          7490 => x"b4",
          7491 => x"11",
          7492 => x"05",
          7493 => x"f1",
          7494 => x"ec",
          7495 => x"38",
          7496 => x"33",
          7497 => x"2e",
          7498 => x"89",
          7499 => x"80",
          7500 => x"89",
          7501 => x"78",
          7502 => x"38",
          7503 => x"08",
          7504 => x"82",
          7505 => x"59",
          7506 => x"88",
          7507 => x"a8",
          7508 => x"39",
          7509 => x"33",
          7510 => x"2e",
          7511 => x"89",
          7512 => x"9a",
          7513 => x"de",
          7514 => x"80",
          7515 => x"82",
          7516 => x"44",
          7517 => x"89",
          7518 => x"80",
          7519 => x"3d",
          7520 => x"53",
          7521 => x"51",
          7522 => x"3f",
          7523 => x"08",
          7524 => x"82",
          7525 => x"59",
          7526 => x"89",
          7527 => x"9c",
          7528 => x"cc",
          7529 => x"e1",
          7530 => x"80",
          7531 => x"82",
          7532 => x"43",
          7533 => x"89",
          7534 => x"78",
          7535 => x"38",
          7536 => x"08",
          7537 => x"82",
          7538 => x"59",
          7539 => x"88",
          7540 => x"b4",
          7541 => x"39",
          7542 => x"33",
          7543 => x"2e",
          7544 => x"89",
          7545 => x"88",
          7546 => x"c8",
          7547 => x"43",
          7548 => x"f8",
          7549 => x"84",
          7550 => x"fe",
          7551 => x"8c",
          7552 => x"2e",
          7553 => x"62",
          7554 => x"88",
          7555 => x"81",
          7556 => x"32",
          7557 => x"72",
          7558 => x"70",
          7559 => x"51",
          7560 => x"80",
          7561 => x"7a",
          7562 => x"38",
          7563 => x"86",
          7564 => x"f5",
          7565 => x"55",
          7566 => x"53",
          7567 => x"51",
          7568 => x"82",
          7569 => x"fe",
          7570 => x"f9",
          7571 => x"3d",
          7572 => x"53",
          7573 => x"51",
          7574 => x"3f",
          7575 => x"08",
          7576 => x"b0",
          7577 => x"fe",
          7578 => x"ff",
          7579 => x"fe",
          7580 => x"82",
          7581 => x"80",
          7582 => x"63",
          7583 => x"cb",
          7584 => x"34",
          7585 => x"44",
          7586 => x"fc",
          7587 => x"84",
          7588 => x"fc",
          7589 => x"8c",
          7590 => x"38",
          7591 => x"63",
          7592 => x"52",
          7593 => x"51",
          7594 => x"3f",
          7595 => x"79",
          7596 => x"ba",
          7597 => x"79",
          7598 => x"ae",
          7599 => x"38",
          7600 => x"a0",
          7601 => x"fe",
          7602 => x"ff",
          7603 => x"fe",
          7604 => x"82",
          7605 => x"80",
          7606 => x"63",
          7607 => x"cb",
          7608 => x"34",
          7609 => x"44",
          7610 => x"82",
          7611 => x"fe",
          7612 => x"ff",
          7613 => x"3d",
          7614 => x"53",
          7615 => x"51",
          7616 => x"3f",
          7617 => x"08",
          7618 => x"88",
          7619 => x"fe",
          7620 => x"ff",
          7621 => x"fe",
          7622 => x"82",
          7623 => x"80",
          7624 => x"60",
          7625 => x"05",
          7626 => x"82",
          7627 => x"78",
          7628 => x"fe",
          7629 => x"ff",
          7630 => x"fe",
          7631 => x"82",
          7632 => x"df",
          7633 => x"39",
          7634 => x"54",
          7635 => x"98",
          7636 => x"c0",
          7637 => x"52",
          7638 => x"fa",
          7639 => x"45",
          7640 => x"78",
          7641 => x"ac",
          7642 => x"26",
          7643 => x"82",
          7644 => x"39",
          7645 => x"f0",
          7646 => x"84",
          7647 => x"fc",
          7648 => x"8c",
          7649 => x"2e",
          7650 => x"59",
          7651 => x"22",
          7652 => x"05",
          7653 => x"41",
          7654 => x"82",
          7655 => x"fe",
          7656 => x"ff",
          7657 => x"3d",
          7658 => x"53",
          7659 => x"51",
          7660 => x"3f",
          7661 => x"08",
          7662 => x"d8",
          7663 => x"fe",
          7664 => x"ff",
          7665 => x"fe",
          7666 => x"82",
          7667 => x"80",
          7668 => x"60",
          7669 => x"59",
          7670 => x"41",
          7671 => x"f0",
          7672 => x"84",
          7673 => x"fc",
          7674 => x"8c",
          7675 => x"38",
          7676 => x"60",
          7677 => x"52",
          7678 => x"51",
          7679 => x"3f",
          7680 => x"79",
          7681 => x"e6",
          7682 => x"79",
          7683 => x"ae",
          7684 => x"38",
          7685 => x"9c",
          7686 => x"fe",
          7687 => x"ff",
          7688 => x"fe",
          7689 => x"82",
          7690 => x"80",
          7691 => x"60",
          7692 => x"59",
          7693 => x"41",
          7694 => x"82",
          7695 => x"fe",
          7696 => x"ff",
          7697 => x"3d",
          7698 => x"53",
          7699 => x"51",
          7700 => x"3f",
          7701 => x"08",
          7702 => x"b8",
          7703 => x"82",
          7704 => x"fe",
          7705 => x"63",
          7706 => x"b4",
          7707 => x"11",
          7708 => x"05",
          7709 => x"91",
          7710 => x"ec",
          7711 => x"f5",
          7712 => x"52",
          7713 => x"51",
          7714 => x"3f",
          7715 => x"2d",
          7716 => x"08",
          7717 => x"fc",
          7718 => x"ec",
          7719 => x"87",
          7720 => x"f6",
          7721 => x"ec",
          7722 => x"84",
          7723 => x"80",
          7724 => x"e1",
          7725 => x"39",
          7726 => x"51",
          7727 => x"3f",
          7728 => x"a5",
          7729 => x"98",
          7730 => x"39",
          7731 => x"51",
          7732 => x"2e",
          7733 => x"7d",
          7734 => x"78",
          7735 => x"d8",
          7736 => x"ff",
          7737 => x"fe",
          7738 => x"82",
          7739 => x"5c",
          7740 => x"82",
          7741 => x"7a",
          7742 => x"38",
          7743 => x"8c",
          7744 => x"39",
          7745 => x"b0",
          7746 => x"39",
          7747 => x"56",
          7748 => x"88",
          7749 => x"53",
          7750 => x"52",
          7751 => x"b0",
          7752 => x"f6",
          7753 => x"39",
          7754 => x"52",
          7755 => x"b0",
          7756 => x"f5",
          7757 => x"39",
          7758 => x"88",
          7759 => x"53",
          7760 => x"52",
          7761 => x"b0",
          7762 => x"f5",
          7763 => x"39",
          7764 => x"53",
          7765 => x"52",
          7766 => x"b0",
          7767 => x"f5",
          7768 => x"89",
          7769 => x"8d",
          7770 => x"56",
          7771 => x"46",
          7772 => x"80",
          7773 => x"80",
          7774 => x"80",
          7775 => x"ff",
          7776 => x"eb",
          7777 => x"8c",
          7778 => x"8c",
          7779 => x"70",
          7780 => x"07",
          7781 => x"5b",
          7782 => x"5a",
          7783 => x"83",
          7784 => x"78",
          7785 => x"78",
          7786 => x"38",
          7787 => x"81",
          7788 => x"59",
          7789 => x"38",
          7790 => x"7d",
          7791 => x"59",
          7792 => x"7e",
          7793 => x"81",
          7794 => x"38",
          7795 => x"51",
          7796 => x"3f",
          7797 => x"fc",
          7798 => x"0b",
          7799 => x"34",
          7800 => x"8c",
          7801 => x"55",
          7802 => x"52",
          7803 => x"d6",
          7804 => x"8c",
          7805 => x"2b",
          7806 => x"53",
          7807 => x"52",
          7808 => x"d6",
          7809 => x"82",
          7810 => x"07",
          7811 => x"c0",
          7812 => x"08",
          7813 => x"84",
          7814 => x"51",
          7815 => x"3f",
          7816 => x"08",
          7817 => x"08",
          7818 => x"84",
          7819 => x"51",
          7820 => x"3f",
          7821 => x"ec",
          7822 => x"0c",
          7823 => x"0b",
          7824 => x"84",
          7825 => x"83",
          7826 => x"94",
          7827 => x"d3",
          7828 => x"8c",
          7829 => x"d6",
          7830 => x"8d",
          7831 => x"e3",
          7832 => x"ec",
          7833 => x"88",
          7834 => x"ed",
          7835 => x"88",
          7836 => x"ed",
          7837 => x"e1",
          7838 => x"ec",
          7839 => x"51",
          7840 => x"f0",
          7841 => x"04",
          7842 => x"93",
          7843 => x"99",
          7844 => x"9f",
          7845 => x"a5",
          7846 => x"ab",
          7847 => x"04",
          7848 => x"88",
          7849 => x"8f",
          7850 => x"96",
          7851 => x"9d",
          7852 => x"a4",
          7853 => x"ab",
          7854 => x"b2",
          7855 => x"b9",
          7856 => x"c0",
          7857 => x"c7",
          7858 => x"ce",
          7859 => x"d4",
          7860 => x"da",
          7861 => x"e0",
          7862 => x"e6",
          7863 => x"ec",
          7864 => x"f2",
          7865 => x"f8",
          7866 => x"fe",
          7867 => x"25",
          7868 => x"64",
          7869 => x"3a",
          7870 => x"25",
          7871 => x"64",
          7872 => x"00",
          7873 => x"20",
          7874 => x"66",
          7875 => x"72",
          7876 => x"6f",
          7877 => x"00",
          7878 => x"72",
          7879 => x"53",
          7880 => x"63",
          7881 => x"69",
          7882 => x"00",
          7883 => x"65",
          7884 => x"65",
          7885 => x"6d",
          7886 => x"6d",
          7887 => x"65",
          7888 => x"00",
          7889 => x"20",
          7890 => x"53",
          7891 => x"4d",
          7892 => x"25",
          7893 => x"3a",
          7894 => x"58",
          7895 => x"00",
          7896 => x"20",
          7897 => x"41",
          7898 => x"20",
          7899 => x"25",
          7900 => x"3a",
          7901 => x"58",
          7902 => x"00",
          7903 => x"20",
          7904 => x"4e",
          7905 => x"41",
          7906 => x"25",
          7907 => x"3a",
          7908 => x"58",
          7909 => x"00",
          7910 => x"20",
          7911 => x"4d",
          7912 => x"20",
          7913 => x"25",
          7914 => x"3a",
          7915 => x"58",
          7916 => x"00",
          7917 => x"20",
          7918 => x"20",
          7919 => x"20",
          7920 => x"25",
          7921 => x"3a",
          7922 => x"58",
          7923 => x"00",
          7924 => x"20",
          7925 => x"43",
          7926 => x"20",
          7927 => x"44",
          7928 => x"63",
          7929 => x"3d",
          7930 => x"64",
          7931 => x"00",
          7932 => x"20",
          7933 => x"45",
          7934 => x"20",
          7935 => x"54",
          7936 => x"72",
          7937 => x"3d",
          7938 => x"64",
          7939 => x"00",
          7940 => x"20",
          7941 => x"52",
          7942 => x"52",
          7943 => x"43",
          7944 => x"6e",
          7945 => x"3d",
          7946 => x"64",
          7947 => x"00",
          7948 => x"20",
          7949 => x"48",
          7950 => x"45",
          7951 => x"53",
          7952 => x"00",
          7953 => x"20",
          7954 => x"49",
          7955 => x"00",
          7956 => x"20",
          7957 => x"54",
          7958 => x"00",
          7959 => x"20",
          7960 => x"0a",
          7961 => x"00",
          7962 => x"20",
          7963 => x"0a",
          7964 => x"00",
          7965 => x"72",
          7966 => x"65",
          7967 => x"00",
          7968 => x"20",
          7969 => x"20",
          7970 => x"65",
          7971 => x"65",
          7972 => x"72",
          7973 => x"64",
          7974 => x"73",
          7975 => x"25",
          7976 => x"0a",
          7977 => x"00",
          7978 => x"20",
          7979 => x"20",
          7980 => x"6f",
          7981 => x"53",
          7982 => x"74",
          7983 => x"64",
          7984 => x"73",
          7985 => x"25",
          7986 => x"0a",
          7987 => x"00",
          7988 => x"20",
          7989 => x"63",
          7990 => x"74",
          7991 => x"20",
          7992 => x"72",
          7993 => x"20",
          7994 => x"20",
          7995 => x"25",
          7996 => x"0a",
          7997 => x"00",
          7998 => x"63",
          7999 => x"00",
          8000 => x"20",
          8001 => x"20",
          8002 => x"20",
          8003 => x"20",
          8004 => x"20",
          8005 => x"20",
          8006 => x"20",
          8007 => x"25",
          8008 => x"0a",
          8009 => x"00",
          8010 => x"20",
          8011 => x"74",
          8012 => x"43",
          8013 => x"6b",
          8014 => x"65",
          8015 => x"20",
          8016 => x"20",
          8017 => x"25",
          8018 => x"30",
          8019 => x"48",
          8020 => x"00",
          8021 => x"20",
          8022 => x"41",
          8023 => x"6c",
          8024 => x"20",
          8025 => x"71",
          8026 => x"20",
          8027 => x"20",
          8028 => x"25",
          8029 => x"30",
          8030 => x"48",
          8031 => x"00",
          8032 => x"20",
          8033 => x"68",
          8034 => x"65",
          8035 => x"52",
          8036 => x"43",
          8037 => x"6b",
          8038 => x"65",
          8039 => x"25",
          8040 => x"30",
          8041 => x"48",
          8042 => x"00",
          8043 => x"6c",
          8044 => x"00",
          8045 => x"69",
          8046 => x"00",
          8047 => x"78",
          8048 => x"00",
          8049 => x"00",
          8050 => x"6d",
          8051 => x"00",
          8052 => x"6e",
          8053 => x"00",
          8054 => x"00",
          8055 => x"2c",
          8056 => x"3d",
          8057 => x"5d",
          8058 => x"00",
          8059 => x"00",
          8060 => x"33",
          8061 => x"00",
          8062 => x"4d",
          8063 => x"53",
          8064 => x"00",
          8065 => x"4e",
          8066 => x"20",
          8067 => x"46",
          8068 => x"32",
          8069 => x"00",
          8070 => x"4e",
          8071 => x"20",
          8072 => x"46",
          8073 => x"20",
          8074 => x"00",
          8075 => x"d8",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"41",
          8080 => x"80",
          8081 => x"49",
          8082 => x"8f",
          8083 => x"4f",
          8084 => x"55",
          8085 => x"9b",
          8086 => x"9f",
          8087 => x"55",
          8088 => x"a7",
          8089 => x"ab",
          8090 => x"af",
          8091 => x"b3",
          8092 => x"b7",
          8093 => x"bb",
          8094 => x"bf",
          8095 => x"c3",
          8096 => x"c7",
          8097 => x"cb",
          8098 => x"cf",
          8099 => x"d3",
          8100 => x"d7",
          8101 => x"db",
          8102 => x"df",
          8103 => x"e3",
          8104 => x"e7",
          8105 => x"eb",
          8106 => x"ef",
          8107 => x"f3",
          8108 => x"f7",
          8109 => x"fb",
          8110 => x"ff",
          8111 => x"3b",
          8112 => x"2f",
          8113 => x"3a",
          8114 => x"7c",
          8115 => x"00",
          8116 => x"04",
          8117 => x"40",
          8118 => x"00",
          8119 => x"00",
          8120 => x"02",
          8121 => x"08",
          8122 => x"20",
          8123 => x"00",
          8124 => x"69",
          8125 => x"00",
          8126 => x"63",
          8127 => x"00",
          8128 => x"69",
          8129 => x"00",
          8130 => x"61",
          8131 => x"00",
          8132 => x"65",
          8133 => x"00",
          8134 => x"65",
          8135 => x"00",
          8136 => x"70",
          8137 => x"00",
          8138 => x"66",
          8139 => x"00",
          8140 => x"6d",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"6c",
          8150 => x"00",
          8151 => x"00",
          8152 => x"74",
          8153 => x"00",
          8154 => x"65",
          8155 => x"00",
          8156 => x"6f",
          8157 => x"00",
          8158 => x"74",
          8159 => x"00",
          8160 => x"73",
          8161 => x"00",
          8162 => x"6b",
          8163 => x"72",
          8164 => x"00",
          8165 => x"65",
          8166 => x"6c",
          8167 => x"72",
          8168 => x"0a",
          8169 => x"00",
          8170 => x"6b",
          8171 => x"74",
          8172 => x"61",
          8173 => x"0a",
          8174 => x"00",
          8175 => x"66",
          8176 => x"20",
          8177 => x"6e",
          8178 => x"00",
          8179 => x"70",
          8180 => x"20",
          8181 => x"6e",
          8182 => x"00",
          8183 => x"61",
          8184 => x"20",
          8185 => x"65",
          8186 => x"65",
          8187 => x"00",
          8188 => x"65",
          8189 => x"64",
          8190 => x"65",
          8191 => x"00",
          8192 => x"65",
          8193 => x"72",
          8194 => x"79",
          8195 => x"69",
          8196 => x"2e",
          8197 => x"00",
          8198 => x"65",
          8199 => x"6e",
          8200 => x"20",
          8201 => x"61",
          8202 => x"2e",
          8203 => x"00",
          8204 => x"69",
          8205 => x"72",
          8206 => x"20",
          8207 => x"74",
          8208 => x"65",
          8209 => x"00",
          8210 => x"76",
          8211 => x"75",
          8212 => x"72",
          8213 => x"20",
          8214 => x"61",
          8215 => x"2e",
          8216 => x"00",
          8217 => x"6b",
          8218 => x"74",
          8219 => x"61",
          8220 => x"64",
          8221 => x"00",
          8222 => x"63",
          8223 => x"61",
          8224 => x"6c",
          8225 => x"69",
          8226 => x"79",
          8227 => x"6d",
          8228 => x"75",
          8229 => x"6f",
          8230 => x"69",
          8231 => x"0a",
          8232 => x"00",
          8233 => x"6d",
          8234 => x"61",
          8235 => x"74",
          8236 => x"0a",
          8237 => x"00",
          8238 => x"65",
          8239 => x"2c",
          8240 => x"65",
          8241 => x"69",
          8242 => x"63",
          8243 => x"65",
          8244 => x"64",
          8245 => x"00",
          8246 => x"65",
          8247 => x"20",
          8248 => x"6b",
          8249 => x"0a",
          8250 => x"00",
          8251 => x"75",
          8252 => x"63",
          8253 => x"74",
          8254 => x"6d",
          8255 => x"2e",
          8256 => x"00",
          8257 => x"20",
          8258 => x"79",
          8259 => x"65",
          8260 => x"69",
          8261 => x"2e",
          8262 => x"00",
          8263 => x"61",
          8264 => x"65",
          8265 => x"69",
          8266 => x"72",
          8267 => x"74",
          8268 => x"00",
          8269 => x"63",
          8270 => x"2e",
          8271 => x"00",
          8272 => x"6e",
          8273 => x"20",
          8274 => x"6f",
          8275 => x"00",
          8276 => x"75",
          8277 => x"74",
          8278 => x"25",
          8279 => x"74",
          8280 => x"75",
          8281 => x"74",
          8282 => x"73",
          8283 => x"0a",
          8284 => x"00",
          8285 => x"64",
          8286 => x"00",
          8287 => x"58",
          8288 => x"00",
          8289 => x"00",
          8290 => x"58",
          8291 => x"00",
          8292 => x"20",
          8293 => x"20",
          8294 => x"00",
          8295 => x"58",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"20",
          8302 => x"28",
          8303 => x"00",
          8304 => x"30",
          8305 => x"30",
          8306 => x"00",
          8307 => x"30",
          8308 => x"00",
          8309 => x"55",
          8310 => x"65",
          8311 => x"30",
          8312 => x"20",
          8313 => x"25",
          8314 => x"2a",
          8315 => x"00",
          8316 => x"20",
          8317 => x"65",
          8318 => x"70",
          8319 => x"61",
          8320 => x"65",
          8321 => x"00",
          8322 => x"65",
          8323 => x"6e",
          8324 => x"72",
          8325 => x"0a",
          8326 => x"00",
          8327 => x"20",
          8328 => x"65",
          8329 => x"70",
          8330 => x"00",
          8331 => x"54",
          8332 => x"44",
          8333 => x"74",
          8334 => x"75",
          8335 => x"00",
          8336 => x"54",
          8337 => x"52",
          8338 => x"74",
          8339 => x"75",
          8340 => x"00",
          8341 => x"54",
          8342 => x"58",
          8343 => x"74",
          8344 => x"75",
          8345 => x"00",
          8346 => x"54",
          8347 => x"58",
          8348 => x"74",
          8349 => x"75",
          8350 => x"00",
          8351 => x"54",
          8352 => x"58",
          8353 => x"74",
          8354 => x"75",
          8355 => x"00",
          8356 => x"54",
          8357 => x"58",
          8358 => x"74",
          8359 => x"75",
          8360 => x"00",
          8361 => x"74",
          8362 => x"20",
          8363 => x"74",
          8364 => x"72",
          8365 => x"0a",
          8366 => x"00",
          8367 => x"62",
          8368 => x"67",
          8369 => x"6d",
          8370 => x"2e",
          8371 => x"00",
          8372 => x"6f",
          8373 => x"63",
          8374 => x"74",
          8375 => x"00",
          8376 => x"00",
          8377 => x"6c",
          8378 => x"74",
          8379 => x"6e",
          8380 => x"61",
          8381 => x"65",
          8382 => x"20",
          8383 => x"64",
          8384 => x"20",
          8385 => x"61",
          8386 => x"69",
          8387 => x"20",
          8388 => x"75",
          8389 => x"79",
          8390 => x"00",
          8391 => x"00",
          8392 => x"61",
          8393 => x"67",
          8394 => x"2e",
          8395 => x"00",
          8396 => x"79",
          8397 => x"2e",
          8398 => x"00",
          8399 => x"70",
          8400 => x"6e",
          8401 => x"2e",
          8402 => x"00",
          8403 => x"6c",
          8404 => x"30",
          8405 => x"2d",
          8406 => x"38",
          8407 => x"25",
          8408 => x"29",
          8409 => x"00",
          8410 => x"70",
          8411 => x"6d",
          8412 => x"0a",
          8413 => x"00",
          8414 => x"6d",
          8415 => x"74",
          8416 => x"00",
          8417 => x"58",
          8418 => x"32",
          8419 => x"00",
          8420 => x"0a",
          8421 => x"00",
          8422 => x"58",
          8423 => x"34",
          8424 => x"00",
          8425 => x"58",
          8426 => x"38",
          8427 => x"00",
          8428 => x"63",
          8429 => x"6e",
          8430 => x"6f",
          8431 => x"40",
          8432 => x"38",
          8433 => x"2e",
          8434 => x"00",
          8435 => x"6c",
          8436 => x"20",
          8437 => x"65",
          8438 => x"25",
          8439 => x"20",
          8440 => x"0a",
          8441 => x"00",
          8442 => x"6c",
          8443 => x"74",
          8444 => x"65",
          8445 => x"6f",
          8446 => x"28",
          8447 => x"2e",
          8448 => x"00",
          8449 => x"74",
          8450 => x"69",
          8451 => x"61",
          8452 => x"69",
          8453 => x"69",
          8454 => x"2e",
          8455 => x"00",
          8456 => x"64",
          8457 => x"62",
          8458 => x"69",
          8459 => x"2e",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"5c",
          8464 => x"25",
          8465 => x"73",
          8466 => x"00",
          8467 => x"5c",
          8468 => x"25",
          8469 => x"00",
          8470 => x"5c",
          8471 => x"00",
          8472 => x"20",
          8473 => x"6d",
          8474 => x"2e",
          8475 => x"00",
          8476 => x"6e",
          8477 => x"2e",
          8478 => x"00",
          8479 => x"62",
          8480 => x"67",
          8481 => x"74",
          8482 => x"75",
          8483 => x"2e",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"ff",
          8488 => x"00",
          8489 => x"ff",
          8490 => x"00",
          8491 => x"ff",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"ff",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"01",
          8505 => x"01",
          8506 => x"01",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"f0",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"f8",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"08",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"10",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"18",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"20",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"28",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"30",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"38",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"3c",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"40",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"44",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"48",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"4c",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"50",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"54",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"5c",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"60",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"68",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"70",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"78",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"80",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"0b",
            10 => x"80",
            11 => x"0c",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"88",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"0b",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"00",
           267 => x"ff",
           268 => x"06",
           269 => x"83",
           270 => x"10",
           271 => x"fc",
           272 => x"51",
           273 => x"80",
           274 => x"ff",
           275 => x"06",
           276 => x"52",
           277 => x"0a",
           278 => x"38",
           279 => x"51",
           280 => x"70",
           281 => x"8e",
           282 => x"70",
           283 => x"0c",
           284 => x"88",
           285 => x"fe",
           286 => x"04",
           287 => x"00",
           288 => x"00",
           289 => x"08",
           290 => x"fd",
           291 => x"53",
           292 => x"05",
           293 => x"08",
           294 => x"51",
           295 => x"88",
           296 => x"0c",
           297 => x"0d",
           298 => x"94",
           299 => x"0c",
           300 => x"81",
           301 => x"8c",
           302 => x"94",
           303 => x"08",
           304 => x"3f",
           305 => x"88",
           306 => x"3d",
           307 => x"04",
           308 => x"94",
           309 => x"0d",
           310 => x"08",
           311 => x"94",
           312 => x"08",
           313 => x"38",
           314 => x"05",
           315 => x"08",
           316 => x"80",
           317 => x"f4",
           318 => x"08",
           319 => x"88",
           320 => x"94",
           321 => x"0c",
           322 => x"05",
           323 => x"fc",
           324 => x"08",
           325 => x"80",
           326 => x"94",
           327 => x"08",
           328 => x"8c",
           329 => x"0b",
           330 => x"05",
           331 => x"fc",
           332 => x"38",
           333 => x"08",
           334 => x"94",
           335 => x"08",
           336 => x"05",
           337 => x"94",
           338 => x"08",
           339 => x"88",
           340 => x"81",
           341 => x"08",
           342 => x"f8",
           343 => x"94",
           344 => x"08",
           345 => x"38",
           346 => x"05",
           347 => x"08",
           348 => x"94",
           349 => x"08",
           350 => x"54",
           351 => x"94",
           352 => x"08",
           353 => x"fb",
           354 => x"0b",
           355 => x"05",
           356 => x"88",
           357 => x"25",
           358 => x"08",
           359 => x"30",
           360 => x"05",
           361 => x"94",
           362 => x"0c",
           363 => x"05",
           364 => x"8c",
           365 => x"8c",
           366 => x"94",
           367 => x"0c",
           368 => x"08",
           369 => x"52",
           370 => x"05",
           371 => x"3f",
           372 => x"94",
           373 => x"0c",
           374 => x"fc",
           375 => x"2e",
           376 => x"08",
           377 => x"30",
           378 => x"05",
           379 => x"f8",
           380 => x"88",
           381 => x"3d",
           382 => x"04",
           383 => x"94",
           384 => x"0d",
           385 => x"08",
           386 => x"80",
           387 => x"f8",
           388 => x"08",
           389 => x"94",
           390 => x"08",
           391 => x"94",
           392 => x"08",
           393 => x"38",
           394 => x"08",
           395 => x"24",
           396 => x"08",
           397 => x"10",
           398 => x"05",
           399 => x"fc",
           400 => x"94",
           401 => x"0c",
           402 => x"08",
           403 => x"80",
           404 => x"38",
           405 => x"05",
           406 => x"88",
           407 => x"a1",
           408 => x"88",
           409 => x"08",
           410 => x"31",
           411 => x"05",
           412 => x"f8",
           413 => x"08",
           414 => x"07",
           415 => x"05",
           416 => x"fc",
           417 => x"2a",
           418 => x"05",
           419 => x"8c",
           420 => x"2a",
           421 => x"05",
           422 => x"39",
           423 => x"05",
           424 => x"8f",
           425 => x"88",
           426 => x"94",
           427 => x"0c",
           428 => x"94",
           429 => x"08",
           430 => x"f4",
           431 => x"94",
           432 => x"08",
           433 => x"3d",
           434 => x"04",
           435 => x"81",
           436 => x"c0",
           437 => x"81",
           438 => x"92",
           439 => x"0b",
           440 => x"8c",
           441 => x"92",
           442 => x"82",
           443 => x"70",
           444 => x"38",
           445 => x"8c",
           446 => x"e9",
           447 => x"92",
           448 => x"80",
           449 => x"71",
           450 => x"c0",
           451 => x"51",
           452 => x"88",
           453 => x"0b",
           454 => x"34",
           455 => x"9f",
           456 => x"0c",
           457 => x"04",
           458 => x"78",
           459 => x"58",
           460 => x"0b",
           461 => x"f0",
           462 => x"52",
           463 => x"70",
           464 => x"81",
           465 => x"38",
           466 => x"c0",
           467 => x"79",
           468 => x"80",
           469 => x"87",
           470 => x"0c",
           471 => x"8c",
           472 => x"2a",
           473 => x"51",
           474 => x"80",
           475 => x"87",
           476 => x"08",
           477 => x"06",
           478 => x"52",
           479 => x"80",
           480 => x"70",
           481 => x"38",
           482 => x"81",
           483 => x"ff",
           484 => x"15",
           485 => x"06",
           486 => x"2e",
           487 => x"c0",
           488 => x"51",
           489 => x"38",
           490 => x"8c",
           491 => x"95",
           492 => x"87",
           493 => x"0c",
           494 => x"8c",
           495 => x"06",
           496 => x"f4",
           497 => x"fc",
           498 => x"52",
           499 => x"2e",
           500 => x"8f",
           501 => x"98",
           502 => x"70",
           503 => x"81",
           504 => x"81",
           505 => x"0c",
           506 => x"04",
           507 => x"74",
           508 => x"71",
           509 => x"2b",
           510 => x"53",
           511 => x"0d",
           512 => x"0d",
           513 => x"33",
           514 => x"71",
           515 => x"88",
           516 => x"14",
           517 => x"07",
           518 => x"33",
           519 => x"0c",
           520 => x"56",
           521 => x"3d",
           522 => x"3d",
           523 => x"0b",
           524 => x"08",
           525 => x"77",
           526 => x"38",
           527 => x"08",
           528 => x"38",
           529 => x"74",
           530 => x"38",
           531 => x"ae",
           532 => x"39",
           533 => x"10",
           534 => x"53",
           535 => x"8c",
           536 => x"52",
           537 => x"52",
           538 => x"3f",
           539 => x"38",
           540 => x"f8",
           541 => x"83",
           542 => x"55",
           543 => x"54",
           544 => x"83",
           545 => x"76",
           546 => x"17",
           547 => x"88",
           548 => x"55",
           549 => x"88",
           550 => x"74",
           551 => x"3f",
           552 => x"0a",
           553 => x"39",
           554 => x"88",
           555 => x"0d",
           556 => x"0d",
           557 => x"9f",
           558 => x"19",
           559 => x"fe",
           560 => x"54",
           561 => x"73",
           562 => x"82",
           563 => x"71",
           564 => x"08",
           565 => x"75",
           566 => x"3d",
           567 => x"3d",
           568 => x"80",
           569 => x"0b",
           570 => x"70",
           571 => x"53",
           572 => x"09",
           573 => x"38",
           574 => x"fd",
           575 => x"08",
           576 => x"9a",
           577 => x"e4",
           578 => x"83",
           579 => x"73",
           580 => x"85",
           581 => x"fc",
           582 => x"0b",
           583 => x"f4",
           584 => x"80",
           585 => x"15",
           586 => x"81",
           587 => x"88",
           588 => x"26",
           589 => x"52",
           590 => x"90",
           591 => x"52",
           592 => x"09",
           593 => x"38",
           594 => x"53",
           595 => x"0c",
           596 => x"8b",
           597 => x"fe",
           598 => x"08",
           599 => x"90",
           600 => x"71",
           601 => x"80",
           602 => x"0c",
           603 => x"04",
           604 => x"78",
           605 => x"9f",
           606 => x"22",
           607 => x"83",
           608 => x"57",
           609 => x"73",
           610 => x"38",
           611 => x"53",
           612 => x"83",
           613 => x"39",
           614 => x"52",
           615 => x"38",
           616 => x"16",
           617 => x"08",
           618 => x"38",
           619 => x"17",
           620 => x"73",
           621 => x"38",
           622 => x"16",
           623 => x"74",
           624 => x"52",
           625 => x"72",
           626 => x"3f",
           627 => x"88",
           628 => x"38",
           629 => x"08",
           630 => x"27",
           631 => x"08",
           632 => x"88",
           633 => x"c9",
           634 => x"90",
           635 => x"75",
           636 => x"71",
           637 => x"3d",
           638 => x"3d",
           639 => x"64",
           640 => x"75",
           641 => x"a0",
           642 => x"06",
           643 => x"16",
           644 => x"ef",
           645 => x"33",
           646 => x"af",
           647 => x"06",
           648 => x"16",
           649 => x"88",
           650 => x"70",
           651 => x"74",
           652 => x"38",
           653 => x"df",
           654 => x"56",
           655 => x"82",
           656 => x"3d",
           657 => x"70",
           658 => x"8a",
           659 => x"70",
           660 => x"34",
           661 => x"74",
           662 => x"81",
           663 => x"80",
           664 => x"88",
           665 => x"5a",
           666 => x"70",
           667 => x"60",
           668 => x"70",
           669 => x"30",
           670 => x"71",
           671 => x"51",
           672 => x"53",
           673 => x"74",
           674 => x"76",
           675 => x"81",
           676 => x"81",
           677 => x"27",
           678 => x"74",
           679 => x"38",
           680 => x"70",
           681 => x"32",
           682 => x"73",
           683 => x"53",
           684 => x"56",
           685 => x"88",
           686 => x"ff",
           687 => x"81",
           688 => x"ff",
           689 => x"53",
           690 => x"76",
           691 => x"98",
           692 => x"7f",
           693 => x"76",
           694 => x"38",
           695 => x"8b",
           696 => x"51",
           697 => x"88",
           698 => x"38",
           699 => x"22",
           700 => x"83",
           701 => x"55",
           702 => x"52",
           703 => x"a8",
           704 => x"57",
           705 => x"fb",
           706 => x"55",
           707 => x"80",
           708 => x"1d",
           709 => x"2a",
           710 => x"51",
           711 => x"b2",
           712 => x"84",
           713 => x"08",
           714 => x"58",
           715 => x"77",
           716 => x"38",
           717 => x"05",
           718 => x"70",
           719 => x"33",
           720 => x"52",
           721 => x"80",
           722 => x"86",
           723 => x"2e",
           724 => x"51",
           725 => x"ff",
           726 => x"08",
           727 => x"b4",
           728 => x"76",
           729 => x"08",
           730 => x"51",
           731 => x"38",
           732 => x"70",
           733 => x"81",
           734 => x"56",
           735 => x"83",
           736 => x"81",
           737 => x"7c",
           738 => x"3f",
           739 => x"1d",
           740 => x"39",
           741 => x"90",
           742 => x"f9",
           743 => x"7b",
           744 => x"54",
           745 => x"77",
           746 => x"f6",
           747 => x"56",
           748 => x"e7",
           749 => x"f8",
           750 => x"08",
           751 => x"06",
           752 => x"74",
           753 => x"2e",
           754 => x"80",
           755 => x"54",
           756 => x"52",
           757 => x"d0",
           758 => x"56",
           759 => x"38",
           760 => x"88",
           761 => x"83",
           762 => x"55",
           763 => x"c6",
           764 => x"82",
           765 => x"53",
           766 => x"51",
           767 => x"88",
           768 => x"08",
           769 => x"51",
           770 => x"88",
           771 => x"ff",
           772 => x"81",
           773 => x"83",
           774 => x"75",
           775 => x"3d",
           776 => x"3d",
           777 => x"80",
           778 => x"0b",
           779 => x"f5",
           780 => x"08",
           781 => x"82",
           782 => x"f2",
           783 => x"53",
           784 => x"53",
           785 => x"d3",
           786 => x"81",
           787 => x"76",
           788 => x"81",
           789 => x"90",
           790 => x"53",
           791 => x"51",
           792 => x"88",
           793 => x"8d",
           794 => x"74",
           795 => x"38",
           796 => x"05",
           797 => x"3f",
           798 => x"08",
           799 => x"5a",
           800 => x"88",
           801 => x"06",
           802 => x"2e",
           803 => x"86",
           804 => x"82",
           805 => x"80",
           806 => x"86",
           807 => x"39",
           808 => x"53",
           809 => x"51",
           810 => x"81",
           811 => x"81",
           812 => x"3d",
           813 => x"f6",
           814 => x"08",
           815 => x"06",
           816 => x"38",
           817 => x"05",
           818 => x"3f",
           819 => x"02",
           820 => x"78",
           821 => x"88",
           822 => x"70",
           823 => x"5b",
           824 => x"88",
           825 => x"ff",
           826 => x"8c",
           827 => x"3d",
           828 => x"34",
           829 => x"05",
           830 => x"3f",
           831 => x"1a",
           832 => x"e2",
           833 => x"e4",
           834 => x"83",
           835 => x"56",
           836 => x"95",
           837 => x"51",
           838 => x"88",
           839 => x"51",
           840 => x"88",
           841 => x"ff",
           842 => x"31",
           843 => x"1b",
           844 => x"2a",
           845 => x"56",
           846 => x"55",
           847 => x"55",
           848 => x"88",
           849 => x"70",
           850 => x"88",
           851 => x"05",
           852 => x"83",
           853 => x"83",
           854 => x"83",
           855 => x"27",
           856 => x"57",
           857 => x"56",
           858 => x"80",
           859 => x"79",
           860 => x"2e",
           861 => x"90",
           862 => x"fb",
           863 => x"81",
           864 => x"90",
           865 => x"39",
           866 => x"18",
           867 => x"79",
           868 => x"06",
           869 => x"19",
           870 => x"05",
           871 => x"55",
           872 => x"1a",
           873 => x"0b",
           874 => x"0c",
           875 => x"88",
           876 => x"0d",
           877 => x"0d",
           878 => x"9f",
           879 => x"85",
           880 => x"2e",
           881 => x"80",
           882 => x"34",
           883 => x"11",
           884 => x"89",
           885 => x"57",
           886 => x"f8",
           887 => x"08",
           888 => x"80",
           889 => x"3d",
           890 => x"80",
           891 => x"02",
           892 => x"70",
           893 => x"81",
           894 => x"57",
           895 => x"85",
           896 => x"a1",
           897 => x"f5",
           898 => x"08",
           899 => x"98",
           900 => x"51",
           901 => x"88",
           902 => x"0c",
           903 => x"0c",
           904 => x"16",
           905 => x"0c",
           906 => x"04",
           907 => x"7d",
           908 => x"0b",
           909 => x"08",
           910 => x"58",
           911 => x"85",
           912 => x"2e",
           913 => x"81",
           914 => x"06",
           915 => x"74",
           916 => x"c3",
           917 => x"74",
           918 => x"86",
           919 => x"81",
           920 => x"57",
           921 => x"9c",
           922 => x"17",
           923 => x"74",
           924 => x"38",
           925 => x"80",
           926 => x"38",
           927 => x"70",
           928 => x"56",
           929 => x"c7",
           930 => x"33",
           931 => x"89",
           932 => x"81",
           933 => x"55",
           934 => x"76",
           935 => x"16",
           936 => x"39",
           937 => x"51",
           938 => x"88",
           939 => x"75",
           940 => x"38",
           941 => x"0c",
           942 => x"51",
           943 => x"88",
           944 => x"08",
           945 => x"8f",
           946 => x"1a",
           947 => x"98",
           948 => x"ff",
           949 => x"71",
           950 => x"77",
           951 => x"38",
           952 => x"54",
           953 => x"83",
           954 => x"a8",
           955 => x"78",
           956 => x"3f",
           957 => x"e5",
           958 => x"08",
           959 => x"0c",
           960 => x"7b",
           961 => x"0c",
           962 => x"2e",
           963 => x"74",
           964 => x"e2",
           965 => x"76",
           966 => x"3d",
           967 => x"3d",
           968 => x"94",
           969 => x"87",
           970 => x"73",
           971 => x"3f",
           972 => x"2b",
           973 => x"8c",
           974 => x"87",
           975 => x"74",
           976 => x"3f",
           977 => x"07",
           978 => x"8c",
           979 => x"94",
           980 => x"87",
           981 => x"73",
           982 => x"3f",
           983 => x"2b",
           984 => x"9c",
           985 => x"87",
           986 => x"74",
           987 => x"3f",
           988 => x"07",
           989 => x"9c",
           990 => x"83",
           991 => x"94",
           992 => x"80",
           993 => x"c0",
           994 => x"9f",
           995 => x"92",
           996 => x"b8",
           997 => x"51",
           998 => x"88",
           999 => x"a0",
          1000 => x"08",
          1001 => x"88",
          1002 => x"3d",
          1003 => x"84",
          1004 => x"51",
          1005 => x"88",
          1006 => x"75",
          1007 => x"2e",
          1008 => x"15",
          1009 => x"a0",
          1010 => x"04",
          1011 => x"39",
          1012 => x"ff",
          1013 => x"ff",
          1014 => x"00",
          1015 => x"ff",
          1016 => x"4f",
          1017 => x"4e",
          1018 => x"4f",
          1019 => x"00",
          1020 => x"00",
          2048 => x"80",
          2049 => x"0b",
          2050 => x"95",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"80",
          2057 => x"0b",
          2058 => x"85",
          2059 => x"80",
          2060 => x"0b",
          2061 => x"a5",
          2062 => x"80",
          2063 => x"0b",
          2064 => x"c5",
          2065 => x"80",
          2066 => x"0b",
          2067 => x"e5",
          2068 => x"80",
          2069 => x"0b",
          2070 => x"85",
          2071 => x"80",
          2072 => x"0b",
          2073 => x"a5",
          2074 => x"80",
          2075 => x"0b",
          2076 => x"c5",
          2077 => x"80",
          2078 => x"0b",
          2079 => x"e5",
          2080 => x"80",
          2081 => x"0b",
          2082 => x"85",
          2083 => x"80",
          2084 => x"0b",
          2085 => x"a5",
          2086 => x"80",
          2087 => x"0b",
          2088 => x"c5",
          2089 => x"80",
          2090 => x"0b",
          2091 => x"e5",
          2092 => x"80",
          2093 => x"0b",
          2094 => x"85",
          2095 => x"80",
          2096 => x"0b",
          2097 => x"a5",
          2098 => x"80",
          2099 => x"0b",
          2100 => x"c5",
          2101 => x"80",
          2102 => x"0b",
          2103 => x"e5",
          2104 => x"80",
          2105 => x"0b",
          2106 => x"85",
          2107 => x"80",
          2108 => x"0b",
          2109 => x"a5",
          2110 => x"80",
          2111 => x"0b",
          2112 => x"c5",
          2113 => x"80",
          2114 => x"0b",
          2115 => x"e5",
          2116 => x"80",
          2117 => x"0b",
          2118 => x"85",
          2119 => x"80",
          2120 => x"0b",
          2121 => x"a5",
          2122 => x"80",
          2123 => x"0b",
          2124 => x"c5",
          2125 => x"80",
          2126 => x"0b",
          2127 => x"e5",
          2128 => x"80",
          2129 => x"0b",
          2130 => x"85",
          2131 => x"00",
          2132 => x"00",
          2133 => x"00",
          2134 => x"00",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"c4",
          2177 => x"8c",
          2178 => x"d4",
          2179 => x"8c",
          2180 => x"80",
          2181 => x"8c",
          2182 => x"e1",
          2183 => x"8c",
          2184 => x"80",
          2185 => x"8c",
          2186 => x"e2",
          2187 => x"8c",
          2188 => x"80",
          2189 => x"8c",
          2190 => x"e2",
          2191 => x"8c",
          2192 => x"80",
          2193 => x"8c",
          2194 => x"e8",
          2195 => x"8c",
          2196 => x"80",
          2197 => x"8c",
          2198 => x"e9",
          2199 => x"8c",
          2200 => x"80",
          2201 => x"8c",
          2202 => x"e2",
          2203 => x"8c",
          2204 => x"80",
          2205 => x"8c",
          2206 => x"ea",
          2207 => x"8c",
          2208 => x"80",
          2209 => x"8c",
          2210 => x"eb",
          2211 => x"8c",
          2212 => x"80",
          2213 => x"8c",
          2214 => x"e8",
          2215 => x"8c",
          2216 => x"80",
          2217 => x"8c",
          2218 => x"e8",
          2219 => x"8c",
          2220 => x"80",
          2221 => x"8c",
          2222 => x"e8",
          2223 => x"8c",
          2224 => x"80",
          2225 => x"8c",
          2226 => x"d6",
          2227 => x"8c",
          2228 => x"80",
          2229 => x"8c",
          2230 => x"d7",
          2231 => x"8c",
          2232 => x"80",
          2233 => x"8c",
          2234 => x"cf",
          2235 => x"8c",
          2236 => x"80",
          2237 => x"8c",
          2238 => x"d1",
          2239 => x"8c",
          2240 => x"80",
          2241 => x"8c",
          2242 => x"d2",
          2243 => x"8c",
          2244 => x"80",
          2245 => x"8c",
          2246 => x"9e",
          2247 => x"8c",
          2248 => x"80",
          2249 => x"8c",
          2250 => x"ab",
          2251 => x"8c",
          2252 => x"80",
          2253 => x"8c",
          2254 => x"a3",
          2255 => x"8c",
          2256 => x"80",
          2257 => x"8c",
          2258 => x"a6",
          2259 => x"8c",
          2260 => x"80",
          2261 => x"8c",
          2262 => x"b0",
          2263 => x"8c",
          2264 => x"80",
          2265 => x"8c",
          2266 => x"b9",
          2267 => x"8c",
          2268 => x"80",
          2269 => x"8c",
          2270 => x"aa",
          2271 => x"8c",
          2272 => x"80",
          2273 => x"8c",
          2274 => x"b3",
          2275 => x"8c",
          2276 => x"80",
          2277 => x"8c",
          2278 => x"b4",
          2279 => x"8c",
          2280 => x"80",
          2281 => x"8c",
          2282 => x"b5",
          2283 => x"8c",
          2284 => x"80",
          2285 => x"8c",
          2286 => x"bc",
          2287 => x"8c",
          2288 => x"80",
          2289 => x"8c",
          2290 => x"ba",
          2291 => x"8c",
          2292 => x"80",
          2293 => x"8c",
          2294 => x"bf",
          2295 => x"8c",
          2296 => x"80",
          2297 => x"8c",
          2298 => x"b6",
          2299 => x"8c",
          2300 => x"80",
          2301 => x"8c",
          2302 => x"c2",
          2303 => x"8c",
          2304 => x"80",
          2305 => x"8c",
          2306 => x"c3",
          2307 => x"8c",
          2308 => x"80",
          2309 => x"8c",
          2310 => x"ac",
          2311 => x"8c",
          2312 => x"80",
          2313 => x"8c",
          2314 => x"ab",
          2315 => x"8c",
          2316 => x"80",
          2317 => x"8c",
          2318 => x"ad",
          2319 => x"8c",
          2320 => x"80",
          2321 => x"8c",
          2322 => x"b6",
          2323 => x"8c",
          2324 => x"80",
          2325 => x"8c",
          2326 => x"c4",
          2327 => x"8c",
          2328 => x"80",
          2329 => x"8c",
          2330 => x"c6",
          2331 => x"8c",
          2332 => x"80",
          2333 => x"8c",
          2334 => x"ca",
          2335 => x"8c",
          2336 => x"80",
          2337 => x"8c",
          2338 => x"9d",
          2339 => x"8c",
          2340 => x"80",
          2341 => x"8c",
          2342 => x"cc",
          2343 => x"8c",
          2344 => x"80",
          2345 => x"8c",
          2346 => x"ef",
          2347 => x"8c",
          2348 => x"80",
          2349 => x"8c",
          2350 => x"f0",
          2351 => x"8c",
          2352 => x"80",
          2353 => x"8c",
          2354 => x"f2",
          2355 => x"8c",
          2356 => x"80",
          2357 => x"8c",
          2358 => x"d0",
          2359 => x"8c",
          2360 => x"80",
          2361 => x"8c",
          2362 => x"d0",
          2363 => x"8c",
          2364 => x"80",
          2365 => x"8c",
          2366 => x"d3",
          2367 => x"8c",
          2368 => x"80",
          2369 => x"8c",
          2370 => x"da",
          2371 => x"8c",
          2372 => x"80",
          2373 => x"8c",
          2374 => x"a4",
          2375 => x"38",
          2376 => x"84",
          2377 => x"0b",
          2378 => x"98",
          2379 => x"80",
          2380 => x"d7",
          2381 => x"82",
          2382 => x"02",
          2383 => x"0c",
          2384 => x"80",
          2385 => x"f8",
          2386 => x"08",
          2387 => x"f8",
          2388 => x"08",
          2389 => x"3f",
          2390 => x"08",
          2391 => x"ec",
          2392 => x"3d",
          2393 => x"f8",
          2394 => x"8c",
          2395 => x"82",
          2396 => x"fd",
          2397 => x"53",
          2398 => x"08",
          2399 => x"52",
          2400 => x"08",
          2401 => x"51",
          2402 => x"8c",
          2403 => x"82",
          2404 => x"54",
          2405 => x"82",
          2406 => x"04",
          2407 => x"08",
          2408 => x"f8",
          2409 => x"0d",
          2410 => x"8c",
          2411 => x"05",
          2412 => x"82",
          2413 => x"f8",
          2414 => x"8c",
          2415 => x"05",
          2416 => x"f8",
          2417 => x"08",
          2418 => x"82",
          2419 => x"fc",
          2420 => x"2e",
          2421 => x"0b",
          2422 => x"08",
          2423 => x"24",
          2424 => x"8c",
          2425 => x"05",
          2426 => x"8c",
          2427 => x"05",
          2428 => x"f8",
          2429 => x"08",
          2430 => x"f8",
          2431 => x"0c",
          2432 => x"82",
          2433 => x"fc",
          2434 => x"2e",
          2435 => x"82",
          2436 => x"8c",
          2437 => x"8c",
          2438 => x"05",
          2439 => x"38",
          2440 => x"08",
          2441 => x"82",
          2442 => x"8c",
          2443 => x"82",
          2444 => x"88",
          2445 => x"8c",
          2446 => x"05",
          2447 => x"f8",
          2448 => x"08",
          2449 => x"f8",
          2450 => x"0c",
          2451 => x"08",
          2452 => x"81",
          2453 => x"f8",
          2454 => x"0c",
          2455 => x"08",
          2456 => x"81",
          2457 => x"f8",
          2458 => x"0c",
          2459 => x"82",
          2460 => x"90",
          2461 => x"2e",
          2462 => x"8c",
          2463 => x"05",
          2464 => x"8c",
          2465 => x"05",
          2466 => x"39",
          2467 => x"08",
          2468 => x"70",
          2469 => x"08",
          2470 => x"51",
          2471 => x"08",
          2472 => x"82",
          2473 => x"85",
          2474 => x"8c",
          2475 => x"fc",
          2476 => x"79",
          2477 => x"05",
          2478 => x"57",
          2479 => x"83",
          2480 => x"38",
          2481 => x"51",
          2482 => x"a4",
          2483 => x"52",
          2484 => x"93",
          2485 => x"70",
          2486 => x"34",
          2487 => x"71",
          2488 => x"81",
          2489 => x"74",
          2490 => x"0c",
          2491 => x"04",
          2492 => x"2b",
          2493 => x"71",
          2494 => x"51",
          2495 => x"72",
          2496 => x"72",
          2497 => x"05",
          2498 => x"71",
          2499 => x"53",
          2500 => x"70",
          2501 => x"0c",
          2502 => x"84",
          2503 => x"f0",
          2504 => x"8f",
          2505 => x"83",
          2506 => x"38",
          2507 => x"84",
          2508 => x"fc",
          2509 => x"83",
          2510 => x"70",
          2511 => x"39",
          2512 => x"77",
          2513 => x"07",
          2514 => x"54",
          2515 => x"38",
          2516 => x"08",
          2517 => x"71",
          2518 => x"80",
          2519 => x"75",
          2520 => x"33",
          2521 => x"06",
          2522 => x"80",
          2523 => x"72",
          2524 => x"75",
          2525 => x"06",
          2526 => x"12",
          2527 => x"33",
          2528 => x"06",
          2529 => x"52",
          2530 => x"72",
          2531 => x"81",
          2532 => x"81",
          2533 => x"71",
          2534 => x"ec",
          2535 => x"87",
          2536 => x"71",
          2537 => x"fb",
          2538 => x"06",
          2539 => x"82",
          2540 => x"51",
          2541 => x"97",
          2542 => x"84",
          2543 => x"54",
          2544 => x"75",
          2545 => x"38",
          2546 => x"52",
          2547 => x"80",
          2548 => x"ec",
          2549 => x"0d",
          2550 => x"0d",
          2551 => x"53",
          2552 => x"52",
          2553 => x"82",
          2554 => x"81",
          2555 => x"07",
          2556 => x"52",
          2557 => x"e8",
          2558 => x"8c",
          2559 => x"3d",
          2560 => x"3d",
          2561 => x"08",
          2562 => x"56",
          2563 => x"80",
          2564 => x"33",
          2565 => x"2e",
          2566 => x"86",
          2567 => x"52",
          2568 => x"53",
          2569 => x"13",
          2570 => x"33",
          2571 => x"06",
          2572 => x"70",
          2573 => x"38",
          2574 => x"80",
          2575 => x"74",
          2576 => x"81",
          2577 => x"70",
          2578 => x"81",
          2579 => x"80",
          2580 => x"05",
          2581 => x"76",
          2582 => x"70",
          2583 => x"0c",
          2584 => x"04",
          2585 => x"76",
          2586 => x"80",
          2587 => x"86",
          2588 => x"52",
          2589 => x"84",
          2590 => x"ec",
          2591 => x"80",
          2592 => x"74",
          2593 => x"8c",
          2594 => x"3d",
          2595 => x"3d",
          2596 => x"11",
          2597 => x"52",
          2598 => x"70",
          2599 => x"98",
          2600 => x"33",
          2601 => x"82",
          2602 => x"26",
          2603 => x"84",
          2604 => x"83",
          2605 => x"26",
          2606 => x"85",
          2607 => x"84",
          2608 => x"26",
          2609 => x"86",
          2610 => x"85",
          2611 => x"26",
          2612 => x"88",
          2613 => x"86",
          2614 => x"e7",
          2615 => x"38",
          2616 => x"54",
          2617 => x"87",
          2618 => x"cc",
          2619 => x"87",
          2620 => x"0c",
          2621 => x"c0",
          2622 => x"82",
          2623 => x"c0",
          2624 => x"83",
          2625 => x"c0",
          2626 => x"84",
          2627 => x"c0",
          2628 => x"85",
          2629 => x"c0",
          2630 => x"86",
          2631 => x"c0",
          2632 => x"74",
          2633 => x"a4",
          2634 => x"c0",
          2635 => x"80",
          2636 => x"98",
          2637 => x"52",
          2638 => x"ec",
          2639 => x"0d",
          2640 => x"0d",
          2641 => x"c0",
          2642 => x"81",
          2643 => x"c0",
          2644 => x"5e",
          2645 => x"87",
          2646 => x"08",
          2647 => x"1c",
          2648 => x"98",
          2649 => x"79",
          2650 => x"87",
          2651 => x"08",
          2652 => x"1c",
          2653 => x"98",
          2654 => x"79",
          2655 => x"87",
          2656 => x"08",
          2657 => x"1c",
          2658 => x"98",
          2659 => x"7b",
          2660 => x"87",
          2661 => x"08",
          2662 => x"1c",
          2663 => x"0c",
          2664 => x"ff",
          2665 => x"83",
          2666 => x"58",
          2667 => x"57",
          2668 => x"56",
          2669 => x"55",
          2670 => x"54",
          2671 => x"53",
          2672 => x"ff",
          2673 => x"f5",
          2674 => x"c9",
          2675 => x"0d",
          2676 => x"0d",
          2677 => x"33",
          2678 => x"9f",
          2679 => x"52",
          2680 => x"82",
          2681 => x"83",
          2682 => x"fb",
          2683 => x"0b",
          2684 => x"94",
          2685 => x"ff",
          2686 => x"56",
          2687 => x"84",
          2688 => x"2e",
          2689 => x"c0",
          2690 => x"70",
          2691 => x"2a",
          2692 => x"53",
          2693 => x"80",
          2694 => x"71",
          2695 => x"81",
          2696 => x"70",
          2697 => x"81",
          2698 => x"06",
          2699 => x"80",
          2700 => x"71",
          2701 => x"81",
          2702 => x"70",
          2703 => x"73",
          2704 => x"51",
          2705 => x"80",
          2706 => x"2e",
          2707 => x"c0",
          2708 => x"75",
          2709 => x"82",
          2710 => x"87",
          2711 => x"fb",
          2712 => x"9f",
          2713 => x"0b",
          2714 => x"33",
          2715 => x"06",
          2716 => x"87",
          2717 => x"51",
          2718 => x"86",
          2719 => x"94",
          2720 => x"08",
          2721 => x"70",
          2722 => x"54",
          2723 => x"2e",
          2724 => x"91",
          2725 => x"06",
          2726 => x"d7",
          2727 => x"32",
          2728 => x"51",
          2729 => x"2e",
          2730 => x"93",
          2731 => x"06",
          2732 => x"ff",
          2733 => x"81",
          2734 => x"87",
          2735 => x"52",
          2736 => x"86",
          2737 => x"94",
          2738 => x"72",
          2739 => x"0d",
          2740 => x"0d",
          2741 => x"74",
          2742 => x"ff",
          2743 => x"57",
          2744 => x"80",
          2745 => x"81",
          2746 => x"15",
          2747 => x"89",
          2748 => x"81",
          2749 => x"57",
          2750 => x"c0",
          2751 => x"75",
          2752 => x"38",
          2753 => x"94",
          2754 => x"70",
          2755 => x"81",
          2756 => x"52",
          2757 => x"8c",
          2758 => x"2a",
          2759 => x"51",
          2760 => x"38",
          2761 => x"70",
          2762 => x"51",
          2763 => x"8d",
          2764 => x"2a",
          2765 => x"51",
          2766 => x"be",
          2767 => x"ff",
          2768 => x"c0",
          2769 => x"70",
          2770 => x"38",
          2771 => x"90",
          2772 => x"0c",
          2773 => x"33",
          2774 => x"06",
          2775 => x"70",
          2776 => x"76",
          2777 => x"0c",
          2778 => x"04",
          2779 => x"0b",
          2780 => x"94",
          2781 => x"ff",
          2782 => x"87",
          2783 => x"51",
          2784 => x"86",
          2785 => x"94",
          2786 => x"08",
          2787 => x"70",
          2788 => x"51",
          2789 => x"2e",
          2790 => x"81",
          2791 => x"87",
          2792 => x"52",
          2793 => x"86",
          2794 => x"94",
          2795 => x"08",
          2796 => x"06",
          2797 => x"0c",
          2798 => x"0d",
          2799 => x"0d",
          2800 => x"89",
          2801 => x"81",
          2802 => x"53",
          2803 => x"84",
          2804 => x"2e",
          2805 => x"c0",
          2806 => x"71",
          2807 => x"2a",
          2808 => x"51",
          2809 => x"52",
          2810 => x"a0",
          2811 => x"ff",
          2812 => x"c0",
          2813 => x"70",
          2814 => x"38",
          2815 => x"90",
          2816 => x"70",
          2817 => x"98",
          2818 => x"51",
          2819 => x"ec",
          2820 => x"0d",
          2821 => x"0d",
          2822 => x"80",
          2823 => x"2a",
          2824 => x"51",
          2825 => x"84",
          2826 => x"c0",
          2827 => x"82",
          2828 => x"87",
          2829 => x"08",
          2830 => x"0c",
          2831 => x"94",
          2832 => x"a0",
          2833 => x"9e",
          2834 => x"89",
          2835 => x"c0",
          2836 => x"82",
          2837 => x"87",
          2838 => x"08",
          2839 => x"0c",
          2840 => x"ac",
          2841 => x"b0",
          2842 => x"9e",
          2843 => x"89",
          2844 => x"c0",
          2845 => x"82",
          2846 => x"87",
          2847 => x"08",
          2848 => x"0c",
          2849 => x"bc",
          2850 => x"c0",
          2851 => x"9e",
          2852 => x"89",
          2853 => x"c0",
          2854 => x"82",
          2855 => x"87",
          2856 => x"08",
          2857 => x"89",
          2858 => x"c0",
          2859 => x"82",
          2860 => x"87",
          2861 => x"08",
          2862 => x"0c",
          2863 => x"8c",
          2864 => x"d8",
          2865 => x"82",
          2866 => x"80",
          2867 => x"9e",
          2868 => x"84",
          2869 => x"51",
          2870 => x"80",
          2871 => x"81",
          2872 => x"89",
          2873 => x"0b",
          2874 => x"90",
          2875 => x"80",
          2876 => x"52",
          2877 => x"2e",
          2878 => x"52",
          2879 => x"de",
          2880 => x"87",
          2881 => x"08",
          2882 => x"0a",
          2883 => x"52",
          2884 => x"83",
          2885 => x"71",
          2886 => x"34",
          2887 => x"c0",
          2888 => x"70",
          2889 => x"06",
          2890 => x"70",
          2891 => x"38",
          2892 => x"82",
          2893 => x"80",
          2894 => x"9e",
          2895 => x"a0",
          2896 => x"51",
          2897 => x"80",
          2898 => x"81",
          2899 => x"89",
          2900 => x"0b",
          2901 => x"90",
          2902 => x"80",
          2903 => x"52",
          2904 => x"2e",
          2905 => x"52",
          2906 => x"e2",
          2907 => x"87",
          2908 => x"08",
          2909 => x"80",
          2910 => x"52",
          2911 => x"83",
          2912 => x"71",
          2913 => x"34",
          2914 => x"c0",
          2915 => x"70",
          2916 => x"06",
          2917 => x"70",
          2918 => x"38",
          2919 => x"82",
          2920 => x"80",
          2921 => x"9e",
          2922 => x"81",
          2923 => x"51",
          2924 => x"80",
          2925 => x"81",
          2926 => x"89",
          2927 => x"0b",
          2928 => x"90",
          2929 => x"c0",
          2930 => x"52",
          2931 => x"2e",
          2932 => x"52",
          2933 => x"e6",
          2934 => x"87",
          2935 => x"08",
          2936 => x"06",
          2937 => x"70",
          2938 => x"38",
          2939 => x"82",
          2940 => x"87",
          2941 => x"08",
          2942 => x"06",
          2943 => x"51",
          2944 => x"82",
          2945 => x"80",
          2946 => x"9e",
          2947 => x"84",
          2948 => x"52",
          2949 => x"2e",
          2950 => x"52",
          2951 => x"e9",
          2952 => x"9e",
          2953 => x"83",
          2954 => x"84",
          2955 => x"51",
          2956 => x"ea",
          2957 => x"87",
          2958 => x"08",
          2959 => x"51",
          2960 => x"80",
          2961 => x"81",
          2962 => x"89",
          2963 => x"c0",
          2964 => x"70",
          2965 => x"51",
          2966 => x"ec",
          2967 => x"0d",
          2968 => x"0d",
          2969 => x"51",
          2970 => x"82",
          2971 => x"54",
          2972 => x"88",
          2973 => x"98",
          2974 => x"3f",
          2975 => x"51",
          2976 => x"82",
          2977 => x"54",
          2978 => x"93",
          2979 => x"b8",
          2980 => x"bc",
          2981 => x"52",
          2982 => x"51",
          2983 => x"82",
          2984 => x"54",
          2985 => x"93",
          2986 => x"b0",
          2987 => x"b4",
          2988 => x"52",
          2989 => x"51",
          2990 => x"82",
          2991 => x"54",
          2992 => x"93",
          2993 => x"98",
          2994 => x"9c",
          2995 => x"52",
          2996 => x"51",
          2997 => x"82",
          2998 => x"54",
          2999 => x"93",
          3000 => x"a0",
          3001 => x"a4",
          3002 => x"52",
          3003 => x"51",
          3004 => x"82",
          3005 => x"54",
          3006 => x"93",
          3007 => x"a8",
          3008 => x"ac",
          3009 => x"52",
          3010 => x"51",
          3011 => x"82",
          3012 => x"54",
          3013 => x"8d",
          3014 => x"e8",
          3015 => x"f7",
          3016 => x"f1",
          3017 => x"eb",
          3018 => x"80",
          3019 => x"82",
          3020 => x"52",
          3021 => x"51",
          3022 => x"82",
          3023 => x"54",
          3024 => x"8d",
          3025 => x"ea",
          3026 => x"f8",
          3027 => x"c5",
          3028 => x"dd",
          3029 => x"80",
          3030 => x"81",
          3031 => x"83",
          3032 => x"89",
          3033 => x"73",
          3034 => x"38",
          3035 => x"51",
          3036 => x"82",
          3037 => x"54",
          3038 => x"88",
          3039 => x"d0",
          3040 => x"3f",
          3041 => x"33",
          3042 => x"2e",
          3043 => x"f8",
          3044 => x"9d",
          3045 => x"e6",
          3046 => x"80",
          3047 => x"81",
          3048 => x"83",
          3049 => x"f8",
          3050 => x"85",
          3051 => x"c0",
          3052 => x"f9",
          3053 => x"dd",
          3054 => x"c4",
          3055 => x"f9",
          3056 => x"d1",
          3057 => x"c8",
          3058 => x"f9",
          3059 => x"c5",
          3060 => x"f8",
          3061 => x"3f",
          3062 => x"22",
          3063 => x"80",
          3064 => x"3f",
          3065 => x"08",
          3066 => x"c0",
          3067 => x"ea",
          3068 => x"8c",
          3069 => x"84",
          3070 => x"71",
          3071 => x"82",
          3072 => x"52",
          3073 => x"51",
          3074 => x"82",
          3075 => x"54",
          3076 => x"a8",
          3077 => x"d4",
          3078 => x"84",
          3079 => x"51",
          3080 => x"82",
          3081 => x"bd",
          3082 => x"76",
          3083 => x"54",
          3084 => x"08",
          3085 => x"d4",
          3086 => x"3f",
          3087 => x"33",
          3088 => x"2e",
          3089 => x"89",
          3090 => x"bd",
          3091 => x"75",
          3092 => x"3f",
          3093 => x"08",
          3094 => x"29",
          3095 => x"54",
          3096 => x"ec",
          3097 => x"fb",
          3098 => x"a9",
          3099 => x"e4",
          3100 => x"3f",
          3101 => x"04",
          3102 => x"02",
          3103 => x"ff",
          3104 => x"84",
          3105 => x"71",
          3106 => x"0b",
          3107 => x"05",
          3108 => x"04",
          3109 => x"51",
          3110 => x"fb",
          3111 => x"39",
          3112 => x"51",
          3113 => x"fb",
          3114 => x"39",
          3115 => x"51",
          3116 => x"fb",
          3117 => x"f9",
          3118 => x"0d",
          3119 => x"80",
          3120 => x"0b",
          3121 => x"84",
          3122 => x"89",
          3123 => x"c0",
          3124 => x"04",
          3125 => x"02",
          3126 => x"53",
          3127 => x"09",
          3128 => x"38",
          3129 => x"3f",
          3130 => x"08",
          3131 => x"2e",
          3132 => x"72",
          3133 => x"84",
          3134 => x"82",
          3135 => x"8f",
          3136 => x"fc",
          3137 => x"80",
          3138 => x"72",
          3139 => x"84",
          3140 => x"fe",
          3141 => x"97",
          3142 => x"8c",
          3143 => x"82",
          3144 => x"54",
          3145 => x"3f",
          3146 => x"fc",
          3147 => x"0d",
          3148 => x"0d",
          3149 => x"33",
          3150 => x"06",
          3151 => x"80",
          3152 => x"72",
          3153 => x"51",
          3154 => x"ff",
          3155 => x"39",
          3156 => x"04",
          3157 => x"77",
          3158 => x"08",
          3159 => x"fc",
          3160 => x"73",
          3161 => x"ff",
          3162 => x"71",
          3163 => x"38",
          3164 => x"06",
          3165 => x"54",
          3166 => x"e7",
          3167 => x"8c",
          3168 => x"3d",
          3169 => x"3d",
          3170 => x"59",
          3171 => x"81",
          3172 => x"56",
          3173 => x"84",
          3174 => x"a5",
          3175 => x"06",
          3176 => x"80",
          3177 => x"81",
          3178 => x"58",
          3179 => x"b0",
          3180 => x"06",
          3181 => x"5a",
          3182 => x"ad",
          3183 => x"06",
          3184 => x"5a",
          3185 => x"05",
          3186 => x"75",
          3187 => x"81",
          3188 => x"77",
          3189 => x"08",
          3190 => x"05",
          3191 => x"5d",
          3192 => x"39",
          3193 => x"72",
          3194 => x"38",
          3195 => x"7b",
          3196 => x"05",
          3197 => x"70",
          3198 => x"33",
          3199 => x"39",
          3200 => x"32",
          3201 => x"72",
          3202 => x"78",
          3203 => x"70",
          3204 => x"07",
          3205 => x"07",
          3206 => x"51",
          3207 => x"80",
          3208 => x"79",
          3209 => x"70",
          3210 => x"33",
          3211 => x"80",
          3212 => x"38",
          3213 => x"e0",
          3214 => x"38",
          3215 => x"81",
          3216 => x"53",
          3217 => x"2e",
          3218 => x"73",
          3219 => x"a2",
          3220 => x"c3",
          3221 => x"38",
          3222 => x"24",
          3223 => x"80",
          3224 => x"8c",
          3225 => x"39",
          3226 => x"2e",
          3227 => x"81",
          3228 => x"80",
          3229 => x"80",
          3230 => x"d5",
          3231 => x"73",
          3232 => x"8e",
          3233 => x"39",
          3234 => x"2e",
          3235 => x"80",
          3236 => x"84",
          3237 => x"56",
          3238 => x"74",
          3239 => x"72",
          3240 => x"38",
          3241 => x"15",
          3242 => x"54",
          3243 => x"38",
          3244 => x"56",
          3245 => x"81",
          3246 => x"72",
          3247 => x"38",
          3248 => x"90",
          3249 => x"06",
          3250 => x"2e",
          3251 => x"51",
          3252 => x"74",
          3253 => x"53",
          3254 => x"fd",
          3255 => x"51",
          3256 => x"ef",
          3257 => x"19",
          3258 => x"53",
          3259 => x"39",
          3260 => x"39",
          3261 => x"39",
          3262 => x"39",
          3263 => x"39",
          3264 => x"d0",
          3265 => x"39",
          3266 => x"70",
          3267 => x"53",
          3268 => x"88",
          3269 => x"19",
          3270 => x"39",
          3271 => x"54",
          3272 => x"74",
          3273 => x"70",
          3274 => x"07",
          3275 => x"55",
          3276 => x"80",
          3277 => x"72",
          3278 => x"38",
          3279 => x"90",
          3280 => x"80",
          3281 => x"5e",
          3282 => x"74",
          3283 => x"3f",
          3284 => x"08",
          3285 => x"7c",
          3286 => x"54",
          3287 => x"82",
          3288 => x"55",
          3289 => x"92",
          3290 => x"53",
          3291 => x"2e",
          3292 => x"14",
          3293 => x"ff",
          3294 => x"14",
          3295 => x"70",
          3296 => x"34",
          3297 => x"30",
          3298 => x"9f",
          3299 => x"57",
          3300 => x"85",
          3301 => x"b1",
          3302 => x"2a",
          3303 => x"51",
          3304 => x"2e",
          3305 => x"3d",
          3306 => x"05",
          3307 => x"34",
          3308 => x"76",
          3309 => x"54",
          3310 => x"72",
          3311 => x"54",
          3312 => x"70",
          3313 => x"56",
          3314 => x"81",
          3315 => x"7b",
          3316 => x"73",
          3317 => x"3f",
          3318 => x"53",
          3319 => x"74",
          3320 => x"53",
          3321 => x"eb",
          3322 => x"77",
          3323 => x"53",
          3324 => x"14",
          3325 => x"54",
          3326 => x"3f",
          3327 => x"74",
          3328 => x"53",
          3329 => x"fb",
          3330 => x"51",
          3331 => x"ef",
          3332 => x"0d",
          3333 => x"0d",
          3334 => x"70",
          3335 => x"08",
          3336 => x"51",
          3337 => x"85",
          3338 => x"fe",
          3339 => x"82",
          3340 => x"85",
          3341 => x"52",
          3342 => x"ca",
          3343 => x"84",
          3344 => x"73",
          3345 => x"82",
          3346 => x"84",
          3347 => x"fd",
          3348 => x"8c",
          3349 => x"82",
          3350 => x"87",
          3351 => x"53",
          3352 => x"fa",
          3353 => x"82",
          3354 => x"85",
          3355 => x"fb",
          3356 => x"79",
          3357 => x"08",
          3358 => x"57",
          3359 => x"71",
          3360 => x"e0",
          3361 => x"80",
          3362 => x"2d",
          3363 => x"08",
          3364 => x"53",
          3365 => x"80",
          3366 => x"8d",
          3367 => x"72",
          3368 => x"30",
          3369 => x"51",
          3370 => x"80",
          3371 => x"71",
          3372 => x"38",
          3373 => x"97",
          3374 => x"25",
          3375 => x"16",
          3376 => x"25",
          3377 => x"14",
          3378 => x"34",
          3379 => x"72",
          3380 => x"3f",
          3381 => x"73",
          3382 => x"72",
          3383 => x"f7",
          3384 => x"53",
          3385 => x"ec",
          3386 => x"0d",
          3387 => x"0d",
          3388 => x"08",
          3389 => x"80",
          3390 => x"76",
          3391 => x"ef",
          3392 => x"8d",
          3393 => x"3d",
          3394 => x"3d",
          3395 => x"5a",
          3396 => x"7a",
          3397 => x"08",
          3398 => x"53",
          3399 => x"09",
          3400 => x"38",
          3401 => x"0c",
          3402 => x"ad",
          3403 => x"06",
          3404 => x"76",
          3405 => x"0c",
          3406 => x"33",
          3407 => x"73",
          3408 => x"81",
          3409 => x"38",
          3410 => x"05",
          3411 => x"08",
          3412 => x"53",
          3413 => x"2e",
          3414 => x"57",
          3415 => x"2e",
          3416 => x"39",
          3417 => x"13",
          3418 => x"08",
          3419 => x"53",
          3420 => x"55",
          3421 => x"80",
          3422 => x"14",
          3423 => x"88",
          3424 => x"27",
          3425 => x"eb",
          3426 => x"53",
          3427 => x"89",
          3428 => x"38",
          3429 => x"55",
          3430 => x"8a",
          3431 => x"a0",
          3432 => x"c2",
          3433 => x"74",
          3434 => x"e0",
          3435 => x"ff",
          3436 => x"d0",
          3437 => x"ff",
          3438 => x"90",
          3439 => x"38",
          3440 => x"81",
          3441 => x"53",
          3442 => x"ca",
          3443 => x"27",
          3444 => x"77",
          3445 => x"08",
          3446 => x"0c",
          3447 => x"33",
          3448 => x"ff",
          3449 => x"80",
          3450 => x"74",
          3451 => x"79",
          3452 => x"74",
          3453 => x"0c",
          3454 => x"04",
          3455 => x"7a",
          3456 => x"80",
          3457 => x"58",
          3458 => x"33",
          3459 => x"a0",
          3460 => x"06",
          3461 => x"13",
          3462 => x"39",
          3463 => x"09",
          3464 => x"38",
          3465 => x"11",
          3466 => x"08",
          3467 => x"54",
          3468 => x"2e",
          3469 => x"80",
          3470 => x"08",
          3471 => x"0c",
          3472 => x"33",
          3473 => x"80",
          3474 => x"38",
          3475 => x"80",
          3476 => x"38",
          3477 => x"57",
          3478 => x"0c",
          3479 => x"33",
          3480 => x"39",
          3481 => x"74",
          3482 => x"38",
          3483 => x"80",
          3484 => x"89",
          3485 => x"38",
          3486 => x"d0",
          3487 => x"55",
          3488 => x"80",
          3489 => x"39",
          3490 => x"d9",
          3491 => x"80",
          3492 => x"27",
          3493 => x"80",
          3494 => x"89",
          3495 => x"70",
          3496 => x"55",
          3497 => x"70",
          3498 => x"55",
          3499 => x"27",
          3500 => x"14",
          3501 => x"06",
          3502 => x"74",
          3503 => x"73",
          3504 => x"38",
          3505 => x"14",
          3506 => x"05",
          3507 => x"08",
          3508 => x"54",
          3509 => x"39",
          3510 => x"84",
          3511 => x"55",
          3512 => x"81",
          3513 => x"8c",
          3514 => x"3d",
          3515 => x"3d",
          3516 => x"05",
          3517 => x"52",
          3518 => x"87",
          3519 => x"f4",
          3520 => x"71",
          3521 => x"0c",
          3522 => x"04",
          3523 => x"02",
          3524 => x"02",
          3525 => x"05",
          3526 => x"83",
          3527 => x"26",
          3528 => x"72",
          3529 => x"c0",
          3530 => x"53",
          3531 => x"74",
          3532 => x"38",
          3533 => x"73",
          3534 => x"c0",
          3535 => x"51",
          3536 => x"85",
          3537 => x"98",
          3538 => x"52",
          3539 => x"82",
          3540 => x"70",
          3541 => x"38",
          3542 => x"8c",
          3543 => x"ec",
          3544 => x"fc",
          3545 => x"52",
          3546 => x"87",
          3547 => x"08",
          3548 => x"2e",
          3549 => x"82",
          3550 => x"34",
          3551 => x"13",
          3552 => x"82",
          3553 => x"86",
          3554 => x"f3",
          3555 => x"62",
          3556 => x"05",
          3557 => x"57",
          3558 => x"83",
          3559 => x"fe",
          3560 => x"8c",
          3561 => x"06",
          3562 => x"71",
          3563 => x"71",
          3564 => x"2b",
          3565 => x"80",
          3566 => x"92",
          3567 => x"c0",
          3568 => x"41",
          3569 => x"5a",
          3570 => x"87",
          3571 => x"0c",
          3572 => x"84",
          3573 => x"08",
          3574 => x"70",
          3575 => x"53",
          3576 => x"2e",
          3577 => x"08",
          3578 => x"70",
          3579 => x"34",
          3580 => x"80",
          3581 => x"53",
          3582 => x"2e",
          3583 => x"53",
          3584 => x"26",
          3585 => x"80",
          3586 => x"87",
          3587 => x"08",
          3588 => x"38",
          3589 => x"8c",
          3590 => x"80",
          3591 => x"78",
          3592 => x"99",
          3593 => x"0c",
          3594 => x"8c",
          3595 => x"08",
          3596 => x"51",
          3597 => x"38",
          3598 => x"8d",
          3599 => x"17",
          3600 => x"81",
          3601 => x"53",
          3602 => x"2e",
          3603 => x"fc",
          3604 => x"52",
          3605 => x"7d",
          3606 => x"ed",
          3607 => x"80",
          3608 => x"71",
          3609 => x"38",
          3610 => x"53",
          3611 => x"ec",
          3612 => x"0d",
          3613 => x"0d",
          3614 => x"02",
          3615 => x"05",
          3616 => x"58",
          3617 => x"80",
          3618 => x"fc",
          3619 => x"8c",
          3620 => x"06",
          3621 => x"71",
          3622 => x"81",
          3623 => x"38",
          3624 => x"2b",
          3625 => x"80",
          3626 => x"92",
          3627 => x"c0",
          3628 => x"40",
          3629 => x"5a",
          3630 => x"c0",
          3631 => x"76",
          3632 => x"76",
          3633 => x"75",
          3634 => x"2a",
          3635 => x"51",
          3636 => x"80",
          3637 => x"7a",
          3638 => x"5c",
          3639 => x"81",
          3640 => x"81",
          3641 => x"06",
          3642 => x"80",
          3643 => x"87",
          3644 => x"08",
          3645 => x"38",
          3646 => x"8c",
          3647 => x"80",
          3648 => x"77",
          3649 => x"99",
          3650 => x"0c",
          3651 => x"8c",
          3652 => x"08",
          3653 => x"51",
          3654 => x"38",
          3655 => x"8d",
          3656 => x"70",
          3657 => x"84",
          3658 => x"5b",
          3659 => x"2e",
          3660 => x"fc",
          3661 => x"52",
          3662 => x"7d",
          3663 => x"f8",
          3664 => x"80",
          3665 => x"71",
          3666 => x"38",
          3667 => x"53",
          3668 => x"ec",
          3669 => x"0d",
          3670 => x"0d",
          3671 => x"05",
          3672 => x"02",
          3673 => x"05",
          3674 => x"54",
          3675 => x"fe",
          3676 => x"ec",
          3677 => x"53",
          3678 => x"80",
          3679 => x"0b",
          3680 => x"8c",
          3681 => x"71",
          3682 => x"dc",
          3683 => x"24",
          3684 => x"84",
          3685 => x"92",
          3686 => x"54",
          3687 => x"8d",
          3688 => x"39",
          3689 => x"80",
          3690 => x"cb",
          3691 => x"70",
          3692 => x"81",
          3693 => x"52",
          3694 => x"8a",
          3695 => x"98",
          3696 => x"71",
          3697 => x"c0",
          3698 => x"52",
          3699 => x"81",
          3700 => x"c0",
          3701 => x"53",
          3702 => x"82",
          3703 => x"71",
          3704 => x"39",
          3705 => x"39",
          3706 => x"77",
          3707 => x"81",
          3708 => x"72",
          3709 => x"84",
          3710 => x"73",
          3711 => x"0c",
          3712 => x"04",
          3713 => x"74",
          3714 => x"71",
          3715 => x"2b",
          3716 => x"ec",
          3717 => x"84",
          3718 => x"fd",
          3719 => x"83",
          3720 => x"12",
          3721 => x"2b",
          3722 => x"07",
          3723 => x"70",
          3724 => x"2b",
          3725 => x"07",
          3726 => x"0c",
          3727 => x"56",
          3728 => x"3d",
          3729 => x"3d",
          3730 => x"84",
          3731 => x"22",
          3732 => x"72",
          3733 => x"54",
          3734 => x"2a",
          3735 => x"34",
          3736 => x"04",
          3737 => x"73",
          3738 => x"70",
          3739 => x"05",
          3740 => x"88",
          3741 => x"72",
          3742 => x"54",
          3743 => x"2a",
          3744 => x"70",
          3745 => x"34",
          3746 => x"51",
          3747 => x"83",
          3748 => x"fe",
          3749 => x"75",
          3750 => x"51",
          3751 => x"92",
          3752 => x"81",
          3753 => x"73",
          3754 => x"55",
          3755 => x"51",
          3756 => x"3d",
          3757 => x"3d",
          3758 => x"76",
          3759 => x"72",
          3760 => x"05",
          3761 => x"11",
          3762 => x"38",
          3763 => x"04",
          3764 => x"78",
          3765 => x"56",
          3766 => x"81",
          3767 => x"74",
          3768 => x"56",
          3769 => x"31",
          3770 => x"52",
          3771 => x"80",
          3772 => x"71",
          3773 => x"38",
          3774 => x"ec",
          3775 => x"0d",
          3776 => x"0d",
          3777 => x"51",
          3778 => x"73",
          3779 => x"81",
          3780 => x"33",
          3781 => x"38",
          3782 => x"8c",
          3783 => x"3d",
          3784 => x"0b",
          3785 => x"0c",
          3786 => x"82",
          3787 => x"04",
          3788 => x"7b",
          3789 => x"83",
          3790 => x"5a",
          3791 => x"80",
          3792 => x"54",
          3793 => x"53",
          3794 => x"53",
          3795 => x"52",
          3796 => x"3f",
          3797 => x"08",
          3798 => x"81",
          3799 => x"82",
          3800 => x"83",
          3801 => x"16",
          3802 => x"18",
          3803 => x"18",
          3804 => x"58",
          3805 => x"9f",
          3806 => x"33",
          3807 => x"2e",
          3808 => x"93",
          3809 => x"76",
          3810 => x"52",
          3811 => x"51",
          3812 => x"83",
          3813 => x"79",
          3814 => x"0c",
          3815 => x"04",
          3816 => x"78",
          3817 => x"80",
          3818 => x"17",
          3819 => x"38",
          3820 => x"fc",
          3821 => x"ec",
          3822 => x"8c",
          3823 => x"38",
          3824 => x"53",
          3825 => x"81",
          3826 => x"f7",
          3827 => x"8c",
          3828 => x"2e",
          3829 => x"55",
          3830 => x"b0",
          3831 => x"82",
          3832 => x"88",
          3833 => x"f8",
          3834 => x"70",
          3835 => x"c0",
          3836 => x"ec",
          3837 => x"8c",
          3838 => x"91",
          3839 => x"55",
          3840 => x"09",
          3841 => x"f0",
          3842 => x"33",
          3843 => x"2e",
          3844 => x"80",
          3845 => x"80",
          3846 => x"ec",
          3847 => x"17",
          3848 => x"fd",
          3849 => x"d4",
          3850 => x"b2",
          3851 => x"96",
          3852 => x"85",
          3853 => x"75",
          3854 => x"3f",
          3855 => x"e4",
          3856 => x"98",
          3857 => x"9c",
          3858 => x"08",
          3859 => x"17",
          3860 => x"3f",
          3861 => x"52",
          3862 => x"51",
          3863 => x"a0",
          3864 => x"05",
          3865 => x"0c",
          3866 => x"75",
          3867 => x"33",
          3868 => x"3f",
          3869 => x"34",
          3870 => x"52",
          3871 => x"51",
          3872 => x"82",
          3873 => x"80",
          3874 => x"81",
          3875 => x"8c",
          3876 => x"3d",
          3877 => x"3d",
          3878 => x"1a",
          3879 => x"fe",
          3880 => x"54",
          3881 => x"73",
          3882 => x"8a",
          3883 => x"71",
          3884 => x"08",
          3885 => x"75",
          3886 => x"0c",
          3887 => x"04",
          3888 => x"7a",
          3889 => x"56",
          3890 => x"77",
          3891 => x"38",
          3892 => x"08",
          3893 => x"38",
          3894 => x"54",
          3895 => x"2e",
          3896 => x"72",
          3897 => x"38",
          3898 => x"8d",
          3899 => x"39",
          3900 => x"81",
          3901 => x"b6",
          3902 => x"2a",
          3903 => x"2a",
          3904 => x"05",
          3905 => x"55",
          3906 => x"82",
          3907 => x"81",
          3908 => x"83",
          3909 => x"b4",
          3910 => x"17",
          3911 => x"a4",
          3912 => x"55",
          3913 => x"57",
          3914 => x"3f",
          3915 => x"08",
          3916 => x"74",
          3917 => x"14",
          3918 => x"70",
          3919 => x"07",
          3920 => x"71",
          3921 => x"52",
          3922 => x"72",
          3923 => x"75",
          3924 => x"58",
          3925 => x"76",
          3926 => x"15",
          3927 => x"73",
          3928 => x"3f",
          3929 => x"08",
          3930 => x"76",
          3931 => x"06",
          3932 => x"05",
          3933 => x"3f",
          3934 => x"08",
          3935 => x"06",
          3936 => x"76",
          3937 => x"15",
          3938 => x"73",
          3939 => x"3f",
          3940 => x"08",
          3941 => x"82",
          3942 => x"06",
          3943 => x"05",
          3944 => x"3f",
          3945 => x"08",
          3946 => x"58",
          3947 => x"58",
          3948 => x"ec",
          3949 => x"0d",
          3950 => x"0d",
          3951 => x"5a",
          3952 => x"59",
          3953 => x"82",
          3954 => x"98",
          3955 => x"82",
          3956 => x"33",
          3957 => x"2e",
          3958 => x"72",
          3959 => x"38",
          3960 => x"8d",
          3961 => x"39",
          3962 => x"81",
          3963 => x"f7",
          3964 => x"2a",
          3965 => x"2a",
          3966 => x"05",
          3967 => x"55",
          3968 => x"82",
          3969 => x"59",
          3970 => x"08",
          3971 => x"74",
          3972 => x"16",
          3973 => x"16",
          3974 => x"59",
          3975 => x"53",
          3976 => x"8f",
          3977 => x"2b",
          3978 => x"74",
          3979 => x"71",
          3980 => x"72",
          3981 => x"0b",
          3982 => x"74",
          3983 => x"17",
          3984 => x"75",
          3985 => x"3f",
          3986 => x"08",
          3987 => x"ec",
          3988 => x"38",
          3989 => x"06",
          3990 => x"78",
          3991 => x"54",
          3992 => x"77",
          3993 => x"33",
          3994 => x"71",
          3995 => x"51",
          3996 => x"34",
          3997 => x"76",
          3998 => x"17",
          3999 => x"75",
          4000 => x"3f",
          4001 => x"08",
          4002 => x"ec",
          4003 => x"38",
          4004 => x"ff",
          4005 => x"10",
          4006 => x"76",
          4007 => x"51",
          4008 => x"be",
          4009 => x"2a",
          4010 => x"05",
          4011 => x"f9",
          4012 => x"8c",
          4013 => x"82",
          4014 => x"ab",
          4015 => x"0a",
          4016 => x"2b",
          4017 => x"70",
          4018 => x"70",
          4019 => x"54",
          4020 => x"82",
          4021 => x"8f",
          4022 => x"07",
          4023 => x"f7",
          4024 => x"0b",
          4025 => x"78",
          4026 => x"0c",
          4027 => x"04",
          4028 => x"7a",
          4029 => x"08",
          4030 => x"59",
          4031 => x"a4",
          4032 => x"17",
          4033 => x"38",
          4034 => x"aa",
          4035 => x"73",
          4036 => x"fd",
          4037 => x"8c",
          4038 => x"82",
          4039 => x"80",
          4040 => x"39",
          4041 => x"eb",
          4042 => x"80",
          4043 => x"8c",
          4044 => x"80",
          4045 => x"52",
          4046 => x"84",
          4047 => x"ec",
          4048 => x"8c",
          4049 => x"2e",
          4050 => x"82",
          4051 => x"81",
          4052 => x"82",
          4053 => x"ff",
          4054 => x"80",
          4055 => x"75",
          4056 => x"3f",
          4057 => x"08",
          4058 => x"16",
          4059 => x"90",
          4060 => x"55",
          4061 => x"27",
          4062 => x"15",
          4063 => x"84",
          4064 => x"07",
          4065 => x"17",
          4066 => x"76",
          4067 => x"a6",
          4068 => x"73",
          4069 => x"0c",
          4070 => x"04",
          4071 => x"7c",
          4072 => x"59",
          4073 => x"95",
          4074 => x"08",
          4075 => x"2e",
          4076 => x"17",
          4077 => x"b2",
          4078 => x"ae",
          4079 => x"7a",
          4080 => x"3f",
          4081 => x"82",
          4082 => x"27",
          4083 => x"82",
          4084 => x"55",
          4085 => x"08",
          4086 => x"d2",
          4087 => x"08",
          4088 => x"08",
          4089 => x"38",
          4090 => x"17",
          4091 => x"54",
          4092 => x"82",
          4093 => x"7a",
          4094 => x"06",
          4095 => x"81",
          4096 => x"17",
          4097 => x"83",
          4098 => x"75",
          4099 => x"f9",
          4100 => x"59",
          4101 => x"08",
          4102 => x"81",
          4103 => x"82",
          4104 => x"59",
          4105 => x"08",
          4106 => x"70",
          4107 => x"25",
          4108 => x"82",
          4109 => x"54",
          4110 => x"55",
          4111 => x"38",
          4112 => x"08",
          4113 => x"38",
          4114 => x"54",
          4115 => x"90",
          4116 => x"18",
          4117 => x"38",
          4118 => x"39",
          4119 => x"38",
          4120 => x"16",
          4121 => x"08",
          4122 => x"38",
          4123 => x"78",
          4124 => x"38",
          4125 => x"51",
          4126 => x"82",
          4127 => x"80",
          4128 => x"80",
          4129 => x"ec",
          4130 => x"09",
          4131 => x"38",
          4132 => x"08",
          4133 => x"ec",
          4134 => x"30",
          4135 => x"80",
          4136 => x"07",
          4137 => x"55",
          4138 => x"38",
          4139 => x"09",
          4140 => x"ae",
          4141 => x"80",
          4142 => x"53",
          4143 => x"51",
          4144 => x"82",
          4145 => x"82",
          4146 => x"30",
          4147 => x"ec",
          4148 => x"25",
          4149 => x"79",
          4150 => x"38",
          4151 => x"8f",
          4152 => x"79",
          4153 => x"f9",
          4154 => x"8c",
          4155 => x"74",
          4156 => x"8c",
          4157 => x"17",
          4158 => x"90",
          4159 => x"54",
          4160 => x"86",
          4161 => x"90",
          4162 => x"17",
          4163 => x"54",
          4164 => x"34",
          4165 => x"56",
          4166 => x"90",
          4167 => x"80",
          4168 => x"82",
          4169 => x"55",
          4170 => x"56",
          4171 => x"82",
          4172 => x"8c",
          4173 => x"f8",
          4174 => x"70",
          4175 => x"f0",
          4176 => x"ec",
          4177 => x"56",
          4178 => x"08",
          4179 => x"7b",
          4180 => x"f6",
          4181 => x"8c",
          4182 => x"8c",
          4183 => x"17",
          4184 => x"80",
          4185 => x"b4",
          4186 => x"57",
          4187 => x"77",
          4188 => x"81",
          4189 => x"15",
          4190 => x"78",
          4191 => x"81",
          4192 => x"53",
          4193 => x"15",
          4194 => x"e9",
          4195 => x"ec",
          4196 => x"df",
          4197 => x"22",
          4198 => x"30",
          4199 => x"70",
          4200 => x"51",
          4201 => x"82",
          4202 => x"8a",
          4203 => x"f8",
          4204 => x"7c",
          4205 => x"56",
          4206 => x"80",
          4207 => x"f1",
          4208 => x"06",
          4209 => x"e9",
          4210 => x"18",
          4211 => x"08",
          4212 => x"38",
          4213 => x"82",
          4214 => x"38",
          4215 => x"54",
          4216 => x"74",
          4217 => x"82",
          4218 => x"22",
          4219 => x"79",
          4220 => x"38",
          4221 => x"98",
          4222 => x"cd",
          4223 => x"22",
          4224 => x"54",
          4225 => x"26",
          4226 => x"52",
          4227 => x"b0",
          4228 => x"ec",
          4229 => x"8c",
          4230 => x"2e",
          4231 => x"0b",
          4232 => x"08",
          4233 => x"98",
          4234 => x"8c",
          4235 => x"85",
          4236 => x"bd",
          4237 => x"31",
          4238 => x"73",
          4239 => x"f4",
          4240 => x"8c",
          4241 => x"18",
          4242 => x"18",
          4243 => x"08",
          4244 => x"72",
          4245 => x"38",
          4246 => x"58",
          4247 => x"89",
          4248 => x"18",
          4249 => x"ff",
          4250 => x"05",
          4251 => x"80",
          4252 => x"8c",
          4253 => x"3d",
          4254 => x"3d",
          4255 => x"08",
          4256 => x"a0",
          4257 => x"54",
          4258 => x"77",
          4259 => x"80",
          4260 => x"0c",
          4261 => x"53",
          4262 => x"80",
          4263 => x"38",
          4264 => x"06",
          4265 => x"b5",
          4266 => x"98",
          4267 => x"14",
          4268 => x"92",
          4269 => x"2a",
          4270 => x"56",
          4271 => x"26",
          4272 => x"80",
          4273 => x"16",
          4274 => x"77",
          4275 => x"53",
          4276 => x"38",
          4277 => x"51",
          4278 => x"82",
          4279 => x"53",
          4280 => x"0b",
          4281 => x"08",
          4282 => x"38",
          4283 => x"8c",
          4284 => x"2e",
          4285 => x"98",
          4286 => x"8c",
          4287 => x"80",
          4288 => x"8a",
          4289 => x"15",
          4290 => x"80",
          4291 => x"14",
          4292 => x"51",
          4293 => x"82",
          4294 => x"53",
          4295 => x"8c",
          4296 => x"2e",
          4297 => x"82",
          4298 => x"ec",
          4299 => x"ba",
          4300 => x"82",
          4301 => x"ff",
          4302 => x"82",
          4303 => x"52",
          4304 => x"f3",
          4305 => x"ec",
          4306 => x"72",
          4307 => x"72",
          4308 => x"f2",
          4309 => x"8c",
          4310 => x"15",
          4311 => x"15",
          4312 => x"b4",
          4313 => x"0c",
          4314 => x"82",
          4315 => x"8a",
          4316 => x"f7",
          4317 => x"7d",
          4318 => x"5b",
          4319 => x"76",
          4320 => x"3f",
          4321 => x"08",
          4322 => x"ec",
          4323 => x"38",
          4324 => x"08",
          4325 => x"08",
          4326 => x"f0",
          4327 => x"8c",
          4328 => x"82",
          4329 => x"80",
          4330 => x"8c",
          4331 => x"18",
          4332 => x"51",
          4333 => x"81",
          4334 => x"81",
          4335 => x"81",
          4336 => x"ec",
          4337 => x"83",
          4338 => x"77",
          4339 => x"72",
          4340 => x"38",
          4341 => x"75",
          4342 => x"81",
          4343 => x"a5",
          4344 => x"ec",
          4345 => x"52",
          4346 => x"8e",
          4347 => x"ec",
          4348 => x"8c",
          4349 => x"2e",
          4350 => x"73",
          4351 => x"81",
          4352 => x"87",
          4353 => x"8c",
          4354 => x"3d",
          4355 => x"3d",
          4356 => x"11",
          4357 => x"ec",
          4358 => x"ec",
          4359 => x"ff",
          4360 => x"33",
          4361 => x"71",
          4362 => x"81",
          4363 => x"94",
          4364 => x"d0",
          4365 => x"ec",
          4366 => x"73",
          4367 => x"82",
          4368 => x"85",
          4369 => x"fc",
          4370 => x"79",
          4371 => x"ff",
          4372 => x"12",
          4373 => x"eb",
          4374 => x"70",
          4375 => x"72",
          4376 => x"81",
          4377 => x"73",
          4378 => x"94",
          4379 => x"d6",
          4380 => x"0d",
          4381 => x"0d",
          4382 => x"55",
          4383 => x"5a",
          4384 => x"08",
          4385 => x"8a",
          4386 => x"08",
          4387 => x"ee",
          4388 => x"8c",
          4389 => x"82",
          4390 => x"80",
          4391 => x"15",
          4392 => x"55",
          4393 => x"38",
          4394 => x"e6",
          4395 => x"33",
          4396 => x"70",
          4397 => x"58",
          4398 => x"86",
          4399 => x"8c",
          4400 => x"73",
          4401 => x"83",
          4402 => x"73",
          4403 => x"38",
          4404 => x"06",
          4405 => x"80",
          4406 => x"75",
          4407 => x"38",
          4408 => x"08",
          4409 => x"54",
          4410 => x"2e",
          4411 => x"83",
          4412 => x"73",
          4413 => x"38",
          4414 => x"51",
          4415 => x"82",
          4416 => x"58",
          4417 => x"08",
          4418 => x"15",
          4419 => x"38",
          4420 => x"0b",
          4421 => x"77",
          4422 => x"0c",
          4423 => x"04",
          4424 => x"77",
          4425 => x"54",
          4426 => x"51",
          4427 => x"82",
          4428 => x"55",
          4429 => x"08",
          4430 => x"14",
          4431 => x"51",
          4432 => x"82",
          4433 => x"55",
          4434 => x"08",
          4435 => x"53",
          4436 => x"08",
          4437 => x"08",
          4438 => x"3f",
          4439 => x"14",
          4440 => x"08",
          4441 => x"3f",
          4442 => x"17",
          4443 => x"8c",
          4444 => x"3d",
          4445 => x"3d",
          4446 => x"08",
          4447 => x"54",
          4448 => x"53",
          4449 => x"82",
          4450 => x"8d",
          4451 => x"08",
          4452 => x"34",
          4453 => x"15",
          4454 => x"0d",
          4455 => x"0d",
          4456 => x"57",
          4457 => x"17",
          4458 => x"08",
          4459 => x"82",
          4460 => x"89",
          4461 => x"55",
          4462 => x"14",
          4463 => x"16",
          4464 => x"71",
          4465 => x"38",
          4466 => x"09",
          4467 => x"38",
          4468 => x"73",
          4469 => x"81",
          4470 => x"ae",
          4471 => x"05",
          4472 => x"15",
          4473 => x"70",
          4474 => x"34",
          4475 => x"8a",
          4476 => x"38",
          4477 => x"05",
          4478 => x"81",
          4479 => x"17",
          4480 => x"12",
          4481 => x"34",
          4482 => x"9c",
          4483 => x"e8",
          4484 => x"8c",
          4485 => x"0c",
          4486 => x"e7",
          4487 => x"8c",
          4488 => x"17",
          4489 => x"51",
          4490 => x"82",
          4491 => x"84",
          4492 => x"3d",
          4493 => x"3d",
          4494 => x"08",
          4495 => x"61",
          4496 => x"55",
          4497 => x"2e",
          4498 => x"55",
          4499 => x"2e",
          4500 => x"80",
          4501 => x"94",
          4502 => x"1c",
          4503 => x"81",
          4504 => x"61",
          4505 => x"56",
          4506 => x"2e",
          4507 => x"83",
          4508 => x"73",
          4509 => x"70",
          4510 => x"25",
          4511 => x"51",
          4512 => x"38",
          4513 => x"0c",
          4514 => x"51",
          4515 => x"26",
          4516 => x"80",
          4517 => x"34",
          4518 => x"51",
          4519 => x"82",
          4520 => x"55",
          4521 => x"91",
          4522 => x"1d",
          4523 => x"8b",
          4524 => x"79",
          4525 => x"3f",
          4526 => x"57",
          4527 => x"55",
          4528 => x"2e",
          4529 => x"80",
          4530 => x"18",
          4531 => x"1a",
          4532 => x"70",
          4533 => x"2a",
          4534 => x"07",
          4535 => x"5a",
          4536 => x"8c",
          4537 => x"54",
          4538 => x"81",
          4539 => x"39",
          4540 => x"70",
          4541 => x"2a",
          4542 => x"75",
          4543 => x"8c",
          4544 => x"2e",
          4545 => x"a0",
          4546 => x"38",
          4547 => x"0c",
          4548 => x"76",
          4549 => x"38",
          4550 => x"b8",
          4551 => x"70",
          4552 => x"5a",
          4553 => x"76",
          4554 => x"38",
          4555 => x"70",
          4556 => x"dc",
          4557 => x"72",
          4558 => x"80",
          4559 => x"51",
          4560 => x"73",
          4561 => x"38",
          4562 => x"18",
          4563 => x"1a",
          4564 => x"55",
          4565 => x"2e",
          4566 => x"83",
          4567 => x"73",
          4568 => x"70",
          4569 => x"25",
          4570 => x"51",
          4571 => x"38",
          4572 => x"75",
          4573 => x"81",
          4574 => x"81",
          4575 => x"27",
          4576 => x"73",
          4577 => x"38",
          4578 => x"70",
          4579 => x"32",
          4580 => x"80",
          4581 => x"2a",
          4582 => x"56",
          4583 => x"81",
          4584 => x"57",
          4585 => x"f5",
          4586 => x"2b",
          4587 => x"25",
          4588 => x"80",
          4589 => x"fc",
          4590 => x"57",
          4591 => x"e6",
          4592 => x"8c",
          4593 => x"2e",
          4594 => x"18",
          4595 => x"1a",
          4596 => x"56",
          4597 => x"3f",
          4598 => x"08",
          4599 => x"e8",
          4600 => x"54",
          4601 => x"80",
          4602 => x"17",
          4603 => x"34",
          4604 => x"11",
          4605 => x"74",
          4606 => x"75",
          4607 => x"dc",
          4608 => x"3f",
          4609 => x"08",
          4610 => x"9f",
          4611 => x"99",
          4612 => x"e0",
          4613 => x"ff",
          4614 => x"79",
          4615 => x"74",
          4616 => x"57",
          4617 => x"77",
          4618 => x"76",
          4619 => x"38",
          4620 => x"73",
          4621 => x"09",
          4622 => x"38",
          4623 => x"84",
          4624 => x"27",
          4625 => x"39",
          4626 => x"f2",
          4627 => x"80",
          4628 => x"54",
          4629 => x"34",
          4630 => x"58",
          4631 => x"f2",
          4632 => x"8c",
          4633 => x"82",
          4634 => x"80",
          4635 => x"1b",
          4636 => x"51",
          4637 => x"82",
          4638 => x"56",
          4639 => x"08",
          4640 => x"9c",
          4641 => x"33",
          4642 => x"80",
          4643 => x"38",
          4644 => x"bf",
          4645 => x"86",
          4646 => x"15",
          4647 => x"2a",
          4648 => x"51",
          4649 => x"92",
          4650 => x"79",
          4651 => x"e4",
          4652 => x"8c",
          4653 => x"2e",
          4654 => x"52",
          4655 => x"ba",
          4656 => x"39",
          4657 => x"33",
          4658 => x"80",
          4659 => x"74",
          4660 => x"81",
          4661 => x"38",
          4662 => x"70",
          4663 => x"82",
          4664 => x"54",
          4665 => x"96",
          4666 => x"06",
          4667 => x"2e",
          4668 => x"ff",
          4669 => x"1c",
          4670 => x"80",
          4671 => x"81",
          4672 => x"ba",
          4673 => x"b6",
          4674 => x"2a",
          4675 => x"51",
          4676 => x"38",
          4677 => x"70",
          4678 => x"81",
          4679 => x"55",
          4680 => x"e1",
          4681 => x"08",
          4682 => x"1d",
          4683 => x"7c",
          4684 => x"3f",
          4685 => x"08",
          4686 => x"fa",
          4687 => x"82",
          4688 => x"8f",
          4689 => x"f6",
          4690 => x"5b",
          4691 => x"70",
          4692 => x"59",
          4693 => x"73",
          4694 => x"c6",
          4695 => x"81",
          4696 => x"70",
          4697 => x"52",
          4698 => x"8d",
          4699 => x"38",
          4700 => x"09",
          4701 => x"a5",
          4702 => x"d0",
          4703 => x"ff",
          4704 => x"53",
          4705 => x"91",
          4706 => x"73",
          4707 => x"d0",
          4708 => x"71",
          4709 => x"f7",
          4710 => x"81",
          4711 => x"55",
          4712 => x"55",
          4713 => x"81",
          4714 => x"74",
          4715 => x"56",
          4716 => x"12",
          4717 => x"70",
          4718 => x"38",
          4719 => x"81",
          4720 => x"51",
          4721 => x"51",
          4722 => x"89",
          4723 => x"70",
          4724 => x"53",
          4725 => x"70",
          4726 => x"51",
          4727 => x"09",
          4728 => x"38",
          4729 => x"38",
          4730 => x"77",
          4731 => x"70",
          4732 => x"2a",
          4733 => x"07",
          4734 => x"51",
          4735 => x"8f",
          4736 => x"84",
          4737 => x"83",
          4738 => x"94",
          4739 => x"74",
          4740 => x"38",
          4741 => x"0c",
          4742 => x"86",
          4743 => x"9c",
          4744 => x"82",
          4745 => x"8c",
          4746 => x"fa",
          4747 => x"56",
          4748 => x"17",
          4749 => x"b0",
          4750 => x"52",
          4751 => x"e0",
          4752 => x"82",
          4753 => x"81",
          4754 => x"b2",
          4755 => x"b4",
          4756 => x"ec",
          4757 => x"ff",
          4758 => x"55",
          4759 => x"d5",
          4760 => x"06",
          4761 => x"80",
          4762 => x"33",
          4763 => x"81",
          4764 => x"81",
          4765 => x"81",
          4766 => x"eb",
          4767 => x"70",
          4768 => x"07",
          4769 => x"73",
          4770 => x"81",
          4771 => x"81",
          4772 => x"83",
          4773 => x"ec",
          4774 => x"16",
          4775 => x"3f",
          4776 => x"08",
          4777 => x"ec",
          4778 => x"9d",
          4779 => x"81",
          4780 => x"81",
          4781 => x"e0",
          4782 => x"8c",
          4783 => x"82",
          4784 => x"80",
          4785 => x"82",
          4786 => x"8c",
          4787 => x"3d",
          4788 => x"3d",
          4789 => x"84",
          4790 => x"05",
          4791 => x"80",
          4792 => x"51",
          4793 => x"82",
          4794 => x"58",
          4795 => x"0b",
          4796 => x"08",
          4797 => x"38",
          4798 => x"08",
          4799 => x"8d",
          4800 => x"08",
          4801 => x"56",
          4802 => x"86",
          4803 => x"75",
          4804 => x"fe",
          4805 => x"54",
          4806 => x"2e",
          4807 => x"14",
          4808 => x"ca",
          4809 => x"ec",
          4810 => x"06",
          4811 => x"54",
          4812 => x"38",
          4813 => x"86",
          4814 => x"82",
          4815 => x"06",
          4816 => x"56",
          4817 => x"38",
          4818 => x"80",
          4819 => x"81",
          4820 => x"52",
          4821 => x"51",
          4822 => x"82",
          4823 => x"81",
          4824 => x"81",
          4825 => x"83",
          4826 => x"87",
          4827 => x"2e",
          4828 => x"82",
          4829 => x"06",
          4830 => x"56",
          4831 => x"38",
          4832 => x"74",
          4833 => x"a3",
          4834 => x"ec",
          4835 => x"06",
          4836 => x"2e",
          4837 => x"80",
          4838 => x"3d",
          4839 => x"83",
          4840 => x"15",
          4841 => x"53",
          4842 => x"8d",
          4843 => x"15",
          4844 => x"3f",
          4845 => x"08",
          4846 => x"70",
          4847 => x"0c",
          4848 => x"16",
          4849 => x"80",
          4850 => x"80",
          4851 => x"54",
          4852 => x"84",
          4853 => x"5b",
          4854 => x"80",
          4855 => x"7a",
          4856 => x"fc",
          4857 => x"8c",
          4858 => x"ff",
          4859 => x"77",
          4860 => x"81",
          4861 => x"76",
          4862 => x"81",
          4863 => x"2e",
          4864 => x"8d",
          4865 => x"26",
          4866 => x"bf",
          4867 => x"f4",
          4868 => x"ec",
          4869 => x"ff",
          4870 => x"84",
          4871 => x"81",
          4872 => x"38",
          4873 => x"51",
          4874 => x"82",
          4875 => x"83",
          4876 => x"58",
          4877 => x"80",
          4878 => x"db",
          4879 => x"8c",
          4880 => x"77",
          4881 => x"80",
          4882 => x"82",
          4883 => x"c4",
          4884 => x"11",
          4885 => x"06",
          4886 => x"8d",
          4887 => x"26",
          4888 => x"74",
          4889 => x"78",
          4890 => x"c1",
          4891 => x"59",
          4892 => x"15",
          4893 => x"2e",
          4894 => x"13",
          4895 => x"72",
          4896 => x"38",
          4897 => x"eb",
          4898 => x"14",
          4899 => x"3f",
          4900 => x"08",
          4901 => x"ec",
          4902 => x"23",
          4903 => x"57",
          4904 => x"83",
          4905 => x"c7",
          4906 => x"d8",
          4907 => x"ec",
          4908 => x"ff",
          4909 => x"8d",
          4910 => x"14",
          4911 => x"3f",
          4912 => x"08",
          4913 => x"14",
          4914 => x"3f",
          4915 => x"08",
          4916 => x"06",
          4917 => x"72",
          4918 => x"97",
          4919 => x"22",
          4920 => x"84",
          4921 => x"5a",
          4922 => x"83",
          4923 => x"14",
          4924 => x"79",
          4925 => x"b0",
          4926 => x"8c",
          4927 => x"82",
          4928 => x"80",
          4929 => x"38",
          4930 => x"08",
          4931 => x"ff",
          4932 => x"38",
          4933 => x"83",
          4934 => x"83",
          4935 => x"74",
          4936 => x"85",
          4937 => x"89",
          4938 => x"76",
          4939 => x"c3",
          4940 => x"70",
          4941 => x"7b",
          4942 => x"73",
          4943 => x"17",
          4944 => x"ac",
          4945 => x"55",
          4946 => x"09",
          4947 => x"38",
          4948 => x"51",
          4949 => x"82",
          4950 => x"83",
          4951 => x"53",
          4952 => x"82",
          4953 => x"82",
          4954 => x"e0",
          4955 => x"ab",
          4956 => x"ec",
          4957 => x"0c",
          4958 => x"53",
          4959 => x"56",
          4960 => x"81",
          4961 => x"13",
          4962 => x"74",
          4963 => x"82",
          4964 => x"74",
          4965 => x"81",
          4966 => x"06",
          4967 => x"83",
          4968 => x"2a",
          4969 => x"72",
          4970 => x"26",
          4971 => x"ff",
          4972 => x"0c",
          4973 => x"15",
          4974 => x"0b",
          4975 => x"76",
          4976 => x"81",
          4977 => x"38",
          4978 => x"51",
          4979 => x"82",
          4980 => x"83",
          4981 => x"53",
          4982 => x"09",
          4983 => x"f9",
          4984 => x"52",
          4985 => x"b8",
          4986 => x"ec",
          4987 => x"38",
          4988 => x"08",
          4989 => x"84",
          4990 => x"d8",
          4991 => x"8c",
          4992 => x"ff",
          4993 => x"72",
          4994 => x"2e",
          4995 => x"80",
          4996 => x"14",
          4997 => x"3f",
          4998 => x"08",
          4999 => x"a4",
          5000 => x"81",
          5001 => x"84",
          5002 => x"d7",
          5003 => x"8c",
          5004 => x"8a",
          5005 => x"2e",
          5006 => x"9d",
          5007 => x"14",
          5008 => x"3f",
          5009 => x"08",
          5010 => x"84",
          5011 => x"d7",
          5012 => x"8c",
          5013 => x"15",
          5014 => x"34",
          5015 => x"22",
          5016 => x"72",
          5017 => x"23",
          5018 => x"23",
          5019 => x"15",
          5020 => x"75",
          5021 => x"0c",
          5022 => x"04",
          5023 => x"77",
          5024 => x"73",
          5025 => x"38",
          5026 => x"72",
          5027 => x"38",
          5028 => x"71",
          5029 => x"38",
          5030 => x"84",
          5031 => x"52",
          5032 => x"09",
          5033 => x"38",
          5034 => x"51",
          5035 => x"82",
          5036 => x"81",
          5037 => x"88",
          5038 => x"08",
          5039 => x"39",
          5040 => x"73",
          5041 => x"74",
          5042 => x"0c",
          5043 => x"04",
          5044 => x"02",
          5045 => x"7a",
          5046 => x"fc",
          5047 => x"f4",
          5048 => x"54",
          5049 => x"8c",
          5050 => x"bc",
          5051 => x"ec",
          5052 => x"82",
          5053 => x"70",
          5054 => x"73",
          5055 => x"38",
          5056 => x"78",
          5057 => x"2e",
          5058 => x"74",
          5059 => x"0c",
          5060 => x"80",
          5061 => x"80",
          5062 => x"70",
          5063 => x"51",
          5064 => x"82",
          5065 => x"54",
          5066 => x"ec",
          5067 => x"0d",
          5068 => x"0d",
          5069 => x"05",
          5070 => x"33",
          5071 => x"54",
          5072 => x"84",
          5073 => x"bf",
          5074 => x"98",
          5075 => x"53",
          5076 => x"05",
          5077 => x"fa",
          5078 => x"ec",
          5079 => x"8c",
          5080 => x"a4",
          5081 => x"68",
          5082 => x"70",
          5083 => x"c6",
          5084 => x"ec",
          5085 => x"8c",
          5086 => x"38",
          5087 => x"05",
          5088 => x"2b",
          5089 => x"80",
          5090 => x"86",
          5091 => x"06",
          5092 => x"2e",
          5093 => x"74",
          5094 => x"38",
          5095 => x"09",
          5096 => x"38",
          5097 => x"f8",
          5098 => x"ec",
          5099 => x"39",
          5100 => x"33",
          5101 => x"73",
          5102 => x"77",
          5103 => x"81",
          5104 => x"73",
          5105 => x"38",
          5106 => x"bc",
          5107 => x"07",
          5108 => x"b4",
          5109 => x"2a",
          5110 => x"51",
          5111 => x"2e",
          5112 => x"62",
          5113 => x"e8",
          5114 => x"8c",
          5115 => x"82",
          5116 => x"52",
          5117 => x"51",
          5118 => x"62",
          5119 => x"8b",
          5120 => x"53",
          5121 => x"51",
          5122 => x"80",
          5123 => x"05",
          5124 => x"3f",
          5125 => x"0b",
          5126 => x"75",
          5127 => x"f1",
          5128 => x"11",
          5129 => x"80",
          5130 => x"97",
          5131 => x"51",
          5132 => x"82",
          5133 => x"55",
          5134 => x"08",
          5135 => x"b7",
          5136 => x"c4",
          5137 => x"05",
          5138 => x"2a",
          5139 => x"51",
          5140 => x"80",
          5141 => x"84",
          5142 => x"39",
          5143 => x"70",
          5144 => x"54",
          5145 => x"a9",
          5146 => x"06",
          5147 => x"2e",
          5148 => x"55",
          5149 => x"73",
          5150 => x"d6",
          5151 => x"8c",
          5152 => x"ff",
          5153 => x"0c",
          5154 => x"8c",
          5155 => x"f8",
          5156 => x"2a",
          5157 => x"51",
          5158 => x"2e",
          5159 => x"80",
          5160 => x"7a",
          5161 => x"a0",
          5162 => x"a4",
          5163 => x"53",
          5164 => x"e6",
          5165 => x"8c",
          5166 => x"8c",
          5167 => x"1b",
          5168 => x"05",
          5169 => x"d3",
          5170 => x"ec",
          5171 => x"ec",
          5172 => x"0c",
          5173 => x"56",
          5174 => x"84",
          5175 => x"90",
          5176 => x"0b",
          5177 => x"80",
          5178 => x"0c",
          5179 => x"1a",
          5180 => x"2a",
          5181 => x"51",
          5182 => x"2e",
          5183 => x"82",
          5184 => x"80",
          5185 => x"38",
          5186 => x"08",
          5187 => x"8a",
          5188 => x"89",
          5189 => x"59",
          5190 => x"76",
          5191 => x"d7",
          5192 => x"8c",
          5193 => x"82",
          5194 => x"81",
          5195 => x"82",
          5196 => x"ec",
          5197 => x"09",
          5198 => x"38",
          5199 => x"78",
          5200 => x"30",
          5201 => x"80",
          5202 => x"77",
          5203 => x"38",
          5204 => x"06",
          5205 => x"c3",
          5206 => x"1a",
          5207 => x"38",
          5208 => x"06",
          5209 => x"2e",
          5210 => x"52",
          5211 => x"a6",
          5212 => x"ec",
          5213 => x"82",
          5214 => x"75",
          5215 => x"8c",
          5216 => x"9c",
          5217 => x"39",
          5218 => x"74",
          5219 => x"8c",
          5220 => x"3d",
          5221 => x"3d",
          5222 => x"65",
          5223 => x"5d",
          5224 => x"0c",
          5225 => x"05",
          5226 => x"f9",
          5227 => x"8c",
          5228 => x"82",
          5229 => x"8a",
          5230 => x"33",
          5231 => x"2e",
          5232 => x"56",
          5233 => x"90",
          5234 => x"06",
          5235 => x"74",
          5236 => x"b6",
          5237 => x"82",
          5238 => x"34",
          5239 => x"aa",
          5240 => x"91",
          5241 => x"56",
          5242 => x"8c",
          5243 => x"1a",
          5244 => x"74",
          5245 => x"38",
          5246 => x"80",
          5247 => x"38",
          5248 => x"70",
          5249 => x"56",
          5250 => x"b2",
          5251 => x"11",
          5252 => x"77",
          5253 => x"5b",
          5254 => x"38",
          5255 => x"88",
          5256 => x"8f",
          5257 => x"08",
          5258 => x"d5",
          5259 => x"8c",
          5260 => x"81",
          5261 => x"9f",
          5262 => x"2e",
          5263 => x"74",
          5264 => x"98",
          5265 => x"7e",
          5266 => x"3f",
          5267 => x"08",
          5268 => x"83",
          5269 => x"ec",
          5270 => x"89",
          5271 => x"77",
          5272 => x"d6",
          5273 => x"7f",
          5274 => x"58",
          5275 => x"75",
          5276 => x"75",
          5277 => x"77",
          5278 => x"7c",
          5279 => x"33",
          5280 => x"3f",
          5281 => x"08",
          5282 => x"7e",
          5283 => x"56",
          5284 => x"2e",
          5285 => x"16",
          5286 => x"55",
          5287 => x"94",
          5288 => x"53",
          5289 => x"b0",
          5290 => x"31",
          5291 => x"05",
          5292 => x"3f",
          5293 => x"56",
          5294 => x"9c",
          5295 => x"19",
          5296 => x"06",
          5297 => x"31",
          5298 => x"76",
          5299 => x"7b",
          5300 => x"08",
          5301 => x"d1",
          5302 => x"8c",
          5303 => x"81",
          5304 => x"94",
          5305 => x"ff",
          5306 => x"05",
          5307 => x"cf",
          5308 => x"76",
          5309 => x"17",
          5310 => x"1e",
          5311 => x"18",
          5312 => x"5e",
          5313 => x"39",
          5314 => x"82",
          5315 => x"90",
          5316 => x"f2",
          5317 => x"63",
          5318 => x"40",
          5319 => x"7e",
          5320 => x"fc",
          5321 => x"51",
          5322 => x"82",
          5323 => x"55",
          5324 => x"08",
          5325 => x"18",
          5326 => x"80",
          5327 => x"74",
          5328 => x"39",
          5329 => x"70",
          5330 => x"81",
          5331 => x"56",
          5332 => x"80",
          5333 => x"38",
          5334 => x"0b",
          5335 => x"82",
          5336 => x"39",
          5337 => x"19",
          5338 => x"83",
          5339 => x"18",
          5340 => x"56",
          5341 => x"27",
          5342 => x"09",
          5343 => x"2e",
          5344 => x"94",
          5345 => x"83",
          5346 => x"56",
          5347 => x"38",
          5348 => x"22",
          5349 => x"89",
          5350 => x"55",
          5351 => x"75",
          5352 => x"18",
          5353 => x"9c",
          5354 => x"85",
          5355 => x"08",
          5356 => x"d7",
          5357 => x"8c",
          5358 => x"82",
          5359 => x"80",
          5360 => x"38",
          5361 => x"ff",
          5362 => x"ff",
          5363 => x"38",
          5364 => x"0c",
          5365 => x"85",
          5366 => x"19",
          5367 => x"b0",
          5368 => x"19",
          5369 => x"81",
          5370 => x"74",
          5371 => x"3f",
          5372 => x"08",
          5373 => x"98",
          5374 => x"7e",
          5375 => x"3f",
          5376 => x"08",
          5377 => x"d2",
          5378 => x"ec",
          5379 => x"89",
          5380 => x"78",
          5381 => x"d5",
          5382 => x"7f",
          5383 => x"58",
          5384 => x"75",
          5385 => x"75",
          5386 => x"78",
          5387 => x"7c",
          5388 => x"33",
          5389 => x"3f",
          5390 => x"08",
          5391 => x"7e",
          5392 => x"78",
          5393 => x"74",
          5394 => x"38",
          5395 => x"b0",
          5396 => x"31",
          5397 => x"05",
          5398 => x"51",
          5399 => x"7e",
          5400 => x"83",
          5401 => x"89",
          5402 => x"db",
          5403 => x"08",
          5404 => x"26",
          5405 => x"51",
          5406 => x"82",
          5407 => x"fd",
          5408 => x"77",
          5409 => x"55",
          5410 => x"0c",
          5411 => x"83",
          5412 => x"80",
          5413 => x"55",
          5414 => x"83",
          5415 => x"9c",
          5416 => x"7e",
          5417 => x"3f",
          5418 => x"08",
          5419 => x"75",
          5420 => x"94",
          5421 => x"ff",
          5422 => x"05",
          5423 => x"3f",
          5424 => x"0b",
          5425 => x"7b",
          5426 => x"08",
          5427 => x"76",
          5428 => x"08",
          5429 => x"1c",
          5430 => x"08",
          5431 => x"5c",
          5432 => x"83",
          5433 => x"74",
          5434 => x"fd",
          5435 => x"18",
          5436 => x"07",
          5437 => x"19",
          5438 => x"75",
          5439 => x"0c",
          5440 => x"04",
          5441 => x"7a",
          5442 => x"05",
          5443 => x"56",
          5444 => x"82",
          5445 => x"57",
          5446 => x"08",
          5447 => x"90",
          5448 => x"86",
          5449 => x"06",
          5450 => x"73",
          5451 => x"e9",
          5452 => x"08",
          5453 => x"cc",
          5454 => x"8c",
          5455 => x"82",
          5456 => x"80",
          5457 => x"16",
          5458 => x"33",
          5459 => x"55",
          5460 => x"34",
          5461 => x"53",
          5462 => x"08",
          5463 => x"3f",
          5464 => x"52",
          5465 => x"c9",
          5466 => x"88",
          5467 => x"96",
          5468 => x"f0",
          5469 => x"92",
          5470 => x"ca",
          5471 => x"81",
          5472 => x"34",
          5473 => x"df",
          5474 => x"ec",
          5475 => x"33",
          5476 => x"55",
          5477 => x"17",
          5478 => x"8c",
          5479 => x"3d",
          5480 => x"3d",
          5481 => x"52",
          5482 => x"3f",
          5483 => x"08",
          5484 => x"ec",
          5485 => x"86",
          5486 => x"52",
          5487 => x"bc",
          5488 => x"ec",
          5489 => x"8c",
          5490 => x"38",
          5491 => x"08",
          5492 => x"82",
          5493 => x"86",
          5494 => x"ff",
          5495 => x"3d",
          5496 => x"3f",
          5497 => x"0b",
          5498 => x"08",
          5499 => x"82",
          5500 => x"82",
          5501 => x"80",
          5502 => x"8c",
          5503 => x"3d",
          5504 => x"3d",
          5505 => x"93",
          5506 => x"52",
          5507 => x"e9",
          5508 => x"8c",
          5509 => x"82",
          5510 => x"80",
          5511 => x"58",
          5512 => x"3d",
          5513 => x"e0",
          5514 => x"8c",
          5515 => x"82",
          5516 => x"bc",
          5517 => x"c7",
          5518 => x"98",
          5519 => x"73",
          5520 => x"38",
          5521 => x"12",
          5522 => x"39",
          5523 => x"33",
          5524 => x"70",
          5525 => x"55",
          5526 => x"2e",
          5527 => x"7f",
          5528 => x"54",
          5529 => x"82",
          5530 => x"94",
          5531 => x"39",
          5532 => x"08",
          5533 => x"81",
          5534 => x"85",
          5535 => x"8c",
          5536 => x"3d",
          5537 => x"3d",
          5538 => x"5b",
          5539 => x"34",
          5540 => x"3d",
          5541 => x"52",
          5542 => x"e8",
          5543 => x"8c",
          5544 => x"82",
          5545 => x"82",
          5546 => x"43",
          5547 => x"11",
          5548 => x"58",
          5549 => x"80",
          5550 => x"38",
          5551 => x"3d",
          5552 => x"d5",
          5553 => x"8c",
          5554 => x"82",
          5555 => x"82",
          5556 => x"52",
          5557 => x"c8",
          5558 => x"ec",
          5559 => x"8c",
          5560 => x"c1",
          5561 => x"7b",
          5562 => x"3f",
          5563 => x"08",
          5564 => x"74",
          5565 => x"3f",
          5566 => x"08",
          5567 => x"ec",
          5568 => x"38",
          5569 => x"51",
          5570 => x"82",
          5571 => x"57",
          5572 => x"08",
          5573 => x"52",
          5574 => x"f2",
          5575 => x"8c",
          5576 => x"a6",
          5577 => x"74",
          5578 => x"3f",
          5579 => x"08",
          5580 => x"ec",
          5581 => x"cc",
          5582 => x"2e",
          5583 => x"86",
          5584 => x"81",
          5585 => x"81",
          5586 => x"3d",
          5587 => x"52",
          5588 => x"c9",
          5589 => x"3d",
          5590 => x"11",
          5591 => x"5a",
          5592 => x"2e",
          5593 => x"b9",
          5594 => x"16",
          5595 => x"33",
          5596 => x"73",
          5597 => x"16",
          5598 => x"26",
          5599 => x"75",
          5600 => x"38",
          5601 => x"05",
          5602 => x"6f",
          5603 => x"ff",
          5604 => x"55",
          5605 => x"74",
          5606 => x"38",
          5607 => x"11",
          5608 => x"74",
          5609 => x"39",
          5610 => x"09",
          5611 => x"38",
          5612 => x"11",
          5613 => x"74",
          5614 => x"82",
          5615 => x"70",
          5616 => x"fc",
          5617 => x"08",
          5618 => x"5c",
          5619 => x"73",
          5620 => x"38",
          5621 => x"1a",
          5622 => x"55",
          5623 => x"38",
          5624 => x"73",
          5625 => x"38",
          5626 => x"76",
          5627 => x"74",
          5628 => x"33",
          5629 => x"05",
          5630 => x"15",
          5631 => x"ba",
          5632 => x"05",
          5633 => x"ff",
          5634 => x"06",
          5635 => x"57",
          5636 => x"18",
          5637 => x"54",
          5638 => x"70",
          5639 => x"34",
          5640 => x"ee",
          5641 => x"34",
          5642 => x"ec",
          5643 => x"0d",
          5644 => x"0d",
          5645 => x"3d",
          5646 => x"71",
          5647 => x"ec",
          5648 => x"8c",
          5649 => x"82",
          5650 => x"82",
          5651 => x"15",
          5652 => x"82",
          5653 => x"15",
          5654 => x"76",
          5655 => x"90",
          5656 => x"81",
          5657 => x"06",
          5658 => x"72",
          5659 => x"56",
          5660 => x"54",
          5661 => x"17",
          5662 => x"78",
          5663 => x"38",
          5664 => x"22",
          5665 => x"59",
          5666 => x"78",
          5667 => x"76",
          5668 => x"51",
          5669 => x"3f",
          5670 => x"08",
          5671 => x"54",
          5672 => x"53",
          5673 => x"3f",
          5674 => x"08",
          5675 => x"38",
          5676 => x"75",
          5677 => x"18",
          5678 => x"31",
          5679 => x"57",
          5680 => x"b1",
          5681 => x"08",
          5682 => x"38",
          5683 => x"51",
          5684 => x"82",
          5685 => x"54",
          5686 => x"08",
          5687 => x"9a",
          5688 => x"ec",
          5689 => x"81",
          5690 => x"8c",
          5691 => x"16",
          5692 => x"16",
          5693 => x"2e",
          5694 => x"76",
          5695 => x"dc",
          5696 => x"31",
          5697 => x"18",
          5698 => x"90",
          5699 => x"81",
          5700 => x"06",
          5701 => x"56",
          5702 => x"9a",
          5703 => x"74",
          5704 => x"3f",
          5705 => x"08",
          5706 => x"ec",
          5707 => x"82",
          5708 => x"56",
          5709 => x"52",
          5710 => x"84",
          5711 => x"ec",
          5712 => x"ff",
          5713 => x"81",
          5714 => x"38",
          5715 => x"98",
          5716 => x"a6",
          5717 => x"16",
          5718 => x"39",
          5719 => x"16",
          5720 => x"75",
          5721 => x"53",
          5722 => x"aa",
          5723 => x"79",
          5724 => x"3f",
          5725 => x"08",
          5726 => x"0b",
          5727 => x"82",
          5728 => x"39",
          5729 => x"16",
          5730 => x"bb",
          5731 => x"2a",
          5732 => x"08",
          5733 => x"15",
          5734 => x"15",
          5735 => x"90",
          5736 => x"16",
          5737 => x"33",
          5738 => x"53",
          5739 => x"34",
          5740 => x"06",
          5741 => x"2e",
          5742 => x"9c",
          5743 => x"85",
          5744 => x"16",
          5745 => x"72",
          5746 => x"0c",
          5747 => x"04",
          5748 => x"79",
          5749 => x"75",
          5750 => x"8a",
          5751 => x"89",
          5752 => x"52",
          5753 => x"05",
          5754 => x"3f",
          5755 => x"08",
          5756 => x"ec",
          5757 => x"38",
          5758 => x"7a",
          5759 => x"d8",
          5760 => x"8c",
          5761 => x"82",
          5762 => x"80",
          5763 => x"16",
          5764 => x"2b",
          5765 => x"74",
          5766 => x"86",
          5767 => x"84",
          5768 => x"06",
          5769 => x"73",
          5770 => x"38",
          5771 => x"52",
          5772 => x"da",
          5773 => x"ec",
          5774 => x"0c",
          5775 => x"14",
          5776 => x"23",
          5777 => x"51",
          5778 => x"82",
          5779 => x"55",
          5780 => x"09",
          5781 => x"38",
          5782 => x"39",
          5783 => x"84",
          5784 => x"0c",
          5785 => x"82",
          5786 => x"89",
          5787 => x"fc",
          5788 => x"87",
          5789 => x"53",
          5790 => x"e7",
          5791 => x"8c",
          5792 => x"38",
          5793 => x"08",
          5794 => x"3d",
          5795 => x"3d",
          5796 => x"89",
          5797 => x"54",
          5798 => x"54",
          5799 => x"82",
          5800 => x"53",
          5801 => x"08",
          5802 => x"74",
          5803 => x"8c",
          5804 => x"73",
          5805 => x"3f",
          5806 => x"08",
          5807 => x"39",
          5808 => x"08",
          5809 => x"d3",
          5810 => x"8c",
          5811 => x"82",
          5812 => x"84",
          5813 => x"06",
          5814 => x"53",
          5815 => x"8c",
          5816 => x"38",
          5817 => x"51",
          5818 => x"72",
          5819 => x"cf",
          5820 => x"8c",
          5821 => x"32",
          5822 => x"72",
          5823 => x"70",
          5824 => x"08",
          5825 => x"54",
          5826 => x"8c",
          5827 => x"3d",
          5828 => x"3d",
          5829 => x"80",
          5830 => x"70",
          5831 => x"52",
          5832 => x"3f",
          5833 => x"08",
          5834 => x"ec",
          5835 => x"64",
          5836 => x"d6",
          5837 => x"8c",
          5838 => x"82",
          5839 => x"a0",
          5840 => x"cb",
          5841 => x"98",
          5842 => x"73",
          5843 => x"38",
          5844 => x"39",
          5845 => x"88",
          5846 => x"75",
          5847 => x"3f",
          5848 => x"ec",
          5849 => x"0d",
          5850 => x"0d",
          5851 => x"5c",
          5852 => x"3d",
          5853 => x"93",
          5854 => x"d6",
          5855 => x"ec",
          5856 => x"8c",
          5857 => x"80",
          5858 => x"0c",
          5859 => x"11",
          5860 => x"90",
          5861 => x"56",
          5862 => x"74",
          5863 => x"75",
          5864 => x"e4",
          5865 => x"81",
          5866 => x"5b",
          5867 => x"82",
          5868 => x"75",
          5869 => x"73",
          5870 => x"81",
          5871 => x"82",
          5872 => x"76",
          5873 => x"f0",
          5874 => x"f4",
          5875 => x"ec",
          5876 => x"d1",
          5877 => x"ec",
          5878 => x"ce",
          5879 => x"ec",
          5880 => x"82",
          5881 => x"07",
          5882 => x"05",
          5883 => x"53",
          5884 => x"98",
          5885 => x"26",
          5886 => x"f9",
          5887 => x"08",
          5888 => x"08",
          5889 => x"98",
          5890 => x"81",
          5891 => x"58",
          5892 => x"3f",
          5893 => x"08",
          5894 => x"ec",
          5895 => x"38",
          5896 => x"77",
          5897 => x"5d",
          5898 => x"74",
          5899 => x"81",
          5900 => x"b4",
          5901 => x"bb",
          5902 => x"8c",
          5903 => x"ff",
          5904 => x"30",
          5905 => x"1b",
          5906 => x"5b",
          5907 => x"39",
          5908 => x"ff",
          5909 => x"82",
          5910 => x"f0",
          5911 => x"30",
          5912 => x"1b",
          5913 => x"5b",
          5914 => x"83",
          5915 => x"58",
          5916 => x"92",
          5917 => x"0c",
          5918 => x"12",
          5919 => x"33",
          5920 => x"54",
          5921 => x"34",
          5922 => x"ec",
          5923 => x"0d",
          5924 => x"0d",
          5925 => x"fc",
          5926 => x"52",
          5927 => x"3f",
          5928 => x"08",
          5929 => x"ec",
          5930 => x"38",
          5931 => x"56",
          5932 => x"38",
          5933 => x"70",
          5934 => x"81",
          5935 => x"55",
          5936 => x"80",
          5937 => x"38",
          5938 => x"54",
          5939 => x"08",
          5940 => x"38",
          5941 => x"82",
          5942 => x"53",
          5943 => x"52",
          5944 => x"8c",
          5945 => x"ec",
          5946 => x"19",
          5947 => x"c9",
          5948 => x"08",
          5949 => x"ff",
          5950 => x"82",
          5951 => x"ff",
          5952 => x"06",
          5953 => x"56",
          5954 => x"08",
          5955 => x"81",
          5956 => x"82",
          5957 => x"75",
          5958 => x"54",
          5959 => x"08",
          5960 => x"27",
          5961 => x"17",
          5962 => x"8c",
          5963 => x"76",
          5964 => x"3f",
          5965 => x"08",
          5966 => x"08",
          5967 => x"90",
          5968 => x"c0",
          5969 => x"90",
          5970 => x"80",
          5971 => x"75",
          5972 => x"75",
          5973 => x"8c",
          5974 => x"3d",
          5975 => x"3d",
          5976 => x"a0",
          5977 => x"05",
          5978 => x"51",
          5979 => x"82",
          5980 => x"55",
          5981 => x"08",
          5982 => x"78",
          5983 => x"08",
          5984 => x"70",
          5985 => x"ae",
          5986 => x"ec",
          5987 => x"8c",
          5988 => x"db",
          5989 => x"fb",
          5990 => x"85",
          5991 => x"06",
          5992 => x"86",
          5993 => x"c7",
          5994 => x"2b",
          5995 => x"24",
          5996 => x"02",
          5997 => x"33",
          5998 => x"58",
          5999 => x"76",
          6000 => x"6b",
          6001 => x"cc",
          6002 => x"8c",
          6003 => x"84",
          6004 => x"06",
          6005 => x"73",
          6006 => x"d4",
          6007 => x"82",
          6008 => x"94",
          6009 => x"81",
          6010 => x"5a",
          6011 => x"08",
          6012 => x"8a",
          6013 => x"54",
          6014 => x"82",
          6015 => x"55",
          6016 => x"08",
          6017 => x"82",
          6018 => x"52",
          6019 => x"e5",
          6020 => x"ec",
          6021 => x"8c",
          6022 => x"38",
          6023 => x"cf",
          6024 => x"ec",
          6025 => x"88",
          6026 => x"ec",
          6027 => x"38",
          6028 => x"c2",
          6029 => x"ec",
          6030 => x"ec",
          6031 => x"82",
          6032 => x"07",
          6033 => x"55",
          6034 => x"2e",
          6035 => x"80",
          6036 => x"80",
          6037 => x"77",
          6038 => x"3f",
          6039 => x"08",
          6040 => x"38",
          6041 => x"ba",
          6042 => x"8c",
          6043 => x"74",
          6044 => x"0c",
          6045 => x"04",
          6046 => x"82",
          6047 => x"c0",
          6048 => x"3d",
          6049 => x"3f",
          6050 => x"08",
          6051 => x"ec",
          6052 => x"38",
          6053 => x"52",
          6054 => x"52",
          6055 => x"3f",
          6056 => x"08",
          6057 => x"ec",
          6058 => x"88",
          6059 => x"39",
          6060 => x"08",
          6061 => x"81",
          6062 => x"38",
          6063 => x"05",
          6064 => x"2a",
          6065 => x"55",
          6066 => x"81",
          6067 => x"5a",
          6068 => x"3d",
          6069 => x"c1",
          6070 => x"8c",
          6071 => x"55",
          6072 => x"ec",
          6073 => x"87",
          6074 => x"ec",
          6075 => x"09",
          6076 => x"38",
          6077 => x"8c",
          6078 => x"2e",
          6079 => x"86",
          6080 => x"81",
          6081 => x"81",
          6082 => x"8c",
          6083 => x"78",
          6084 => x"3f",
          6085 => x"08",
          6086 => x"ec",
          6087 => x"38",
          6088 => x"52",
          6089 => x"ff",
          6090 => x"78",
          6091 => x"b4",
          6092 => x"54",
          6093 => x"15",
          6094 => x"b2",
          6095 => x"ca",
          6096 => x"b6",
          6097 => x"53",
          6098 => x"53",
          6099 => x"3f",
          6100 => x"b4",
          6101 => x"d4",
          6102 => x"b6",
          6103 => x"54",
          6104 => x"d5",
          6105 => x"53",
          6106 => x"11",
          6107 => x"d7",
          6108 => x"81",
          6109 => x"34",
          6110 => x"a4",
          6111 => x"ec",
          6112 => x"8c",
          6113 => x"38",
          6114 => x"0a",
          6115 => x"05",
          6116 => x"d0",
          6117 => x"64",
          6118 => x"c9",
          6119 => x"54",
          6120 => x"15",
          6121 => x"81",
          6122 => x"34",
          6123 => x"b8",
          6124 => x"8c",
          6125 => x"8b",
          6126 => x"75",
          6127 => x"ff",
          6128 => x"73",
          6129 => x"0c",
          6130 => x"04",
          6131 => x"a9",
          6132 => x"51",
          6133 => x"82",
          6134 => x"ff",
          6135 => x"a9",
          6136 => x"ee",
          6137 => x"ec",
          6138 => x"8c",
          6139 => x"d3",
          6140 => x"a9",
          6141 => x"9d",
          6142 => x"58",
          6143 => x"82",
          6144 => x"55",
          6145 => x"08",
          6146 => x"02",
          6147 => x"33",
          6148 => x"54",
          6149 => x"82",
          6150 => x"53",
          6151 => x"52",
          6152 => x"88",
          6153 => x"b4",
          6154 => x"53",
          6155 => x"3d",
          6156 => x"ff",
          6157 => x"aa",
          6158 => x"73",
          6159 => x"3f",
          6160 => x"08",
          6161 => x"ec",
          6162 => x"63",
          6163 => x"81",
          6164 => x"65",
          6165 => x"2e",
          6166 => x"55",
          6167 => x"82",
          6168 => x"84",
          6169 => x"06",
          6170 => x"73",
          6171 => x"3f",
          6172 => x"08",
          6173 => x"ec",
          6174 => x"38",
          6175 => x"53",
          6176 => x"95",
          6177 => x"16",
          6178 => x"87",
          6179 => x"05",
          6180 => x"34",
          6181 => x"70",
          6182 => x"81",
          6183 => x"55",
          6184 => x"74",
          6185 => x"73",
          6186 => x"78",
          6187 => x"83",
          6188 => x"16",
          6189 => x"2a",
          6190 => x"51",
          6191 => x"80",
          6192 => x"38",
          6193 => x"80",
          6194 => x"52",
          6195 => x"be",
          6196 => x"ec",
          6197 => x"51",
          6198 => x"3f",
          6199 => x"8c",
          6200 => x"2e",
          6201 => x"82",
          6202 => x"52",
          6203 => x"b5",
          6204 => x"8c",
          6205 => x"80",
          6206 => x"58",
          6207 => x"ec",
          6208 => x"38",
          6209 => x"54",
          6210 => x"09",
          6211 => x"38",
          6212 => x"52",
          6213 => x"af",
          6214 => x"81",
          6215 => x"34",
          6216 => x"8c",
          6217 => x"38",
          6218 => x"ca",
          6219 => x"ec",
          6220 => x"8c",
          6221 => x"38",
          6222 => x"b5",
          6223 => x"8c",
          6224 => x"74",
          6225 => x"0c",
          6226 => x"04",
          6227 => x"02",
          6228 => x"33",
          6229 => x"80",
          6230 => x"57",
          6231 => x"95",
          6232 => x"52",
          6233 => x"d2",
          6234 => x"8c",
          6235 => x"82",
          6236 => x"80",
          6237 => x"5a",
          6238 => x"3d",
          6239 => x"c9",
          6240 => x"8c",
          6241 => x"82",
          6242 => x"b8",
          6243 => x"cf",
          6244 => x"a0",
          6245 => x"55",
          6246 => x"75",
          6247 => x"71",
          6248 => x"33",
          6249 => x"74",
          6250 => x"57",
          6251 => x"8b",
          6252 => x"54",
          6253 => x"15",
          6254 => x"ff",
          6255 => x"82",
          6256 => x"55",
          6257 => x"ec",
          6258 => x"0d",
          6259 => x"0d",
          6260 => x"53",
          6261 => x"05",
          6262 => x"51",
          6263 => x"82",
          6264 => x"55",
          6265 => x"08",
          6266 => x"76",
          6267 => x"93",
          6268 => x"51",
          6269 => x"82",
          6270 => x"55",
          6271 => x"08",
          6272 => x"80",
          6273 => x"81",
          6274 => x"86",
          6275 => x"38",
          6276 => x"86",
          6277 => x"90",
          6278 => x"54",
          6279 => x"ff",
          6280 => x"76",
          6281 => x"83",
          6282 => x"51",
          6283 => x"3f",
          6284 => x"08",
          6285 => x"8c",
          6286 => x"3d",
          6287 => x"3d",
          6288 => x"5c",
          6289 => x"98",
          6290 => x"52",
          6291 => x"d1",
          6292 => x"8c",
          6293 => x"8c",
          6294 => x"70",
          6295 => x"08",
          6296 => x"51",
          6297 => x"80",
          6298 => x"38",
          6299 => x"06",
          6300 => x"80",
          6301 => x"38",
          6302 => x"5f",
          6303 => x"3d",
          6304 => x"ff",
          6305 => x"82",
          6306 => x"57",
          6307 => x"08",
          6308 => x"74",
          6309 => x"c3",
          6310 => x"8c",
          6311 => x"82",
          6312 => x"bf",
          6313 => x"ec",
          6314 => x"ec",
          6315 => x"59",
          6316 => x"81",
          6317 => x"56",
          6318 => x"33",
          6319 => x"16",
          6320 => x"27",
          6321 => x"56",
          6322 => x"80",
          6323 => x"80",
          6324 => x"ff",
          6325 => x"70",
          6326 => x"56",
          6327 => x"e8",
          6328 => x"76",
          6329 => x"81",
          6330 => x"80",
          6331 => x"57",
          6332 => x"78",
          6333 => x"51",
          6334 => x"2e",
          6335 => x"73",
          6336 => x"38",
          6337 => x"08",
          6338 => x"b1",
          6339 => x"8c",
          6340 => x"82",
          6341 => x"a7",
          6342 => x"33",
          6343 => x"c3",
          6344 => x"2e",
          6345 => x"e4",
          6346 => x"2e",
          6347 => x"56",
          6348 => x"05",
          6349 => x"e3",
          6350 => x"ec",
          6351 => x"76",
          6352 => x"0c",
          6353 => x"04",
          6354 => x"82",
          6355 => x"ff",
          6356 => x"9d",
          6357 => x"fa",
          6358 => x"ec",
          6359 => x"ec",
          6360 => x"82",
          6361 => x"83",
          6362 => x"53",
          6363 => x"3d",
          6364 => x"ff",
          6365 => x"73",
          6366 => x"70",
          6367 => x"52",
          6368 => x"9f",
          6369 => x"bc",
          6370 => x"74",
          6371 => x"6d",
          6372 => x"70",
          6373 => x"af",
          6374 => x"8c",
          6375 => x"2e",
          6376 => x"70",
          6377 => x"57",
          6378 => x"fd",
          6379 => x"ec",
          6380 => x"8d",
          6381 => x"2b",
          6382 => x"81",
          6383 => x"86",
          6384 => x"ec",
          6385 => x"9f",
          6386 => x"ff",
          6387 => x"54",
          6388 => x"8a",
          6389 => x"70",
          6390 => x"06",
          6391 => x"ff",
          6392 => x"38",
          6393 => x"15",
          6394 => x"80",
          6395 => x"74",
          6396 => x"bc",
          6397 => x"89",
          6398 => x"ec",
          6399 => x"81",
          6400 => x"88",
          6401 => x"26",
          6402 => x"39",
          6403 => x"86",
          6404 => x"81",
          6405 => x"ff",
          6406 => x"38",
          6407 => x"54",
          6408 => x"81",
          6409 => x"81",
          6410 => x"78",
          6411 => x"5a",
          6412 => x"6d",
          6413 => x"81",
          6414 => x"57",
          6415 => x"9f",
          6416 => x"38",
          6417 => x"54",
          6418 => x"81",
          6419 => x"b1",
          6420 => x"2e",
          6421 => x"a7",
          6422 => x"15",
          6423 => x"54",
          6424 => x"09",
          6425 => x"38",
          6426 => x"76",
          6427 => x"41",
          6428 => x"52",
          6429 => x"52",
          6430 => x"b3",
          6431 => x"ec",
          6432 => x"8c",
          6433 => x"f7",
          6434 => x"74",
          6435 => x"e5",
          6436 => x"ec",
          6437 => x"8c",
          6438 => x"38",
          6439 => x"38",
          6440 => x"74",
          6441 => x"39",
          6442 => x"08",
          6443 => x"81",
          6444 => x"38",
          6445 => x"74",
          6446 => x"38",
          6447 => x"51",
          6448 => x"3f",
          6449 => x"08",
          6450 => x"ec",
          6451 => x"a0",
          6452 => x"ec",
          6453 => x"51",
          6454 => x"3f",
          6455 => x"0b",
          6456 => x"8b",
          6457 => x"67",
          6458 => x"a7",
          6459 => x"81",
          6460 => x"34",
          6461 => x"ad",
          6462 => x"8c",
          6463 => x"73",
          6464 => x"8c",
          6465 => x"3d",
          6466 => x"3d",
          6467 => x"02",
          6468 => x"cb",
          6469 => x"3d",
          6470 => x"72",
          6471 => x"5a",
          6472 => x"82",
          6473 => x"58",
          6474 => x"08",
          6475 => x"91",
          6476 => x"77",
          6477 => x"7c",
          6478 => x"38",
          6479 => x"59",
          6480 => x"90",
          6481 => x"81",
          6482 => x"06",
          6483 => x"73",
          6484 => x"54",
          6485 => x"82",
          6486 => x"39",
          6487 => x"8b",
          6488 => x"11",
          6489 => x"2b",
          6490 => x"54",
          6491 => x"fe",
          6492 => x"ff",
          6493 => x"70",
          6494 => x"07",
          6495 => x"8c",
          6496 => x"8c",
          6497 => x"40",
          6498 => x"55",
          6499 => x"88",
          6500 => x"08",
          6501 => x"38",
          6502 => x"77",
          6503 => x"56",
          6504 => x"51",
          6505 => x"3f",
          6506 => x"55",
          6507 => x"08",
          6508 => x"38",
          6509 => x"8c",
          6510 => x"2e",
          6511 => x"82",
          6512 => x"ff",
          6513 => x"38",
          6514 => x"08",
          6515 => x"16",
          6516 => x"2e",
          6517 => x"87",
          6518 => x"74",
          6519 => x"74",
          6520 => x"81",
          6521 => x"38",
          6522 => x"ff",
          6523 => x"2e",
          6524 => x"7b",
          6525 => x"80",
          6526 => x"81",
          6527 => x"81",
          6528 => x"06",
          6529 => x"56",
          6530 => x"52",
          6531 => x"af",
          6532 => x"8c",
          6533 => x"82",
          6534 => x"80",
          6535 => x"81",
          6536 => x"56",
          6537 => x"d3",
          6538 => x"ff",
          6539 => x"7c",
          6540 => x"55",
          6541 => x"b3",
          6542 => x"1b",
          6543 => x"1b",
          6544 => x"33",
          6545 => x"54",
          6546 => x"34",
          6547 => x"fe",
          6548 => x"08",
          6549 => x"74",
          6550 => x"75",
          6551 => x"16",
          6552 => x"33",
          6553 => x"73",
          6554 => x"77",
          6555 => x"8c",
          6556 => x"3d",
          6557 => x"3d",
          6558 => x"02",
          6559 => x"eb",
          6560 => x"3d",
          6561 => x"59",
          6562 => x"8b",
          6563 => x"82",
          6564 => x"24",
          6565 => x"82",
          6566 => x"84",
          6567 => x"88",
          6568 => x"51",
          6569 => x"2e",
          6570 => x"75",
          6571 => x"ec",
          6572 => x"06",
          6573 => x"7e",
          6574 => x"d0",
          6575 => x"ec",
          6576 => x"06",
          6577 => x"56",
          6578 => x"74",
          6579 => x"76",
          6580 => x"81",
          6581 => x"8a",
          6582 => x"b2",
          6583 => x"fc",
          6584 => x"52",
          6585 => x"a4",
          6586 => x"8c",
          6587 => x"38",
          6588 => x"80",
          6589 => x"74",
          6590 => x"26",
          6591 => x"15",
          6592 => x"74",
          6593 => x"38",
          6594 => x"80",
          6595 => x"84",
          6596 => x"92",
          6597 => x"80",
          6598 => x"38",
          6599 => x"06",
          6600 => x"2e",
          6601 => x"56",
          6602 => x"78",
          6603 => x"89",
          6604 => x"2b",
          6605 => x"43",
          6606 => x"38",
          6607 => x"30",
          6608 => x"77",
          6609 => x"91",
          6610 => x"c2",
          6611 => x"f8",
          6612 => x"52",
          6613 => x"a4",
          6614 => x"56",
          6615 => x"08",
          6616 => x"77",
          6617 => x"77",
          6618 => x"ec",
          6619 => x"45",
          6620 => x"bf",
          6621 => x"8e",
          6622 => x"26",
          6623 => x"74",
          6624 => x"48",
          6625 => x"75",
          6626 => x"38",
          6627 => x"81",
          6628 => x"fa",
          6629 => x"2a",
          6630 => x"56",
          6631 => x"2e",
          6632 => x"87",
          6633 => x"82",
          6634 => x"38",
          6635 => x"55",
          6636 => x"83",
          6637 => x"81",
          6638 => x"56",
          6639 => x"80",
          6640 => x"38",
          6641 => x"83",
          6642 => x"06",
          6643 => x"78",
          6644 => x"91",
          6645 => x"0b",
          6646 => x"22",
          6647 => x"80",
          6648 => x"74",
          6649 => x"38",
          6650 => x"56",
          6651 => x"17",
          6652 => x"57",
          6653 => x"2e",
          6654 => x"75",
          6655 => x"79",
          6656 => x"fe",
          6657 => x"82",
          6658 => x"84",
          6659 => x"05",
          6660 => x"5e",
          6661 => x"80",
          6662 => x"ec",
          6663 => x"8a",
          6664 => x"fd",
          6665 => x"75",
          6666 => x"38",
          6667 => x"78",
          6668 => x"8c",
          6669 => x"0b",
          6670 => x"22",
          6671 => x"80",
          6672 => x"74",
          6673 => x"38",
          6674 => x"56",
          6675 => x"17",
          6676 => x"57",
          6677 => x"2e",
          6678 => x"75",
          6679 => x"79",
          6680 => x"fe",
          6681 => x"82",
          6682 => x"10",
          6683 => x"82",
          6684 => x"9f",
          6685 => x"38",
          6686 => x"8c",
          6687 => x"82",
          6688 => x"05",
          6689 => x"2a",
          6690 => x"56",
          6691 => x"17",
          6692 => x"81",
          6693 => x"60",
          6694 => x"65",
          6695 => x"12",
          6696 => x"30",
          6697 => x"74",
          6698 => x"59",
          6699 => x"7d",
          6700 => x"81",
          6701 => x"76",
          6702 => x"41",
          6703 => x"76",
          6704 => x"90",
          6705 => x"62",
          6706 => x"51",
          6707 => x"26",
          6708 => x"75",
          6709 => x"31",
          6710 => x"65",
          6711 => x"fe",
          6712 => x"82",
          6713 => x"58",
          6714 => x"09",
          6715 => x"38",
          6716 => x"08",
          6717 => x"26",
          6718 => x"78",
          6719 => x"79",
          6720 => x"78",
          6721 => x"86",
          6722 => x"82",
          6723 => x"06",
          6724 => x"83",
          6725 => x"82",
          6726 => x"27",
          6727 => x"8f",
          6728 => x"55",
          6729 => x"26",
          6730 => x"59",
          6731 => x"62",
          6732 => x"74",
          6733 => x"38",
          6734 => x"88",
          6735 => x"ec",
          6736 => x"26",
          6737 => x"86",
          6738 => x"1a",
          6739 => x"79",
          6740 => x"38",
          6741 => x"80",
          6742 => x"2e",
          6743 => x"83",
          6744 => x"9f",
          6745 => x"8b",
          6746 => x"06",
          6747 => x"74",
          6748 => x"84",
          6749 => x"52",
          6750 => x"a2",
          6751 => x"53",
          6752 => x"52",
          6753 => x"a2",
          6754 => x"80",
          6755 => x"51",
          6756 => x"3f",
          6757 => x"34",
          6758 => x"ff",
          6759 => x"1b",
          6760 => x"a2",
          6761 => x"90",
          6762 => x"83",
          6763 => x"70",
          6764 => x"80",
          6765 => x"55",
          6766 => x"ff",
          6767 => x"66",
          6768 => x"ff",
          6769 => x"38",
          6770 => x"ff",
          6771 => x"1b",
          6772 => x"f2",
          6773 => x"74",
          6774 => x"51",
          6775 => x"3f",
          6776 => x"1c",
          6777 => x"98",
          6778 => x"a0",
          6779 => x"ff",
          6780 => x"51",
          6781 => x"3f",
          6782 => x"1b",
          6783 => x"e4",
          6784 => x"2e",
          6785 => x"80",
          6786 => x"88",
          6787 => x"80",
          6788 => x"ff",
          6789 => x"7c",
          6790 => x"51",
          6791 => x"3f",
          6792 => x"1b",
          6793 => x"bc",
          6794 => x"b0",
          6795 => x"a0",
          6796 => x"52",
          6797 => x"ff",
          6798 => x"ff",
          6799 => x"c0",
          6800 => x"0b",
          6801 => x"34",
          6802 => x"fc",
          6803 => x"c7",
          6804 => x"39",
          6805 => x"0a",
          6806 => x"51",
          6807 => x"3f",
          6808 => x"ff",
          6809 => x"1b",
          6810 => x"da",
          6811 => x"0b",
          6812 => x"a9",
          6813 => x"34",
          6814 => x"fc",
          6815 => x"1b",
          6816 => x"8f",
          6817 => x"d5",
          6818 => x"1b",
          6819 => x"ff",
          6820 => x"81",
          6821 => x"7a",
          6822 => x"ff",
          6823 => x"81",
          6824 => x"ec",
          6825 => x"38",
          6826 => x"09",
          6827 => x"ee",
          6828 => x"60",
          6829 => x"7a",
          6830 => x"ff",
          6831 => x"84",
          6832 => x"52",
          6833 => x"9f",
          6834 => x"8b",
          6835 => x"52",
          6836 => x"9f",
          6837 => x"8a",
          6838 => x"52",
          6839 => x"51",
          6840 => x"3f",
          6841 => x"83",
          6842 => x"ff",
          6843 => x"82",
          6844 => x"1b",
          6845 => x"ec",
          6846 => x"d5",
          6847 => x"ff",
          6848 => x"75",
          6849 => x"05",
          6850 => x"7e",
          6851 => x"e5",
          6852 => x"60",
          6853 => x"52",
          6854 => x"9a",
          6855 => x"53",
          6856 => x"51",
          6857 => x"3f",
          6858 => x"58",
          6859 => x"09",
          6860 => x"38",
          6861 => x"51",
          6862 => x"3f",
          6863 => x"1b",
          6864 => x"a0",
          6865 => x"52",
          6866 => x"91",
          6867 => x"ff",
          6868 => x"81",
          6869 => x"f8",
          6870 => x"7a",
          6871 => x"84",
          6872 => x"61",
          6873 => x"26",
          6874 => x"57",
          6875 => x"53",
          6876 => x"51",
          6877 => x"3f",
          6878 => x"08",
          6879 => x"84",
          6880 => x"8c",
          6881 => x"7a",
          6882 => x"aa",
          6883 => x"75",
          6884 => x"56",
          6885 => x"81",
          6886 => x"80",
          6887 => x"38",
          6888 => x"83",
          6889 => x"63",
          6890 => x"74",
          6891 => x"38",
          6892 => x"54",
          6893 => x"52",
          6894 => x"99",
          6895 => x"8c",
          6896 => x"c1",
          6897 => x"75",
          6898 => x"56",
          6899 => x"8c",
          6900 => x"2e",
          6901 => x"56",
          6902 => x"ff",
          6903 => x"84",
          6904 => x"2e",
          6905 => x"56",
          6906 => x"58",
          6907 => x"38",
          6908 => x"77",
          6909 => x"ff",
          6910 => x"82",
          6911 => x"78",
          6912 => x"c2",
          6913 => x"1b",
          6914 => x"34",
          6915 => x"16",
          6916 => x"82",
          6917 => x"83",
          6918 => x"84",
          6919 => x"67",
          6920 => x"fd",
          6921 => x"51",
          6922 => x"3f",
          6923 => x"16",
          6924 => x"ec",
          6925 => x"bf",
          6926 => x"86",
          6927 => x"8c",
          6928 => x"16",
          6929 => x"83",
          6930 => x"ff",
          6931 => x"66",
          6932 => x"1b",
          6933 => x"8c",
          6934 => x"77",
          6935 => x"7e",
          6936 => x"91",
          6937 => x"82",
          6938 => x"a2",
          6939 => x"80",
          6940 => x"ff",
          6941 => x"81",
          6942 => x"ec",
          6943 => x"89",
          6944 => x"8a",
          6945 => x"86",
          6946 => x"ec",
          6947 => x"82",
          6948 => x"99",
          6949 => x"f5",
          6950 => x"60",
          6951 => x"79",
          6952 => x"5a",
          6953 => x"78",
          6954 => x"8d",
          6955 => x"55",
          6956 => x"fc",
          6957 => x"51",
          6958 => x"7a",
          6959 => x"81",
          6960 => x"8c",
          6961 => x"74",
          6962 => x"38",
          6963 => x"81",
          6964 => x"81",
          6965 => x"8a",
          6966 => x"06",
          6967 => x"76",
          6968 => x"76",
          6969 => x"55",
          6970 => x"ec",
          6971 => x"0d",
          6972 => x"0d",
          6973 => x"70",
          6974 => x"74",
          6975 => x"ea",
          6976 => x"74",
          6977 => x"14",
          6978 => x"de",
          6979 => x"55",
          6980 => x"55",
          6981 => x"2e",
          6982 => x"56",
          6983 => x"9f",
          6984 => x"51",
          6985 => x"38",
          6986 => x"09",
          6987 => x"38",
          6988 => x"81",
          6989 => x"72",
          6990 => x"29",
          6991 => x"05",
          6992 => x"70",
          6993 => x"fe",
          6994 => x"82",
          6995 => x"8b",
          6996 => x"33",
          6997 => x"2e",
          6998 => x"81",
          6999 => x"ff",
          7000 => x"96",
          7001 => x"38",
          7002 => x"82",
          7003 => x"88",
          7004 => x"ff",
          7005 => x"52",
          7006 => x"81",
          7007 => x"84",
          7008 => x"9c",
          7009 => x"08",
          7010 => x"88",
          7011 => x"39",
          7012 => x"51",
          7013 => x"81",
          7014 => x"80",
          7015 => x"ff",
          7016 => x"eb",
          7017 => x"cc",
          7018 => x"39",
          7019 => x"51",
          7020 => x"81",
          7021 => x"80",
          7022 => x"80",
          7023 => x"cf",
          7024 => x"98",
          7025 => x"39",
          7026 => x"51",
          7027 => x"82",
          7028 => x"bb",
          7029 => x"e4",
          7030 => x"82",
          7031 => x"af",
          7032 => x"a4",
          7033 => x"82",
          7034 => x"a3",
          7035 => x"d8",
          7036 => x"82",
          7037 => x"97",
          7038 => x"84",
          7039 => x"82",
          7040 => x"8b",
          7041 => x"b4",
          7042 => x"82",
          7043 => x"ff",
          7044 => x"83",
          7045 => x"fb",
          7046 => x"79",
          7047 => x"87",
          7048 => x"38",
          7049 => x"87",
          7050 => x"91",
          7051 => x"52",
          7052 => x"ee",
          7053 => x"8c",
          7054 => x"75",
          7055 => x"f7",
          7056 => x"ec",
          7057 => x"53",
          7058 => x"82",
          7059 => x"8b",
          7060 => x"3d",
          7061 => x"3d",
          7062 => x"84",
          7063 => x"05",
          7064 => x"80",
          7065 => x"70",
          7066 => x"25",
          7067 => x"59",
          7068 => x"87",
          7069 => x"38",
          7070 => x"76",
          7071 => x"ff",
          7072 => x"93",
          7073 => x"ff",
          7074 => x"76",
          7075 => x"70",
          7076 => x"9d",
          7077 => x"ec",
          7078 => x"8c",
          7079 => x"38",
          7080 => x"08",
          7081 => x"88",
          7082 => x"ec",
          7083 => x"3d",
          7084 => x"84",
          7085 => x"52",
          7086 => x"da",
          7087 => x"ec",
          7088 => x"8c",
          7089 => x"38",
          7090 => x"80",
          7091 => x"74",
          7092 => x"59",
          7093 => x"96",
          7094 => x"51",
          7095 => x"76",
          7096 => x"07",
          7097 => x"30",
          7098 => x"72",
          7099 => x"51",
          7100 => x"2e",
          7101 => x"82",
          7102 => x"c0",
          7103 => x"52",
          7104 => x"93",
          7105 => x"75",
          7106 => x"0c",
          7107 => x"04",
          7108 => x"7b",
          7109 => x"b3",
          7110 => x"58",
          7111 => x"53",
          7112 => x"51",
          7113 => x"82",
          7114 => x"a4",
          7115 => x"2e",
          7116 => x"81",
          7117 => x"98",
          7118 => x"7f",
          7119 => x"ec",
          7120 => x"7d",
          7121 => x"82",
          7122 => x"57",
          7123 => x"04",
          7124 => x"ec",
          7125 => x"0d",
          7126 => x"0d",
          7127 => x"02",
          7128 => x"cf",
          7129 => x"73",
          7130 => x"5f",
          7131 => x"5e",
          7132 => x"82",
          7133 => x"ff",
          7134 => x"82",
          7135 => x"ff",
          7136 => x"80",
          7137 => x"27",
          7138 => x"7b",
          7139 => x"38",
          7140 => x"a7",
          7141 => x"39",
          7142 => x"72",
          7143 => x"38",
          7144 => x"82",
          7145 => x"ff",
          7146 => x"89",
          7147 => x"94",
          7148 => x"fd",
          7149 => x"55",
          7150 => x"74",
          7151 => x"7a",
          7152 => x"72",
          7153 => x"82",
          7154 => x"88",
          7155 => x"39",
          7156 => x"51",
          7157 => x"3f",
          7158 => x"a1",
          7159 => x"53",
          7160 => x"8e",
          7161 => x"52",
          7162 => x"51",
          7163 => x"3f",
          7164 => x"83",
          7165 => x"82",
          7166 => x"15",
          7167 => x"ff",
          7168 => x"ff",
          7169 => x"83",
          7170 => x"82",
          7171 => x"55",
          7172 => x"bc",
          7173 => x"70",
          7174 => x"80",
          7175 => x"27",
          7176 => x"56",
          7177 => x"74",
          7178 => x"81",
          7179 => x"06",
          7180 => x"06",
          7181 => x"80",
          7182 => x"73",
          7183 => x"85",
          7184 => x"83",
          7185 => x"ff",
          7186 => x"81",
          7187 => x"39",
          7188 => x"51",
          7189 => x"3f",
          7190 => x"1c",
          7191 => x"f6",
          7192 => x"8c",
          7193 => x"2b",
          7194 => x"51",
          7195 => x"2e",
          7196 => x"ab",
          7197 => x"c5",
          7198 => x"ec",
          7199 => x"70",
          7200 => x"a0",
          7201 => x"72",
          7202 => x"30",
          7203 => x"73",
          7204 => x"51",
          7205 => x"57",
          7206 => x"73",
          7207 => x"76",
          7208 => x"81",
          7209 => x"80",
          7210 => x"7c",
          7211 => x"78",
          7212 => x"38",
          7213 => x"82",
          7214 => x"8f",
          7215 => x"fc",
          7216 => x"9b",
          7217 => x"83",
          7218 => x"83",
          7219 => x"ff",
          7220 => x"82",
          7221 => x"51",
          7222 => x"3f",
          7223 => x"54",
          7224 => x"53",
          7225 => x"33",
          7226 => x"d4",
          7227 => x"a5",
          7228 => x"2e",
          7229 => x"fa",
          7230 => x"3d",
          7231 => x"3d",
          7232 => x"96",
          7233 => x"fe",
          7234 => x"81",
          7235 => x"c1",
          7236 => x"f0",
          7237 => x"b9",
          7238 => x"fe",
          7239 => x"72",
          7240 => x"81",
          7241 => x"71",
          7242 => x"38",
          7243 => x"f1",
          7244 => x"84",
          7245 => x"f3",
          7246 => x"51",
          7247 => x"3f",
          7248 => x"70",
          7249 => x"52",
          7250 => x"95",
          7251 => x"fe",
          7252 => x"82",
          7253 => x"fe",
          7254 => x"80",
          7255 => x"f1",
          7256 => x"2a",
          7257 => x"51",
          7258 => x"2e",
          7259 => x"51",
          7260 => x"3f",
          7261 => x"51",
          7262 => x"3f",
          7263 => x"f0",
          7264 => x"84",
          7265 => x"06",
          7266 => x"80",
          7267 => x"81",
          7268 => x"bd",
          7269 => x"c0",
          7270 => x"b5",
          7271 => x"fe",
          7272 => x"72",
          7273 => x"81",
          7274 => x"71",
          7275 => x"38",
          7276 => x"f0",
          7277 => x"84",
          7278 => x"f2",
          7279 => x"51",
          7280 => x"3f",
          7281 => x"70",
          7282 => x"52",
          7283 => x"95",
          7284 => x"fe",
          7285 => x"82",
          7286 => x"fe",
          7287 => x"80",
          7288 => x"ed",
          7289 => x"2a",
          7290 => x"51",
          7291 => x"2e",
          7292 => x"51",
          7293 => x"3f",
          7294 => x"51",
          7295 => x"3f",
          7296 => x"ef",
          7297 => x"88",
          7298 => x"06",
          7299 => x"80",
          7300 => x"81",
          7301 => x"b9",
          7302 => x"90",
          7303 => x"b1",
          7304 => x"fe",
          7305 => x"fe",
          7306 => x"84",
          7307 => x"fb",
          7308 => x"79",
          7309 => x"56",
          7310 => x"51",
          7311 => x"3f",
          7312 => x"33",
          7313 => x"38",
          7314 => x"85",
          7315 => x"a3",
          7316 => x"b9",
          7317 => x"8c",
          7318 => x"70",
          7319 => x"08",
          7320 => x"82",
          7321 => x"51",
          7322 => x"89",
          7323 => x"89",
          7324 => x"73",
          7325 => x"81",
          7326 => x"82",
          7327 => x"74",
          7328 => x"f4",
          7329 => x"8c",
          7330 => x"2e",
          7331 => x"8c",
          7332 => x"fe",
          7333 => x"8e",
          7334 => x"f0",
          7335 => x"3f",
          7336 => x"89",
          7337 => x"89",
          7338 => x"73",
          7339 => x"81",
          7340 => x"74",
          7341 => x"ff",
          7342 => x"80",
          7343 => x"ec",
          7344 => x"0d",
          7345 => x"0d",
          7346 => x"82",
          7347 => x"5f",
          7348 => x"7c",
          7349 => x"b4",
          7350 => x"ec",
          7351 => x"06",
          7352 => x"2e",
          7353 => x"a2",
          7354 => x"e0",
          7355 => x"70",
          7356 => x"82",
          7357 => x"53",
          7358 => x"8e",
          7359 => x"b7",
          7360 => x"8c",
          7361 => x"2e",
          7362 => x"85",
          7363 => x"c1",
          7364 => x"5f",
          7365 => x"9c",
          7366 => x"95",
          7367 => x"70",
          7368 => x"f8",
          7369 => x"fe",
          7370 => x"3d",
          7371 => x"51",
          7372 => x"82",
          7373 => x"90",
          7374 => x"2c",
          7375 => x"80",
          7376 => x"b3",
          7377 => x"c2",
          7378 => x"78",
          7379 => x"d5",
          7380 => x"24",
          7381 => x"80",
          7382 => x"38",
          7383 => x"80",
          7384 => x"e9",
          7385 => x"c0",
          7386 => x"38",
          7387 => x"24",
          7388 => x"78",
          7389 => x"92",
          7390 => x"39",
          7391 => x"2e",
          7392 => x"78",
          7393 => x"92",
          7394 => x"c3",
          7395 => x"38",
          7396 => x"2e",
          7397 => x"8a",
          7398 => x"81",
          7399 => x"99",
          7400 => x"83",
          7401 => x"78",
          7402 => x"89",
          7403 => x"9d",
          7404 => x"85",
          7405 => x"38",
          7406 => x"b4",
          7407 => x"11",
          7408 => x"05",
          7409 => x"c2",
          7410 => x"ec",
          7411 => x"fe",
          7412 => x"3d",
          7413 => x"53",
          7414 => x"51",
          7415 => x"3f",
          7416 => x"08",
          7417 => x"ad",
          7418 => x"fe",
          7419 => x"ff",
          7420 => x"ff",
          7421 => x"82",
          7422 => x"86",
          7423 => x"ec",
          7424 => x"86",
          7425 => x"fa",
          7426 => x"63",
          7427 => x"7b",
          7428 => x"38",
          7429 => x"7a",
          7430 => x"5c",
          7431 => x"26",
          7432 => x"e1",
          7433 => x"ff",
          7434 => x"ff",
          7435 => x"ff",
          7436 => x"82",
          7437 => x"80",
          7438 => x"38",
          7439 => x"fc",
          7440 => x"84",
          7441 => x"81",
          7442 => x"8c",
          7443 => x"2e",
          7444 => x"b4",
          7445 => x"11",
          7446 => x"05",
          7447 => x"aa",
          7448 => x"ec",
          7449 => x"fd",
          7450 => x"86",
          7451 => x"f9",
          7452 => x"5a",
          7453 => x"81",
          7454 => x"59",
          7455 => x"05",
          7456 => x"34",
          7457 => x"42",
          7458 => x"3d",
          7459 => x"53",
          7460 => x"51",
          7461 => x"3f",
          7462 => x"08",
          7463 => x"f5",
          7464 => x"fe",
          7465 => x"ff",
          7466 => x"ff",
          7467 => x"82",
          7468 => x"80",
          7469 => x"38",
          7470 => x"f8",
          7471 => x"84",
          7472 => x"80",
          7473 => x"8c",
          7474 => x"2e",
          7475 => x"82",
          7476 => x"fe",
          7477 => x"63",
          7478 => x"27",
          7479 => x"70",
          7480 => x"5e",
          7481 => x"7c",
          7482 => x"78",
          7483 => x"79",
          7484 => x"52",
          7485 => x"51",
          7486 => x"3f",
          7487 => x"81",
          7488 => x"d5",
          7489 => x"e4",
          7490 => x"39",
          7491 => x"80",
          7492 => x"84",
          7493 => x"ff",
          7494 => x"8c",
          7495 => x"df",
          7496 => x"e0",
          7497 => x"80",
          7498 => x"82",
          7499 => x"44",
          7500 => x"82",
          7501 => x"59",
          7502 => x"88",
          7503 => x"a0",
          7504 => x"39",
          7505 => x"33",
          7506 => x"2e",
          7507 => x"89",
          7508 => x"ab",
          7509 => x"e3",
          7510 => x"80",
          7511 => x"82",
          7512 => x"44",
          7513 => x"89",
          7514 => x"78",
          7515 => x"38",
          7516 => x"08",
          7517 => x"82",
          7518 => x"fc",
          7519 => x"b4",
          7520 => x"11",
          7521 => x"05",
          7522 => x"fe",
          7523 => x"ec",
          7524 => x"38",
          7525 => x"33",
          7526 => x"2e",
          7527 => x"89",
          7528 => x"80",
          7529 => x"89",
          7530 => x"78",
          7531 => x"38",
          7532 => x"08",
          7533 => x"82",
          7534 => x"59",
          7535 => x"88",
          7536 => x"ac",
          7537 => x"39",
          7538 => x"33",
          7539 => x"2e",
          7540 => x"89",
          7541 => x"99",
          7542 => x"de",
          7543 => x"80",
          7544 => x"82",
          7545 => x"43",
          7546 => x"89",
          7547 => x"05",
          7548 => x"fe",
          7549 => x"ff",
          7550 => x"fe",
          7551 => x"82",
          7552 => x"80",
          7553 => x"80",
          7554 => x"7a",
          7555 => x"38",
          7556 => x"90",
          7557 => x"70",
          7558 => x"2a",
          7559 => x"51",
          7560 => x"78",
          7561 => x"38",
          7562 => x"83",
          7563 => x"82",
          7564 => x"fe",
          7565 => x"a0",
          7566 => x"61",
          7567 => x"63",
          7568 => x"3f",
          7569 => x"51",
          7570 => x"3f",
          7571 => x"b4",
          7572 => x"11",
          7573 => x"05",
          7574 => x"ae",
          7575 => x"ec",
          7576 => x"f9",
          7577 => x"3d",
          7578 => x"53",
          7579 => x"51",
          7580 => x"3f",
          7581 => x"08",
          7582 => x"38",
          7583 => x"80",
          7584 => x"79",
          7585 => x"05",
          7586 => x"fe",
          7587 => x"ff",
          7588 => x"fe",
          7589 => x"82",
          7590 => x"e0",
          7591 => x"39",
          7592 => x"54",
          7593 => x"84",
          7594 => x"e9",
          7595 => x"52",
          7596 => x"fb",
          7597 => x"45",
          7598 => x"78",
          7599 => x"d5",
          7600 => x"27",
          7601 => x"3d",
          7602 => x"53",
          7603 => x"51",
          7604 => x"3f",
          7605 => x"08",
          7606 => x"38",
          7607 => x"80",
          7608 => x"79",
          7609 => x"05",
          7610 => x"39",
          7611 => x"51",
          7612 => x"3f",
          7613 => x"b4",
          7614 => x"11",
          7615 => x"05",
          7616 => x"f8",
          7617 => x"ec",
          7618 => x"f8",
          7619 => x"3d",
          7620 => x"53",
          7621 => x"51",
          7622 => x"3f",
          7623 => x"08",
          7624 => x"38",
          7625 => x"be",
          7626 => x"70",
          7627 => x"23",
          7628 => x"3d",
          7629 => x"53",
          7630 => x"51",
          7631 => x"3f",
          7632 => x"08",
          7633 => x"cd",
          7634 => x"22",
          7635 => x"87",
          7636 => x"f9",
          7637 => x"f8",
          7638 => x"fe",
          7639 => x"79",
          7640 => x"59",
          7641 => x"f7",
          7642 => x"9f",
          7643 => x"60",
          7644 => x"d5",
          7645 => x"fe",
          7646 => x"ff",
          7647 => x"fe",
          7648 => x"82",
          7649 => x"80",
          7650 => x"60",
          7651 => x"05",
          7652 => x"82",
          7653 => x"78",
          7654 => x"39",
          7655 => x"51",
          7656 => x"3f",
          7657 => x"b4",
          7658 => x"11",
          7659 => x"05",
          7660 => x"c8",
          7661 => x"ec",
          7662 => x"f6",
          7663 => x"3d",
          7664 => x"53",
          7665 => x"51",
          7666 => x"3f",
          7667 => x"08",
          7668 => x"38",
          7669 => x"0c",
          7670 => x"05",
          7671 => x"fe",
          7672 => x"ff",
          7673 => x"fe",
          7674 => x"82",
          7675 => x"e4",
          7676 => x"39",
          7677 => x"54",
          7678 => x"a4",
          7679 => x"95",
          7680 => x"52",
          7681 => x"f8",
          7682 => x"45",
          7683 => x"78",
          7684 => x"81",
          7685 => x"27",
          7686 => x"3d",
          7687 => x"53",
          7688 => x"51",
          7689 => x"3f",
          7690 => x"08",
          7691 => x"38",
          7692 => x"0c",
          7693 => x"05",
          7694 => x"39",
          7695 => x"51",
          7696 => x"3f",
          7697 => x"b4",
          7698 => x"11",
          7699 => x"05",
          7700 => x"b6",
          7701 => x"ec",
          7702 => x"f5",
          7703 => x"52",
          7704 => x"51",
          7705 => x"3f",
          7706 => x"04",
          7707 => x"80",
          7708 => x"84",
          7709 => x"f9",
          7710 => x"8c",
          7711 => x"2e",
          7712 => x"63",
          7713 => x"cc",
          7714 => x"89",
          7715 => x"78",
          7716 => x"ec",
          7717 => x"f4",
          7718 => x"8c",
          7719 => x"82",
          7720 => x"fe",
          7721 => x"f4",
          7722 => x"88",
          7723 => x"f1",
          7724 => x"d8",
          7725 => x"dd",
          7726 => x"a0",
          7727 => x"f1",
          7728 => x"ff",
          7729 => x"eb",
          7730 => x"c9",
          7731 => x"33",
          7732 => x"80",
          7733 => x"38",
          7734 => x"59",
          7735 => x"81",
          7736 => x"3d",
          7737 => x"51",
          7738 => x"3f",
          7739 => x"08",
          7740 => x"7a",
          7741 => x"38",
          7742 => x"89",
          7743 => x"2e",
          7744 => x"cd",
          7745 => x"2e",
          7746 => x"c5",
          7747 => x"b4",
          7748 => x"82",
          7749 => x"80",
          7750 => x"bc",
          7751 => x"ff",
          7752 => x"fe",
          7753 => x"bb",
          7754 => x"dc",
          7755 => x"ff",
          7756 => x"fe",
          7757 => x"ab",
          7758 => x"82",
          7759 => x"80",
          7760 => x"cc",
          7761 => x"ff",
          7762 => x"fe",
          7763 => x"93",
          7764 => x"80",
          7765 => x"d8",
          7766 => x"ff",
          7767 => x"fe",
          7768 => x"82",
          7769 => x"82",
          7770 => x"80",
          7771 => x"11",
          7772 => x"55",
          7773 => x"80",
          7774 => x"80",
          7775 => x"3d",
          7776 => x"51",
          7777 => x"82",
          7778 => x"82",
          7779 => x"09",
          7780 => x"72",
          7781 => x"51",
          7782 => x"80",
          7783 => x"26",
          7784 => x"5a",
          7785 => x"59",
          7786 => x"8d",
          7787 => x"70",
          7788 => x"5c",
          7789 => x"bb",
          7790 => x"32",
          7791 => x"07",
          7792 => x"38",
          7793 => x"09",
          7794 => x"c9",
          7795 => x"e0",
          7796 => x"c1",
          7797 => x"39",
          7798 => x"80",
          7799 => x"a0",
          7800 => x"94",
          7801 => x"54",
          7802 => x"80",
          7803 => x"fe",
          7804 => x"82",
          7805 => x"90",
          7806 => x"55",
          7807 => x"80",
          7808 => x"fe",
          7809 => x"72",
          7810 => x"08",
          7811 => x"87",
          7812 => x"70",
          7813 => x"87",
          7814 => x"72",
          7815 => x"97",
          7816 => x"ec",
          7817 => x"75",
          7818 => x"87",
          7819 => x"73",
          7820 => x"83",
          7821 => x"8c",
          7822 => x"75",
          7823 => x"83",
          7824 => x"94",
          7825 => x"80",
          7826 => x"c0",
          7827 => x"80",
          7828 => x"82",
          7829 => x"80",
          7830 => x"82",
          7831 => x"fe",
          7832 => x"fe",
          7833 => x"82",
          7834 => x"fe",
          7835 => x"82",
          7836 => x"fe",
          7837 => x"81",
          7838 => x"fe",
          7839 => x"81",
          7840 => x"3f",
          7841 => x"80",
          7842 => x"30",
          7843 => x"30",
          7844 => x"30",
          7845 => x"30",
          7846 => x"30",
          7847 => x"6e",
          7848 => x"6d",
          7849 => x"6d",
          7850 => x"6d",
          7851 => x"6d",
          7852 => x"6d",
          7853 => x"6d",
          7854 => x"6d",
          7855 => x"6d",
          7856 => x"6d",
          7857 => x"6d",
          7858 => x"6d",
          7859 => x"6d",
          7860 => x"6d",
          7861 => x"6d",
          7862 => x"6d",
          7863 => x"6d",
          7864 => x"6d",
          7865 => x"6d",
          7866 => x"6d",
          7867 => x"2f",
          7868 => x"25",
          7869 => x"64",
          7870 => x"3a",
          7871 => x"25",
          7872 => x"0a",
          7873 => x"43",
          7874 => x"6e",
          7875 => x"75",
          7876 => x"69",
          7877 => x"00",
          7878 => x"66",
          7879 => x"20",
          7880 => x"20",
          7881 => x"66",
          7882 => x"00",
          7883 => x"44",
          7884 => x"63",
          7885 => x"69",
          7886 => x"65",
          7887 => x"74",
          7888 => x"0a",
          7889 => x"20",
          7890 => x"20",
          7891 => x"41",
          7892 => x"28",
          7893 => x"58",
          7894 => x"38",
          7895 => x"0a",
          7896 => x"20",
          7897 => x"52",
          7898 => x"20",
          7899 => x"28",
          7900 => x"58",
          7901 => x"38",
          7902 => x"0a",
          7903 => x"20",
          7904 => x"53",
          7905 => x"52",
          7906 => x"28",
          7907 => x"58",
          7908 => x"38",
          7909 => x"0a",
          7910 => x"20",
          7911 => x"41",
          7912 => x"20",
          7913 => x"28",
          7914 => x"58",
          7915 => x"38",
          7916 => x"0a",
          7917 => x"20",
          7918 => x"4d",
          7919 => x"20",
          7920 => x"28",
          7921 => x"58",
          7922 => x"38",
          7923 => x"0a",
          7924 => x"20",
          7925 => x"20",
          7926 => x"44",
          7927 => x"28",
          7928 => x"69",
          7929 => x"20",
          7930 => x"32",
          7931 => x"0a",
          7932 => x"20",
          7933 => x"4d",
          7934 => x"20",
          7935 => x"28",
          7936 => x"65",
          7937 => x"20",
          7938 => x"32",
          7939 => x"0a",
          7940 => x"20",
          7941 => x"54",
          7942 => x"54",
          7943 => x"28",
          7944 => x"6e",
          7945 => x"73",
          7946 => x"32",
          7947 => x"0a",
          7948 => x"20",
          7949 => x"53",
          7950 => x"4e",
          7951 => x"55",
          7952 => x"00",
          7953 => x"20",
          7954 => x"20",
          7955 => x"0a",
          7956 => x"20",
          7957 => x"43",
          7958 => x"00",
          7959 => x"20",
          7960 => x"32",
          7961 => x"00",
          7962 => x"20",
          7963 => x"49",
          7964 => x"00",
          7965 => x"64",
          7966 => x"73",
          7967 => x"0a",
          7968 => x"20",
          7969 => x"55",
          7970 => x"73",
          7971 => x"56",
          7972 => x"6f",
          7973 => x"64",
          7974 => x"73",
          7975 => x"20",
          7976 => x"58",
          7977 => x"00",
          7978 => x"20",
          7979 => x"55",
          7980 => x"6d",
          7981 => x"20",
          7982 => x"72",
          7983 => x"64",
          7984 => x"73",
          7985 => x"20",
          7986 => x"58",
          7987 => x"00",
          7988 => x"20",
          7989 => x"61",
          7990 => x"53",
          7991 => x"74",
          7992 => x"64",
          7993 => x"73",
          7994 => x"20",
          7995 => x"20",
          7996 => x"58",
          7997 => x"00",
          7998 => x"73",
          7999 => x"00",
          8000 => x"20",
          8001 => x"55",
          8002 => x"20",
          8003 => x"20",
          8004 => x"20",
          8005 => x"20",
          8006 => x"20",
          8007 => x"20",
          8008 => x"58",
          8009 => x"00",
          8010 => x"20",
          8011 => x"73",
          8012 => x"20",
          8013 => x"63",
          8014 => x"72",
          8015 => x"20",
          8016 => x"20",
          8017 => x"20",
          8018 => x"25",
          8019 => x"4d",
          8020 => x"00",
          8021 => x"20",
          8022 => x"52",
          8023 => x"43",
          8024 => x"6b",
          8025 => x"65",
          8026 => x"20",
          8027 => x"20",
          8028 => x"20",
          8029 => x"25",
          8030 => x"4d",
          8031 => x"00",
          8032 => x"20",
          8033 => x"73",
          8034 => x"6e",
          8035 => x"44",
          8036 => x"20",
          8037 => x"63",
          8038 => x"72",
          8039 => x"20",
          8040 => x"25",
          8041 => x"4d",
          8042 => x"00",
          8043 => x"61",
          8044 => x"00",
          8045 => x"64",
          8046 => x"00",
          8047 => x"65",
          8048 => x"00",
          8049 => x"4f",
          8050 => x"4f",
          8051 => x"00",
          8052 => x"6b",
          8053 => x"6e",
          8054 => x"00",
          8055 => x"2b",
          8056 => x"3c",
          8057 => x"5b",
          8058 => x"00",
          8059 => x"54",
          8060 => x"54",
          8061 => x"00",
          8062 => x"90",
          8063 => x"4f",
          8064 => x"30",
          8065 => x"20",
          8066 => x"45",
          8067 => x"20",
          8068 => x"33",
          8069 => x"20",
          8070 => x"20",
          8071 => x"45",
          8072 => x"20",
          8073 => x"20",
          8074 => x"20",
          8075 => x"7d",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"45",
          8080 => x"8f",
          8081 => x"45",
          8082 => x"8e",
          8083 => x"92",
          8084 => x"55",
          8085 => x"9a",
          8086 => x"9e",
          8087 => x"4f",
          8088 => x"a6",
          8089 => x"aa",
          8090 => x"ae",
          8091 => x"b2",
          8092 => x"b6",
          8093 => x"ba",
          8094 => x"be",
          8095 => x"c2",
          8096 => x"c6",
          8097 => x"ca",
          8098 => x"ce",
          8099 => x"d2",
          8100 => x"d6",
          8101 => x"da",
          8102 => x"de",
          8103 => x"e2",
          8104 => x"e6",
          8105 => x"ea",
          8106 => x"ee",
          8107 => x"f2",
          8108 => x"f6",
          8109 => x"fa",
          8110 => x"fe",
          8111 => x"2c",
          8112 => x"5d",
          8113 => x"2a",
          8114 => x"3f",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"02",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"6e",
          8125 => x"00",
          8126 => x"6f",
          8127 => x"00",
          8128 => x"6e",
          8129 => x"00",
          8130 => x"6f",
          8131 => x"00",
          8132 => x"78",
          8133 => x"00",
          8134 => x"6c",
          8135 => x"00",
          8136 => x"6f",
          8137 => x"00",
          8138 => x"69",
          8139 => x"00",
          8140 => x"75",
          8141 => x"00",
          8142 => x"62",
          8143 => x"68",
          8144 => x"77",
          8145 => x"64",
          8146 => x"65",
          8147 => x"64",
          8148 => x"65",
          8149 => x"6c",
          8150 => x"00",
          8151 => x"70",
          8152 => x"73",
          8153 => x"74",
          8154 => x"73",
          8155 => x"00",
          8156 => x"66",
          8157 => x"00",
          8158 => x"73",
          8159 => x"00",
          8160 => x"61",
          8161 => x"00",
          8162 => x"73",
          8163 => x"72",
          8164 => x"0a",
          8165 => x"74",
          8166 => x"61",
          8167 => x"72",
          8168 => x"2e",
          8169 => x"00",
          8170 => x"73",
          8171 => x"6f",
          8172 => x"65",
          8173 => x"2e",
          8174 => x"00",
          8175 => x"20",
          8176 => x"65",
          8177 => x"75",
          8178 => x"0a",
          8179 => x"20",
          8180 => x"68",
          8181 => x"75",
          8182 => x"0a",
          8183 => x"76",
          8184 => x"64",
          8185 => x"6c",
          8186 => x"6d",
          8187 => x"00",
          8188 => x"63",
          8189 => x"20",
          8190 => x"69",
          8191 => x"0a",
          8192 => x"6c",
          8193 => x"6c",
          8194 => x"64",
          8195 => x"78",
          8196 => x"73",
          8197 => x"00",
          8198 => x"6c",
          8199 => x"61",
          8200 => x"65",
          8201 => x"76",
          8202 => x"64",
          8203 => x"00",
          8204 => x"20",
          8205 => x"77",
          8206 => x"65",
          8207 => x"6f",
          8208 => x"74",
          8209 => x"0a",
          8210 => x"69",
          8211 => x"6e",
          8212 => x"65",
          8213 => x"73",
          8214 => x"76",
          8215 => x"64",
          8216 => x"00",
          8217 => x"73",
          8218 => x"6f",
          8219 => x"6e",
          8220 => x"65",
          8221 => x"00",
          8222 => x"20",
          8223 => x"70",
          8224 => x"62",
          8225 => x"66",
          8226 => x"73",
          8227 => x"65",
          8228 => x"6f",
          8229 => x"20",
          8230 => x"64",
          8231 => x"2e",
          8232 => x"00",
          8233 => x"72",
          8234 => x"20",
          8235 => x"72",
          8236 => x"2e",
          8237 => x"00",
          8238 => x"6d",
          8239 => x"74",
          8240 => x"70",
          8241 => x"74",
          8242 => x"20",
          8243 => x"63",
          8244 => x"65",
          8245 => x"00",
          8246 => x"6c",
          8247 => x"73",
          8248 => x"63",
          8249 => x"2e",
          8250 => x"00",
          8251 => x"73",
          8252 => x"69",
          8253 => x"6e",
          8254 => x"65",
          8255 => x"79",
          8256 => x"00",
          8257 => x"6f",
          8258 => x"6e",
          8259 => x"70",
          8260 => x"66",
          8261 => x"73",
          8262 => x"00",
          8263 => x"72",
          8264 => x"74",
          8265 => x"20",
          8266 => x"6f",
          8267 => x"63",
          8268 => x"00",
          8269 => x"63",
          8270 => x"73",
          8271 => x"00",
          8272 => x"6b",
          8273 => x"6e",
          8274 => x"72",
          8275 => x"0a",
          8276 => x"6c",
          8277 => x"79",
          8278 => x"20",
          8279 => x"61",
          8280 => x"6c",
          8281 => x"79",
          8282 => x"2f",
          8283 => x"2e",
          8284 => x"00",
          8285 => x"61",
          8286 => x"00",
          8287 => x"38",
          8288 => x"00",
          8289 => x"20",
          8290 => x"34",
          8291 => x"00",
          8292 => x"20",
          8293 => x"20",
          8294 => x"00",
          8295 => x"32",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"0a",
          8300 => x"53",
          8301 => x"2a",
          8302 => x"20",
          8303 => x"00",
          8304 => x"2f",
          8305 => x"32",
          8306 => x"00",
          8307 => x"2e",
          8308 => x"00",
          8309 => x"50",
          8310 => x"72",
          8311 => x"25",
          8312 => x"29",
          8313 => x"20",
          8314 => x"2a",
          8315 => x"00",
          8316 => x"55",
          8317 => x"74",
          8318 => x"75",
          8319 => x"48",
          8320 => x"6c",
          8321 => x"00",
          8322 => x"6d",
          8323 => x"69",
          8324 => x"72",
          8325 => x"74",
          8326 => x"00",
          8327 => x"32",
          8328 => x"74",
          8329 => x"75",
          8330 => x"00",
          8331 => x"43",
          8332 => x"52",
          8333 => x"6e",
          8334 => x"72",
          8335 => x"0a",
          8336 => x"43",
          8337 => x"57",
          8338 => x"6e",
          8339 => x"72",
          8340 => x"0a",
          8341 => x"52",
          8342 => x"52",
          8343 => x"6e",
          8344 => x"72",
          8345 => x"0a",
          8346 => x"52",
          8347 => x"54",
          8348 => x"6e",
          8349 => x"72",
          8350 => x"0a",
          8351 => x"52",
          8352 => x"52",
          8353 => x"6e",
          8354 => x"72",
          8355 => x"0a",
          8356 => x"52",
          8357 => x"54",
          8358 => x"6e",
          8359 => x"72",
          8360 => x"0a",
          8361 => x"74",
          8362 => x"67",
          8363 => x"20",
          8364 => x"65",
          8365 => x"2e",
          8366 => x"00",
          8367 => x"61",
          8368 => x"6e",
          8369 => x"69",
          8370 => x"2e",
          8371 => x"00",
          8372 => x"74",
          8373 => x"65",
          8374 => x"61",
          8375 => x"00",
          8376 => x"00",
          8377 => x"69",
          8378 => x"20",
          8379 => x"69",
          8380 => x"69",
          8381 => x"73",
          8382 => x"64",
          8383 => x"72",
          8384 => x"2c",
          8385 => x"65",
          8386 => x"20",
          8387 => x"74",
          8388 => x"6e",
          8389 => x"6c",
          8390 => x"00",
          8391 => x"00",
          8392 => x"65",
          8393 => x"6e",
          8394 => x"2e",
          8395 => x"00",
          8396 => x"70",
          8397 => x"67",
          8398 => x"00",
          8399 => x"6d",
          8400 => x"69",
          8401 => x"2e",
          8402 => x"00",
          8403 => x"38",
          8404 => x"25",
          8405 => x"29",
          8406 => x"30",
          8407 => x"28",
          8408 => x"78",
          8409 => x"00",
          8410 => x"6d",
          8411 => x"65",
          8412 => x"79",
          8413 => x"00",
          8414 => x"6f",
          8415 => x"65",
          8416 => x"0a",
          8417 => x"38",
          8418 => x"30",
          8419 => x"00",
          8420 => x"3f",
          8421 => x"00",
          8422 => x"38",
          8423 => x"30",
          8424 => x"00",
          8425 => x"38",
          8426 => x"30",
          8427 => x"00",
          8428 => x"65",
          8429 => x"69",
          8430 => x"63",
          8431 => x"20",
          8432 => x"30",
          8433 => x"2e",
          8434 => x"00",
          8435 => x"6c",
          8436 => x"67",
          8437 => x"64",
          8438 => x"20",
          8439 => x"78",
          8440 => x"2e",
          8441 => x"00",
          8442 => x"6c",
          8443 => x"65",
          8444 => x"6e",
          8445 => x"63",
          8446 => x"20",
          8447 => x"29",
          8448 => x"00",
          8449 => x"73",
          8450 => x"74",
          8451 => x"20",
          8452 => x"6c",
          8453 => x"74",
          8454 => x"2e",
          8455 => x"00",
          8456 => x"6c",
          8457 => x"65",
          8458 => x"74",
          8459 => x"2e",
          8460 => x"00",
          8461 => x"55",
          8462 => x"6e",
          8463 => x"3a",
          8464 => x"5c",
          8465 => x"25",
          8466 => x"00",
          8467 => x"3a",
          8468 => x"5c",
          8469 => x"00",
          8470 => x"3a",
          8471 => x"00",
          8472 => x"64",
          8473 => x"6d",
          8474 => x"64",
          8475 => x"00",
          8476 => x"6e",
          8477 => x"67",
          8478 => x"0a",
          8479 => x"61",
          8480 => x"6e",
          8481 => x"6e",
          8482 => x"72",
          8483 => x"73",
          8484 => x"0a",
          8485 => x"00",
          8486 => x"00",
          8487 => x"7f",
          8488 => x"00",
          8489 => x"7f",
          8490 => x"00",
          8491 => x"7f",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"ff",
          8496 => x"00",
          8497 => x"00",
          8498 => x"78",
          8499 => x"00",
          8500 => x"e1",
          8501 => x"e1",
          8502 => x"e1",
          8503 => x"00",
          8504 => x"01",
          8505 => x"01",
          8506 => x"10",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"7e",
          8512 => x"01",
          8513 => x"00",
          8514 => x"00",
          8515 => x"7e",
          8516 => x"01",
          8517 => x"00",
          8518 => x"00",
          8519 => x"7f",
          8520 => x"03",
          8521 => x"00",
          8522 => x"00",
          8523 => x"7f",
          8524 => x"03",
          8525 => x"00",
          8526 => x"00",
          8527 => x"7f",
          8528 => x"03",
          8529 => x"00",
          8530 => x"00",
          8531 => x"7f",
          8532 => x"04",
          8533 => x"00",
          8534 => x"00",
          8535 => x"7f",
          8536 => x"04",
          8537 => x"00",
          8538 => x"00",
          8539 => x"7f",
          8540 => x"04",
          8541 => x"00",
          8542 => x"00",
          8543 => x"7f",
          8544 => x"04",
          8545 => x"00",
          8546 => x"00",
          8547 => x"7f",
          8548 => x"04",
          8549 => x"00",
          8550 => x"00",
          8551 => x"7f",
          8552 => x"04",
          8553 => x"00",
          8554 => x"00",
          8555 => x"7f",
          8556 => x"04",
          8557 => x"00",
          8558 => x"00",
          8559 => x"7f",
          8560 => x"05",
          8561 => x"00",
          8562 => x"00",
          8563 => x"7f",
          8564 => x"05",
          8565 => x"00",
          8566 => x"00",
          8567 => x"7f",
          8568 => x"05",
          8569 => x"00",
          8570 => x"00",
          8571 => x"7f",
          8572 => x"05",
          8573 => x"00",
          8574 => x"00",
          8575 => x"7f",
          8576 => x"07",
          8577 => x"00",
          8578 => x"00",
          8579 => x"7f",
          8580 => x"07",
          8581 => x"00",
          8582 => x"00",
          8583 => x"7f",
          8584 => x"08",
          8585 => x"00",
          8586 => x"00",
          8587 => x"7f",
          8588 => x"08",
          8589 => x"00",
          8590 => x"00",
          8591 => x"7f",
          8592 => x"08",
          8593 => x"00",
          8594 => x"00",
          8595 => x"7f",
          8596 => x"08",
          8597 => x"00",
          8598 => x"00",
          8599 => x"7f",
          8600 => x"09",
          8601 => x"00",
          8602 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"88",
            11 => x"90",
            12 => x"88",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"ac",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"04",
           267 => x"81",
           268 => x"83",
           269 => x"05",
           270 => x"10",
           271 => x"72",
           272 => x"51",
           273 => x"72",
           274 => x"06",
           275 => x"72",
           276 => x"10",
           277 => x"10",
           278 => x"ed",
           279 => x"53",
           280 => x"f4",
           281 => x"27",
           282 => x"71",
           283 => x"53",
           284 => x"0b",
           285 => x"88",
           286 => x"9d",
           287 => x"04",
           288 => x"04",
           289 => x"94",
           290 => x"0c",
           291 => x"80",
           292 => x"8c",
           293 => x"94",
           294 => x"08",
           295 => x"3f",
           296 => x"88",
           297 => x"3d",
           298 => x"04",
           299 => x"94",
           300 => x"0d",
           301 => x"08",
           302 => x"52",
           303 => x"05",
           304 => x"b9",
           305 => x"70",
           306 => x"85",
           307 => x"0c",
           308 => x"02",
           309 => x"3d",
           310 => x"94",
           311 => x"0c",
           312 => x"05",
           313 => x"ab",
           314 => x"88",
           315 => x"94",
           316 => x"0c",
           317 => x"08",
           318 => x"94",
           319 => x"08",
           320 => x"0b",
           321 => x"05",
           322 => x"f4",
           323 => x"08",
           324 => x"94",
           325 => x"08",
           326 => x"38",
           327 => x"05",
           328 => x"08",
           329 => x"80",
           330 => x"f0",
           331 => x"08",
           332 => x"88",
           333 => x"94",
           334 => x"0c",
           335 => x"05",
           336 => x"fc",
           337 => x"53",
           338 => x"05",
           339 => x"08",
           340 => x"51",
           341 => x"88",
           342 => x"08",
           343 => x"54",
           344 => x"05",
           345 => x"8c",
           346 => x"f8",
           347 => x"94",
           348 => x"0c",
           349 => x"05",
           350 => x"0c",
           351 => x"0d",
           352 => x"94",
           353 => x"0c",
           354 => x"80",
           355 => x"fc",
           356 => x"08",
           357 => x"80",
           358 => x"94",
           359 => x"08",
           360 => x"88",
           361 => x"0b",
           362 => x"05",
           363 => x"8c",
           364 => x"25",
           365 => x"08",
           366 => x"30",
           367 => x"05",
           368 => x"94",
           369 => x"08",
           370 => x"88",
           371 => x"ad",
           372 => x"70",
           373 => x"05",
           374 => x"08",
           375 => x"80",
           376 => x"94",
           377 => x"08",
           378 => x"f8",
           379 => x"08",
           380 => x"70",
           381 => x"87",
           382 => x"0c",
           383 => x"02",
           384 => x"3d",
           385 => x"94",
           386 => x"0c",
           387 => x"08",
           388 => x"94",
           389 => x"08",
           390 => x"05",
           391 => x"38",
           392 => x"05",
           393 => x"a3",
           394 => x"94",
           395 => x"08",
           396 => x"94",
           397 => x"08",
           398 => x"8c",
           399 => x"08",
           400 => x"10",
           401 => x"05",
           402 => x"94",
           403 => x"08",
           404 => x"c9",
           405 => x"8c",
           406 => x"08",
           407 => x"26",
           408 => x"08",
           409 => x"94",
           410 => x"08",
           411 => x"88",
           412 => x"08",
           413 => x"94",
           414 => x"08",
           415 => x"f8",
           416 => x"08",
           417 => x"81",
           418 => x"fc",
           419 => x"08",
           420 => x"81",
           421 => x"8c",
           422 => x"af",
           423 => x"90",
           424 => x"2e",
           425 => x"08",
           426 => x"70",
           427 => x"05",
           428 => x"39",
           429 => x"05",
           430 => x"08",
           431 => x"51",
           432 => x"05",
           433 => x"85",
           434 => x"0c",
           435 => x"0d",
           436 => x"87",
           437 => x"0c",
           438 => x"c0",
           439 => x"85",
           440 => x"98",
           441 => x"c0",
           442 => x"70",
           443 => x"51",
           444 => x"8a",
           445 => x"98",
           446 => x"70",
           447 => x"c0",
           448 => x"fc",
           449 => x"52",
           450 => x"87",
           451 => x"08",
           452 => x"2e",
           453 => x"0b",
           454 => x"f0",
           455 => x"0b",
           456 => x"88",
           457 => x"0d",
           458 => x"0d",
           459 => x"56",
           460 => x"0b",
           461 => x"9f",
           462 => x"06",
           463 => x"52",
           464 => x"09",
           465 => x"9e",
           466 => x"87",
           467 => x"0c",
           468 => x"92",
           469 => x"0b",
           470 => x"8c",
           471 => x"92",
           472 => x"85",
           473 => x"06",
           474 => x"70",
           475 => x"38",
           476 => x"84",
           477 => x"ff",
           478 => x"27",
           479 => x"73",
           480 => x"38",
           481 => x"8b",
           482 => x"70",
           483 => x"34",
           484 => x"81",
           485 => x"a2",
           486 => x"80",
           487 => x"87",
           488 => x"08",
           489 => x"b5",
           490 => x"98",
           491 => x"70",
           492 => x"0b",
           493 => x"8c",
           494 => x"92",
           495 => x"82",
           496 => x"70",
           497 => x"73",
           498 => x"06",
           499 => x"72",
           500 => x"06",
           501 => x"c0",
           502 => x"51",
           503 => x"09",
           504 => x"38",
           505 => x"88",
           506 => x"0d",
           507 => x"0d",
           508 => x"33",
           509 => x"88",
           510 => x"0c",
           511 => x"3d",
           512 => x"3d",
           513 => x"11",
           514 => x"33",
           515 => x"71",
           516 => x"81",
           517 => x"72",
           518 => x"75",
           519 => x"88",
           520 => x"54",
           521 => x"85",
           522 => x"f9",
           523 => x"0b",
           524 => x"f4",
           525 => x"81",
           526 => x"ed",
           527 => x"17",
           528 => x"e5",
           529 => x"55",
           530 => x"89",
           531 => x"2e",
           532 => x"d5",
           533 => x"76",
           534 => x"06",
           535 => x"2a",
           536 => x"05",
           537 => x"70",
           538 => x"bd",
           539 => x"b9",
           540 => x"fe",
           541 => x"08",
           542 => x"06",
           543 => x"84",
           544 => x"2b",
           545 => x"53",
           546 => x"8c",
           547 => x"52",
           548 => x"52",
           549 => x"3f",
           550 => x"38",
           551 => x"e2",
           552 => x"f0",
           553 => x"83",
           554 => x"74",
           555 => x"3d",
           556 => x"3d",
           557 => x"0b",
           558 => x"fe",
           559 => x"08",
           560 => x"56",
           561 => x"74",
           562 => x"38",
           563 => x"75",
           564 => x"16",
           565 => x"53",
           566 => x"87",
           567 => x"fd",
           568 => x"54",
           569 => x"0b",
           570 => x"08",
           571 => x"53",
           572 => x"2e",
           573 => x"8c",
           574 => x"51",
           575 => x"88",
           576 => x"53",
           577 => x"fd",
           578 => x"08",
           579 => x"06",
           580 => x"0c",
           581 => x"04",
           582 => x"76",
           583 => x"9f",
           584 => x"55",
           585 => x"88",
           586 => x"72",
           587 => x"38",
           588 => x"73",
           589 => x"81",
           590 => x"72",
           591 => x"33",
           592 => x"2e",
           593 => x"85",
           594 => x"08",
           595 => x"16",
           596 => x"2e",
           597 => x"51",
           598 => x"88",
           599 => x"39",
           600 => x"52",
           601 => x"0c",
           602 => x"88",
           603 => x"0d",
           604 => x"0d",
           605 => x"0b",
           606 => x"71",
           607 => x"70",
           608 => x"06",
           609 => x"55",
           610 => x"88",
           611 => x"08",
           612 => x"38",
           613 => x"dc",
           614 => x"06",
           615 => x"cf",
           616 => x"90",
           617 => x"15",
           618 => x"8f",
           619 => x"84",
           620 => x"52",
           621 => x"bc",
           622 => x"82",
           623 => x"05",
           624 => x"06",
           625 => x"38",
           626 => x"df",
           627 => x"71",
           628 => x"a0",
           629 => x"88",
           630 => x"08",
           631 => x"88",
           632 => x"0c",
           633 => x"fd",
           634 => x"08",
           635 => x"73",
           636 => x"52",
           637 => x"88",
           638 => x"f2",
           639 => x"62",
           640 => x"5c",
           641 => x"74",
           642 => x"81",
           643 => x"81",
           644 => x"56",
           645 => x"70",
           646 => x"74",
           647 => x"81",
           648 => x"81",
           649 => x"0b",
           650 => x"62",
           651 => x"55",
           652 => x"8f",
           653 => x"fd",
           654 => x"08",
           655 => x"34",
           656 => x"93",
           657 => x"08",
           658 => x"5f",
           659 => x"76",
           660 => x"58",
           661 => x"55",
           662 => x"09",
           663 => x"38",
           664 => x"5b",
           665 => x"5f",
           666 => x"1c",
           667 => x"06",
           668 => x"33",
           669 => x"70",
           670 => x"27",
           671 => x"07",
           672 => x"5b",
           673 => x"55",
           674 => x"38",
           675 => x"09",
           676 => x"38",
           677 => x"7a",
           678 => x"55",
           679 => x"9f",
           680 => x"32",
           681 => x"ae",
           682 => x"70",
           683 => x"2a",
           684 => x"51",
           685 => x"38",
           686 => x"5a",
           687 => x"77",
           688 => x"81",
           689 => x"1c",
           690 => x"55",
           691 => x"ff",
           692 => x"1e",
           693 => x"55",
           694 => x"83",
           695 => x"74",
           696 => x"7b",
           697 => x"3f",
           698 => x"ef",
           699 => x"7b",
           700 => x"2b",
           701 => x"54",
           702 => x"08",
           703 => x"f8",
           704 => x"08",
           705 => x"80",
           706 => x"33",
           707 => x"2e",
           708 => x"8b",
           709 => x"83",
           710 => x"06",
           711 => x"74",
           712 => x"7d",
           713 => x"88",
           714 => x"5b",
           715 => x"58",
           716 => x"9a",
           717 => x"81",
           718 => x"79",
           719 => x"5b",
           720 => x"31",
           721 => x"75",
           722 => x"38",
           723 => x"80",
           724 => x"7b",
           725 => x"3f",
           726 => x"88",
           727 => x"08",
           728 => x"39",
           729 => x"1c",
           730 => x"33",
           731 => x"a5",
           732 => x"33",
           733 => x"70",
           734 => x"56",
           735 => x"38",
           736 => x"39",
           737 => x"39",
           738 => x"d3",
           739 => x"88",
           740 => x"af",
           741 => x"0c",
           742 => x"04",
           743 => x"79",
           744 => x"82",
           745 => x"53",
           746 => x"51",
           747 => x"83",
           748 => x"80",
           749 => x"51",
           750 => x"88",
           751 => x"ff",
           752 => x"56",
           753 => x"d5",
           754 => x"06",
           755 => x"75",
           756 => x"77",
           757 => x"f6",
           758 => x"08",
           759 => x"94",
           760 => x"f8",
           761 => x"08",
           762 => x"06",
           763 => x"82",
           764 => x"38",
           765 => x"d2",
           766 => x"76",
           767 => x"3f",
           768 => x"88",
           769 => x"76",
           770 => x"3f",
           771 => x"ff",
           772 => x"74",
           773 => x"2e",
           774 => x"56",
           775 => x"89",
           776 => x"ed",
           777 => x"59",
           778 => x"0b",
           779 => x"0c",
           780 => x"88",
           781 => x"55",
           782 => x"82",
           783 => x"75",
           784 => x"70",
           785 => x"fe",
           786 => x"08",
           787 => x"57",
           788 => x"09",
           789 => x"38",
           790 => x"be",
           791 => x"75",
           792 => x"3f",
           793 => x"38",
           794 => x"55",
           795 => x"ac",
           796 => x"e4",
           797 => x"8a",
           798 => x"88",
           799 => x"52",
           800 => x"3f",
           801 => x"ff",
           802 => x"83",
           803 => x"06",
           804 => x"56",
           805 => x"76",
           806 => x"38",
           807 => x"8f",
           808 => x"8d",
           809 => x"75",
           810 => x"3f",
           811 => x"08",
           812 => x"95",
           813 => x"51",
           814 => x"88",
           815 => x"ff",
           816 => x"8c",
           817 => x"f3",
           818 => x"b6",
           819 => x"58",
           820 => x"33",
           821 => x"02",
           822 => x"05",
           823 => x"59",
           824 => x"3f",
           825 => x"ff",
           826 => x"05",
           827 => x"8c",
           828 => x"1a",
           829 => x"e0",
           830 => x"f1",
           831 => x"84",
           832 => x"3d",
           833 => x"f5",
           834 => x"08",
           835 => x"06",
           836 => x"38",
           837 => x"05",
           838 => x"3f",
           839 => x"7a",
           840 => x"3f",
           841 => x"ff",
           842 => x"71",
           843 => x"84",
           844 => x"84",
           845 => x"33",
           846 => x"31",
           847 => x"51",
           848 => x"3f",
           849 => x"05",
           850 => x"0c",
           851 => x"8a",
           852 => x"74",
           853 => x"26",
           854 => x"57",
           855 => x"76",
           856 => x"83",
           857 => x"86",
           858 => x"2e",
           859 => x"76",
           860 => x"83",
           861 => x"06",
           862 => x"3d",
           863 => x"f5",
           864 => x"08",
           865 => x"88",
           866 => x"08",
           867 => x"0c",
           868 => x"ff",
           869 => x"08",
           870 => x"2a",
           871 => x"0c",
           872 => x"81",
           873 => x"0b",
           874 => x"f4",
           875 => x"75",
           876 => x"3d",
           877 => x"3d",
           878 => x"0b",
           879 => x"55",
           880 => x"80",
           881 => x"38",
           882 => x"16",
           883 => x"e0",
           884 => x"54",
           885 => x"54",
           886 => x"51",
           887 => x"88",
           888 => x"08",
           889 => x"88",
           890 => x"73",
           891 => x"38",
           892 => x"33",
           893 => x"70",
           894 => x"55",
           895 => x"2e",
           896 => x"54",
           897 => x"51",
           898 => x"88",
           899 => x"0c",
           900 => x"05",
           901 => x"3f",
           902 => x"16",
           903 => x"16",
           904 => x"81",
           905 => x"88",
           906 => x"0d",
           907 => x"0d",
           908 => x"0b",
           909 => x"f4",
           910 => x"5c",
           911 => x"0c",
           912 => x"80",
           913 => x"38",
           914 => x"81",
           915 => x"57",
           916 => x"81",
           917 => x"39",
           918 => x"34",
           919 => x"0b",
           920 => x"81",
           921 => x"39",
           922 => x"98",
           923 => x"55",
           924 => x"83",
           925 => x"77",
           926 => x"9a",
           927 => x"08",
           928 => x"06",
           929 => x"80",
           930 => x"16",
           931 => x"77",
           932 => x"70",
           933 => x"5b",
           934 => x"38",
           935 => x"a0",
           936 => x"8b",
           937 => x"08",
           938 => x"3f",
           939 => x"81",
           940 => x"aa",
           941 => x"17",
           942 => x"08",
           943 => x"3f",
           944 => x"88",
           945 => x"ff",
           946 => x"08",
           947 => x"0c",
           948 => x"83",
           949 => x"80",
           950 => x"55",
           951 => x"83",
           952 => x"74",
           953 => x"08",
           954 => x"53",
           955 => x"52",
           956 => x"b5",
           957 => x"fe",
           958 => x"16",
           959 => x"17",
           960 => x"31",
           961 => x"7c",
           962 => x"80",
           963 => x"38",
           964 => x"fe",
           965 => x"57",
           966 => x"8c",
           967 => x"fb",
           968 => x"c0",
           969 => x"54",
           970 => x"52",
           971 => x"d7",
           972 => x"90",
           973 => x"94",
           974 => x"54",
           975 => x"52",
           976 => x"c3",
           977 => x"08",
           978 => x"94",
           979 => x"c0",
           980 => x"54",
           981 => x"52",
           982 => x"ab",
           983 => x"90",
           984 => x"94",
           985 => x"54",
           986 => x"52",
           987 => x"97",
           988 => x"08",
           989 => x"94",
           990 => x"80",
           991 => x"c0",
           992 => x"8c",
           993 => x"87",
           994 => x"0c",
           995 => x"f9",
           996 => x"08",
           997 => x"e0",
           998 => x"3f",
           999 => x"38",
          1000 => x"88",
          1001 => x"98",
          1002 => x"87",
          1003 => x"53",
          1004 => x"74",
          1005 => x"3f",
          1006 => x"38",
          1007 => x"80",
          1008 => x"73",
          1009 => x"39",
          1010 => x"73",
          1011 => x"fb",
          1012 => x"ff",
          1013 => x"00",
          1014 => x"ff",
          1015 => x"ff",
          1016 => x"4f",
          1017 => x"49",
          1018 => x"52",
          1019 => x"00",
          1020 => x"00",
          2048 => x"0b",
          2049 => x"0b",
          2050 => x"ca",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"0b",
          2057 => x"04",
          2058 => x"c4",
          2059 => x"0b",
          2060 => x"04",
          2061 => x"c4",
          2062 => x"0b",
          2063 => x"04",
          2064 => x"c4",
          2065 => x"0b",
          2066 => x"04",
          2067 => x"c4",
          2068 => x"0b",
          2069 => x"04",
          2070 => x"c5",
          2071 => x"0b",
          2072 => x"04",
          2073 => x"c5",
          2074 => x"0b",
          2075 => x"04",
          2076 => x"c5",
          2077 => x"0b",
          2078 => x"04",
          2079 => x"c5",
          2080 => x"0b",
          2081 => x"04",
          2082 => x"c6",
          2083 => x"0b",
          2084 => x"04",
          2085 => x"c6",
          2086 => x"0b",
          2087 => x"04",
          2088 => x"c6",
          2089 => x"0b",
          2090 => x"04",
          2091 => x"c6",
          2092 => x"0b",
          2093 => x"04",
          2094 => x"c7",
          2095 => x"0b",
          2096 => x"04",
          2097 => x"c7",
          2098 => x"0b",
          2099 => x"04",
          2100 => x"c7",
          2101 => x"0b",
          2102 => x"04",
          2103 => x"c7",
          2104 => x"0b",
          2105 => x"04",
          2106 => x"c8",
          2107 => x"0b",
          2108 => x"04",
          2109 => x"c8",
          2110 => x"0b",
          2111 => x"04",
          2112 => x"c8",
          2113 => x"0b",
          2114 => x"04",
          2115 => x"c8",
          2116 => x"0b",
          2117 => x"04",
          2118 => x"c9",
          2119 => x"0b",
          2120 => x"04",
          2121 => x"c9",
          2122 => x"0b",
          2123 => x"04",
          2124 => x"c9",
          2125 => x"0b",
          2126 => x"04",
          2127 => x"c9",
          2128 => x"0b",
          2129 => x"04",
          2130 => x"ca",
          2131 => x"00",
          2132 => x"00",
          2133 => x"00",
          2134 => x"00",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"80",
          2177 => x"82",
          2178 => x"80",
          2179 => x"82",
          2180 => x"83",
          2181 => x"82",
          2182 => x"80",
          2183 => x"82",
          2184 => x"83",
          2185 => x"82",
          2186 => x"80",
          2187 => x"82",
          2188 => x"83",
          2189 => x"82",
          2190 => x"80",
          2191 => x"82",
          2192 => x"83",
          2193 => x"82",
          2194 => x"80",
          2195 => x"82",
          2196 => x"83",
          2197 => x"82",
          2198 => x"80",
          2199 => x"82",
          2200 => x"83",
          2201 => x"82",
          2202 => x"80",
          2203 => x"82",
          2204 => x"83",
          2205 => x"82",
          2206 => x"80",
          2207 => x"82",
          2208 => x"83",
          2209 => x"82",
          2210 => x"80",
          2211 => x"82",
          2212 => x"83",
          2213 => x"82",
          2214 => x"80",
          2215 => x"82",
          2216 => x"83",
          2217 => x"82",
          2218 => x"80",
          2219 => x"82",
          2220 => x"83",
          2221 => x"82",
          2222 => x"80",
          2223 => x"82",
          2224 => x"83",
          2225 => x"82",
          2226 => x"80",
          2227 => x"82",
          2228 => x"83",
          2229 => x"82",
          2230 => x"80",
          2231 => x"82",
          2232 => x"83",
          2233 => x"82",
          2234 => x"80",
          2235 => x"82",
          2236 => x"83",
          2237 => x"82",
          2238 => x"80",
          2239 => x"82",
          2240 => x"83",
          2241 => x"82",
          2242 => x"80",
          2243 => x"82",
          2244 => x"83",
          2245 => x"82",
          2246 => x"81",
          2247 => x"82",
          2248 => x"83",
          2249 => x"82",
          2250 => x"81",
          2251 => x"82",
          2252 => x"83",
          2253 => x"82",
          2254 => x"81",
          2255 => x"82",
          2256 => x"83",
          2257 => x"82",
          2258 => x"81",
          2259 => x"82",
          2260 => x"83",
          2261 => x"82",
          2262 => x"81",
          2263 => x"82",
          2264 => x"83",
          2265 => x"82",
          2266 => x"81",
          2267 => x"82",
          2268 => x"83",
          2269 => x"82",
          2270 => x"81",
          2271 => x"82",
          2272 => x"83",
          2273 => x"82",
          2274 => x"81",
          2275 => x"82",
          2276 => x"83",
          2277 => x"82",
          2278 => x"81",
          2279 => x"82",
          2280 => x"83",
          2281 => x"82",
          2282 => x"81",
          2283 => x"82",
          2284 => x"83",
          2285 => x"82",
          2286 => x"81",
          2287 => x"82",
          2288 => x"83",
          2289 => x"82",
          2290 => x"81",
          2291 => x"82",
          2292 => x"83",
          2293 => x"82",
          2294 => x"81",
          2295 => x"82",
          2296 => x"83",
          2297 => x"82",
          2298 => x"81",
          2299 => x"82",
          2300 => x"83",
          2301 => x"82",
          2302 => x"81",
          2303 => x"82",
          2304 => x"83",
          2305 => x"82",
          2306 => x"81",
          2307 => x"82",
          2308 => x"83",
          2309 => x"82",
          2310 => x"81",
          2311 => x"82",
          2312 => x"83",
          2313 => x"82",
          2314 => x"81",
          2315 => x"82",
          2316 => x"83",
          2317 => x"82",
          2318 => x"81",
          2319 => x"82",
          2320 => x"83",
          2321 => x"82",
          2322 => x"81",
          2323 => x"82",
          2324 => x"83",
          2325 => x"82",
          2326 => x"81",
          2327 => x"82",
          2328 => x"83",
          2329 => x"82",
          2330 => x"81",
          2331 => x"82",
          2332 => x"83",
          2333 => x"82",
          2334 => x"81",
          2335 => x"82",
          2336 => x"83",
          2337 => x"82",
          2338 => x"81",
          2339 => x"82",
          2340 => x"83",
          2341 => x"82",
          2342 => x"81",
          2343 => x"82",
          2344 => x"83",
          2345 => x"82",
          2346 => x"80",
          2347 => x"82",
          2348 => x"83",
          2349 => x"82",
          2350 => x"80",
          2351 => x"82",
          2352 => x"83",
          2353 => x"82",
          2354 => x"80",
          2355 => x"82",
          2356 => x"83",
          2357 => x"82",
          2358 => x"80",
          2359 => x"82",
          2360 => x"83",
          2361 => x"82",
          2362 => x"80",
          2363 => x"82",
          2364 => x"83",
          2365 => x"82",
          2366 => x"80",
          2367 => x"82",
          2368 => x"83",
          2369 => x"82",
          2370 => x"81",
          2371 => x"82",
          2372 => x"83",
          2373 => x"82",
          2374 => x"82",
          2375 => x"8e",
          2376 => x"70",
          2377 => x"0c",
          2378 => x"ca",
          2379 => x"c4",
          2380 => x"f3",
          2381 => x"04",
          2382 => x"08",
          2383 => x"f8",
          2384 => x"0d",
          2385 => x"8c",
          2386 => x"05",
          2387 => x"8c",
          2388 => x"05",
          2389 => x"c5",
          2390 => x"ec",
          2391 => x"8c",
          2392 => x"85",
          2393 => x"8c",
          2394 => x"82",
          2395 => x"02",
          2396 => x"0c",
          2397 => x"81",
          2398 => x"f8",
          2399 => x"08",
          2400 => x"f8",
          2401 => x"08",
          2402 => x"82",
          2403 => x"70",
          2404 => x"0c",
          2405 => x"0d",
          2406 => x"0c",
          2407 => x"f8",
          2408 => x"8c",
          2409 => x"3d",
          2410 => x"82",
          2411 => x"fc",
          2412 => x"0b",
          2413 => x"08",
          2414 => x"82",
          2415 => x"8c",
          2416 => x"8c",
          2417 => x"05",
          2418 => x"38",
          2419 => x"08",
          2420 => x"80",
          2421 => x"80",
          2422 => x"f8",
          2423 => x"08",
          2424 => x"82",
          2425 => x"8c",
          2426 => x"82",
          2427 => x"8c",
          2428 => x"8c",
          2429 => x"05",
          2430 => x"8c",
          2431 => x"05",
          2432 => x"39",
          2433 => x"08",
          2434 => x"80",
          2435 => x"38",
          2436 => x"08",
          2437 => x"82",
          2438 => x"88",
          2439 => x"ad",
          2440 => x"f8",
          2441 => x"08",
          2442 => x"08",
          2443 => x"31",
          2444 => x"08",
          2445 => x"82",
          2446 => x"f8",
          2447 => x"8c",
          2448 => x"05",
          2449 => x"8c",
          2450 => x"05",
          2451 => x"f8",
          2452 => x"08",
          2453 => x"8c",
          2454 => x"05",
          2455 => x"f8",
          2456 => x"08",
          2457 => x"8c",
          2458 => x"05",
          2459 => x"39",
          2460 => x"08",
          2461 => x"80",
          2462 => x"82",
          2463 => x"88",
          2464 => x"82",
          2465 => x"f4",
          2466 => x"91",
          2467 => x"f8",
          2468 => x"08",
          2469 => x"f8",
          2470 => x"0c",
          2471 => x"f8",
          2472 => x"08",
          2473 => x"0c",
          2474 => x"82",
          2475 => x"04",
          2476 => x"76",
          2477 => x"8c",
          2478 => x"33",
          2479 => x"55",
          2480 => x"8a",
          2481 => x"06",
          2482 => x"2e",
          2483 => x"12",
          2484 => x"2e",
          2485 => x"73",
          2486 => x"55",
          2487 => x"52",
          2488 => x"09",
          2489 => x"38",
          2490 => x"ec",
          2491 => x"0d",
          2492 => x"88",
          2493 => x"70",
          2494 => x"07",
          2495 => x"8f",
          2496 => x"38",
          2497 => x"84",
          2498 => x"72",
          2499 => x"05",
          2500 => x"71",
          2501 => x"53",
          2502 => x"70",
          2503 => x"0c",
          2504 => x"71",
          2505 => x"38",
          2506 => x"90",
          2507 => x"70",
          2508 => x"0c",
          2509 => x"71",
          2510 => x"38",
          2511 => x"8e",
          2512 => x"0d",
          2513 => x"72",
          2514 => x"53",
          2515 => x"93",
          2516 => x"73",
          2517 => x"54",
          2518 => x"2e",
          2519 => x"73",
          2520 => x"71",
          2521 => x"ff",
          2522 => x"70",
          2523 => x"38",
          2524 => x"70",
          2525 => x"81",
          2526 => x"81",
          2527 => x"71",
          2528 => x"ff",
          2529 => x"54",
          2530 => x"38",
          2531 => x"73",
          2532 => x"75",
          2533 => x"71",
          2534 => x"8c",
          2535 => x"52",
          2536 => x"04",
          2537 => x"f7",
          2538 => x"14",
          2539 => x"84",
          2540 => x"06",
          2541 => x"70",
          2542 => x"14",
          2543 => x"08",
          2544 => x"71",
          2545 => x"dc",
          2546 => x"54",
          2547 => x"39",
          2548 => x"8c",
          2549 => x"3d",
          2550 => x"3d",
          2551 => x"83",
          2552 => x"2b",
          2553 => x"3f",
          2554 => x"08",
          2555 => x"72",
          2556 => x"54",
          2557 => x"25",
          2558 => x"82",
          2559 => x"84",
          2560 => x"fb",
          2561 => x"70",
          2562 => x"53",
          2563 => x"2e",
          2564 => x"71",
          2565 => x"a0",
          2566 => x"06",
          2567 => x"12",
          2568 => x"71",
          2569 => x"81",
          2570 => x"73",
          2571 => x"ff",
          2572 => x"55",
          2573 => x"83",
          2574 => x"70",
          2575 => x"38",
          2576 => x"73",
          2577 => x"51",
          2578 => x"09",
          2579 => x"38",
          2580 => x"81",
          2581 => x"72",
          2582 => x"51",
          2583 => x"ec",
          2584 => x"0d",
          2585 => x"0d",
          2586 => x"08",
          2587 => x"38",
          2588 => x"05",
          2589 => x"9b",
          2590 => x"8c",
          2591 => x"38",
          2592 => x"39",
          2593 => x"82",
          2594 => x"86",
          2595 => x"fc",
          2596 => x"82",
          2597 => x"05",
          2598 => x"52",
          2599 => x"81",
          2600 => x"13",
          2601 => x"51",
          2602 => x"9e",
          2603 => x"38",
          2604 => x"51",
          2605 => x"97",
          2606 => x"38",
          2607 => x"51",
          2608 => x"bb",
          2609 => x"38",
          2610 => x"51",
          2611 => x"bb",
          2612 => x"38",
          2613 => x"55",
          2614 => x"87",
          2615 => x"d9",
          2616 => x"22",
          2617 => x"73",
          2618 => x"80",
          2619 => x"0b",
          2620 => x"9c",
          2621 => x"87",
          2622 => x"0c",
          2623 => x"87",
          2624 => x"0c",
          2625 => x"87",
          2626 => x"0c",
          2627 => x"87",
          2628 => x"0c",
          2629 => x"87",
          2630 => x"0c",
          2631 => x"87",
          2632 => x"0c",
          2633 => x"98",
          2634 => x"87",
          2635 => x"0c",
          2636 => x"c0",
          2637 => x"80",
          2638 => x"8c",
          2639 => x"3d",
          2640 => x"3d",
          2641 => x"87",
          2642 => x"5d",
          2643 => x"87",
          2644 => x"08",
          2645 => x"23",
          2646 => x"b8",
          2647 => x"82",
          2648 => x"c0",
          2649 => x"5a",
          2650 => x"34",
          2651 => x"b0",
          2652 => x"84",
          2653 => x"c0",
          2654 => x"5a",
          2655 => x"34",
          2656 => x"a8",
          2657 => x"86",
          2658 => x"c0",
          2659 => x"5c",
          2660 => x"23",
          2661 => x"a0",
          2662 => x"8a",
          2663 => x"7d",
          2664 => x"ff",
          2665 => x"7b",
          2666 => x"06",
          2667 => x"33",
          2668 => x"33",
          2669 => x"33",
          2670 => x"33",
          2671 => x"33",
          2672 => x"ff",
          2673 => x"81",
          2674 => x"94",
          2675 => x"3d",
          2676 => x"3d",
          2677 => x"05",
          2678 => x"70",
          2679 => x"52",
          2680 => x"0b",
          2681 => x"34",
          2682 => x"04",
          2683 => x"77",
          2684 => x"89",
          2685 => x"81",
          2686 => x"55",
          2687 => x"94",
          2688 => x"80",
          2689 => x"87",
          2690 => x"51",
          2691 => x"96",
          2692 => x"06",
          2693 => x"70",
          2694 => x"38",
          2695 => x"70",
          2696 => x"51",
          2697 => x"72",
          2698 => x"81",
          2699 => x"70",
          2700 => x"38",
          2701 => x"70",
          2702 => x"51",
          2703 => x"38",
          2704 => x"06",
          2705 => x"94",
          2706 => x"80",
          2707 => x"87",
          2708 => x"52",
          2709 => x"75",
          2710 => x"0c",
          2711 => x"04",
          2712 => x"02",
          2713 => x"0b",
          2714 => x"94",
          2715 => x"ff",
          2716 => x"56",
          2717 => x"84",
          2718 => x"2e",
          2719 => x"c0",
          2720 => x"70",
          2721 => x"2a",
          2722 => x"53",
          2723 => x"80",
          2724 => x"71",
          2725 => x"81",
          2726 => x"70",
          2727 => x"81",
          2728 => x"06",
          2729 => x"80",
          2730 => x"71",
          2731 => x"81",
          2732 => x"70",
          2733 => x"73",
          2734 => x"51",
          2735 => x"80",
          2736 => x"2e",
          2737 => x"c0",
          2738 => x"75",
          2739 => x"3d",
          2740 => x"3d",
          2741 => x"80",
          2742 => x"81",
          2743 => x"53",
          2744 => x"2e",
          2745 => x"71",
          2746 => x"81",
          2747 => x"82",
          2748 => x"70",
          2749 => x"59",
          2750 => x"87",
          2751 => x"51",
          2752 => x"86",
          2753 => x"94",
          2754 => x"08",
          2755 => x"70",
          2756 => x"54",
          2757 => x"2e",
          2758 => x"91",
          2759 => x"06",
          2760 => x"d7",
          2761 => x"32",
          2762 => x"51",
          2763 => x"2e",
          2764 => x"93",
          2765 => x"06",
          2766 => x"ff",
          2767 => x"81",
          2768 => x"87",
          2769 => x"52",
          2770 => x"86",
          2771 => x"94",
          2772 => x"72",
          2773 => x"74",
          2774 => x"ff",
          2775 => x"57",
          2776 => x"38",
          2777 => x"ec",
          2778 => x"0d",
          2779 => x"0d",
          2780 => x"89",
          2781 => x"81",
          2782 => x"52",
          2783 => x"84",
          2784 => x"2e",
          2785 => x"c0",
          2786 => x"70",
          2787 => x"2a",
          2788 => x"51",
          2789 => x"80",
          2790 => x"71",
          2791 => x"51",
          2792 => x"80",
          2793 => x"2e",
          2794 => x"c0",
          2795 => x"71",
          2796 => x"ff",
          2797 => x"ec",
          2798 => x"3d",
          2799 => x"3d",
          2800 => x"82",
          2801 => x"70",
          2802 => x"52",
          2803 => x"94",
          2804 => x"80",
          2805 => x"87",
          2806 => x"52",
          2807 => x"82",
          2808 => x"06",
          2809 => x"ff",
          2810 => x"2e",
          2811 => x"81",
          2812 => x"87",
          2813 => x"52",
          2814 => x"86",
          2815 => x"94",
          2816 => x"08",
          2817 => x"70",
          2818 => x"53",
          2819 => x"8c",
          2820 => x"3d",
          2821 => x"3d",
          2822 => x"9e",
          2823 => x"9c",
          2824 => x"51",
          2825 => x"2e",
          2826 => x"87",
          2827 => x"08",
          2828 => x"0c",
          2829 => x"a8",
          2830 => x"9c",
          2831 => x"9e",
          2832 => x"89",
          2833 => x"c0",
          2834 => x"82",
          2835 => x"87",
          2836 => x"08",
          2837 => x"0c",
          2838 => x"a0",
          2839 => x"ac",
          2840 => x"9e",
          2841 => x"89",
          2842 => x"c0",
          2843 => x"82",
          2844 => x"87",
          2845 => x"08",
          2846 => x"0c",
          2847 => x"b8",
          2848 => x"bc",
          2849 => x"9e",
          2850 => x"89",
          2851 => x"c0",
          2852 => x"82",
          2853 => x"87",
          2854 => x"08",
          2855 => x"0c",
          2856 => x"80",
          2857 => x"82",
          2858 => x"87",
          2859 => x"08",
          2860 => x"0c",
          2861 => x"88",
          2862 => x"d4",
          2863 => x"9e",
          2864 => x"89",
          2865 => x"0b",
          2866 => x"34",
          2867 => x"c0",
          2868 => x"70",
          2869 => x"06",
          2870 => x"70",
          2871 => x"38",
          2872 => x"82",
          2873 => x"80",
          2874 => x"9e",
          2875 => x"88",
          2876 => x"51",
          2877 => x"80",
          2878 => x"81",
          2879 => x"89",
          2880 => x"0b",
          2881 => x"90",
          2882 => x"80",
          2883 => x"52",
          2884 => x"2e",
          2885 => x"52",
          2886 => x"df",
          2887 => x"87",
          2888 => x"08",
          2889 => x"80",
          2890 => x"52",
          2891 => x"83",
          2892 => x"71",
          2893 => x"34",
          2894 => x"c0",
          2895 => x"70",
          2896 => x"06",
          2897 => x"70",
          2898 => x"38",
          2899 => x"82",
          2900 => x"80",
          2901 => x"9e",
          2902 => x"90",
          2903 => x"51",
          2904 => x"80",
          2905 => x"81",
          2906 => x"89",
          2907 => x"0b",
          2908 => x"90",
          2909 => x"80",
          2910 => x"52",
          2911 => x"2e",
          2912 => x"52",
          2913 => x"e3",
          2914 => x"87",
          2915 => x"08",
          2916 => x"80",
          2917 => x"52",
          2918 => x"83",
          2919 => x"71",
          2920 => x"34",
          2921 => x"c0",
          2922 => x"70",
          2923 => x"06",
          2924 => x"70",
          2925 => x"38",
          2926 => x"82",
          2927 => x"80",
          2928 => x"9e",
          2929 => x"80",
          2930 => x"51",
          2931 => x"80",
          2932 => x"81",
          2933 => x"89",
          2934 => x"0b",
          2935 => x"90",
          2936 => x"80",
          2937 => x"52",
          2938 => x"83",
          2939 => x"71",
          2940 => x"34",
          2941 => x"90",
          2942 => x"80",
          2943 => x"2a",
          2944 => x"70",
          2945 => x"34",
          2946 => x"c0",
          2947 => x"70",
          2948 => x"51",
          2949 => x"80",
          2950 => x"81",
          2951 => x"89",
          2952 => x"c0",
          2953 => x"70",
          2954 => x"70",
          2955 => x"51",
          2956 => x"89",
          2957 => x"0b",
          2958 => x"90",
          2959 => x"06",
          2960 => x"70",
          2961 => x"38",
          2962 => x"82",
          2963 => x"87",
          2964 => x"08",
          2965 => x"51",
          2966 => x"89",
          2967 => x"3d",
          2968 => x"3d",
          2969 => x"84",
          2970 => x"3f",
          2971 => x"33",
          2972 => x"2e",
          2973 => x"f6",
          2974 => x"b6",
          2975 => x"ac",
          2976 => x"3f",
          2977 => x"33",
          2978 => x"2e",
          2979 => x"89",
          2980 => x"89",
          2981 => x"54",
          2982 => x"c4",
          2983 => x"3f",
          2984 => x"33",
          2985 => x"2e",
          2986 => x"89",
          2987 => x"89",
          2988 => x"54",
          2989 => x"e0",
          2990 => x"3f",
          2991 => x"33",
          2992 => x"2e",
          2993 => x"89",
          2994 => x"89",
          2995 => x"54",
          2996 => x"fc",
          2997 => x"3f",
          2998 => x"33",
          2999 => x"2e",
          3000 => x"89",
          3001 => x"89",
          3002 => x"54",
          3003 => x"98",
          3004 => x"3f",
          3005 => x"33",
          3006 => x"2e",
          3007 => x"89",
          3008 => x"89",
          3009 => x"54",
          3010 => x"b4",
          3011 => x"3f",
          3012 => x"33",
          3013 => x"2e",
          3014 => x"89",
          3015 => x"81",
          3016 => x"89",
          3017 => x"89",
          3018 => x"73",
          3019 => x"38",
          3020 => x"33",
          3021 => x"f0",
          3022 => x"3f",
          3023 => x"33",
          3024 => x"2e",
          3025 => x"89",
          3026 => x"81",
          3027 => x"89",
          3028 => x"89",
          3029 => x"73",
          3030 => x"38",
          3031 => x"51",
          3032 => x"82",
          3033 => x"54",
          3034 => x"88",
          3035 => x"c4",
          3036 => x"3f",
          3037 => x"33",
          3038 => x"2e",
          3039 => x"f8",
          3040 => x"ae",
          3041 => x"e5",
          3042 => x"80",
          3043 => x"81",
          3044 => x"83",
          3045 => x"89",
          3046 => x"73",
          3047 => x"38",
          3048 => x"51",
          3049 => x"81",
          3050 => x"83",
          3051 => x"89",
          3052 => x"81",
          3053 => x"88",
          3054 => x"89",
          3055 => x"81",
          3056 => x"88",
          3057 => x"89",
          3058 => x"81",
          3059 => x"88",
          3060 => x"f9",
          3061 => x"da",
          3062 => x"cc",
          3063 => x"fa",
          3064 => x"b2",
          3065 => x"d0",
          3066 => x"84",
          3067 => x"51",
          3068 => x"82",
          3069 => x"bd",
          3070 => x"76",
          3071 => x"54",
          3072 => x"08",
          3073 => x"a8",
          3074 => x"3f",
          3075 => x"33",
          3076 => x"2e",
          3077 => x"89",
          3078 => x"bd",
          3079 => x"75",
          3080 => x"3f",
          3081 => x"08",
          3082 => x"29",
          3083 => x"54",
          3084 => x"ec",
          3085 => x"fa",
          3086 => x"da",
          3087 => x"de",
          3088 => x"80",
          3089 => x"82",
          3090 => x"56",
          3091 => x"52",
          3092 => x"e4",
          3093 => x"ec",
          3094 => x"c0",
          3095 => x"31",
          3096 => x"8c",
          3097 => x"81",
          3098 => x"87",
          3099 => x"86",
          3100 => x"be",
          3101 => x"0d",
          3102 => x"0d",
          3103 => x"33",
          3104 => x"71",
          3105 => x"38",
          3106 => x"0b",
          3107 => x"88",
          3108 => x"08",
          3109 => x"ac",
          3110 => x"81",
          3111 => x"97",
          3112 => x"bc",
          3113 => x"81",
          3114 => x"8b",
          3115 => x"c8",
          3116 => x"81",
          3117 => x"80",
          3118 => x"3d",
          3119 => x"88",
          3120 => x"80",
          3121 => x"96",
          3122 => x"82",
          3123 => x"87",
          3124 => x"0c",
          3125 => x"0d",
          3126 => x"33",
          3127 => x"2e",
          3128 => x"85",
          3129 => x"ed",
          3130 => x"84",
          3131 => x"80",
          3132 => x"72",
          3133 => x"8d",
          3134 => x"05",
          3135 => x"0c",
          3136 => x"8c",
          3137 => x"71",
          3138 => x"38",
          3139 => x"2d",
          3140 => x"04",
          3141 => x"02",
          3142 => x"82",
          3143 => x"76",
          3144 => x"0c",
          3145 => x"ad",
          3146 => x"8c",
          3147 => x"3d",
          3148 => x"3d",
          3149 => x"73",
          3150 => x"ff",
          3151 => x"71",
          3152 => x"38",
          3153 => x"06",
          3154 => x"54",
          3155 => x"e7",
          3156 => x"0d",
          3157 => x"0d",
          3158 => x"fc",
          3159 => x"8c",
          3160 => x"54",
          3161 => x"81",
          3162 => x"53",
          3163 => x"8e",
          3164 => x"ff",
          3165 => x"14",
          3166 => x"3f",
          3167 => x"82",
          3168 => x"86",
          3169 => x"ec",
          3170 => x"68",
          3171 => x"70",
          3172 => x"33",
          3173 => x"2e",
          3174 => x"75",
          3175 => x"81",
          3176 => x"38",
          3177 => x"70",
          3178 => x"33",
          3179 => x"75",
          3180 => x"81",
          3181 => x"81",
          3182 => x"75",
          3183 => x"81",
          3184 => x"82",
          3185 => x"81",
          3186 => x"56",
          3187 => x"09",
          3188 => x"38",
          3189 => x"71",
          3190 => x"81",
          3191 => x"59",
          3192 => x"9d",
          3193 => x"53",
          3194 => x"95",
          3195 => x"29",
          3196 => x"76",
          3197 => x"79",
          3198 => x"5b",
          3199 => x"e5",
          3200 => x"ec",
          3201 => x"70",
          3202 => x"25",
          3203 => x"32",
          3204 => x"72",
          3205 => x"73",
          3206 => x"58",
          3207 => x"73",
          3208 => x"38",
          3209 => x"79",
          3210 => x"5b",
          3211 => x"75",
          3212 => x"de",
          3213 => x"80",
          3214 => x"89",
          3215 => x"70",
          3216 => x"55",
          3217 => x"cf",
          3218 => x"38",
          3219 => x"24",
          3220 => x"80",
          3221 => x"8e",
          3222 => x"c3",
          3223 => x"73",
          3224 => x"81",
          3225 => x"99",
          3226 => x"c4",
          3227 => x"38",
          3228 => x"73",
          3229 => x"81",
          3230 => x"80",
          3231 => x"38",
          3232 => x"2e",
          3233 => x"f9",
          3234 => x"d8",
          3235 => x"38",
          3236 => x"77",
          3237 => x"08",
          3238 => x"80",
          3239 => x"55",
          3240 => x"8d",
          3241 => x"70",
          3242 => x"51",
          3243 => x"f5",
          3244 => x"2a",
          3245 => x"74",
          3246 => x"53",
          3247 => x"8f",
          3248 => x"fc",
          3249 => x"81",
          3250 => x"80",
          3251 => x"73",
          3252 => x"3f",
          3253 => x"56",
          3254 => x"27",
          3255 => x"a0",
          3256 => x"3f",
          3257 => x"84",
          3258 => x"33",
          3259 => x"93",
          3260 => x"95",
          3261 => x"91",
          3262 => x"8d",
          3263 => x"89",
          3264 => x"fb",
          3265 => x"86",
          3266 => x"2a",
          3267 => x"51",
          3268 => x"2e",
          3269 => x"84",
          3270 => x"86",
          3271 => x"78",
          3272 => x"08",
          3273 => x"32",
          3274 => x"72",
          3275 => x"51",
          3276 => x"74",
          3277 => x"38",
          3278 => x"88",
          3279 => x"7a",
          3280 => x"55",
          3281 => x"3d",
          3282 => x"52",
          3283 => x"9b",
          3284 => x"ec",
          3285 => x"06",
          3286 => x"52",
          3287 => x"3f",
          3288 => x"08",
          3289 => x"27",
          3290 => x"14",
          3291 => x"f8",
          3292 => x"87",
          3293 => x"81",
          3294 => x"b0",
          3295 => x"7d",
          3296 => x"5f",
          3297 => x"75",
          3298 => x"07",
          3299 => x"54",
          3300 => x"26",
          3301 => x"ff",
          3302 => x"84",
          3303 => x"06",
          3304 => x"80",
          3305 => x"96",
          3306 => x"e0",
          3307 => x"73",
          3308 => x"57",
          3309 => x"06",
          3310 => x"54",
          3311 => x"a0",
          3312 => x"2a",
          3313 => x"54",
          3314 => x"38",
          3315 => x"76",
          3316 => x"38",
          3317 => x"fd",
          3318 => x"06",
          3319 => x"38",
          3320 => x"56",
          3321 => x"26",
          3322 => x"3d",
          3323 => x"05",
          3324 => x"ff",
          3325 => x"53",
          3326 => x"d9",
          3327 => x"38",
          3328 => x"56",
          3329 => x"27",
          3330 => x"a0",
          3331 => x"3f",
          3332 => x"3d",
          3333 => x"3d",
          3334 => x"70",
          3335 => x"52",
          3336 => x"73",
          3337 => x"3f",
          3338 => x"04",
          3339 => x"74",
          3340 => x"0c",
          3341 => x"05",
          3342 => x"fa",
          3343 => x"8d",
          3344 => x"80",
          3345 => x"0b",
          3346 => x"0c",
          3347 => x"04",
          3348 => x"82",
          3349 => x"76",
          3350 => x"0c",
          3351 => x"05",
          3352 => x"53",
          3353 => x"72",
          3354 => x"0c",
          3355 => x"04",
          3356 => x"77",
          3357 => x"80",
          3358 => x"54",
          3359 => x"54",
          3360 => x"80",
          3361 => x"8d",
          3362 => x"71",
          3363 => x"ec",
          3364 => x"06",
          3365 => x"2e",
          3366 => x"72",
          3367 => x"38",
          3368 => x"70",
          3369 => x"25",
          3370 => x"73",
          3371 => x"38",
          3372 => x"86",
          3373 => x"54",
          3374 => x"73",
          3375 => x"ff",
          3376 => x"72",
          3377 => x"74",
          3378 => x"72",
          3379 => x"54",
          3380 => x"81",
          3381 => x"39",
          3382 => x"80",
          3383 => x"51",
          3384 => x"81",
          3385 => x"8c",
          3386 => x"3d",
          3387 => x"3d",
          3388 => x"80",
          3389 => x"8d",
          3390 => x"53",
          3391 => x"fe",
          3392 => x"82",
          3393 => x"84",
          3394 => x"f8",
          3395 => x"7c",
          3396 => x"70",
          3397 => x"75",
          3398 => x"55",
          3399 => x"2e",
          3400 => x"87",
          3401 => x"76",
          3402 => x"73",
          3403 => x"81",
          3404 => x"81",
          3405 => x"77",
          3406 => x"70",
          3407 => x"58",
          3408 => x"09",
          3409 => x"c2",
          3410 => x"81",
          3411 => x"75",
          3412 => x"55",
          3413 => x"e2",
          3414 => x"90",
          3415 => x"f8",
          3416 => x"8f",
          3417 => x"81",
          3418 => x"75",
          3419 => x"55",
          3420 => x"81",
          3421 => x"27",
          3422 => x"d0",
          3423 => x"55",
          3424 => x"73",
          3425 => x"80",
          3426 => x"14",
          3427 => x"72",
          3428 => x"e0",
          3429 => x"80",
          3430 => x"39",
          3431 => x"55",
          3432 => x"80",
          3433 => x"e0",
          3434 => x"38",
          3435 => x"81",
          3436 => x"53",
          3437 => x"81",
          3438 => x"53",
          3439 => x"8e",
          3440 => x"70",
          3441 => x"55",
          3442 => x"27",
          3443 => x"77",
          3444 => x"74",
          3445 => x"76",
          3446 => x"77",
          3447 => x"70",
          3448 => x"55",
          3449 => x"77",
          3450 => x"38",
          3451 => x"74",
          3452 => x"55",
          3453 => x"ec",
          3454 => x"0d",
          3455 => x"0d",
          3456 => x"56",
          3457 => x"0c",
          3458 => x"70",
          3459 => x"73",
          3460 => x"81",
          3461 => x"81",
          3462 => x"ed",
          3463 => x"2e",
          3464 => x"8e",
          3465 => x"08",
          3466 => x"76",
          3467 => x"56",
          3468 => x"b0",
          3469 => x"06",
          3470 => x"75",
          3471 => x"76",
          3472 => x"70",
          3473 => x"73",
          3474 => x"8b",
          3475 => x"73",
          3476 => x"85",
          3477 => x"82",
          3478 => x"76",
          3479 => x"70",
          3480 => x"ac",
          3481 => x"a0",
          3482 => x"fa",
          3483 => x"53",
          3484 => x"57",
          3485 => x"98",
          3486 => x"39",
          3487 => x"80",
          3488 => x"26",
          3489 => x"86",
          3490 => x"80",
          3491 => x"57",
          3492 => x"74",
          3493 => x"38",
          3494 => x"27",
          3495 => x"14",
          3496 => x"06",
          3497 => x"14",
          3498 => x"06",
          3499 => x"74",
          3500 => x"f9",
          3501 => x"ff",
          3502 => x"89",
          3503 => x"38",
          3504 => x"c5",
          3505 => x"29",
          3506 => x"81",
          3507 => x"76",
          3508 => x"56",
          3509 => x"ba",
          3510 => x"2e",
          3511 => x"30",
          3512 => x"0c",
          3513 => x"82",
          3514 => x"8a",
          3515 => x"ff",
          3516 => x"8f",
          3517 => x"81",
          3518 => x"26",
          3519 => x"89",
          3520 => x"52",
          3521 => x"ec",
          3522 => x"0d",
          3523 => x"0d",
          3524 => x"33",
          3525 => x"9f",
          3526 => x"53",
          3527 => x"81",
          3528 => x"38",
          3529 => x"87",
          3530 => x"11",
          3531 => x"54",
          3532 => x"84",
          3533 => x"54",
          3534 => x"87",
          3535 => x"11",
          3536 => x"0c",
          3537 => x"c0",
          3538 => x"70",
          3539 => x"70",
          3540 => x"51",
          3541 => x"8a",
          3542 => x"98",
          3543 => x"70",
          3544 => x"08",
          3545 => x"06",
          3546 => x"38",
          3547 => x"8c",
          3548 => x"80",
          3549 => x"71",
          3550 => x"14",
          3551 => x"f4",
          3552 => x"70",
          3553 => x"0c",
          3554 => x"04",
          3555 => x"60",
          3556 => x"8c",
          3557 => x"33",
          3558 => x"5b",
          3559 => x"5a",
          3560 => x"82",
          3561 => x"81",
          3562 => x"52",
          3563 => x"38",
          3564 => x"84",
          3565 => x"92",
          3566 => x"c0",
          3567 => x"87",
          3568 => x"13",
          3569 => x"57",
          3570 => x"0b",
          3571 => x"8c",
          3572 => x"0c",
          3573 => x"75",
          3574 => x"2a",
          3575 => x"51",
          3576 => x"80",
          3577 => x"7b",
          3578 => x"7b",
          3579 => x"5d",
          3580 => x"59",
          3581 => x"06",
          3582 => x"73",
          3583 => x"81",
          3584 => x"ff",
          3585 => x"72",
          3586 => x"38",
          3587 => x"8c",
          3588 => x"c3",
          3589 => x"98",
          3590 => x"71",
          3591 => x"38",
          3592 => x"2e",
          3593 => x"76",
          3594 => x"92",
          3595 => x"72",
          3596 => x"06",
          3597 => x"f7",
          3598 => x"5a",
          3599 => x"80",
          3600 => x"70",
          3601 => x"5a",
          3602 => x"80",
          3603 => x"73",
          3604 => x"06",
          3605 => x"38",
          3606 => x"fe",
          3607 => x"fc",
          3608 => x"52",
          3609 => x"83",
          3610 => x"71",
          3611 => x"8c",
          3612 => x"3d",
          3613 => x"3d",
          3614 => x"64",
          3615 => x"bf",
          3616 => x"40",
          3617 => x"59",
          3618 => x"58",
          3619 => x"82",
          3620 => x"81",
          3621 => x"52",
          3622 => x"09",
          3623 => x"b1",
          3624 => x"84",
          3625 => x"92",
          3626 => x"c0",
          3627 => x"87",
          3628 => x"13",
          3629 => x"56",
          3630 => x"87",
          3631 => x"0c",
          3632 => x"82",
          3633 => x"58",
          3634 => x"84",
          3635 => x"06",
          3636 => x"71",
          3637 => x"38",
          3638 => x"05",
          3639 => x"0c",
          3640 => x"73",
          3641 => x"81",
          3642 => x"71",
          3643 => x"38",
          3644 => x"8c",
          3645 => x"d0",
          3646 => x"98",
          3647 => x"71",
          3648 => x"38",
          3649 => x"2e",
          3650 => x"76",
          3651 => x"92",
          3652 => x"72",
          3653 => x"06",
          3654 => x"f7",
          3655 => x"59",
          3656 => x"1a",
          3657 => x"06",
          3658 => x"59",
          3659 => x"80",
          3660 => x"73",
          3661 => x"06",
          3662 => x"38",
          3663 => x"fe",
          3664 => x"fc",
          3665 => x"52",
          3666 => x"83",
          3667 => x"71",
          3668 => x"8c",
          3669 => x"3d",
          3670 => x"3d",
          3671 => x"84",
          3672 => x"33",
          3673 => x"a7",
          3674 => x"54",
          3675 => x"fa",
          3676 => x"8c",
          3677 => x"06",
          3678 => x"72",
          3679 => x"85",
          3680 => x"98",
          3681 => x"56",
          3682 => x"80",
          3683 => x"76",
          3684 => x"74",
          3685 => x"c0",
          3686 => x"54",
          3687 => x"2e",
          3688 => x"d4",
          3689 => x"2e",
          3690 => x"80",
          3691 => x"08",
          3692 => x"70",
          3693 => x"51",
          3694 => x"2e",
          3695 => x"c0",
          3696 => x"52",
          3697 => x"87",
          3698 => x"08",
          3699 => x"38",
          3700 => x"87",
          3701 => x"14",
          3702 => x"70",
          3703 => x"52",
          3704 => x"96",
          3705 => x"92",
          3706 => x"0a",
          3707 => x"39",
          3708 => x"0c",
          3709 => x"39",
          3710 => x"54",
          3711 => x"ec",
          3712 => x"0d",
          3713 => x"0d",
          3714 => x"33",
          3715 => x"88",
          3716 => x"8c",
          3717 => x"51",
          3718 => x"04",
          3719 => x"75",
          3720 => x"82",
          3721 => x"90",
          3722 => x"2b",
          3723 => x"33",
          3724 => x"88",
          3725 => x"71",
          3726 => x"ec",
          3727 => x"54",
          3728 => x"85",
          3729 => x"ff",
          3730 => x"02",
          3731 => x"05",
          3732 => x"70",
          3733 => x"05",
          3734 => x"88",
          3735 => x"72",
          3736 => x"0d",
          3737 => x"0d",
          3738 => x"52",
          3739 => x"81",
          3740 => x"70",
          3741 => x"70",
          3742 => x"05",
          3743 => x"88",
          3744 => x"72",
          3745 => x"54",
          3746 => x"2a",
          3747 => x"34",
          3748 => x"04",
          3749 => x"76",
          3750 => x"54",
          3751 => x"2e",
          3752 => x"70",
          3753 => x"33",
          3754 => x"05",
          3755 => x"11",
          3756 => x"84",
          3757 => x"fe",
          3758 => x"77",
          3759 => x"53",
          3760 => x"81",
          3761 => x"ff",
          3762 => x"f4",
          3763 => x"0d",
          3764 => x"0d",
          3765 => x"56",
          3766 => x"70",
          3767 => x"33",
          3768 => x"05",
          3769 => x"71",
          3770 => x"56",
          3771 => x"72",
          3772 => x"38",
          3773 => x"e2",
          3774 => x"8c",
          3775 => x"3d",
          3776 => x"3d",
          3777 => x"54",
          3778 => x"71",
          3779 => x"38",
          3780 => x"70",
          3781 => x"f3",
          3782 => x"82",
          3783 => x"84",
          3784 => x"80",
          3785 => x"ec",
          3786 => x"0b",
          3787 => x"0c",
          3788 => x"0d",
          3789 => x"0b",
          3790 => x"56",
          3791 => x"2e",
          3792 => x"81",
          3793 => x"08",
          3794 => x"70",
          3795 => x"33",
          3796 => x"a2",
          3797 => x"ec",
          3798 => x"09",
          3799 => x"38",
          3800 => x"08",
          3801 => x"b0",
          3802 => x"a4",
          3803 => x"9c",
          3804 => x"56",
          3805 => x"27",
          3806 => x"16",
          3807 => x"82",
          3808 => x"06",
          3809 => x"54",
          3810 => x"78",
          3811 => x"33",
          3812 => x"3f",
          3813 => x"5a",
          3814 => x"ec",
          3815 => x"0d",
          3816 => x"0d",
          3817 => x"56",
          3818 => x"b0",
          3819 => x"af",
          3820 => x"fe",
          3821 => x"8c",
          3822 => x"82",
          3823 => x"9f",
          3824 => x"74",
          3825 => x"52",
          3826 => x"51",
          3827 => x"82",
          3828 => x"80",
          3829 => x"ff",
          3830 => x"74",
          3831 => x"76",
          3832 => x"0c",
          3833 => x"04",
          3834 => x"7a",
          3835 => x"fe",
          3836 => x"8c",
          3837 => x"82",
          3838 => x"81",
          3839 => x"33",
          3840 => x"2e",
          3841 => x"80",
          3842 => x"17",
          3843 => x"81",
          3844 => x"06",
          3845 => x"84",
          3846 => x"8c",
          3847 => x"b4",
          3848 => x"56",
          3849 => x"82",
          3850 => x"84",
          3851 => x"fc",
          3852 => x"8b",
          3853 => x"52",
          3854 => x"a9",
          3855 => x"85",
          3856 => x"84",
          3857 => x"fc",
          3858 => x"17",
          3859 => x"9c",
          3860 => x"91",
          3861 => x"08",
          3862 => x"17",
          3863 => x"3f",
          3864 => x"81",
          3865 => x"19",
          3866 => x"53",
          3867 => x"17",
          3868 => x"82",
          3869 => x"18",
          3870 => x"80",
          3871 => x"33",
          3872 => x"3f",
          3873 => x"08",
          3874 => x"38",
          3875 => x"82",
          3876 => x"8a",
          3877 => x"fb",
          3878 => x"fe",
          3879 => x"08",
          3880 => x"56",
          3881 => x"74",
          3882 => x"38",
          3883 => x"75",
          3884 => x"16",
          3885 => x"53",
          3886 => x"ec",
          3887 => x"0d",
          3888 => x"0d",
          3889 => x"08",
          3890 => x"81",
          3891 => x"df",
          3892 => x"15",
          3893 => x"d7",
          3894 => x"33",
          3895 => x"82",
          3896 => x"38",
          3897 => x"89",
          3898 => x"2e",
          3899 => x"bf",
          3900 => x"2e",
          3901 => x"81",
          3902 => x"81",
          3903 => x"89",
          3904 => x"08",
          3905 => x"52",
          3906 => x"3f",
          3907 => x"08",
          3908 => x"74",
          3909 => x"14",
          3910 => x"81",
          3911 => x"2a",
          3912 => x"05",
          3913 => x"57",
          3914 => x"f5",
          3915 => x"ec",
          3916 => x"38",
          3917 => x"06",
          3918 => x"33",
          3919 => x"78",
          3920 => x"06",
          3921 => x"5c",
          3922 => x"53",
          3923 => x"38",
          3924 => x"06",
          3925 => x"39",
          3926 => x"a4",
          3927 => x"52",
          3928 => x"bd",
          3929 => x"ec",
          3930 => x"38",
          3931 => x"fe",
          3932 => x"b4",
          3933 => x"8d",
          3934 => x"ec",
          3935 => x"ff",
          3936 => x"39",
          3937 => x"a4",
          3938 => x"52",
          3939 => x"91",
          3940 => x"ec",
          3941 => x"76",
          3942 => x"fc",
          3943 => x"b4",
          3944 => x"f8",
          3945 => x"ec",
          3946 => x"06",
          3947 => x"81",
          3948 => x"8c",
          3949 => x"3d",
          3950 => x"3d",
          3951 => x"7e",
          3952 => x"82",
          3953 => x"27",
          3954 => x"76",
          3955 => x"27",
          3956 => x"75",
          3957 => x"79",
          3958 => x"38",
          3959 => x"89",
          3960 => x"2e",
          3961 => x"80",
          3962 => x"2e",
          3963 => x"81",
          3964 => x"81",
          3965 => x"89",
          3966 => x"08",
          3967 => x"52",
          3968 => x"3f",
          3969 => x"08",
          3970 => x"ec",
          3971 => x"38",
          3972 => x"06",
          3973 => x"81",
          3974 => x"06",
          3975 => x"77",
          3976 => x"2e",
          3977 => x"84",
          3978 => x"06",
          3979 => x"06",
          3980 => x"53",
          3981 => x"81",
          3982 => x"34",
          3983 => x"a4",
          3984 => x"52",
          3985 => x"d9",
          3986 => x"ec",
          3987 => x"8c",
          3988 => x"94",
          3989 => x"ff",
          3990 => x"05",
          3991 => x"54",
          3992 => x"38",
          3993 => x"74",
          3994 => x"06",
          3995 => x"07",
          3996 => x"74",
          3997 => x"39",
          3998 => x"a4",
          3999 => x"52",
          4000 => x"9d",
          4001 => x"ec",
          4002 => x"8c",
          4003 => x"d8",
          4004 => x"ff",
          4005 => x"76",
          4006 => x"06",
          4007 => x"05",
          4008 => x"3f",
          4009 => x"87",
          4010 => x"08",
          4011 => x"51",
          4012 => x"82",
          4013 => x"59",
          4014 => x"08",
          4015 => x"f0",
          4016 => x"82",
          4017 => x"06",
          4018 => x"05",
          4019 => x"54",
          4020 => x"3f",
          4021 => x"08",
          4022 => x"74",
          4023 => x"51",
          4024 => x"81",
          4025 => x"34",
          4026 => x"ec",
          4027 => x"0d",
          4028 => x"0d",
          4029 => x"72",
          4030 => x"56",
          4031 => x"27",
          4032 => x"98",
          4033 => x"9d",
          4034 => x"2e",
          4035 => x"53",
          4036 => x"51",
          4037 => x"82",
          4038 => x"54",
          4039 => x"08",
          4040 => x"93",
          4041 => x"80",
          4042 => x"54",
          4043 => x"82",
          4044 => x"54",
          4045 => x"74",
          4046 => x"fb",
          4047 => x"8c",
          4048 => x"82",
          4049 => x"80",
          4050 => x"38",
          4051 => x"08",
          4052 => x"38",
          4053 => x"08",
          4054 => x"38",
          4055 => x"52",
          4056 => x"d6",
          4057 => x"ec",
          4058 => x"98",
          4059 => x"11",
          4060 => x"57",
          4061 => x"74",
          4062 => x"81",
          4063 => x"0c",
          4064 => x"81",
          4065 => x"84",
          4066 => x"55",
          4067 => x"ff",
          4068 => x"54",
          4069 => x"ec",
          4070 => x"0d",
          4071 => x"0d",
          4072 => x"08",
          4073 => x"79",
          4074 => x"17",
          4075 => x"80",
          4076 => x"98",
          4077 => x"26",
          4078 => x"58",
          4079 => x"52",
          4080 => x"fd",
          4081 => x"74",
          4082 => x"08",
          4083 => x"38",
          4084 => x"08",
          4085 => x"ec",
          4086 => x"82",
          4087 => x"17",
          4088 => x"ec",
          4089 => x"c7",
          4090 => x"90",
          4091 => x"56",
          4092 => x"2e",
          4093 => x"77",
          4094 => x"81",
          4095 => x"38",
          4096 => x"98",
          4097 => x"26",
          4098 => x"56",
          4099 => x"51",
          4100 => x"80",
          4101 => x"ec",
          4102 => x"09",
          4103 => x"38",
          4104 => x"08",
          4105 => x"ec",
          4106 => x"30",
          4107 => x"80",
          4108 => x"07",
          4109 => x"08",
          4110 => x"55",
          4111 => x"ef",
          4112 => x"ec",
          4113 => x"95",
          4114 => x"08",
          4115 => x"27",
          4116 => x"98",
          4117 => x"89",
          4118 => x"85",
          4119 => x"db",
          4120 => x"81",
          4121 => x"17",
          4122 => x"89",
          4123 => x"75",
          4124 => x"ac",
          4125 => x"7a",
          4126 => x"3f",
          4127 => x"08",
          4128 => x"38",
          4129 => x"8c",
          4130 => x"2e",
          4131 => x"86",
          4132 => x"ec",
          4133 => x"8c",
          4134 => x"70",
          4135 => x"07",
          4136 => x"7c",
          4137 => x"55",
          4138 => x"f8",
          4139 => x"2e",
          4140 => x"ff",
          4141 => x"55",
          4142 => x"ff",
          4143 => x"76",
          4144 => x"3f",
          4145 => x"08",
          4146 => x"08",
          4147 => x"8c",
          4148 => x"80",
          4149 => x"55",
          4150 => x"94",
          4151 => x"2e",
          4152 => x"53",
          4153 => x"51",
          4154 => x"82",
          4155 => x"55",
          4156 => x"75",
          4157 => x"98",
          4158 => x"05",
          4159 => x"56",
          4160 => x"26",
          4161 => x"15",
          4162 => x"84",
          4163 => x"07",
          4164 => x"18",
          4165 => x"ff",
          4166 => x"2e",
          4167 => x"39",
          4168 => x"39",
          4169 => x"08",
          4170 => x"81",
          4171 => x"74",
          4172 => x"0c",
          4173 => x"04",
          4174 => x"7a",
          4175 => x"f3",
          4176 => x"8c",
          4177 => x"81",
          4178 => x"ec",
          4179 => x"38",
          4180 => x"51",
          4181 => x"82",
          4182 => x"82",
          4183 => x"b0",
          4184 => x"84",
          4185 => x"52",
          4186 => x"52",
          4187 => x"3f",
          4188 => x"39",
          4189 => x"8a",
          4190 => x"75",
          4191 => x"38",
          4192 => x"19",
          4193 => x"81",
          4194 => x"ed",
          4195 => x"8c",
          4196 => x"2e",
          4197 => x"15",
          4198 => x"70",
          4199 => x"07",
          4200 => x"53",
          4201 => x"75",
          4202 => x"0c",
          4203 => x"04",
          4204 => x"7a",
          4205 => x"58",
          4206 => x"f0",
          4207 => x"80",
          4208 => x"9f",
          4209 => x"80",
          4210 => x"90",
          4211 => x"17",
          4212 => x"aa",
          4213 => x"53",
          4214 => x"88",
          4215 => x"08",
          4216 => x"38",
          4217 => x"53",
          4218 => x"17",
          4219 => x"72",
          4220 => x"fe",
          4221 => x"08",
          4222 => x"80",
          4223 => x"16",
          4224 => x"2b",
          4225 => x"75",
          4226 => x"73",
          4227 => x"f5",
          4228 => x"8c",
          4229 => x"82",
          4230 => x"ff",
          4231 => x"81",
          4232 => x"ec",
          4233 => x"38",
          4234 => x"82",
          4235 => x"26",
          4236 => x"58",
          4237 => x"73",
          4238 => x"39",
          4239 => x"51",
          4240 => x"82",
          4241 => x"98",
          4242 => x"94",
          4243 => x"17",
          4244 => x"58",
          4245 => x"9a",
          4246 => x"81",
          4247 => x"74",
          4248 => x"98",
          4249 => x"83",
          4250 => x"b4",
          4251 => x"0c",
          4252 => x"82",
          4253 => x"8a",
          4254 => x"f8",
          4255 => x"70",
          4256 => x"08",
          4257 => x"57",
          4258 => x"0a",
          4259 => x"38",
          4260 => x"15",
          4261 => x"08",
          4262 => x"72",
          4263 => x"cb",
          4264 => x"ff",
          4265 => x"81",
          4266 => x"13",
          4267 => x"94",
          4268 => x"74",
          4269 => x"85",
          4270 => x"22",
          4271 => x"73",
          4272 => x"38",
          4273 => x"8a",
          4274 => x"05",
          4275 => x"06",
          4276 => x"8a",
          4277 => x"73",
          4278 => x"3f",
          4279 => x"08",
          4280 => x"81",
          4281 => x"ec",
          4282 => x"ff",
          4283 => x"82",
          4284 => x"ff",
          4285 => x"38",
          4286 => x"82",
          4287 => x"26",
          4288 => x"7b",
          4289 => x"98",
          4290 => x"55",
          4291 => x"94",
          4292 => x"73",
          4293 => x"3f",
          4294 => x"08",
          4295 => x"82",
          4296 => x"80",
          4297 => x"38",
          4298 => x"8c",
          4299 => x"2e",
          4300 => x"55",
          4301 => x"08",
          4302 => x"38",
          4303 => x"08",
          4304 => x"fb",
          4305 => x"8c",
          4306 => x"38",
          4307 => x"0c",
          4308 => x"51",
          4309 => x"82",
          4310 => x"98",
          4311 => x"90",
          4312 => x"16",
          4313 => x"15",
          4314 => x"74",
          4315 => x"0c",
          4316 => x"04",
          4317 => x"7b",
          4318 => x"5b",
          4319 => x"52",
          4320 => x"ac",
          4321 => x"ec",
          4322 => x"8c",
          4323 => x"ec",
          4324 => x"ec",
          4325 => x"17",
          4326 => x"51",
          4327 => x"82",
          4328 => x"54",
          4329 => x"08",
          4330 => x"82",
          4331 => x"9c",
          4332 => x"33",
          4333 => x"72",
          4334 => x"09",
          4335 => x"38",
          4336 => x"8c",
          4337 => x"72",
          4338 => x"55",
          4339 => x"53",
          4340 => x"8e",
          4341 => x"56",
          4342 => x"09",
          4343 => x"38",
          4344 => x"8c",
          4345 => x"81",
          4346 => x"fd",
          4347 => x"8c",
          4348 => x"82",
          4349 => x"80",
          4350 => x"38",
          4351 => x"09",
          4352 => x"38",
          4353 => x"82",
          4354 => x"8b",
          4355 => x"fd",
          4356 => x"9a",
          4357 => x"eb",
          4358 => x"8c",
          4359 => x"ff",
          4360 => x"70",
          4361 => x"53",
          4362 => x"09",
          4363 => x"38",
          4364 => x"eb",
          4365 => x"8c",
          4366 => x"2b",
          4367 => x"72",
          4368 => x"0c",
          4369 => x"04",
          4370 => x"77",
          4371 => x"ff",
          4372 => x"9a",
          4373 => x"55",
          4374 => x"76",
          4375 => x"53",
          4376 => x"09",
          4377 => x"38",
          4378 => x"52",
          4379 => x"eb",
          4380 => x"3d",
          4381 => x"3d",
          4382 => x"5b",
          4383 => x"08",
          4384 => x"15",
          4385 => x"81",
          4386 => x"15",
          4387 => x"51",
          4388 => x"82",
          4389 => x"58",
          4390 => x"08",
          4391 => x"9c",
          4392 => x"33",
          4393 => x"86",
          4394 => x"80",
          4395 => x"13",
          4396 => x"06",
          4397 => x"06",
          4398 => x"72",
          4399 => x"82",
          4400 => x"53",
          4401 => x"2e",
          4402 => x"53",
          4403 => x"a9",
          4404 => x"74",
          4405 => x"72",
          4406 => x"38",
          4407 => x"99",
          4408 => x"ec",
          4409 => x"06",
          4410 => x"88",
          4411 => x"06",
          4412 => x"54",
          4413 => x"a0",
          4414 => x"74",
          4415 => x"3f",
          4416 => x"08",
          4417 => x"ec",
          4418 => x"98",
          4419 => x"fa",
          4420 => x"80",
          4421 => x"0c",
          4422 => x"ec",
          4423 => x"0d",
          4424 => x"0d",
          4425 => x"57",
          4426 => x"73",
          4427 => x"3f",
          4428 => x"08",
          4429 => x"ec",
          4430 => x"98",
          4431 => x"75",
          4432 => x"3f",
          4433 => x"08",
          4434 => x"ec",
          4435 => x"a0",
          4436 => x"ec",
          4437 => x"14",
          4438 => x"db",
          4439 => x"a0",
          4440 => x"14",
          4441 => x"ac",
          4442 => x"83",
          4443 => x"82",
          4444 => x"87",
          4445 => x"fd",
          4446 => x"70",
          4447 => x"08",
          4448 => x"55",
          4449 => x"3f",
          4450 => x"08",
          4451 => x"13",
          4452 => x"73",
          4453 => x"83",
          4454 => x"3d",
          4455 => x"3d",
          4456 => x"57",
          4457 => x"89",
          4458 => x"17",
          4459 => x"81",
          4460 => x"70",
          4461 => x"55",
          4462 => x"08",
          4463 => x"81",
          4464 => x"52",
          4465 => x"a8",
          4466 => x"2e",
          4467 => x"84",
          4468 => x"52",
          4469 => x"09",
          4470 => x"38",
          4471 => x"81",
          4472 => x"81",
          4473 => x"73",
          4474 => x"55",
          4475 => x"55",
          4476 => x"c5",
          4477 => x"88",
          4478 => x"0b",
          4479 => x"9c",
          4480 => x"8b",
          4481 => x"17",
          4482 => x"08",
          4483 => x"52",
          4484 => x"82",
          4485 => x"76",
          4486 => x"51",
          4487 => x"82",
          4488 => x"86",
          4489 => x"12",
          4490 => x"3f",
          4491 => x"08",
          4492 => x"88",
          4493 => x"f3",
          4494 => x"70",
          4495 => x"80",
          4496 => x"51",
          4497 => x"af",
          4498 => x"81",
          4499 => x"dc",
          4500 => x"74",
          4501 => x"38",
          4502 => x"88",
          4503 => x"39",
          4504 => x"80",
          4505 => x"56",
          4506 => x"af",
          4507 => x"06",
          4508 => x"56",
          4509 => x"32",
          4510 => x"80",
          4511 => x"51",
          4512 => x"dc",
          4513 => x"1c",
          4514 => x"33",
          4515 => x"9f",
          4516 => x"ff",
          4517 => x"1c",
          4518 => x"7a",
          4519 => x"3f",
          4520 => x"08",
          4521 => x"39",
          4522 => x"a0",
          4523 => x"5e",
          4524 => x"52",
          4525 => x"ff",
          4526 => x"59",
          4527 => x"33",
          4528 => x"ae",
          4529 => x"06",
          4530 => x"78",
          4531 => x"81",
          4532 => x"32",
          4533 => x"9f",
          4534 => x"26",
          4535 => x"53",
          4536 => x"73",
          4537 => x"17",
          4538 => x"34",
          4539 => x"db",
          4540 => x"32",
          4541 => x"9f",
          4542 => x"54",
          4543 => x"2e",
          4544 => x"80",
          4545 => x"75",
          4546 => x"bd",
          4547 => x"7e",
          4548 => x"a0",
          4549 => x"bd",
          4550 => x"82",
          4551 => x"18",
          4552 => x"1a",
          4553 => x"a0",
          4554 => x"fc",
          4555 => x"32",
          4556 => x"80",
          4557 => x"30",
          4558 => x"71",
          4559 => x"51",
          4560 => x"55",
          4561 => x"ac",
          4562 => x"81",
          4563 => x"78",
          4564 => x"51",
          4565 => x"af",
          4566 => x"06",
          4567 => x"55",
          4568 => x"32",
          4569 => x"80",
          4570 => x"51",
          4571 => x"db",
          4572 => x"39",
          4573 => x"09",
          4574 => x"38",
          4575 => x"7c",
          4576 => x"54",
          4577 => x"a2",
          4578 => x"32",
          4579 => x"ae",
          4580 => x"72",
          4581 => x"9f",
          4582 => x"51",
          4583 => x"74",
          4584 => x"88",
          4585 => x"fe",
          4586 => x"98",
          4587 => x"80",
          4588 => x"75",
          4589 => x"81",
          4590 => x"33",
          4591 => x"51",
          4592 => x"82",
          4593 => x"80",
          4594 => x"78",
          4595 => x"81",
          4596 => x"5a",
          4597 => x"d2",
          4598 => x"ec",
          4599 => x"80",
          4600 => x"1c",
          4601 => x"27",
          4602 => x"79",
          4603 => x"74",
          4604 => x"7a",
          4605 => x"74",
          4606 => x"39",
          4607 => x"fb",
          4608 => x"fe",
          4609 => x"ec",
          4610 => x"ff",
          4611 => x"73",
          4612 => x"38",
          4613 => x"81",
          4614 => x"54",
          4615 => x"75",
          4616 => x"17",
          4617 => x"39",
          4618 => x"0c",
          4619 => x"99",
          4620 => x"54",
          4621 => x"2e",
          4622 => x"84",
          4623 => x"34",
          4624 => x"76",
          4625 => x"8b",
          4626 => x"81",
          4627 => x"56",
          4628 => x"80",
          4629 => x"1b",
          4630 => x"08",
          4631 => x"51",
          4632 => x"82",
          4633 => x"56",
          4634 => x"08",
          4635 => x"98",
          4636 => x"76",
          4637 => x"3f",
          4638 => x"08",
          4639 => x"ec",
          4640 => x"38",
          4641 => x"70",
          4642 => x"73",
          4643 => x"be",
          4644 => x"33",
          4645 => x"73",
          4646 => x"8b",
          4647 => x"83",
          4648 => x"06",
          4649 => x"73",
          4650 => x"53",
          4651 => x"51",
          4652 => x"82",
          4653 => x"80",
          4654 => x"75",
          4655 => x"f3",
          4656 => x"9f",
          4657 => x"1c",
          4658 => x"74",
          4659 => x"38",
          4660 => x"09",
          4661 => x"e7",
          4662 => x"2a",
          4663 => x"77",
          4664 => x"51",
          4665 => x"2e",
          4666 => x"81",
          4667 => x"80",
          4668 => x"38",
          4669 => x"ab",
          4670 => x"55",
          4671 => x"75",
          4672 => x"73",
          4673 => x"55",
          4674 => x"82",
          4675 => x"06",
          4676 => x"ab",
          4677 => x"33",
          4678 => x"70",
          4679 => x"55",
          4680 => x"2e",
          4681 => x"1b",
          4682 => x"06",
          4683 => x"52",
          4684 => x"db",
          4685 => x"ec",
          4686 => x"0c",
          4687 => x"74",
          4688 => x"0c",
          4689 => x"04",
          4690 => x"7c",
          4691 => x"08",
          4692 => x"55",
          4693 => x"59",
          4694 => x"81",
          4695 => x"70",
          4696 => x"33",
          4697 => x"52",
          4698 => x"2e",
          4699 => x"ee",
          4700 => x"2e",
          4701 => x"81",
          4702 => x"33",
          4703 => x"81",
          4704 => x"52",
          4705 => x"26",
          4706 => x"14",
          4707 => x"06",
          4708 => x"52",
          4709 => x"80",
          4710 => x"0b",
          4711 => x"59",
          4712 => x"7a",
          4713 => x"70",
          4714 => x"33",
          4715 => x"05",
          4716 => x"9f",
          4717 => x"53",
          4718 => x"89",
          4719 => x"70",
          4720 => x"54",
          4721 => x"12",
          4722 => x"26",
          4723 => x"12",
          4724 => x"06",
          4725 => x"30",
          4726 => x"51",
          4727 => x"2e",
          4728 => x"85",
          4729 => x"be",
          4730 => x"74",
          4731 => x"30",
          4732 => x"9f",
          4733 => x"2a",
          4734 => x"54",
          4735 => x"2e",
          4736 => x"15",
          4737 => x"55",
          4738 => x"ff",
          4739 => x"39",
          4740 => x"86",
          4741 => x"7c",
          4742 => x"51",
          4743 => x"8d",
          4744 => x"70",
          4745 => x"0c",
          4746 => x"04",
          4747 => x"78",
          4748 => x"83",
          4749 => x"0b",
          4750 => x"79",
          4751 => x"e2",
          4752 => x"55",
          4753 => x"08",
          4754 => x"84",
          4755 => x"df",
          4756 => x"8c",
          4757 => x"ff",
          4758 => x"83",
          4759 => x"d4",
          4760 => x"81",
          4761 => x"38",
          4762 => x"17",
          4763 => x"74",
          4764 => x"09",
          4765 => x"38",
          4766 => x"81",
          4767 => x"30",
          4768 => x"79",
          4769 => x"54",
          4770 => x"74",
          4771 => x"09",
          4772 => x"38",
          4773 => x"fb",
          4774 => x"ea",
          4775 => x"b1",
          4776 => x"ec",
          4777 => x"8c",
          4778 => x"2e",
          4779 => x"53",
          4780 => x"52",
          4781 => x"51",
          4782 => x"82",
          4783 => x"55",
          4784 => x"08",
          4785 => x"38",
          4786 => x"82",
          4787 => x"88",
          4788 => x"f2",
          4789 => x"02",
          4790 => x"cb",
          4791 => x"55",
          4792 => x"60",
          4793 => x"3f",
          4794 => x"08",
          4795 => x"80",
          4796 => x"ec",
          4797 => x"fc",
          4798 => x"ec",
          4799 => x"82",
          4800 => x"70",
          4801 => x"8c",
          4802 => x"2e",
          4803 => x"73",
          4804 => x"81",
          4805 => x"33",
          4806 => x"80",
          4807 => x"81",
          4808 => x"d7",
          4809 => x"8c",
          4810 => x"ff",
          4811 => x"06",
          4812 => x"98",
          4813 => x"2e",
          4814 => x"74",
          4815 => x"81",
          4816 => x"8a",
          4817 => x"ac",
          4818 => x"39",
          4819 => x"77",
          4820 => x"81",
          4821 => x"33",
          4822 => x"3f",
          4823 => x"08",
          4824 => x"70",
          4825 => x"55",
          4826 => x"86",
          4827 => x"80",
          4828 => x"74",
          4829 => x"81",
          4830 => x"8a",
          4831 => x"f4",
          4832 => x"53",
          4833 => x"fd",
          4834 => x"8c",
          4835 => x"ff",
          4836 => x"82",
          4837 => x"06",
          4838 => x"8c",
          4839 => x"58",
          4840 => x"f6",
          4841 => x"58",
          4842 => x"2e",
          4843 => x"fa",
          4844 => x"e8",
          4845 => x"ec",
          4846 => x"78",
          4847 => x"5a",
          4848 => x"90",
          4849 => x"75",
          4850 => x"38",
          4851 => x"3d",
          4852 => x"70",
          4853 => x"08",
          4854 => x"7a",
          4855 => x"38",
          4856 => x"51",
          4857 => x"82",
          4858 => x"81",
          4859 => x"81",
          4860 => x"38",
          4861 => x"83",
          4862 => x"38",
          4863 => x"84",
          4864 => x"38",
          4865 => x"81",
          4866 => x"38",
          4867 => x"db",
          4868 => x"8c",
          4869 => x"ff",
          4870 => x"72",
          4871 => x"09",
          4872 => x"d0",
          4873 => x"14",
          4874 => x"3f",
          4875 => x"08",
          4876 => x"06",
          4877 => x"38",
          4878 => x"51",
          4879 => x"82",
          4880 => x"58",
          4881 => x"0c",
          4882 => x"33",
          4883 => x"80",
          4884 => x"ff",
          4885 => x"ff",
          4886 => x"55",
          4887 => x"81",
          4888 => x"38",
          4889 => x"06",
          4890 => x"80",
          4891 => x"52",
          4892 => x"8a",
          4893 => x"80",
          4894 => x"ff",
          4895 => x"53",
          4896 => x"86",
          4897 => x"83",
          4898 => x"c5",
          4899 => x"f5",
          4900 => x"ec",
          4901 => x"8c",
          4902 => x"15",
          4903 => x"06",
          4904 => x"76",
          4905 => x"80",
          4906 => x"da",
          4907 => x"8c",
          4908 => x"ff",
          4909 => x"74",
          4910 => x"d4",
          4911 => x"dc",
          4912 => x"ec",
          4913 => x"c2",
          4914 => x"b9",
          4915 => x"ec",
          4916 => x"ff",
          4917 => x"56",
          4918 => x"83",
          4919 => x"14",
          4920 => x"71",
          4921 => x"5a",
          4922 => x"26",
          4923 => x"8a",
          4924 => x"74",
          4925 => x"ff",
          4926 => x"82",
          4927 => x"55",
          4928 => x"08",
          4929 => x"ec",
          4930 => x"ec",
          4931 => x"ff",
          4932 => x"83",
          4933 => x"74",
          4934 => x"26",
          4935 => x"57",
          4936 => x"26",
          4937 => x"57",
          4938 => x"56",
          4939 => x"82",
          4940 => x"15",
          4941 => x"0c",
          4942 => x"0c",
          4943 => x"a4",
          4944 => x"1d",
          4945 => x"54",
          4946 => x"2e",
          4947 => x"af",
          4948 => x"14",
          4949 => x"3f",
          4950 => x"08",
          4951 => x"06",
          4952 => x"72",
          4953 => x"79",
          4954 => x"80",
          4955 => x"d9",
          4956 => x"8c",
          4957 => x"15",
          4958 => x"2b",
          4959 => x"8d",
          4960 => x"2e",
          4961 => x"77",
          4962 => x"0c",
          4963 => x"76",
          4964 => x"38",
          4965 => x"70",
          4966 => x"81",
          4967 => x"53",
          4968 => x"89",
          4969 => x"56",
          4970 => x"08",
          4971 => x"38",
          4972 => x"15",
          4973 => x"8c",
          4974 => x"80",
          4975 => x"34",
          4976 => x"09",
          4977 => x"92",
          4978 => x"14",
          4979 => x"3f",
          4980 => x"08",
          4981 => x"06",
          4982 => x"2e",
          4983 => x"80",
          4984 => x"1b",
          4985 => x"db",
          4986 => x"8c",
          4987 => x"ea",
          4988 => x"ec",
          4989 => x"34",
          4990 => x"51",
          4991 => x"82",
          4992 => x"83",
          4993 => x"53",
          4994 => x"d5",
          4995 => x"06",
          4996 => x"b4",
          4997 => x"84",
          4998 => x"ec",
          4999 => x"85",
          5000 => x"09",
          5001 => x"38",
          5002 => x"51",
          5003 => x"82",
          5004 => x"86",
          5005 => x"f2",
          5006 => x"06",
          5007 => x"9c",
          5008 => x"d8",
          5009 => x"ec",
          5010 => x"0c",
          5011 => x"51",
          5012 => x"82",
          5013 => x"8c",
          5014 => x"74",
          5015 => x"98",
          5016 => x"53",
          5017 => x"98",
          5018 => x"15",
          5019 => x"94",
          5020 => x"56",
          5021 => x"ec",
          5022 => x"0d",
          5023 => x"0d",
          5024 => x"55",
          5025 => x"b9",
          5026 => x"53",
          5027 => x"b1",
          5028 => x"52",
          5029 => x"a9",
          5030 => x"22",
          5031 => x"57",
          5032 => x"2e",
          5033 => x"99",
          5034 => x"33",
          5035 => x"3f",
          5036 => x"08",
          5037 => x"71",
          5038 => x"74",
          5039 => x"83",
          5040 => x"78",
          5041 => x"52",
          5042 => x"ec",
          5043 => x"0d",
          5044 => x"0d",
          5045 => x"33",
          5046 => x"3d",
          5047 => x"56",
          5048 => x"8b",
          5049 => x"82",
          5050 => x"24",
          5051 => x"8c",
          5052 => x"29",
          5053 => x"05",
          5054 => x"55",
          5055 => x"84",
          5056 => x"34",
          5057 => x"80",
          5058 => x"80",
          5059 => x"75",
          5060 => x"75",
          5061 => x"38",
          5062 => x"3d",
          5063 => x"05",
          5064 => x"3f",
          5065 => x"08",
          5066 => x"8c",
          5067 => x"3d",
          5068 => x"3d",
          5069 => x"84",
          5070 => x"05",
          5071 => x"89",
          5072 => x"2e",
          5073 => x"77",
          5074 => x"54",
          5075 => x"05",
          5076 => x"84",
          5077 => x"f6",
          5078 => x"8c",
          5079 => x"82",
          5080 => x"84",
          5081 => x"5c",
          5082 => x"3d",
          5083 => x"ed",
          5084 => x"8c",
          5085 => x"82",
          5086 => x"92",
          5087 => x"d7",
          5088 => x"98",
          5089 => x"73",
          5090 => x"38",
          5091 => x"9c",
          5092 => x"80",
          5093 => x"38",
          5094 => x"95",
          5095 => x"2e",
          5096 => x"aa",
          5097 => x"ea",
          5098 => x"8c",
          5099 => x"9e",
          5100 => x"05",
          5101 => x"54",
          5102 => x"38",
          5103 => x"70",
          5104 => x"54",
          5105 => x"8e",
          5106 => x"83",
          5107 => x"88",
          5108 => x"83",
          5109 => x"83",
          5110 => x"06",
          5111 => x"80",
          5112 => x"38",
          5113 => x"51",
          5114 => x"82",
          5115 => x"56",
          5116 => x"0a",
          5117 => x"05",
          5118 => x"3f",
          5119 => x"0b",
          5120 => x"80",
          5121 => x"7a",
          5122 => x"3f",
          5123 => x"9c",
          5124 => x"d1",
          5125 => x"81",
          5126 => x"34",
          5127 => x"80",
          5128 => x"b0",
          5129 => x"54",
          5130 => x"52",
          5131 => x"05",
          5132 => x"3f",
          5133 => x"08",
          5134 => x"ec",
          5135 => x"38",
          5136 => x"82",
          5137 => x"b2",
          5138 => x"84",
          5139 => x"06",
          5140 => x"73",
          5141 => x"38",
          5142 => x"ad",
          5143 => x"2a",
          5144 => x"51",
          5145 => x"2e",
          5146 => x"81",
          5147 => x"80",
          5148 => x"87",
          5149 => x"39",
          5150 => x"51",
          5151 => x"82",
          5152 => x"7b",
          5153 => x"12",
          5154 => x"82",
          5155 => x"81",
          5156 => x"83",
          5157 => x"06",
          5158 => x"80",
          5159 => x"77",
          5160 => x"58",
          5161 => x"08",
          5162 => x"63",
          5163 => x"63",
          5164 => x"57",
          5165 => x"82",
          5166 => x"82",
          5167 => x"88",
          5168 => x"9c",
          5169 => x"d2",
          5170 => x"8c",
          5171 => x"8c",
          5172 => x"1b",
          5173 => x"0c",
          5174 => x"22",
          5175 => x"77",
          5176 => x"80",
          5177 => x"34",
          5178 => x"1a",
          5179 => x"94",
          5180 => x"85",
          5181 => x"06",
          5182 => x"80",
          5183 => x"38",
          5184 => x"08",
          5185 => x"84",
          5186 => x"ec",
          5187 => x"0c",
          5188 => x"70",
          5189 => x"52",
          5190 => x"39",
          5191 => x"51",
          5192 => x"82",
          5193 => x"57",
          5194 => x"08",
          5195 => x"38",
          5196 => x"8c",
          5197 => x"2e",
          5198 => x"83",
          5199 => x"75",
          5200 => x"74",
          5201 => x"07",
          5202 => x"54",
          5203 => x"8a",
          5204 => x"75",
          5205 => x"73",
          5206 => x"98",
          5207 => x"a9",
          5208 => x"ff",
          5209 => x"80",
          5210 => x"76",
          5211 => x"d6",
          5212 => x"8c",
          5213 => x"38",
          5214 => x"39",
          5215 => x"82",
          5216 => x"05",
          5217 => x"84",
          5218 => x"0c",
          5219 => x"82",
          5220 => x"97",
          5221 => x"f2",
          5222 => x"63",
          5223 => x"40",
          5224 => x"7e",
          5225 => x"fc",
          5226 => x"51",
          5227 => x"82",
          5228 => x"55",
          5229 => x"08",
          5230 => x"19",
          5231 => x"80",
          5232 => x"74",
          5233 => x"39",
          5234 => x"81",
          5235 => x"56",
          5236 => x"82",
          5237 => x"39",
          5238 => x"1a",
          5239 => x"82",
          5240 => x"0b",
          5241 => x"81",
          5242 => x"39",
          5243 => x"94",
          5244 => x"55",
          5245 => x"83",
          5246 => x"7b",
          5247 => x"89",
          5248 => x"08",
          5249 => x"06",
          5250 => x"81",
          5251 => x"8a",
          5252 => x"05",
          5253 => x"06",
          5254 => x"a8",
          5255 => x"38",
          5256 => x"55",
          5257 => x"19",
          5258 => x"51",
          5259 => x"82",
          5260 => x"55",
          5261 => x"ff",
          5262 => x"ff",
          5263 => x"38",
          5264 => x"0c",
          5265 => x"52",
          5266 => x"cb",
          5267 => x"ec",
          5268 => x"ff",
          5269 => x"8c",
          5270 => x"7c",
          5271 => x"57",
          5272 => x"80",
          5273 => x"1a",
          5274 => x"22",
          5275 => x"75",
          5276 => x"38",
          5277 => x"58",
          5278 => x"53",
          5279 => x"1b",
          5280 => x"88",
          5281 => x"ec",
          5282 => x"38",
          5283 => x"33",
          5284 => x"80",
          5285 => x"b0",
          5286 => x"31",
          5287 => x"27",
          5288 => x"80",
          5289 => x"52",
          5290 => x"77",
          5291 => x"7d",
          5292 => x"e0",
          5293 => x"2b",
          5294 => x"76",
          5295 => x"94",
          5296 => x"ff",
          5297 => x"71",
          5298 => x"7b",
          5299 => x"38",
          5300 => x"19",
          5301 => x"51",
          5302 => x"82",
          5303 => x"fe",
          5304 => x"53",
          5305 => x"83",
          5306 => x"b4",
          5307 => x"51",
          5308 => x"7b",
          5309 => x"08",
          5310 => x"76",
          5311 => x"08",
          5312 => x"0c",
          5313 => x"f3",
          5314 => x"75",
          5315 => x"0c",
          5316 => x"04",
          5317 => x"60",
          5318 => x"40",
          5319 => x"80",
          5320 => x"3d",
          5321 => x"77",
          5322 => x"3f",
          5323 => x"08",
          5324 => x"ec",
          5325 => x"91",
          5326 => x"74",
          5327 => x"38",
          5328 => x"b8",
          5329 => x"33",
          5330 => x"70",
          5331 => x"56",
          5332 => x"74",
          5333 => x"a4",
          5334 => x"82",
          5335 => x"34",
          5336 => x"98",
          5337 => x"91",
          5338 => x"56",
          5339 => x"94",
          5340 => x"11",
          5341 => x"76",
          5342 => x"75",
          5343 => x"80",
          5344 => x"38",
          5345 => x"70",
          5346 => x"56",
          5347 => x"fd",
          5348 => x"11",
          5349 => x"77",
          5350 => x"5c",
          5351 => x"38",
          5352 => x"88",
          5353 => x"74",
          5354 => x"52",
          5355 => x"18",
          5356 => x"51",
          5357 => x"82",
          5358 => x"55",
          5359 => x"08",
          5360 => x"ab",
          5361 => x"2e",
          5362 => x"74",
          5363 => x"95",
          5364 => x"19",
          5365 => x"08",
          5366 => x"88",
          5367 => x"55",
          5368 => x"9c",
          5369 => x"09",
          5370 => x"38",
          5371 => x"c1",
          5372 => x"ec",
          5373 => x"38",
          5374 => x"52",
          5375 => x"97",
          5376 => x"ec",
          5377 => x"fe",
          5378 => x"8c",
          5379 => x"7c",
          5380 => x"57",
          5381 => x"80",
          5382 => x"1b",
          5383 => x"22",
          5384 => x"75",
          5385 => x"38",
          5386 => x"59",
          5387 => x"53",
          5388 => x"1a",
          5389 => x"be",
          5390 => x"ec",
          5391 => x"38",
          5392 => x"08",
          5393 => x"56",
          5394 => x"9b",
          5395 => x"53",
          5396 => x"77",
          5397 => x"7d",
          5398 => x"16",
          5399 => x"3f",
          5400 => x"0b",
          5401 => x"78",
          5402 => x"80",
          5403 => x"18",
          5404 => x"08",
          5405 => x"7e",
          5406 => x"3f",
          5407 => x"08",
          5408 => x"7e",
          5409 => x"0c",
          5410 => x"19",
          5411 => x"08",
          5412 => x"84",
          5413 => x"57",
          5414 => x"27",
          5415 => x"56",
          5416 => x"52",
          5417 => x"f9",
          5418 => x"ec",
          5419 => x"38",
          5420 => x"52",
          5421 => x"83",
          5422 => x"b4",
          5423 => x"d4",
          5424 => x"81",
          5425 => x"34",
          5426 => x"7e",
          5427 => x"0c",
          5428 => x"1a",
          5429 => x"94",
          5430 => x"1b",
          5431 => x"5e",
          5432 => x"27",
          5433 => x"55",
          5434 => x"0c",
          5435 => x"90",
          5436 => x"c0",
          5437 => x"90",
          5438 => x"56",
          5439 => x"ec",
          5440 => x"0d",
          5441 => x"0d",
          5442 => x"fc",
          5443 => x"52",
          5444 => x"3f",
          5445 => x"08",
          5446 => x"ec",
          5447 => x"38",
          5448 => x"70",
          5449 => x"81",
          5450 => x"55",
          5451 => x"80",
          5452 => x"16",
          5453 => x"51",
          5454 => x"82",
          5455 => x"57",
          5456 => x"08",
          5457 => x"a4",
          5458 => x"11",
          5459 => x"55",
          5460 => x"16",
          5461 => x"08",
          5462 => x"75",
          5463 => x"e8",
          5464 => x"08",
          5465 => x"51",
          5466 => x"82",
          5467 => x"52",
          5468 => x"c9",
          5469 => x"52",
          5470 => x"c9",
          5471 => x"54",
          5472 => x"15",
          5473 => x"cc",
          5474 => x"8c",
          5475 => x"17",
          5476 => x"06",
          5477 => x"90",
          5478 => x"82",
          5479 => x"8a",
          5480 => x"fc",
          5481 => x"70",
          5482 => x"d9",
          5483 => x"ec",
          5484 => x"8c",
          5485 => x"38",
          5486 => x"05",
          5487 => x"f1",
          5488 => x"8c",
          5489 => x"82",
          5490 => x"87",
          5491 => x"ec",
          5492 => x"72",
          5493 => x"0c",
          5494 => x"04",
          5495 => x"84",
          5496 => x"e4",
          5497 => x"80",
          5498 => x"ec",
          5499 => x"38",
          5500 => x"08",
          5501 => x"34",
          5502 => x"82",
          5503 => x"83",
          5504 => x"ef",
          5505 => x"53",
          5506 => x"05",
          5507 => x"51",
          5508 => x"82",
          5509 => x"55",
          5510 => x"08",
          5511 => x"76",
          5512 => x"93",
          5513 => x"51",
          5514 => x"82",
          5515 => x"55",
          5516 => x"08",
          5517 => x"80",
          5518 => x"70",
          5519 => x"56",
          5520 => x"89",
          5521 => x"94",
          5522 => x"b2",
          5523 => x"05",
          5524 => x"2a",
          5525 => x"51",
          5526 => x"80",
          5527 => x"76",
          5528 => x"52",
          5529 => x"3f",
          5530 => x"08",
          5531 => x"8e",
          5532 => x"ec",
          5533 => x"09",
          5534 => x"38",
          5535 => x"82",
          5536 => x"93",
          5537 => x"e4",
          5538 => x"6f",
          5539 => x"7a",
          5540 => x"9e",
          5541 => x"05",
          5542 => x"51",
          5543 => x"82",
          5544 => x"57",
          5545 => x"08",
          5546 => x"7b",
          5547 => x"94",
          5548 => x"55",
          5549 => x"73",
          5550 => x"ed",
          5551 => x"93",
          5552 => x"55",
          5553 => x"82",
          5554 => x"57",
          5555 => x"08",
          5556 => x"68",
          5557 => x"c9",
          5558 => x"8c",
          5559 => x"82",
          5560 => x"82",
          5561 => x"52",
          5562 => x"a3",
          5563 => x"ec",
          5564 => x"52",
          5565 => x"b8",
          5566 => x"ec",
          5567 => x"8c",
          5568 => x"a2",
          5569 => x"74",
          5570 => x"3f",
          5571 => x"08",
          5572 => x"ec",
          5573 => x"69",
          5574 => x"d9",
          5575 => x"82",
          5576 => x"2e",
          5577 => x"52",
          5578 => x"cf",
          5579 => x"ec",
          5580 => x"8c",
          5581 => x"2e",
          5582 => x"84",
          5583 => x"06",
          5584 => x"57",
          5585 => x"76",
          5586 => x"9e",
          5587 => x"05",
          5588 => x"dc",
          5589 => x"90",
          5590 => x"81",
          5591 => x"56",
          5592 => x"80",
          5593 => x"02",
          5594 => x"81",
          5595 => x"70",
          5596 => x"56",
          5597 => x"81",
          5598 => x"78",
          5599 => x"38",
          5600 => x"99",
          5601 => x"81",
          5602 => x"18",
          5603 => x"18",
          5604 => x"58",
          5605 => x"33",
          5606 => x"ee",
          5607 => x"6f",
          5608 => x"af",
          5609 => x"8d",
          5610 => x"2e",
          5611 => x"8a",
          5612 => x"6f",
          5613 => x"af",
          5614 => x"0b",
          5615 => x"33",
          5616 => x"81",
          5617 => x"70",
          5618 => x"52",
          5619 => x"56",
          5620 => x"8d",
          5621 => x"70",
          5622 => x"51",
          5623 => x"f5",
          5624 => x"54",
          5625 => x"a7",
          5626 => x"74",
          5627 => x"38",
          5628 => x"73",
          5629 => x"81",
          5630 => x"81",
          5631 => x"39",
          5632 => x"81",
          5633 => x"74",
          5634 => x"81",
          5635 => x"91",
          5636 => x"6e",
          5637 => x"59",
          5638 => x"7a",
          5639 => x"5c",
          5640 => x"26",
          5641 => x"7a",
          5642 => x"8c",
          5643 => x"3d",
          5644 => x"3d",
          5645 => x"8d",
          5646 => x"54",
          5647 => x"55",
          5648 => x"82",
          5649 => x"53",
          5650 => x"08",
          5651 => x"91",
          5652 => x"72",
          5653 => x"8c",
          5654 => x"73",
          5655 => x"38",
          5656 => x"70",
          5657 => x"81",
          5658 => x"57",
          5659 => x"73",
          5660 => x"08",
          5661 => x"94",
          5662 => x"75",
          5663 => x"97",
          5664 => x"11",
          5665 => x"2b",
          5666 => x"73",
          5667 => x"38",
          5668 => x"16",
          5669 => x"a0",
          5670 => x"ec",
          5671 => x"78",
          5672 => x"55",
          5673 => x"90",
          5674 => x"ec",
          5675 => x"96",
          5676 => x"70",
          5677 => x"94",
          5678 => x"71",
          5679 => x"08",
          5680 => x"53",
          5681 => x"15",
          5682 => x"a6",
          5683 => x"74",
          5684 => x"3f",
          5685 => x"08",
          5686 => x"ec",
          5687 => x"81",
          5688 => x"8c",
          5689 => x"2e",
          5690 => x"82",
          5691 => x"88",
          5692 => x"98",
          5693 => x"80",
          5694 => x"38",
          5695 => x"80",
          5696 => x"77",
          5697 => x"08",
          5698 => x"0c",
          5699 => x"70",
          5700 => x"81",
          5701 => x"5a",
          5702 => x"2e",
          5703 => x"52",
          5704 => x"f9",
          5705 => x"ec",
          5706 => x"8c",
          5707 => x"38",
          5708 => x"08",
          5709 => x"73",
          5710 => x"c7",
          5711 => x"8c",
          5712 => x"73",
          5713 => x"38",
          5714 => x"af",
          5715 => x"73",
          5716 => x"27",
          5717 => x"98",
          5718 => x"a0",
          5719 => x"08",
          5720 => x"0c",
          5721 => x"06",
          5722 => x"2e",
          5723 => x"52",
          5724 => x"a3",
          5725 => x"ec",
          5726 => x"82",
          5727 => x"34",
          5728 => x"c4",
          5729 => x"91",
          5730 => x"53",
          5731 => x"89",
          5732 => x"ec",
          5733 => x"94",
          5734 => x"8c",
          5735 => x"27",
          5736 => x"8c",
          5737 => x"15",
          5738 => x"07",
          5739 => x"16",
          5740 => x"ff",
          5741 => x"80",
          5742 => x"77",
          5743 => x"2e",
          5744 => x"9c",
          5745 => x"53",
          5746 => x"ec",
          5747 => x"0d",
          5748 => x"0d",
          5749 => x"54",
          5750 => x"81",
          5751 => x"53",
          5752 => x"05",
          5753 => x"84",
          5754 => x"e7",
          5755 => x"ec",
          5756 => x"8c",
          5757 => x"ea",
          5758 => x"0c",
          5759 => x"51",
          5760 => x"82",
          5761 => x"55",
          5762 => x"08",
          5763 => x"ab",
          5764 => x"98",
          5765 => x"80",
          5766 => x"38",
          5767 => x"70",
          5768 => x"81",
          5769 => x"57",
          5770 => x"ad",
          5771 => x"08",
          5772 => x"d3",
          5773 => x"8c",
          5774 => x"17",
          5775 => x"86",
          5776 => x"17",
          5777 => x"75",
          5778 => x"3f",
          5779 => x"08",
          5780 => x"2e",
          5781 => x"85",
          5782 => x"86",
          5783 => x"2e",
          5784 => x"76",
          5785 => x"73",
          5786 => x"0c",
          5787 => x"04",
          5788 => x"76",
          5789 => x"05",
          5790 => x"53",
          5791 => x"82",
          5792 => x"87",
          5793 => x"ec",
          5794 => x"86",
          5795 => x"fb",
          5796 => x"79",
          5797 => x"05",
          5798 => x"56",
          5799 => x"3f",
          5800 => x"08",
          5801 => x"ec",
          5802 => x"38",
          5803 => x"82",
          5804 => x"52",
          5805 => x"f8",
          5806 => x"ec",
          5807 => x"ca",
          5808 => x"ec",
          5809 => x"51",
          5810 => x"82",
          5811 => x"53",
          5812 => x"08",
          5813 => x"81",
          5814 => x"80",
          5815 => x"82",
          5816 => x"a6",
          5817 => x"73",
          5818 => x"3f",
          5819 => x"51",
          5820 => x"82",
          5821 => x"84",
          5822 => x"70",
          5823 => x"2c",
          5824 => x"ec",
          5825 => x"51",
          5826 => x"82",
          5827 => x"87",
          5828 => x"ee",
          5829 => x"57",
          5830 => x"3d",
          5831 => x"3d",
          5832 => x"af",
          5833 => x"ec",
          5834 => x"8c",
          5835 => x"38",
          5836 => x"51",
          5837 => x"82",
          5838 => x"55",
          5839 => x"08",
          5840 => x"80",
          5841 => x"70",
          5842 => x"58",
          5843 => x"85",
          5844 => x"8d",
          5845 => x"2e",
          5846 => x"52",
          5847 => x"be",
          5848 => x"8c",
          5849 => x"3d",
          5850 => x"3d",
          5851 => x"55",
          5852 => x"92",
          5853 => x"52",
          5854 => x"de",
          5855 => x"8c",
          5856 => x"82",
          5857 => x"82",
          5858 => x"74",
          5859 => x"98",
          5860 => x"11",
          5861 => x"59",
          5862 => x"75",
          5863 => x"38",
          5864 => x"81",
          5865 => x"5b",
          5866 => x"82",
          5867 => x"39",
          5868 => x"08",
          5869 => x"59",
          5870 => x"09",
          5871 => x"38",
          5872 => x"57",
          5873 => x"3d",
          5874 => x"c1",
          5875 => x"8c",
          5876 => x"2e",
          5877 => x"8c",
          5878 => x"2e",
          5879 => x"8c",
          5880 => x"70",
          5881 => x"08",
          5882 => x"7a",
          5883 => x"7f",
          5884 => x"54",
          5885 => x"77",
          5886 => x"80",
          5887 => x"15",
          5888 => x"ec",
          5889 => x"75",
          5890 => x"52",
          5891 => x"52",
          5892 => x"8d",
          5893 => x"ec",
          5894 => x"8c",
          5895 => x"d6",
          5896 => x"33",
          5897 => x"1a",
          5898 => x"54",
          5899 => x"09",
          5900 => x"38",
          5901 => x"ff",
          5902 => x"82",
          5903 => x"83",
          5904 => x"70",
          5905 => x"25",
          5906 => x"59",
          5907 => x"9b",
          5908 => x"51",
          5909 => x"3f",
          5910 => x"08",
          5911 => x"70",
          5912 => x"25",
          5913 => x"59",
          5914 => x"75",
          5915 => x"7a",
          5916 => x"ff",
          5917 => x"7c",
          5918 => x"90",
          5919 => x"11",
          5920 => x"56",
          5921 => x"15",
          5922 => x"8c",
          5923 => x"3d",
          5924 => x"3d",
          5925 => x"3d",
          5926 => x"70",
          5927 => x"dd",
          5928 => x"ec",
          5929 => x"8c",
          5930 => x"a8",
          5931 => x"33",
          5932 => x"a0",
          5933 => x"33",
          5934 => x"70",
          5935 => x"55",
          5936 => x"73",
          5937 => x"8e",
          5938 => x"08",
          5939 => x"18",
          5940 => x"80",
          5941 => x"38",
          5942 => x"08",
          5943 => x"08",
          5944 => x"c4",
          5945 => x"8c",
          5946 => x"88",
          5947 => x"80",
          5948 => x"17",
          5949 => x"51",
          5950 => x"3f",
          5951 => x"08",
          5952 => x"81",
          5953 => x"81",
          5954 => x"ec",
          5955 => x"09",
          5956 => x"38",
          5957 => x"39",
          5958 => x"77",
          5959 => x"ec",
          5960 => x"08",
          5961 => x"98",
          5962 => x"82",
          5963 => x"52",
          5964 => x"bd",
          5965 => x"ec",
          5966 => x"17",
          5967 => x"0c",
          5968 => x"80",
          5969 => x"73",
          5970 => x"75",
          5971 => x"38",
          5972 => x"34",
          5973 => x"82",
          5974 => x"89",
          5975 => x"e2",
          5976 => x"53",
          5977 => x"a4",
          5978 => x"3d",
          5979 => x"3f",
          5980 => x"08",
          5981 => x"ec",
          5982 => x"38",
          5983 => x"3d",
          5984 => x"3d",
          5985 => x"d1",
          5986 => x"8c",
          5987 => x"82",
          5988 => x"81",
          5989 => x"80",
          5990 => x"70",
          5991 => x"81",
          5992 => x"56",
          5993 => x"81",
          5994 => x"98",
          5995 => x"74",
          5996 => x"38",
          5997 => x"05",
          5998 => x"06",
          5999 => x"55",
          6000 => x"38",
          6001 => x"51",
          6002 => x"82",
          6003 => x"74",
          6004 => x"81",
          6005 => x"56",
          6006 => x"80",
          6007 => x"54",
          6008 => x"08",
          6009 => x"2e",
          6010 => x"73",
          6011 => x"ec",
          6012 => x"52",
          6013 => x"52",
          6014 => x"3f",
          6015 => x"08",
          6016 => x"ec",
          6017 => x"38",
          6018 => x"08",
          6019 => x"cc",
          6020 => x"8c",
          6021 => x"82",
          6022 => x"86",
          6023 => x"80",
          6024 => x"8c",
          6025 => x"2e",
          6026 => x"8c",
          6027 => x"c0",
          6028 => x"ce",
          6029 => x"8c",
          6030 => x"8c",
          6031 => x"70",
          6032 => x"08",
          6033 => x"51",
          6034 => x"80",
          6035 => x"73",
          6036 => x"38",
          6037 => x"52",
          6038 => x"95",
          6039 => x"ec",
          6040 => x"8c",
          6041 => x"ff",
          6042 => x"82",
          6043 => x"55",
          6044 => x"ec",
          6045 => x"0d",
          6046 => x"0d",
          6047 => x"3d",
          6048 => x"9a",
          6049 => x"cb",
          6050 => x"ec",
          6051 => x"8c",
          6052 => x"b0",
          6053 => x"69",
          6054 => x"70",
          6055 => x"97",
          6056 => x"ec",
          6057 => x"8c",
          6058 => x"38",
          6059 => x"94",
          6060 => x"ec",
          6061 => x"09",
          6062 => x"88",
          6063 => x"df",
          6064 => x"85",
          6065 => x"51",
          6066 => x"74",
          6067 => x"78",
          6068 => x"8a",
          6069 => x"57",
          6070 => x"82",
          6071 => x"75",
          6072 => x"8c",
          6073 => x"38",
          6074 => x"8c",
          6075 => x"2e",
          6076 => x"83",
          6077 => x"82",
          6078 => x"ff",
          6079 => x"06",
          6080 => x"54",
          6081 => x"73",
          6082 => x"82",
          6083 => x"52",
          6084 => x"a4",
          6085 => x"ec",
          6086 => x"8c",
          6087 => x"9a",
          6088 => x"a0",
          6089 => x"51",
          6090 => x"3f",
          6091 => x"0b",
          6092 => x"78",
          6093 => x"bf",
          6094 => x"88",
          6095 => x"80",
          6096 => x"ff",
          6097 => x"75",
          6098 => x"11",
          6099 => x"f8",
          6100 => x"78",
          6101 => x"80",
          6102 => x"ff",
          6103 => x"78",
          6104 => x"80",
          6105 => x"7f",
          6106 => x"d4",
          6107 => x"c9",
          6108 => x"54",
          6109 => x"15",
          6110 => x"cb",
          6111 => x"8c",
          6112 => x"82",
          6113 => x"b2",
          6114 => x"b2",
          6115 => x"96",
          6116 => x"b5",
          6117 => x"53",
          6118 => x"51",
          6119 => x"64",
          6120 => x"8b",
          6121 => x"54",
          6122 => x"15",
          6123 => x"ff",
          6124 => x"82",
          6125 => x"54",
          6126 => x"53",
          6127 => x"51",
          6128 => x"3f",
          6129 => x"ec",
          6130 => x"0d",
          6131 => x"0d",
          6132 => x"05",
          6133 => x"3f",
          6134 => x"3d",
          6135 => x"52",
          6136 => x"d5",
          6137 => x"8c",
          6138 => x"82",
          6139 => x"82",
          6140 => x"4d",
          6141 => x"52",
          6142 => x"52",
          6143 => x"3f",
          6144 => x"08",
          6145 => x"ec",
          6146 => x"38",
          6147 => x"05",
          6148 => x"06",
          6149 => x"73",
          6150 => x"a0",
          6151 => x"08",
          6152 => x"ff",
          6153 => x"ff",
          6154 => x"ac",
          6155 => x"92",
          6156 => x"54",
          6157 => x"3f",
          6158 => x"52",
          6159 => x"f7",
          6160 => x"ec",
          6161 => x"8c",
          6162 => x"38",
          6163 => x"09",
          6164 => x"38",
          6165 => x"08",
          6166 => x"88",
          6167 => x"39",
          6168 => x"08",
          6169 => x"81",
          6170 => x"38",
          6171 => x"b1",
          6172 => x"ec",
          6173 => x"8c",
          6174 => x"c8",
          6175 => x"93",
          6176 => x"ff",
          6177 => x"8d",
          6178 => x"b4",
          6179 => x"af",
          6180 => x"17",
          6181 => x"33",
          6182 => x"70",
          6183 => x"55",
          6184 => x"38",
          6185 => x"54",
          6186 => x"34",
          6187 => x"0b",
          6188 => x"8b",
          6189 => x"84",
          6190 => x"06",
          6191 => x"73",
          6192 => x"e5",
          6193 => x"2e",
          6194 => x"75",
          6195 => x"c6",
          6196 => x"8c",
          6197 => x"78",
          6198 => x"bb",
          6199 => x"82",
          6200 => x"80",
          6201 => x"38",
          6202 => x"08",
          6203 => x"ff",
          6204 => x"82",
          6205 => x"79",
          6206 => x"58",
          6207 => x"8c",
          6208 => x"c0",
          6209 => x"33",
          6210 => x"2e",
          6211 => x"99",
          6212 => x"75",
          6213 => x"c6",
          6214 => x"54",
          6215 => x"15",
          6216 => x"82",
          6217 => x"9c",
          6218 => x"c8",
          6219 => x"8c",
          6220 => x"82",
          6221 => x"8c",
          6222 => x"ff",
          6223 => x"82",
          6224 => x"55",
          6225 => x"ec",
          6226 => x"0d",
          6227 => x"0d",
          6228 => x"05",
          6229 => x"05",
          6230 => x"33",
          6231 => x"53",
          6232 => x"05",
          6233 => x"51",
          6234 => x"82",
          6235 => x"55",
          6236 => x"08",
          6237 => x"78",
          6238 => x"95",
          6239 => x"51",
          6240 => x"82",
          6241 => x"55",
          6242 => x"08",
          6243 => x"80",
          6244 => x"81",
          6245 => x"86",
          6246 => x"38",
          6247 => x"61",
          6248 => x"12",
          6249 => x"7a",
          6250 => x"51",
          6251 => x"74",
          6252 => x"78",
          6253 => x"83",
          6254 => x"51",
          6255 => x"3f",
          6256 => x"08",
          6257 => x"8c",
          6258 => x"3d",
          6259 => x"3d",
          6260 => x"82",
          6261 => x"d0",
          6262 => x"3d",
          6263 => x"3f",
          6264 => x"08",
          6265 => x"ec",
          6266 => x"38",
          6267 => x"52",
          6268 => x"05",
          6269 => x"3f",
          6270 => x"08",
          6271 => x"ec",
          6272 => x"02",
          6273 => x"33",
          6274 => x"54",
          6275 => x"a6",
          6276 => x"22",
          6277 => x"71",
          6278 => x"53",
          6279 => x"51",
          6280 => x"3f",
          6281 => x"0b",
          6282 => x"76",
          6283 => x"b8",
          6284 => x"ec",
          6285 => x"82",
          6286 => x"93",
          6287 => x"ea",
          6288 => x"6b",
          6289 => x"53",
          6290 => x"05",
          6291 => x"51",
          6292 => x"82",
          6293 => x"82",
          6294 => x"30",
          6295 => x"ec",
          6296 => x"25",
          6297 => x"79",
          6298 => x"85",
          6299 => x"75",
          6300 => x"73",
          6301 => x"f9",
          6302 => x"80",
          6303 => x"8d",
          6304 => x"54",
          6305 => x"3f",
          6306 => x"08",
          6307 => x"ec",
          6308 => x"38",
          6309 => x"51",
          6310 => x"82",
          6311 => x"57",
          6312 => x"08",
          6313 => x"8c",
          6314 => x"8c",
          6315 => x"5b",
          6316 => x"18",
          6317 => x"18",
          6318 => x"74",
          6319 => x"81",
          6320 => x"78",
          6321 => x"8b",
          6322 => x"54",
          6323 => x"75",
          6324 => x"38",
          6325 => x"1b",
          6326 => x"55",
          6327 => x"2e",
          6328 => x"39",
          6329 => x"09",
          6330 => x"38",
          6331 => x"80",
          6332 => x"70",
          6333 => x"25",
          6334 => x"80",
          6335 => x"38",
          6336 => x"bc",
          6337 => x"11",
          6338 => x"ff",
          6339 => x"82",
          6340 => x"57",
          6341 => x"08",
          6342 => x"70",
          6343 => x"80",
          6344 => x"83",
          6345 => x"80",
          6346 => x"84",
          6347 => x"a7",
          6348 => x"b4",
          6349 => x"ad",
          6350 => x"8c",
          6351 => x"0c",
          6352 => x"ec",
          6353 => x"0d",
          6354 => x"0d",
          6355 => x"3d",
          6356 => x"52",
          6357 => x"ce",
          6358 => x"8c",
          6359 => x"8c",
          6360 => x"54",
          6361 => x"08",
          6362 => x"8b",
          6363 => x"8b",
          6364 => x"59",
          6365 => x"3f",
          6366 => x"33",
          6367 => x"06",
          6368 => x"57",
          6369 => x"81",
          6370 => x"58",
          6371 => x"06",
          6372 => x"4e",
          6373 => x"ff",
          6374 => x"82",
          6375 => x"80",
          6376 => x"6c",
          6377 => x"53",
          6378 => x"ae",
          6379 => x"8c",
          6380 => x"2e",
          6381 => x"88",
          6382 => x"6d",
          6383 => x"55",
          6384 => x"8c",
          6385 => x"ff",
          6386 => x"83",
          6387 => x"51",
          6388 => x"26",
          6389 => x"15",
          6390 => x"ff",
          6391 => x"80",
          6392 => x"87",
          6393 => x"bc",
          6394 => x"74",
          6395 => x"38",
          6396 => x"fd",
          6397 => x"ae",
          6398 => x"8c",
          6399 => x"38",
          6400 => x"27",
          6401 => x"89",
          6402 => x"8b",
          6403 => x"27",
          6404 => x"55",
          6405 => x"81",
          6406 => x"8f",
          6407 => x"2a",
          6408 => x"70",
          6409 => x"34",
          6410 => x"74",
          6411 => x"05",
          6412 => x"17",
          6413 => x"70",
          6414 => x"52",
          6415 => x"73",
          6416 => x"c8",
          6417 => x"33",
          6418 => x"73",
          6419 => x"81",
          6420 => x"80",
          6421 => x"02",
          6422 => x"76",
          6423 => x"51",
          6424 => x"2e",
          6425 => x"87",
          6426 => x"57",
          6427 => x"79",
          6428 => x"80",
          6429 => x"70",
          6430 => x"ba",
          6431 => x"8c",
          6432 => x"82",
          6433 => x"80",
          6434 => x"52",
          6435 => x"bf",
          6436 => x"8c",
          6437 => x"82",
          6438 => x"8d",
          6439 => x"c4",
          6440 => x"e5",
          6441 => x"c6",
          6442 => x"ec",
          6443 => x"09",
          6444 => x"cc",
          6445 => x"76",
          6446 => x"c4",
          6447 => x"74",
          6448 => x"b0",
          6449 => x"ec",
          6450 => x"8c",
          6451 => x"38",
          6452 => x"8c",
          6453 => x"67",
          6454 => x"db",
          6455 => x"88",
          6456 => x"34",
          6457 => x"52",
          6458 => x"ab",
          6459 => x"54",
          6460 => x"15",
          6461 => x"ff",
          6462 => x"82",
          6463 => x"54",
          6464 => x"82",
          6465 => x"9c",
          6466 => x"f2",
          6467 => x"62",
          6468 => x"80",
          6469 => x"93",
          6470 => x"55",
          6471 => x"5e",
          6472 => x"3f",
          6473 => x"08",
          6474 => x"ec",
          6475 => x"38",
          6476 => x"58",
          6477 => x"38",
          6478 => x"97",
          6479 => x"08",
          6480 => x"38",
          6481 => x"70",
          6482 => x"81",
          6483 => x"55",
          6484 => x"87",
          6485 => x"39",
          6486 => x"90",
          6487 => x"82",
          6488 => x"8a",
          6489 => x"89",
          6490 => x"7f",
          6491 => x"56",
          6492 => x"3f",
          6493 => x"06",
          6494 => x"72",
          6495 => x"82",
          6496 => x"05",
          6497 => x"7c",
          6498 => x"55",
          6499 => x"27",
          6500 => x"16",
          6501 => x"83",
          6502 => x"76",
          6503 => x"80",
          6504 => x"79",
          6505 => x"99",
          6506 => x"7f",
          6507 => x"14",
          6508 => x"83",
          6509 => x"82",
          6510 => x"81",
          6511 => x"38",
          6512 => x"08",
          6513 => x"95",
          6514 => x"ec",
          6515 => x"81",
          6516 => x"7b",
          6517 => x"06",
          6518 => x"39",
          6519 => x"56",
          6520 => x"09",
          6521 => x"b9",
          6522 => x"80",
          6523 => x"80",
          6524 => x"78",
          6525 => x"7a",
          6526 => x"38",
          6527 => x"73",
          6528 => x"81",
          6529 => x"ff",
          6530 => x"74",
          6531 => x"ff",
          6532 => x"82",
          6533 => x"58",
          6534 => x"08",
          6535 => x"74",
          6536 => x"16",
          6537 => x"73",
          6538 => x"39",
          6539 => x"7e",
          6540 => x"0c",
          6541 => x"2e",
          6542 => x"88",
          6543 => x"8c",
          6544 => x"1a",
          6545 => x"07",
          6546 => x"1b",
          6547 => x"08",
          6548 => x"16",
          6549 => x"75",
          6550 => x"38",
          6551 => x"90",
          6552 => x"15",
          6553 => x"54",
          6554 => x"34",
          6555 => x"82",
          6556 => x"90",
          6557 => x"e9",
          6558 => x"6d",
          6559 => x"80",
          6560 => x"9d",
          6561 => x"5c",
          6562 => x"3f",
          6563 => x"0b",
          6564 => x"08",
          6565 => x"38",
          6566 => x"08",
          6567 => x"8d",
          6568 => x"08",
          6569 => x"80",
          6570 => x"80",
          6571 => x"8c",
          6572 => x"ff",
          6573 => x"52",
          6574 => x"a0",
          6575 => x"8c",
          6576 => x"ff",
          6577 => x"06",
          6578 => x"56",
          6579 => x"38",
          6580 => x"70",
          6581 => x"55",
          6582 => x"8b",
          6583 => x"3d",
          6584 => x"83",
          6585 => x"ff",
          6586 => x"82",
          6587 => x"99",
          6588 => x"74",
          6589 => x"38",
          6590 => x"80",
          6591 => x"ff",
          6592 => x"55",
          6593 => x"83",
          6594 => x"78",
          6595 => x"38",
          6596 => x"26",
          6597 => x"81",
          6598 => x"8b",
          6599 => x"79",
          6600 => x"80",
          6601 => x"93",
          6602 => x"39",
          6603 => x"6e",
          6604 => x"89",
          6605 => x"48",
          6606 => x"83",
          6607 => x"61",
          6608 => x"25",
          6609 => x"55",
          6610 => x"8a",
          6611 => x"3d",
          6612 => x"81",
          6613 => x"ff",
          6614 => x"81",
          6615 => x"ec",
          6616 => x"38",
          6617 => x"70",
          6618 => x"8c",
          6619 => x"56",
          6620 => x"38",
          6621 => x"55",
          6622 => x"75",
          6623 => x"38",
          6624 => x"70",
          6625 => x"ff",
          6626 => x"83",
          6627 => x"78",
          6628 => x"89",
          6629 => x"81",
          6630 => x"06",
          6631 => x"80",
          6632 => x"77",
          6633 => x"74",
          6634 => x"8d",
          6635 => x"06",
          6636 => x"2e",
          6637 => x"77",
          6638 => x"93",
          6639 => x"74",
          6640 => x"cb",
          6641 => x"7d",
          6642 => x"81",
          6643 => x"38",
          6644 => x"66",
          6645 => x"81",
          6646 => x"e0",
          6647 => x"74",
          6648 => x"38",
          6649 => x"98",
          6650 => x"e0",
          6651 => x"82",
          6652 => x"57",
          6653 => x"80",
          6654 => x"76",
          6655 => x"38",
          6656 => x"51",
          6657 => x"3f",
          6658 => x"08",
          6659 => x"87",
          6660 => x"2a",
          6661 => x"5c",
          6662 => x"8c",
          6663 => x"80",
          6664 => x"44",
          6665 => x"0a",
          6666 => x"ec",
          6667 => x"39",
          6668 => x"66",
          6669 => x"81",
          6670 => x"d0",
          6671 => x"74",
          6672 => x"38",
          6673 => x"98",
          6674 => x"d0",
          6675 => x"82",
          6676 => x"57",
          6677 => x"80",
          6678 => x"76",
          6679 => x"38",
          6680 => x"51",
          6681 => x"3f",
          6682 => x"08",
          6683 => x"57",
          6684 => x"08",
          6685 => x"96",
          6686 => x"82",
          6687 => x"10",
          6688 => x"08",
          6689 => x"72",
          6690 => x"59",
          6691 => x"ff",
          6692 => x"5d",
          6693 => x"44",
          6694 => x"11",
          6695 => x"70",
          6696 => x"71",
          6697 => x"06",
          6698 => x"52",
          6699 => x"40",
          6700 => x"09",
          6701 => x"38",
          6702 => x"18",
          6703 => x"39",
          6704 => x"79",
          6705 => x"70",
          6706 => x"58",
          6707 => x"76",
          6708 => x"38",
          6709 => x"7d",
          6710 => x"70",
          6711 => x"55",
          6712 => x"3f",
          6713 => x"08",
          6714 => x"2e",
          6715 => x"9b",
          6716 => x"ec",
          6717 => x"f5",
          6718 => x"38",
          6719 => x"38",
          6720 => x"59",
          6721 => x"38",
          6722 => x"7d",
          6723 => x"81",
          6724 => x"38",
          6725 => x"0b",
          6726 => x"08",
          6727 => x"78",
          6728 => x"1a",
          6729 => x"c0",
          6730 => x"74",
          6731 => x"39",
          6732 => x"55",
          6733 => x"8f",
          6734 => x"fd",
          6735 => x"8c",
          6736 => x"f5",
          6737 => x"78",
          6738 => x"79",
          6739 => x"80",
          6740 => x"f1",
          6741 => x"39",
          6742 => x"81",
          6743 => x"06",
          6744 => x"55",
          6745 => x"27",
          6746 => x"81",
          6747 => x"56",
          6748 => x"38",
          6749 => x"80",
          6750 => x"ff",
          6751 => x"8b",
          6752 => x"f8",
          6753 => x"ff",
          6754 => x"84",
          6755 => x"1b",
          6756 => x"b3",
          6757 => x"1c",
          6758 => x"ff",
          6759 => x"8e",
          6760 => x"a1",
          6761 => x"0b",
          6762 => x"7d",
          6763 => x"30",
          6764 => x"84",
          6765 => x"51",
          6766 => x"51",
          6767 => x"3f",
          6768 => x"83",
          6769 => x"90",
          6770 => x"ff",
          6771 => x"93",
          6772 => x"a0",
          6773 => x"39",
          6774 => x"1b",
          6775 => x"85",
          6776 => x"95",
          6777 => x"52",
          6778 => x"ff",
          6779 => x"81",
          6780 => x"1b",
          6781 => x"cf",
          6782 => x"9c",
          6783 => x"a0",
          6784 => x"83",
          6785 => x"06",
          6786 => x"82",
          6787 => x"52",
          6788 => x"51",
          6789 => x"3f",
          6790 => x"1b",
          6791 => x"c5",
          6792 => x"ac",
          6793 => x"a0",
          6794 => x"52",
          6795 => x"ff",
          6796 => x"86",
          6797 => x"51",
          6798 => x"3f",
          6799 => x"80",
          6800 => x"a9",
          6801 => x"1c",
          6802 => x"81",
          6803 => x"80",
          6804 => x"ae",
          6805 => x"b2",
          6806 => x"1b",
          6807 => x"85",
          6808 => x"ff",
          6809 => x"96",
          6810 => x"9f",
          6811 => x"80",
          6812 => x"34",
          6813 => x"1c",
          6814 => x"81",
          6815 => x"ab",
          6816 => x"a0",
          6817 => x"d4",
          6818 => x"fe",
          6819 => x"59",
          6820 => x"3f",
          6821 => x"53",
          6822 => x"51",
          6823 => x"3f",
          6824 => x"8c",
          6825 => x"e7",
          6826 => x"2e",
          6827 => x"80",
          6828 => x"54",
          6829 => x"53",
          6830 => x"51",
          6831 => x"3f",
          6832 => x"80",
          6833 => x"ff",
          6834 => x"84",
          6835 => x"d2",
          6836 => x"ff",
          6837 => x"86",
          6838 => x"f2",
          6839 => x"1b",
          6840 => x"81",
          6841 => x"52",
          6842 => x"51",
          6843 => x"3f",
          6844 => x"ec",
          6845 => x"9e",
          6846 => x"d4",
          6847 => x"51",
          6848 => x"3f",
          6849 => x"87",
          6850 => x"52",
          6851 => x"9a",
          6852 => x"54",
          6853 => x"7a",
          6854 => x"ff",
          6855 => x"65",
          6856 => x"7a",
          6857 => x"8f",
          6858 => x"80",
          6859 => x"2e",
          6860 => x"9a",
          6861 => x"7a",
          6862 => x"a9",
          6863 => x"84",
          6864 => x"9e",
          6865 => x"0a",
          6866 => x"51",
          6867 => x"ff",
          6868 => x"7d",
          6869 => x"38",
          6870 => x"52",
          6871 => x"9e",
          6872 => x"55",
          6873 => x"62",
          6874 => x"74",
          6875 => x"75",
          6876 => x"7e",
          6877 => x"fe",
          6878 => x"ec",
          6879 => x"38",
          6880 => x"82",
          6881 => x"52",
          6882 => x"9e",
          6883 => x"16",
          6884 => x"56",
          6885 => x"38",
          6886 => x"77",
          6887 => x"8d",
          6888 => x"7d",
          6889 => x"38",
          6890 => x"57",
          6891 => x"83",
          6892 => x"76",
          6893 => x"7a",
          6894 => x"ff",
          6895 => x"82",
          6896 => x"81",
          6897 => x"16",
          6898 => x"56",
          6899 => x"38",
          6900 => x"83",
          6901 => x"86",
          6902 => x"ff",
          6903 => x"38",
          6904 => x"82",
          6905 => x"81",
          6906 => x"06",
          6907 => x"fe",
          6908 => x"53",
          6909 => x"51",
          6910 => x"3f",
          6911 => x"52",
          6912 => x"9c",
          6913 => x"be",
          6914 => x"75",
          6915 => x"81",
          6916 => x"0b",
          6917 => x"77",
          6918 => x"75",
          6919 => x"60",
          6920 => x"80",
          6921 => x"75",
          6922 => x"8c",
          6923 => x"85",
          6924 => x"8c",
          6925 => x"2a",
          6926 => x"75",
          6927 => x"82",
          6928 => x"87",
          6929 => x"52",
          6930 => x"51",
          6931 => x"3f",
          6932 => x"ca",
          6933 => x"9c",
          6934 => x"54",
          6935 => x"52",
          6936 => x"98",
          6937 => x"56",
          6938 => x"08",
          6939 => x"53",
          6940 => x"51",
          6941 => x"3f",
          6942 => x"8c",
          6943 => x"38",
          6944 => x"56",
          6945 => x"56",
          6946 => x"8c",
          6947 => x"75",
          6948 => x"0c",
          6949 => x"04",
          6950 => x"7d",
          6951 => x"80",
          6952 => x"05",
          6953 => x"76",
          6954 => x"38",
          6955 => x"11",
          6956 => x"53",
          6957 => x"79",
          6958 => x"3f",
          6959 => x"09",
          6960 => x"38",
          6961 => x"55",
          6962 => x"db",
          6963 => x"70",
          6964 => x"34",
          6965 => x"74",
          6966 => x"81",
          6967 => x"80",
          6968 => x"55",
          6969 => x"76",
          6970 => x"8c",
          6971 => x"3d",
          6972 => x"3d",
          6973 => x"08",
          6974 => x"57",
          6975 => x"80",
          6976 => x"39",
          6977 => x"85",
          6978 => x"80",
          6979 => x"15",
          6980 => x"33",
          6981 => x"a0",
          6982 => x"81",
          6983 => x"70",
          6984 => x"06",
          6985 => x"e6",
          6986 => x"2e",
          6987 => x"88",
          6988 => x"70",
          6989 => x"34",
          6990 => x"90",
          6991 => x"fc",
          6992 => x"53",
          6993 => x"54",
          6994 => x"3f",
          6995 => x"08",
          6996 => x"14",
          6997 => x"81",
          6998 => x"38",
          6999 => x"81",
          7000 => x"53",
          7001 => x"d2",
          7002 => x"72",
          7003 => x"0c",
          7004 => x"04",
          7005 => x"73",
          7006 => x"26",
          7007 => x"71",
          7008 => x"f5",
          7009 => x"71",
          7010 => x"ff",
          7011 => x"80",
          7012 => x"94",
          7013 => x"39",
          7014 => x"51",
          7015 => x"81",
          7016 => x"80",
          7017 => x"ff",
          7018 => x"e4",
          7019 => x"dc",
          7020 => x"39",
          7021 => x"51",
          7022 => x"82",
          7023 => x"80",
          7024 => x"80",
          7025 => x"c8",
          7026 => x"b0",
          7027 => x"39",
          7028 => x"51",
          7029 => x"80",
          7030 => x"39",
          7031 => x"51",
          7032 => x"81",
          7033 => x"39",
          7034 => x"51",
          7035 => x"81",
          7036 => x"39",
          7037 => x"51",
          7038 => x"82",
          7039 => x"39",
          7040 => x"51",
          7041 => x"82",
          7042 => x"39",
          7043 => x"51",
          7044 => x"3f",
          7045 => x"04",
          7046 => x"77",
          7047 => x"74",
          7048 => x"8a",
          7049 => x"75",
          7050 => x"51",
          7051 => x"e8",
          7052 => x"fe",
          7053 => x"82",
          7054 => x"52",
          7055 => x"ed",
          7056 => x"8c",
          7057 => x"79",
          7058 => x"82",
          7059 => x"ff",
          7060 => x"87",
          7061 => x"ec",
          7062 => x"02",
          7063 => x"e3",
          7064 => x"57",
          7065 => x"30",
          7066 => x"73",
          7067 => x"59",
          7068 => x"77",
          7069 => x"83",
          7070 => x"74",
          7071 => x"81",
          7072 => x"55",
          7073 => x"80",
          7074 => x"53",
          7075 => x"3d",
          7076 => x"c1",
          7077 => x"8c",
          7078 => x"82",
          7079 => x"b8",
          7080 => x"ec",
          7081 => x"98",
          7082 => x"8c",
          7083 => x"96",
          7084 => x"54",
          7085 => x"77",
          7086 => x"c5",
          7087 => x"8c",
          7088 => x"82",
          7089 => x"90",
          7090 => x"74",
          7091 => x"38",
          7092 => x"19",
          7093 => x"39",
          7094 => x"05",
          7095 => x"3f",
          7096 => x"78",
          7097 => x"7b",
          7098 => x"2a",
          7099 => x"57",
          7100 => x"80",
          7101 => x"82",
          7102 => x"87",
          7103 => x"08",
          7104 => x"fe",
          7105 => x"56",
          7106 => x"ec",
          7107 => x"0d",
          7108 => x"0d",
          7109 => x"05",
          7110 => x"57",
          7111 => x"80",
          7112 => x"79",
          7113 => x"3f",
          7114 => x"08",
          7115 => x"80",
          7116 => x"75",
          7117 => x"38",
          7118 => x"55",
          7119 => x"8c",
          7120 => x"52",
          7121 => x"2d",
          7122 => x"08",
          7123 => x"77",
          7124 => x"8c",
          7125 => x"3d",
          7126 => x"3d",
          7127 => x"63",
          7128 => x"80",
          7129 => x"73",
          7130 => x"41",
          7131 => x"5e",
          7132 => x"52",
          7133 => x"51",
          7134 => x"3f",
          7135 => x"51",
          7136 => x"3f",
          7137 => x"79",
          7138 => x"38",
          7139 => x"89",
          7140 => x"2e",
          7141 => x"c6",
          7142 => x"53",
          7143 => x"8e",
          7144 => x"52",
          7145 => x"51",
          7146 => x"3f",
          7147 => x"83",
          7148 => x"82",
          7149 => x"15",
          7150 => x"39",
          7151 => x"72",
          7152 => x"38",
          7153 => x"82",
          7154 => x"ff",
          7155 => x"89",
          7156 => x"90",
          7157 => x"da",
          7158 => x"55",
          7159 => x"18",
          7160 => x"27",
          7161 => x"33",
          7162 => x"9c",
          7163 => x"a6",
          7164 => x"82",
          7165 => x"ff",
          7166 => x"81",
          7167 => x"51",
          7168 => x"3f",
          7169 => x"82",
          7170 => x"ff",
          7171 => x"80",
          7172 => x"27",
          7173 => x"18",
          7174 => x"53",
          7175 => x"7a",
          7176 => x"81",
          7177 => x"9f",
          7178 => x"38",
          7179 => x"73",
          7180 => x"ff",
          7181 => x"72",
          7182 => x"38",
          7183 => x"26",
          7184 => x"51",
          7185 => x"51",
          7186 => x"3f",
          7187 => x"c1",
          7188 => x"ac",
          7189 => x"da",
          7190 => x"79",
          7191 => x"fe",
          7192 => x"82",
          7193 => x"98",
          7194 => x"2c",
          7195 => x"a0",
          7196 => x"06",
          7197 => x"f6",
          7198 => x"8c",
          7199 => x"2b",
          7200 => x"70",
          7201 => x"30",
          7202 => x"70",
          7203 => x"07",
          7204 => x"06",
          7205 => x"59",
          7206 => x"80",
          7207 => x"38",
          7208 => x"09",
          7209 => x"38",
          7210 => x"39",
          7211 => x"72",
          7212 => x"be",
          7213 => x"72",
          7214 => x"0c",
          7215 => x"04",
          7216 => x"02",
          7217 => x"82",
          7218 => x"82",
          7219 => x"55",
          7220 => x"3f",
          7221 => x"22",
          7222 => x"9d",
          7223 => x"c0",
          7224 => x"cc",
          7225 => x"cd",
          7226 => x"83",
          7227 => x"86",
          7228 => x"80",
          7229 => x"fe",
          7230 => x"86",
          7231 => x"fe",
          7232 => x"c0",
          7233 => x"53",
          7234 => x"3f",
          7235 => x"f1",
          7236 => x"83",
          7237 => x"f3",
          7238 => x"51",
          7239 => x"3f",
          7240 => x"70",
          7241 => x"52",
          7242 => x"95",
          7243 => x"fe",
          7244 => x"82",
          7245 => x"fe",
          7246 => x"80",
          7247 => x"92",
          7248 => x"2a",
          7249 => x"51",
          7250 => x"2e",
          7251 => x"51",
          7252 => x"3f",
          7253 => x"51",
          7254 => x"3f",
          7255 => x"f0",
          7256 => x"83",
          7257 => x"06",
          7258 => x"80",
          7259 => x"81",
          7260 => x"de",
          7261 => x"ac",
          7262 => x"d6",
          7263 => x"fe",
          7264 => x"72",
          7265 => x"81",
          7266 => x"71",
          7267 => x"38",
          7268 => x"f0",
          7269 => x"84",
          7270 => x"f2",
          7271 => x"51",
          7272 => x"3f",
          7273 => x"70",
          7274 => x"52",
          7275 => x"95",
          7276 => x"fe",
          7277 => x"82",
          7278 => x"fe",
          7279 => x"80",
          7280 => x"8e",
          7281 => x"2a",
          7282 => x"51",
          7283 => x"2e",
          7284 => x"51",
          7285 => x"3f",
          7286 => x"51",
          7287 => x"3f",
          7288 => x"ef",
          7289 => x"87",
          7290 => x"06",
          7291 => x"80",
          7292 => x"81",
          7293 => x"da",
          7294 => x"fc",
          7295 => x"d2",
          7296 => x"fe",
          7297 => x"72",
          7298 => x"81",
          7299 => x"71",
          7300 => x"38",
          7301 => x"ef",
          7302 => x"85",
          7303 => x"f1",
          7304 => x"51",
          7305 => x"3f",
          7306 => x"3f",
          7307 => x"04",
          7308 => x"77",
          7309 => x"56",
          7310 => x"75",
          7311 => x"f0",
          7312 => x"f8",
          7313 => x"a7",
          7314 => x"82",
          7315 => x"82",
          7316 => x"ff",
          7317 => x"82",
          7318 => x"30",
          7319 => x"ec",
          7320 => x"25",
          7321 => x"51",
          7322 => x"82",
          7323 => x"82",
          7324 => x"54",
          7325 => x"09",
          7326 => x"38",
          7327 => x"53",
          7328 => x"51",
          7329 => x"82",
          7330 => x"80",
          7331 => x"82",
          7332 => x"51",
          7333 => x"3f",
          7334 => x"a3",
          7335 => x"83",
          7336 => x"82",
          7337 => x"82",
          7338 => x"54",
          7339 => x"09",
          7340 => x"38",
          7341 => x"51",
          7342 => x"3f",
          7343 => x"8c",
          7344 => x"3d",
          7345 => x"3d",
          7346 => x"71",
          7347 => x"0c",
          7348 => x"52",
          7349 => x"88",
          7350 => x"8c",
          7351 => x"ff",
          7352 => x"7d",
          7353 => x"06",
          7354 => x"85",
          7355 => x"3d",
          7356 => x"ff",
          7357 => x"7c",
          7358 => x"82",
          7359 => x"ff",
          7360 => x"82",
          7361 => x"7d",
          7362 => x"82",
          7363 => x"8d",
          7364 => x"70",
          7365 => x"86",
          7366 => x"fc",
          7367 => x"3d",
          7368 => x"80",
          7369 => x"51",
          7370 => x"b4",
          7371 => x"05",
          7372 => x"3f",
          7373 => x"08",
          7374 => x"90",
          7375 => x"78",
          7376 => x"87",
          7377 => x"80",
          7378 => x"38",
          7379 => x"81",
          7380 => x"bd",
          7381 => x"78",
          7382 => x"ba",
          7383 => x"2e",
          7384 => x"8a",
          7385 => x"80",
          7386 => x"a1",
          7387 => x"c0",
          7388 => x"38",
          7389 => x"82",
          7390 => x"d2",
          7391 => x"f9",
          7392 => x"38",
          7393 => x"24",
          7394 => x"80",
          7395 => x"98",
          7396 => x"f8",
          7397 => x"38",
          7398 => x"78",
          7399 => x"8a",
          7400 => x"81",
          7401 => x"38",
          7402 => x"2e",
          7403 => x"8a",
          7404 => x"81",
          7405 => x"8f",
          7406 => x"39",
          7407 => x"80",
          7408 => x"84",
          7409 => x"82",
          7410 => x"8c",
          7411 => x"2e",
          7412 => x"b4",
          7413 => x"11",
          7414 => x"05",
          7415 => x"ab",
          7416 => x"ec",
          7417 => x"fe",
          7418 => x"3d",
          7419 => x"53",
          7420 => x"51",
          7421 => x"3f",
          7422 => x"08",
          7423 => x"8c",
          7424 => x"82",
          7425 => x"fe",
          7426 => x"63",
          7427 => x"79",
          7428 => x"f2",
          7429 => x"78",
          7430 => x"05",
          7431 => x"7a",
          7432 => x"81",
          7433 => x"3d",
          7434 => x"53",
          7435 => x"51",
          7436 => x"3f",
          7437 => x"08",
          7438 => x"da",
          7439 => x"fe",
          7440 => x"ff",
          7441 => x"ff",
          7442 => x"82",
          7443 => x"80",
          7444 => x"38",
          7445 => x"f8",
          7446 => x"84",
          7447 => x"81",
          7448 => x"8c",
          7449 => x"2e",
          7450 => x"82",
          7451 => x"fe",
          7452 => x"63",
          7453 => x"27",
          7454 => x"61",
          7455 => x"81",
          7456 => x"79",
          7457 => x"05",
          7458 => x"b4",
          7459 => x"11",
          7460 => x"05",
          7461 => x"f3",
          7462 => x"ec",
          7463 => x"fc",
          7464 => x"3d",
          7465 => x"53",
          7466 => x"51",
          7467 => x"3f",
          7468 => x"08",
          7469 => x"de",
          7470 => x"fe",
          7471 => x"ff",
          7472 => x"ff",
          7473 => x"82",
          7474 => x"80",
          7475 => x"38",
          7476 => x"51",
          7477 => x"3f",
          7478 => x"63",
          7479 => x"61",
          7480 => x"33",
          7481 => x"78",
          7482 => x"38",
          7483 => x"54",
          7484 => x"79",
          7485 => x"cc",
          7486 => x"9a",
          7487 => x"62",
          7488 => x"5a",
          7489 => x"86",
          7490 => x"bd",
          7491 => x"ff",
          7492 => x"ff",
          7493 => x"fe",
          7494 => x"82",
          7495 => x"80",
          7496 => x"89",
          7497 => x"78",
          7498 => x"38",
          7499 => x"08",
          7500 => x"39",
          7501 => x"33",
          7502 => x"2e",
          7503 => x"89",
          7504 => x"bc",
          7505 => x"e2",
          7506 => x"80",
          7507 => x"82",
          7508 => x"44",
          7509 => x"89",
          7510 => x"78",
          7511 => x"38",
          7512 => x"08",
          7513 => x"82",
          7514 => x"59",
          7515 => x"88",
          7516 => x"b8",
          7517 => x"39",
          7518 => x"08",
          7519 => x"44",
          7520 => x"fc",
          7521 => x"84",
          7522 => x"fe",
          7523 => x"8c",
          7524 => x"de",
          7525 => x"e0",
          7526 => x"80",
          7527 => x"82",
          7528 => x"43",
          7529 => x"82",
          7530 => x"59",
          7531 => x"88",
          7532 => x"a4",
          7533 => x"39",
          7534 => x"33",
          7535 => x"2e",
          7536 => x"89",
          7537 => x"aa",
          7538 => x"e3",
          7539 => x"80",
          7540 => x"82",
          7541 => x"43",
          7542 => x"89",
          7543 => x"78",
          7544 => x"38",
          7545 => x"08",
          7546 => x"82",
          7547 => x"88",
          7548 => x"3d",
          7549 => x"53",
          7550 => x"51",
          7551 => x"3f",
          7552 => x"08",
          7553 => x"38",
          7554 => x"5c",
          7555 => x"83",
          7556 => x"7a",
          7557 => x"30",
          7558 => x"9f",
          7559 => x"06",
          7560 => x"5a",
          7561 => x"88",
          7562 => x"2e",
          7563 => x"42",
          7564 => x"51",
          7565 => x"3f",
          7566 => x"54",
          7567 => x"52",
          7568 => x"96",
          7569 => x"f8",
          7570 => x"e6",
          7571 => x"39",
          7572 => x"80",
          7573 => x"84",
          7574 => x"fd",
          7575 => x"8c",
          7576 => x"2e",
          7577 => x"b4",
          7578 => x"11",
          7579 => x"05",
          7580 => x"97",
          7581 => x"ec",
          7582 => x"a5",
          7583 => x"02",
          7584 => x"33",
          7585 => x"81",
          7586 => x"3d",
          7587 => x"53",
          7588 => x"51",
          7589 => x"3f",
          7590 => x"08",
          7591 => x"f6",
          7592 => x"33",
          7593 => x"87",
          7594 => x"fa",
          7595 => x"f8",
          7596 => x"fe",
          7597 => x"79",
          7598 => x"59",
          7599 => x"f8",
          7600 => x"79",
          7601 => x"b4",
          7602 => x"11",
          7603 => x"05",
          7604 => x"b7",
          7605 => x"ec",
          7606 => x"91",
          7607 => x"02",
          7608 => x"33",
          7609 => x"81",
          7610 => x"b5",
          7611 => x"90",
          7612 => x"be",
          7613 => x"39",
          7614 => x"f4",
          7615 => x"84",
          7616 => x"fd",
          7617 => x"8c",
          7618 => x"2e",
          7619 => x"b4",
          7620 => x"11",
          7621 => x"05",
          7622 => x"e1",
          7623 => x"ec",
          7624 => x"a6",
          7625 => x"02",
          7626 => x"79",
          7627 => x"5b",
          7628 => x"b4",
          7629 => x"11",
          7630 => x"05",
          7631 => x"bd",
          7632 => x"ec",
          7633 => x"f7",
          7634 => x"70",
          7635 => x"82",
          7636 => x"fe",
          7637 => x"80",
          7638 => x"51",
          7639 => x"3f",
          7640 => x"33",
          7641 => x"2e",
          7642 => x"78",
          7643 => x"38",
          7644 => x"41",
          7645 => x"3d",
          7646 => x"53",
          7647 => x"51",
          7648 => x"3f",
          7649 => x"08",
          7650 => x"38",
          7651 => x"be",
          7652 => x"70",
          7653 => x"23",
          7654 => x"ae",
          7655 => x"90",
          7656 => x"8e",
          7657 => x"39",
          7658 => x"f4",
          7659 => x"84",
          7660 => x"fc",
          7661 => x"8c",
          7662 => x"2e",
          7663 => x"b4",
          7664 => x"11",
          7665 => x"05",
          7666 => x"b1",
          7667 => x"ec",
          7668 => x"a1",
          7669 => x"71",
          7670 => x"84",
          7671 => x"3d",
          7672 => x"53",
          7673 => x"51",
          7674 => x"3f",
          7675 => x"08",
          7676 => x"a2",
          7677 => x"08",
          7678 => x"87",
          7679 => x"f8",
          7680 => x"f8",
          7681 => x"fe",
          7682 => x"79",
          7683 => x"59",
          7684 => x"f6",
          7685 => x"79",
          7686 => x"b4",
          7687 => x"11",
          7688 => x"05",
          7689 => x"d5",
          7690 => x"ec",
          7691 => x"8d",
          7692 => x"71",
          7693 => x"84",
          7694 => x"b9",
          7695 => x"90",
          7696 => x"ee",
          7697 => x"39",
          7698 => x"80",
          7699 => x"84",
          7700 => x"f9",
          7701 => x"8c",
          7702 => x"2e",
          7703 => x"63",
          7704 => x"b0",
          7705 => x"ae",
          7706 => x"78",
          7707 => x"ff",
          7708 => x"ff",
          7709 => x"fe",
          7710 => x"82",
          7711 => x"80",
          7712 => x"38",
          7713 => x"87",
          7714 => x"f7",
          7715 => x"59",
          7716 => x"8c",
          7717 => x"2e",
          7718 => x"82",
          7719 => x"52",
          7720 => x"51",
          7721 => x"3f",
          7722 => x"82",
          7723 => x"fe",
          7724 => x"fe",
          7725 => x"f4",
          7726 => x"88",
          7727 => x"f0",
          7728 => x"59",
          7729 => x"fe",
          7730 => x"f4",
          7731 => x"70",
          7732 => x"78",
          7733 => x"be",
          7734 => x"06",
          7735 => x"2e",
          7736 => x"b4",
          7737 => x"05",
          7738 => x"97",
          7739 => x"ec",
          7740 => x"5b",
          7741 => x"b2",
          7742 => x"24",
          7743 => x"81",
          7744 => x"80",
          7745 => x"83",
          7746 => x"80",
          7747 => x"88",
          7748 => x"55",
          7749 => x"54",
          7750 => x"88",
          7751 => x"3d",
          7752 => x"51",
          7753 => x"3f",
          7754 => x"88",
          7755 => x"3d",
          7756 => x"51",
          7757 => x"3f",
          7758 => x"55",
          7759 => x"54",
          7760 => x"88",
          7761 => x"3d",
          7762 => x"51",
          7763 => x"3f",
          7764 => x"54",
          7765 => x"88",
          7766 => x"3d",
          7767 => x"51",
          7768 => x"3f",
          7769 => x"58",
          7770 => x"57",
          7771 => x"81",
          7772 => x"05",
          7773 => x"83",
          7774 => x"83",
          7775 => x"b4",
          7776 => x"05",
          7777 => x"3f",
          7778 => x"08",
          7779 => x"08",
          7780 => x"70",
          7781 => x"25",
          7782 => x"5f",
          7783 => x"83",
          7784 => x"81",
          7785 => x"06",
          7786 => x"2e",
          7787 => x"1b",
          7788 => x"06",
          7789 => x"fe",
          7790 => x"81",
          7791 => x"32",
          7792 => x"8a",
          7793 => x"2e",
          7794 => x"f2",
          7795 => x"88",
          7796 => x"f4",
          7797 => x"be",
          7798 => x"0d",
          7799 => x"8d",
          7800 => x"c0",
          7801 => x"08",
          7802 => x"84",
          7803 => x"51",
          7804 => x"3f",
          7805 => x"08",
          7806 => x"08",
          7807 => x"84",
          7808 => x"51",
          7809 => x"3f",
          7810 => x"ec",
          7811 => x"0c",
          7812 => x"9c",
          7813 => x"55",
          7814 => x"52",
          7815 => x"d6",
          7816 => x"8c",
          7817 => x"2b",
          7818 => x"53",
          7819 => x"52",
          7820 => x"d6",
          7821 => x"82",
          7822 => x"07",
          7823 => x"80",
          7824 => x"c0",
          7825 => x"8c",
          7826 => x"87",
          7827 => x"0c",
          7828 => x"0b",
          7829 => x"0c",
          7830 => x"0b",
          7831 => x"0c",
          7832 => x"3f",
          7833 => x"3f",
          7834 => x"51",
          7835 => x"3f",
          7836 => x"51",
          7837 => x"3f",
          7838 => x"51",
          7839 => x"3f",
          7840 => x"bc",
          7841 => x"3f",
          7842 => x"00",
          7843 => x"00",
          7844 => x"00",
          7845 => x"00",
          7846 => x"00",
          7847 => x"00",
          7848 => x"00",
          7849 => x"00",
          7850 => x"00",
          7851 => x"00",
          7852 => x"00",
          7853 => x"00",
          7854 => x"00",
          7855 => x"00",
          7856 => x"00",
          7857 => x"00",
          7858 => x"00",
          7859 => x"00",
          7860 => x"00",
          7861 => x"00",
          7862 => x"00",
          7863 => x"00",
          7864 => x"00",
          7865 => x"00",
          7866 => x"00",
          7867 => x"64",
          7868 => x"2f",
          7869 => x"25",
          7870 => x"64",
          7871 => x"2e",
          7872 => x"64",
          7873 => x"6f",
          7874 => x"6f",
          7875 => x"67",
          7876 => x"74",
          7877 => x"00",
          7878 => x"28",
          7879 => x"6d",
          7880 => x"43",
          7881 => x"6e",
          7882 => x"29",
          7883 => x"0a",
          7884 => x"69",
          7885 => x"20",
          7886 => x"6c",
          7887 => x"6e",
          7888 => x"3a",
          7889 => x"20",
          7890 => x"42",
          7891 => x"52",
          7892 => x"20",
          7893 => x"38",
          7894 => x"30",
          7895 => x"2e",
          7896 => x"20",
          7897 => x"44",
          7898 => x"20",
          7899 => x"20",
          7900 => x"38",
          7901 => x"30",
          7902 => x"2e",
          7903 => x"20",
          7904 => x"4e",
          7905 => x"42",
          7906 => x"20",
          7907 => x"38",
          7908 => x"30",
          7909 => x"2e",
          7910 => x"20",
          7911 => x"52",
          7912 => x"20",
          7913 => x"20",
          7914 => x"38",
          7915 => x"30",
          7916 => x"2e",
          7917 => x"20",
          7918 => x"41",
          7919 => x"20",
          7920 => x"20",
          7921 => x"38",
          7922 => x"30",
          7923 => x"2e",
          7924 => x"20",
          7925 => x"44",
          7926 => x"52",
          7927 => x"20",
          7928 => x"76",
          7929 => x"73",
          7930 => x"30",
          7931 => x"2e",
          7932 => x"20",
          7933 => x"49",
          7934 => x"31",
          7935 => x"20",
          7936 => x"6d",
          7937 => x"20",
          7938 => x"30",
          7939 => x"2e",
          7940 => x"20",
          7941 => x"4e",
          7942 => x"43",
          7943 => x"20",
          7944 => x"61",
          7945 => x"6c",
          7946 => x"30",
          7947 => x"2e",
          7948 => x"20",
          7949 => x"49",
          7950 => x"4f",
          7951 => x"42",
          7952 => x"00",
          7953 => x"20",
          7954 => x"42",
          7955 => x"43",
          7956 => x"20",
          7957 => x"4f",
          7958 => x"0a",
          7959 => x"20",
          7960 => x"53",
          7961 => x"00",
          7962 => x"20",
          7963 => x"50",
          7964 => x"00",
          7965 => x"64",
          7966 => x"73",
          7967 => x"3a",
          7968 => x"20",
          7969 => x"50",
          7970 => x"65",
          7971 => x"20",
          7972 => x"74",
          7973 => x"41",
          7974 => x"65",
          7975 => x"3d",
          7976 => x"38",
          7977 => x"00",
          7978 => x"20",
          7979 => x"50",
          7980 => x"65",
          7981 => x"79",
          7982 => x"61",
          7983 => x"41",
          7984 => x"65",
          7985 => x"3d",
          7986 => x"38",
          7987 => x"00",
          7988 => x"20",
          7989 => x"74",
          7990 => x"20",
          7991 => x"72",
          7992 => x"64",
          7993 => x"73",
          7994 => x"20",
          7995 => x"3d",
          7996 => x"38",
          7997 => x"00",
          7998 => x"69",
          7999 => x"0a",
          8000 => x"20",
          8001 => x"50",
          8002 => x"64",
          8003 => x"20",
          8004 => x"20",
          8005 => x"20",
          8006 => x"20",
          8007 => x"3d",
          8008 => x"34",
          8009 => x"00",
          8010 => x"20",
          8011 => x"79",
          8012 => x"6d",
          8013 => x"6f",
          8014 => x"46",
          8015 => x"20",
          8016 => x"20",
          8017 => x"3d",
          8018 => x"2e",
          8019 => x"64",
          8020 => x"0a",
          8021 => x"20",
          8022 => x"44",
          8023 => x"20",
          8024 => x"63",
          8025 => x"72",
          8026 => x"20",
          8027 => x"20",
          8028 => x"3d",
          8029 => x"2e",
          8030 => x"64",
          8031 => x"0a",
          8032 => x"20",
          8033 => x"69",
          8034 => x"6f",
          8035 => x"53",
          8036 => x"4d",
          8037 => x"6f",
          8038 => x"46",
          8039 => x"3d",
          8040 => x"2e",
          8041 => x"64",
          8042 => x"0a",
          8043 => x"6d",
          8044 => x"00",
          8045 => x"65",
          8046 => x"6d",
          8047 => x"6c",
          8048 => x"00",
          8049 => x"56",
          8050 => x"56",
          8051 => x"6e",
          8052 => x"6e",
          8053 => x"77",
          8054 => x"44",
          8055 => x"2a",
          8056 => x"3b",
          8057 => x"3f",
          8058 => x"7f",
          8059 => x"41",
          8060 => x"41",
          8061 => x"00",
          8062 => x"fe",
          8063 => x"44",
          8064 => x"2e",
          8065 => x"4f",
          8066 => x"4d",
          8067 => x"20",
          8068 => x"54",
          8069 => x"20",
          8070 => x"4f",
          8071 => x"4d",
          8072 => x"20",
          8073 => x"54",
          8074 => x"20",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"9a",
          8080 => x"41",
          8081 => x"45",
          8082 => x"49",
          8083 => x"92",
          8084 => x"4f",
          8085 => x"99",
          8086 => x"9d",
          8087 => x"49",
          8088 => x"a5",
          8089 => x"a9",
          8090 => x"ad",
          8091 => x"b1",
          8092 => x"b5",
          8093 => x"b9",
          8094 => x"bd",
          8095 => x"c1",
          8096 => x"c5",
          8097 => x"c9",
          8098 => x"cd",
          8099 => x"d1",
          8100 => x"d5",
          8101 => x"d9",
          8102 => x"dd",
          8103 => x"e1",
          8104 => x"e5",
          8105 => x"e9",
          8106 => x"ed",
          8107 => x"f1",
          8108 => x"f5",
          8109 => x"f9",
          8110 => x"fd",
          8111 => x"2e",
          8112 => x"5b",
          8113 => x"22",
          8114 => x"3e",
          8115 => x"00",
          8116 => x"01",
          8117 => x"10",
          8118 => x"00",
          8119 => x"00",
          8120 => x"01",
          8121 => x"04",
          8122 => x"10",
          8123 => x"00",
          8124 => x"69",
          8125 => x"00",
          8126 => x"69",
          8127 => x"6c",
          8128 => x"69",
          8129 => x"00",
          8130 => x"6c",
          8131 => x"00",
          8132 => x"65",
          8133 => x"00",
          8134 => x"63",
          8135 => x"72",
          8136 => x"63",
          8137 => x"00",
          8138 => x"64",
          8139 => x"00",
          8140 => x"64",
          8141 => x"00",
          8142 => x"65",
          8143 => x"65",
          8144 => x"65",
          8145 => x"69",
          8146 => x"69",
          8147 => x"66",
          8148 => x"66",
          8149 => x"61",
          8150 => x"00",
          8151 => x"6d",
          8152 => x"65",
          8153 => x"72",
          8154 => x"65",
          8155 => x"00",
          8156 => x"6e",
          8157 => x"00",
          8158 => x"65",
          8159 => x"00",
          8160 => x"62",
          8161 => x"63",
          8162 => x"69",
          8163 => x"45",
          8164 => x"72",
          8165 => x"6e",
          8166 => x"6e",
          8167 => x"65",
          8168 => x"72",
          8169 => x"00",
          8170 => x"69",
          8171 => x"6e",
          8172 => x"72",
          8173 => x"79",
          8174 => x"00",
          8175 => x"6f",
          8176 => x"6c",
          8177 => x"6f",
          8178 => x"2e",
          8179 => x"6f",
          8180 => x"74",
          8181 => x"6f",
          8182 => x"2e",
          8183 => x"6e",
          8184 => x"69",
          8185 => x"69",
          8186 => x"61",
          8187 => x"0a",
          8188 => x"63",
          8189 => x"73",
          8190 => x"6e",
          8191 => x"2e",
          8192 => x"69",
          8193 => x"61",
          8194 => x"61",
          8195 => x"65",
          8196 => x"74",
          8197 => x"00",
          8198 => x"69",
          8199 => x"68",
          8200 => x"6c",
          8201 => x"6e",
          8202 => x"69",
          8203 => x"00",
          8204 => x"44",
          8205 => x"20",
          8206 => x"74",
          8207 => x"72",
          8208 => x"63",
          8209 => x"2e",
          8210 => x"72",
          8211 => x"20",
          8212 => x"62",
          8213 => x"69",
          8214 => x"6e",
          8215 => x"69",
          8216 => x"00",
          8217 => x"69",
          8218 => x"6e",
          8219 => x"65",
          8220 => x"6c",
          8221 => x"0a",
          8222 => x"6f",
          8223 => x"6d",
          8224 => x"69",
          8225 => x"20",
          8226 => x"65",
          8227 => x"74",
          8228 => x"66",
          8229 => x"64",
          8230 => x"20",
          8231 => x"6b",
          8232 => x"00",
          8233 => x"6f",
          8234 => x"74",
          8235 => x"6f",
          8236 => x"64",
          8237 => x"00",
          8238 => x"69",
          8239 => x"75",
          8240 => x"6f",
          8241 => x"61",
          8242 => x"6e",
          8243 => x"6e",
          8244 => x"6c",
          8245 => x"0a",
          8246 => x"69",
          8247 => x"69",
          8248 => x"6f",
          8249 => x"64",
          8250 => x"00",
          8251 => x"6e",
          8252 => x"66",
          8253 => x"65",
          8254 => x"6d",
          8255 => x"72",
          8256 => x"00",
          8257 => x"6f",
          8258 => x"61",
          8259 => x"6f",
          8260 => x"20",
          8261 => x"65",
          8262 => x"00",
          8263 => x"61",
          8264 => x"65",
          8265 => x"73",
          8266 => x"63",
          8267 => x"65",
          8268 => x"0a",
          8269 => x"75",
          8270 => x"73",
          8271 => x"00",
          8272 => x"6e",
          8273 => x"77",
          8274 => x"72",
          8275 => x"2e",
          8276 => x"25",
          8277 => x"62",
          8278 => x"73",
          8279 => x"20",
          8280 => x"25",
          8281 => x"62",
          8282 => x"73",
          8283 => x"63",
          8284 => x"00",
          8285 => x"65",
          8286 => x"00",
          8287 => x"30",
          8288 => x"00",
          8289 => x"20",
          8290 => x"30",
          8291 => x"00",
          8292 => x"20",
          8293 => x"20",
          8294 => x"00",
          8295 => x"30",
          8296 => x"00",
          8297 => x"20",
          8298 => x"7c",
          8299 => x"0d",
          8300 => x"4f",
          8301 => x"2a",
          8302 => x"73",
          8303 => x"00",
          8304 => x"30",
          8305 => x"2f",
          8306 => x"30",
          8307 => x"31",
          8308 => x"00",
          8309 => x"5a",
          8310 => x"20",
          8311 => x"20",
          8312 => x"78",
          8313 => x"73",
          8314 => x"20",
          8315 => x"0a",
          8316 => x"50",
          8317 => x"6e",
          8318 => x"72",
          8319 => x"20",
          8320 => x"64",
          8321 => x"0a",
          8322 => x"69",
          8323 => x"20",
          8324 => x"65",
          8325 => x"70",
          8326 => x"00",
          8327 => x"53",
          8328 => x"6e",
          8329 => x"72",
          8330 => x"0a",
          8331 => x"4f",
          8332 => x"20",
          8333 => x"69",
          8334 => x"72",
          8335 => x"74",
          8336 => x"4f",
          8337 => x"20",
          8338 => x"69",
          8339 => x"72",
          8340 => x"74",
          8341 => x"41",
          8342 => x"20",
          8343 => x"69",
          8344 => x"72",
          8345 => x"74",
          8346 => x"41",
          8347 => x"20",
          8348 => x"69",
          8349 => x"72",
          8350 => x"74",
          8351 => x"41",
          8352 => x"20",
          8353 => x"69",
          8354 => x"72",
          8355 => x"74",
          8356 => x"41",
          8357 => x"20",
          8358 => x"69",
          8359 => x"72",
          8360 => x"74",
          8361 => x"65",
          8362 => x"6e",
          8363 => x"70",
          8364 => x"6d",
          8365 => x"2e",
          8366 => x"00",
          8367 => x"6e",
          8368 => x"69",
          8369 => x"74",
          8370 => x"72",
          8371 => x"0a",
          8372 => x"75",
          8373 => x"78",
          8374 => x"62",
          8375 => x"00",
          8376 => x"3a",
          8377 => x"61",
          8378 => x"64",
          8379 => x"20",
          8380 => x"74",
          8381 => x"69",
          8382 => x"73",
          8383 => x"61",
          8384 => x"30",
          8385 => x"6c",
          8386 => x"65",
          8387 => x"69",
          8388 => x"61",
          8389 => x"6c",
          8390 => x"0a",
          8391 => x"20",
          8392 => x"6c",
          8393 => x"69",
          8394 => x"2e",
          8395 => x"00",
          8396 => x"6f",
          8397 => x"6e",
          8398 => x"2e",
          8399 => x"6f",
          8400 => x"72",
          8401 => x"2e",
          8402 => x"00",
          8403 => x"30",
          8404 => x"28",
          8405 => x"78",
          8406 => x"25",
          8407 => x"78",
          8408 => x"38",
          8409 => x"00",
          8410 => x"75",
          8411 => x"4d",
          8412 => x"72",
          8413 => x"00",
          8414 => x"43",
          8415 => x"6c",
          8416 => x"2e",
          8417 => x"30",
          8418 => x"25",
          8419 => x"2d",
          8420 => x"3f",
          8421 => x"00",
          8422 => x"30",
          8423 => x"25",
          8424 => x"2d",
          8425 => x"30",
          8426 => x"25",
          8427 => x"2d",
          8428 => x"78",
          8429 => x"74",
          8430 => x"20",
          8431 => x"65",
          8432 => x"25",
          8433 => x"20",
          8434 => x"0a",
          8435 => x"61",
          8436 => x"6e",
          8437 => x"6f",
          8438 => x"40",
          8439 => x"38",
          8440 => x"2e",
          8441 => x"00",
          8442 => x"61",
          8443 => x"72",
          8444 => x"72",
          8445 => x"20",
          8446 => x"65",
          8447 => x"64",
          8448 => x"00",
          8449 => x"65",
          8450 => x"72",
          8451 => x"67",
          8452 => x"70",
          8453 => x"61",
          8454 => x"6e",
          8455 => x"0a",
          8456 => x"6f",
          8457 => x"72",
          8458 => x"6f",
          8459 => x"67",
          8460 => x"0a",
          8461 => x"50",
          8462 => x"69",
          8463 => x"64",
          8464 => x"73",
          8465 => x"2e",
          8466 => x"00",
          8467 => x"64",
          8468 => x"73",
          8469 => x"00",
          8470 => x"64",
          8471 => x"73",
          8472 => x"61",
          8473 => x"6f",
          8474 => x"6e",
          8475 => x"00",
          8476 => x"75",
          8477 => x"6e",
          8478 => x"2e",
          8479 => x"6e",
          8480 => x"69",
          8481 => x"69",
          8482 => x"72",
          8483 => x"74",
          8484 => x"2e",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"01",
          8491 => x"00",
          8492 => x"01",
          8493 => x"81",
          8494 => x"00",
          8495 => x"7f",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"f5",
          8501 => x"f5",
          8502 => x"f5",
          8503 => x"00",
          8504 => x"01",
          8505 => x"01",
          8506 => x"01",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"02",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"04",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"14",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"2b",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"30",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"3c",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"3d",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"3f",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"40",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"41",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"42",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"43",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"50",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"51",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"54",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"55",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"79",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"78",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"82",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"83",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"85",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"87",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"8c",
          8601 => x"00",
          8602 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"e0",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"0b",
            11 => x"2d",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"c4",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"d0",
           163 => x"10",
           164 => x"06",
           165 => x"88",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"cf",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"81",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"04",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"51",
           267 => x"73",
           268 => x"73",
           269 => x"81",
           270 => x"10",
           271 => x"07",
           272 => x"0c",
           273 => x"72",
           274 => x"81",
           275 => x"09",
           276 => x"71",
           277 => x"0a",
           278 => x"72",
           279 => x"51",
           280 => x"9f",
           281 => x"a4",
           282 => x"80",
           283 => x"05",
           284 => x"0b",
           285 => x"04",
           286 => x"9e",
           287 => x"80",
           288 => x"fe",
           289 => x"00",
           290 => x"94",
           291 => x"0d",
           292 => x"08",
           293 => x"52",
           294 => x"05",
           295 => x"de",
           296 => x"70",
           297 => x"85",
           298 => x"0c",
           299 => x"02",
           300 => x"3d",
           301 => x"94",
           302 => x"08",
           303 => x"88",
           304 => x"82",
           305 => x"08",
           306 => x"54",
           307 => x"94",
           308 => x"08",
           309 => x"f9",
           310 => x"0b",
           311 => x"05",
           312 => x"88",
           313 => x"25",
           314 => x"08",
           315 => x"30",
           316 => x"05",
           317 => x"94",
           318 => x"0c",
           319 => x"05",
           320 => x"81",
           321 => x"f4",
           322 => x"08",
           323 => x"94",
           324 => x"0c",
           325 => x"05",
           326 => x"ab",
           327 => x"8c",
           328 => x"94",
           329 => x"0c",
           330 => x"08",
           331 => x"94",
           332 => x"08",
           333 => x"0b",
           334 => x"05",
           335 => x"f0",
           336 => x"08",
           337 => x"80",
           338 => x"8c",
           339 => x"94",
           340 => x"08",
           341 => x"3f",
           342 => x"94",
           343 => x"0c",
           344 => x"fc",
           345 => x"2e",
           346 => x"08",
           347 => x"30",
           348 => x"05",
           349 => x"f8",
           350 => x"88",
           351 => x"3d",
           352 => x"04",
           353 => x"94",
           354 => x"0d",
           355 => x"08",
           356 => x"94",
           357 => x"08",
           358 => x"38",
           359 => x"05",
           360 => x"08",
           361 => x"81",
           362 => x"fc",
           363 => x"08",
           364 => x"80",
           365 => x"94",
           366 => x"08",
           367 => x"8c",
           368 => x"53",
           369 => x"05",
           370 => x"08",
           371 => x"51",
           372 => x"08",
           373 => x"f8",
           374 => x"94",
           375 => x"08",
           376 => x"38",
           377 => x"05",
           378 => x"08",
           379 => x"94",
           380 => x"08",
           381 => x"54",
           382 => x"94",
           383 => x"08",
           384 => x"fd",
           385 => x"0b",
           386 => x"05",
           387 => x"94",
           388 => x"0c",
           389 => x"05",
           390 => x"88",
           391 => x"ac",
           392 => x"fc",
           393 => x"2e",
           394 => x"0b",
           395 => x"05",
           396 => x"38",
           397 => x"05",
           398 => x"08",
           399 => x"94",
           400 => x"08",
           401 => x"fc",
           402 => x"39",
           403 => x"05",
           404 => x"80",
           405 => x"08",
           406 => x"94",
           407 => x"08",
           408 => x"94",
           409 => x"08",
           410 => x"05",
           411 => x"08",
           412 => x"94",
           413 => x"08",
           414 => x"05",
           415 => x"08",
           416 => x"94",
           417 => x"08",
           418 => x"08",
           419 => x"94",
           420 => x"08",
           421 => x"08",
           422 => x"ff",
           423 => x"08",
           424 => x"80",
           425 => x"94",
           426 => x"08",
           427 => x"f4",
           428 => x"8d",
           429 => x"f8",
           430 => x"94",
           431 => x"0c",
           432 => x"f4",
           433 => x"0c",
           434 => x"94",
           435 => x"3d",
           436 => x"0b",
           437 => x"8c",
           438 => x"87",
           439 => x"0c",
           440 => x"c0",
           441 => x"87",
           442 => x"08",
           443 => x"51",
           444 => x"2e",
           445 => x"c0",
           446 => x"51",
           447 => x"87",
           448 => x"08",
           449 => x"06",
           450 => x"38",
           451 => x"8c",
           452 => x"80",
           453 => x"71",
           454 => x"9f",
           455 => x"0b",
           456 => x"33",
           457 => x"3d",
           458 => x"3d",
           459 => x"7d",
           460 => x"80",
           461 => x"0b",
           462 => x"81",
           463 => x"82",
           464 => x"2e",
           465 => x"81",
           466 => x"0b",
           467 => x"8c",
           468 => x"c0",
           469 => x"84",
           470 => x"92",
           471 => x"c0",
           472 => x"70",
           473 => x"81",
           474 => x"53",
           475 => x"a7",
           476 => x"92",
           477 => x"81",
           478 => x"79",
           479 => x"51",
           480 => x"90",
           481 => x"2e",
           482 => x"76",
           483 => x"58",
           484 => x"54",
           485 => x"72",
           486 => x"70",
           487 => x"38",
           488 => x"8c",
           489 => x"ff",
           490 => x"c0",
           491 => x"51",
           492 => x"81",
           493 => x"92",
           494 => x"c0",
           495 => x"70",
           496 => x"51",
           497 => x"80",
           498 => x"80",
           499 => x"70",
           500 => x"81",
           501 => x"87",
           502 => x"08",
           503 => x"2e",
           504 => x"83",
           505 => x"71",
           506 => x"3d",
           507 => x"3d",
           508 => x"11",
           509 => x"71",
           510 => x"88",
           511 => x"84",
           512 => x"fd",
           513 => x"83",
           514 => x"12",
           515 => x"2b",
           516 => x"07",
           517 => x"70",
           518 => x"2b",
           519 => x"07",
           520 => x"53",
           521 => x"52",
           522 => x"04",
           523 => x"79",
           524 => x"9f",
           525 => x"57",
           526 => x"80",
           527 => x"88",
           528 => x"80",
           529 => x"33",
           530 => x"2e",
           531 => x"83",
           532 => x"80",
           533 => x"54",
           534 => x"fe",
           535 => x"88",
           536 => x"08",
           537 => x"3d",
           538 => x"fd",
           539 => x"08",
           540 => x"51",
           541 => x"88",
           542 => x"ff",
           543 => x"39",
           544 => x"82",
           545 => x"06",
           546 => x"2a",
           547 => x"05",
           548 => x"70",
           549 => x"92",
           550 => x"8e",
           551 => x"fe",
           552 => x"08",
           553 => x"55",
           554 => x"55",
           555 => x"89",
           556 => x"fb",
           557 => x"0b",
           558 => x"08",
           559 => x"12",
           560 => x"55",
           561 => x"56",
           562 => x"8d",
           563 => x"33",
           564 => x"94",
           565 => x"57",
           566 => x"0c",
           567 => x"04",
           568 => x"75",
           569 => x"0b",
           570 => x"f4",
           571 => x"51",
           572 => x"83",
           573 => x"06",
           574 => x"14",
           575 => x"3f",
           576 => x"2b",
           577 => x"51",
           578 => x"88",
           579 => x"ff",
           580 => x"88",
           581 => x"0d",
           582 => x"0d",
           583 => x"0b",
           584 => x"55",
           585 => x"23",
           586 => x"53",
           587 => x"88",
           588 => x"08",
           589 => x"38",
           590 => x"39",
           591 => x"73",
           592 => x"83",
           593 => x"06",
           594 => x"14",
           595 => x"8c",
           596 => x"80",
           597 => x"72",
           598 => x"3f",
           599 => x"85",
           600 => x"08",
           601 => x"16",
           602 => x"71",
           603 => x"3d",
           604 => x"3d",
           605 => x"0b",
           606 => x"08",
           607 => x"05",
           608 => x"ff",
           609 => x"57",
           610 => x"2e",
           611 => x"15",
           612 => x"86",
           613 => x"80",
           614 => x"8f",
           615 => x"80",
           616 => x"13",
           617 => x"8c",
           618 => x"72",
           619 => x"0b",
           620 => x"57",
           621 => x"27",
           622 => x"39",
           623 => x"ff",
           624 => x"2a",
           625 => x"a8",
           626 => x"fc",
           627 => x"52",
           628 => x"27",
           629 => x"52",
           630 => x"17",
           631 => x"38",
           632 => x"16",
           633 => x"51",
           634 => x"88",
           635 => x"0c",
           636 => x"80",
           637 => x"0c",
           638 => x"04",
           639 => x"60",
           640 => x"5e",
           641 => x"55",
           642 => x"09",
           643 => x"38",
           644 => x"44",
           645 => x"62",
           646 => x"56",
           647 => x"09",
           648 => x"38",
           649 => x"80",
           650 => x"0c",
           651 => x"51",
           652 => x"26",
           653 => x"51",
           654 => x"88",
           655 => x"7d",
           656 => x"39",
           657 => x"1d",
           658 => x"5a",
           659 => x"a0",
           660 => x"05",
           661 => x"15",
           662 => x"2e",
           663 => x"ef",
           664 => x"59",
           665 => x"08",
           666 => x"81",
           667 => x"ff",
           668 => x"70",
           669 => x"32",
           670 => x"73",
           671 => x"25",
           672 => x"52",
           673 => x"57",
           674 => x"c7",
           675 => x"2e",
           676 => x"83",
           677 => x"77",
           678 => x"07",
           679 => x"2e",
           680 => x"88",
           681 => x"78",
           682 => x"30",
           683 => x"9f",
           684 => x"57",
           685 => x"9b",
           686 => x"8b",
           687 => x"39",
           688 => x"70",
           689 => x"72",
           690 => x"57",
           691 => x"34",
           692 => x"7a",
           693 => x"80",
           694 => x"26",
           695 => x"55",
           696 => x"34",
           697 => x"b1",
           698 => x"80",
           699 => x"54",
           700 => x"85",
           701 => x"06",
           702 => x"1c",
           703 => x"51",
           704 => x"88",
           705 => x"08",
           706 => x"7c",
           707 => x"80",
           708 => x"38",
           709 => x"70",
           710 => x"81",
           711 => x"56",
           712 => x"8b",
           713 => x"08",
           714 => x"5b",
           715 => x"18",
           716 => x"2e",
           717 => x"70",
           718 => x"33",
           719 => x"05",
           720 => x"71",
           721 => x"56",
           722 => x"e2",
           723 => x"75",
           724 => x"38",
           725 => x"9a",
           726 => x"39",
           727 => x"88",
           728 => x"83",
           729 => x"84",
           730 => x"11",
           731 => x"74",
           732 => x"1d",
           733 => x"2a",
           734 => x"51",
           735 => x"89",
           736 => x"92",
           737 => x"8e",
           738 => x"fa",
           739 => x"08",
           740 => x"fd",
           741 => x"88",
           742 => x"0d",
           743 => x"0d",
           744 => x"57",
           745 => x"fe",
           746 => x"76",
           747 => x"3f",
           748 => x"08",
           749 => x"76",
           750 => x"3f",
           751 => x"ff",
           752 => x"82",
           753 => x"d4",
           754 => x"81",
           755 => x"38",
           756 => x"53",
           757 => x"51",
           758 => x"88",
           759 => x"08",
           760 => x"51",
           761 => x"88",
           762 => x"ff",
           763 => x"81",
           764 => x"a9",
           765 => x"80",
           766 => x"52",
           767 => x"aa",
           768 => x"56",
           769 => x"38",
           770 => x"e2",
           771 => x"83",
           772 => x"55",
           773 => x"c6",
           774 => x"81",
           775 => x"0c",
           776 => x"04",
           777 => x"65",
           778 => x"0b",
           779 => x"f4",
           780 => x"3f",
           781 => x"06",
           782 => x"74",
           783 => x"74",
           784 => x"3d",
           785 => x"5a",
           786 => x"88",
           787 => x"06",
           788 => x"2e",
           789 => x"b3",
           790 => x"83",
           791 => x"52",
           792 => x"c6",
           793 => x"ab",
           794 => x"33",
           795 => x"2e",
           796 => x"3d",
           797 => x"f7",
           798 => x"08",
           799 => x"76",
           800 => x"99",
           801 => x"81",
           802 => x"76",
           803 => x"81",
           804 => x"81",
           805 => x"39",
           806 => x"86",
           807 => x"82",
           808 => x"54",
           809 => x"52",
           810 => x"fe",
           811 => x"88",
           812 => x"38",
           813 => x"05",
           814 => x"3f",
           815 => x"ff",
           816 => x"77",
           817 => x"3d",
           818 => x"f6",
           819 => x"08",
           820 => x"05",
           821 => x"29",
           822 => x"ad",
           823 => x"52",
           824 => x"8a",
           825 => x"83",
           826 => x"7a",
           827 => x"0c",
           828 => x"82",
           829 => x"3d",
           830 => x"f5",
           831 => x"08",
           832 => x"95",
           833 => x"51",
           834 => x"88",
           835 => x"ff",
           836 => x"8c",
           837 => x"ef",
           838 => x"e7",
           839 => x"56",
           840 => x"ca",
           841 => x"83",
           842 => x"76",
           843 => x"31",
           844 => x"70",
           845 => x"1d",
           846 => x"71",
           847 => x"5c",
           848 => x"c4",
           849 => x"82",
           850 => x"1b",
           851 => x"e0",
           852 => x"56",
           853 => x"fe",
           854 => x"82",
           855 => x"f6",
           856 => x"38",
           857 => x"39",
           858 => x"80",
           859 => x"38",
           860 => x"76",
           861 => x"81",
           862 => x"95",
           863 => x"51",
           864 => x"88",
           865 => x"0c",
           866 => x"19",
           867 => x"1a",
           868 => x"ff",
           869 => x"1a",
           870 => x"84",
           871 => x"1b",
           872 => x"0b",
           873 => x"78",
           874 => x"9f",
           875 => x"56",
           876 => x"95",
           877 => x"ea",
           878 => x"0b",
           879 => x"08",
           880 => x"74",
           881 => x"df",
           882 => x"81",
           883 => x"3d",
           884 => x"69",
           885 => x"70",
           886 => x"05",
           887 => x"3f",
           888 => x"88",
           889 => x"38",
           890 => x"54",
           891 => x"93",
           892 => x"05",
           893 => x"2a",
           894 => x"51",
           895 => x"80",
           896 => x"83",
           897 => x"75",
           898 => x"3f",
           899 => x"16",
           900 => x"dc",
           901 => x"eb",
           902 => x"9c",
           903 => x"98",
           904 => x"0b",
           905 => x"73",
           906 => x"3d",
           907 => x"3d",
           908 => x"7e",
           909 => x"9f",
           910 => x"5b",
           911 => x"7b",
           912 => x"75",
           913 => x"d1",
           914 => x"33",
           915 => x"84",
           916 => x"2e",
           917 => x"91",
           918 => x"17",
           919 => x"80",
           920 => x"34",
           921 => x"b1",
           922 => x"08",
           923 => x"31",
           924 => x"27",
           925 => x"58",
           926 => x"81",
           927 => x"16",
           928 => x"ff",
           929 => x"74",
           930 => x"82",
           931 => x"05",
           932 => x"06",
           933 => x"06",
           934 => x"9e",
           935 => x"38",
           936 => x"55",
           937 => x"16",
           938 => x"80",
           939 => x"55",
           940 => x"ff",
           941 => x"a4",
           942 => x"16",
           943 => x"f3",
           944 => x"55",
           945 => x"2e",
           946 => x"88",
           947 => x"17",
           948 => x"08",
           949 => x"84",
           950 => x"51",
           951 => x"27",
           952 => x"55",
           953 => x"16",
           954 => x"06",
           955 => x"08",
           956 => x"f0",
           957 => x"08",
           958 => x"98",
           959 => x"98",
           960 => x"75",
           961 => x"16",
           962 => x"78",
           963 => x"e8",
           964 => x"59",
           965 => x"80",
           966 => x"0c",
           967 => x"04",
           968 => x"87",
           969 => x"08",
           970 => x"80",
           971 => x"ea",
           972 => x"08",
           973 => x"c0",
           974 => x"56",
           975 => x"80",
           976 => x"ea",
           977 => x"88",
           978 => x"c0",
           979 => x"87",
           980 => x"08",
           981 => x"80",
           982 => x"ea",
           983 => x"08",
           984 => x"c0",
           985 => x"56",
           986 => x"80",
           987 => x"ea",
           988 => x"88",
           989 => x"c0",
           990 => x"8c",
           991 => x"87",
           992 => x"0c",
           993 => x"0b",
           994 => x"94",
           995 => x"51",
           996 => x"88",
           997 => x"9f",
           998 => x"9b",
           999 => x"ae",
          1000 => x"0b",
          1001 => x"c0",
          1002 => x"55",
          1003 => x"05",
          1004 => x"52",
          1005 => x"f6",
          1006 => x"8d",
          1007 => x"73",
          1008 => x"38",
          1009 => x"e4",
          1010 => x"54",
          1011 => x"54",
          1012 => x"00",
          1013 => x"ff",
          1014 => x"ff",
          1015 => x"ff",
          1016 => x"42",
          1017 => x"54",
          1018 => x"2e",
          1019 => x"00",
          1020 => x"01",
          2048 => x"0b",
          2049 => x"80",
          2050 => x"80",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"0b",
          2057 => x"80",
          2058 => x"80",
          2059 => x"0b",
          2060 => x"95",
          2061 => x"80",
          2062 => x"0b",
          2063 => x"b5",
          2064 => x"80",
          2065 => x"0b",
          2066 => x"d5",
          2067 => x"80",
          2068 => x"0b",
          2069 => x"f5",
          2070 => x"80",
          2071 => x"0b",
          2072 => x"95",
          2073 => x"80",
          2074 => x"0b",
          2075 => x"b5",
          2076 => x"80",
          2077 => x"0b",
          2078 => x"d5",
          2079 => x"80",
          2080 => x"0b",
          2081 => x"f5",
          2082 => x"80",
          2083 => x"0b",
          2084 => x"95",
          2085 => x"80",
          2086 => x"0b",
          2087 => x"b5",
          2088 => x"80",
          2089 => x"0b",
          2090 => x"d5",
          2091 => x"80",
          2092 => x"0b",
          2093 => x"f5",
          2094 => x"80",
          2095 => x"0b",
          2096 => x"95",
          2097 => x"80",
          2098 => x"0b",
          2099 => x"b5",
          2100 => x"80",
          2101 => x"0b",
          2102 => x"d5",
          2103 => x"80",
          2104 => x"0b",
          2105 => x"f5",
          2106 => x"80",
          2107 => x"0b",
          2108 => x"95",
          2109 => x"80",
          2110 => x"0b",
          2111 => x"b5",
          2112 => x"80",
          2113 => x"0b",
          2114 => x"d5",
          2115 => x"80",
          2116 => x"0b",
          2117 => x"f5",
          2118 => x"80",
          2119 => x"0b",
          2120 => x"95",
          2121 => x"80",
          2122 => x"0b",
          2123 => x"b5",
          2124 => x"80",
          2125 => x"0b",
          2126 => x"d5",
          2127 => x"80",
          2128 => x"0b",
          2129 => x"f5",
          2130 => x"80",
          2131 => x"00",
          2132 => x"00",
          2133 => x"00",
          2134 => x"00",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"00",
          2177 => x"04",
          2178 => x"0c",
          2179 => x"2d",
          2180 => x"08",
          2181 => x"04",
          2182 => x"0c",
          2183 => x"2d",
          2184 => x"08",
          2185 => x"04",
          2186 => x"0c",
          2187 => x"2d",
          2188 => x"08",
          2189 => x"04",
          2190 => x"0c",
          2191 => x"2d",
          2192 => x"08",
          2193 => x"04",
          2194 => x"0c",
          2195 => x"2d",
          2196 => x"08",
          2197 => x"04",
          2198 => x"0c",
          2199 => x"2d",
          2200 => x"08",
          2201 => x"04",
          2202 => x"0c",
          2203 => x"2d",
          2204 => x"08",
          2205 => x"04",
          2206 => x"0c",
          2207 => x"2d",
          2208 => x"08",
          2209 => x"04",
          2210 => x"0c",
          2211 => x"2d",
          2212 => x"08",
          2213 => x"04",
          2214 => x"0c",
          2215 => x"2d",
          2216 => x"08",
          2217 => x"04",
          2218 => x"0c",
          2219 => x"2d",
          2220 => x"08",
          2221 => x"04",
          2222 => x"0c",
          2223 => x"2d",
          2224 => x"08",
          2225 => x"04",
          2226 => x"0c",
          2227 => x"2d",
          2228 => x"08",
          2229 => x"04",
          2230 => x"0c",
          2231 => x"2d",
          2232 => x"08",
          2233 => x"04",
          2234 => x"0c",
          2235 => x"2d",
          2236 => x"08",
          2237 => x"04",
          2238 => x"0c",
          2239 => x"2d",
          2240 => x"08",
          2241 => x"04",
          2242 => x"0c",
          2243 => x"2d",
          2244 => x"08",
          2245 => x"04",
          2246 => x"0c",
          2247 => x"2d",
          2248 => x"08",
          2249 => x"04",
          2250 => x"0c",
          2251 => x"2d",
          2252 => x"08",
          2253 => x"04",
          2254 => x"0c",
          2255 => x"2d",
          2256 => x"08",
          2257 => x"04",
          2258 => x"0c",
          2259 => x"2d",
          2260 => x"08",
          2261 => x"04",
          2262 => x"0c",
          2263 => x"2d",
          2264 => x"08",
          2265 => x"04",
          2266 => x"0c",
          2267 => x"2d",
          2268 => x"08",
          2269 => x"04",
          2270 => x"0c",
          2271 => x"2d",
          2272 => x"08",
          2273 => x"04",
          2274 => x"0c",
          2275 => x"2d",
          2276 => x"08",
          2277 => x"04",
          2278 => x"0c",
          2279 => x"2d",
          2280 => x"08",
          2281 => x"04",
          2282 => x"0c",
          2283 => x"2d",
          2284 => x"08",
          2285 => x"04",
          2286 => x"0c",
          2287 => x"2d",
          2288 => x"08",
          2289 => x"04",
          2290 => x"0c",
          2291 => x"2d",
          2292 => x"08",
          2293 => x"04",
          2294 => x"0c",
          2295 => x"2d",
          2296 => x"08",
          2297 => x"04",
          2298 => x"0c",
          2299 => x"2d",
          2300 => x"08",
          2301 => x"04",
          2302 => x"0c",
          2303 => x"2d",
          2304 => x"08",
          2305 => x"04",
          2306 => x"0c",
          2307 => x"2d",
          2308 => x"08",
          2309 => x"04",
          2310 => x"0c",
          2311 => x"2d",
          2312 => x"08",
          2313 => x"04",
          2314 => x"0c",
          2315 => x"2d",
          2316 => x"08",
          2317 => x"04",
          2318 => x"0c",
          2319 => x"2d",
          2320 => x"08",
          2321 => x"04",
          2322 => x"0c",
          2323 => x"2d",
          2324 => x"08",
          2325 => x"04",
          2326 => x"0c",
          2327 => x"2d",
          2328 => x"08",
          2329 => x"04",
          2330 => x"0c",
          2331 => x"2d",
          2332 => x"08",
          2333 => x"04",
          2334 => x"0c",
          2335 => x"2d",
          2336 => x"08",
          2337 => x"04",
          2338 => x"0c",
          2339 => x"2d",
          2340 => x"08",
          2341 => x"04",
          2342 => x"0c",
          2343 => x"2d",
          2344 => x"08",
          2345 => x"04",
          2346 => x"0c",
          2347 => x"2d",
          2348 => x"08",
          2349 => x"04",
          2350 => x"0c",
          2351 => x"2d",
          2352 => x"08",
          2353 => x"04",
          2354 => x"0c",
          2355 => x"2d",
          2356 => x"08",
          2357 => x"04",
          2358 => x"0c",
          2359 => x"2d",
          2360 => x"08",
          2361 => x"04",
          2362 => x"0c",
          2363 => x"2d",
          2364 => x"08",
          2365 => x"04",
          2366 => x"0c",
          2367 => x"2d",
          2368 => x"08",
          2369 => x"04",
          2370 => x"0c",
          2371 => x"2d",
          2372 => x"08",
          2373 => x"04",
          2374 => x"70",
          2375 => x"27",
          2376 => x"71",
          2377 => x"53",
          2378 => x"80",
          2379 => x"80",
          2380 => x"81",
          2381 => x"3c",
          2382 => x"f8",
          2383 => x"8c",
          2384 => x"3d",
          2385 => x"82",
          2386 => x"8c",
          2387 => x"82",
          2388 => x"88",
          2389 => x"80",
          2390 => x"8c",
          2391 => x"82",
          2392 => x"54",
          2393 => x"82",
          2394 => x"04",
          2395 => x"08",
          2396 => x"f8",
          2397 => x"0d",
          2398 => x"8c",
          2399 => x"05",
          2400 => x"8c",
          2401 => x"05",
          2402 => x"3f",
          2403 => x"08",
          2404 => x"ec",
          2405 => x"3d",
          2406 => x"f8",
          2407 => x"8c",
          2408 => x"82",
          2409 => x"fd",
          2410 => x"0b",
          2411 => x"08",
          2412 => x"80",
          2413 => x"f8",
          2414 => x"0c",
          2415 => x"08",
          2416 => x"82",
          2417 => x"88",
          2418 => x"b9",
          2419 => x"f8",
          2420 => x"08",
          2421 => x"38",
          2422 => x"8c",
          2423 => x"05",
          2424 => x"38",
          2425 => x"08",
          2426 => x"10",
          2427 => x"08",
          2428 => x"82",
          2429 => x"fc",
          2430 => x"82",
          2431 => x"fc",
          2432 => x"b8",
          2433 => x"f8",
          2434 => x"08",
          2435 => x"e1",
          2436 => x"f8",
          2437 => x"08",
          2438 => x"08",
          2439 => x"26",
          2440 => x"8c",
          2441 => x"05",
          2442 => x"f8",
          2443 => x"08",
          2444 => x"f8",
          2445 => x"0c",
          2446 => x"08",
          2447 => x"82",
          2448 => x"fc",
          2449 => x"82",
          2450 => x"f8",
          2451 => x"8c",
          2452 => x"05",
          2453 => x"82",
          2454 => x"fc",
          2455 => x"8c",
          2456 => x"05",
          2457 => x"82",
          2458 => x"8c",
          2459 => x"95",
          2460 => x"f8",
          2461 => x"08",
          2462 => x"38",
          2463 => x"08",
          2464 => x"70",
          2465 => x"08",
          2466 => x"51",
          2467 => x"8c",
          2468 => x"05",
          2469 => x"8c",
          2470 => x"05",
          2471 => x"8c",
          2472 => x"05",
          2473 => x"ec",
          2474 => x"0d",
          2475 => x"0c",
          2476 => x"0d",
          2477 => x"02",
          2478 => x"05",
          2479 => x"53",
          2480 => x"27",
          2481 => x"83",
          2482 => x"80",
          2483 => x"ff",
          2484 => x"ff",
          2485 => x"73",
          2486 => x"05",
          2487 => x"12",
          2488 => x"2e",
          2489 => x"ef",
          2490 => x"8c",
          2491 => x"3d",
          2492 => x"74",
          2493 => x"07",
          2494 => x"2b",
          2495 => x"51",
          2496 => x"a5",
          2497 => x"70",
          2498 => x"0c",
          2499 => x"84",
          2500 => x"72",
          2501 => x"05",
          2502 => x"71",
          2503 => x"53",
          2504 => x"52",
          2505 => x"dd",
          2506 => x"27",
          2507 => x"71",
          2508 => x"53",
          2509 => x"52",
          2510 => x"f2",
          2511 => x"ff",
          2512 => x"3d",
          2513 => x"70",
          2514 => x"06",
          2515 => x"70",
          2516 => x"73",
          2517 => x"56",
          2518 => x"08",
          2519 => x"38",
          2520 => x"52",
          2521 => x"81",
          2522 => x"54",
          2523 => x"9d",
          2524 => x"55",
          2525 => x"09",
          2526 => x"38",
          2527 => x"14",
          2528 => x"81",
          2529 => x"56",
          2530 => x"e5",
          2531 => x"55",
          2532 => x"06",
          2533 => x"06",
          2534 => x"82",
          2535 => x"52",
          2536 => x"0d",
          2537 => x"70",
          2538 => x"ff",
          2539 => x"f8",
          2540 => x"80",
          2541 => x"51",
          2542 => x"84",
          2543 => x"71",
          2544 => x"54",
          2545 => x"2e",
          2546 => x"75",
          2547 => x"94",
          2548 => x"82",
          2549 => x"87",
          2550 => x"fe",
          2551 => x"52",
          2552 => x"88",
          2553 => x"86",
          2554 => x"ec",
          2555 => x"06",
          2556 => x"14",
          2557 => x"80",
          2558 => x"71",
          2559 => x"0c",
          2560 => x"04",
          2561 => x"77",
          2562 => x"53",
          2563 => x"80",
          2564 => x"38",
          2565 => x"70",
          2566 => x"81",
          2567 => x"81",
          2568 => x"39",
          2569 => x"39",
          2570 => x"80",
          2571 => x"81",
          2572 => x"55",
          2573 => x"2e",
          2574 => x"55",
          2575 => x"84",
          2576 => x"38",
          2577 => x"06",
          2578 => x"2e",
          2579 => x"88",
          2580 => x"70",
          2581 => x"34",
          2582 => x"71",
          2583 => x"8c",
          2584 => x"3d",
          2585 => x"3d",
          2586 => x"72",
          2587 => x"91",
          2588 => x"fc",
          2589 => x"51",
          2590 => x"82",
          2591 => x"85",
          2592 => x"83",
          2593 => x"72",
          2594 => x"0c",
          2595 => x"04",
          2596 => x"76",
          2597 => x"ff",
          2598 => x"81",
          2599 => x"26",
          2600 => x"83",
          2601 => x"05",
          2602 => x"70",
          2603 => x"8a",
          2604 => x"33",
          2605 => x"70",
          2606 => x"fe",
          2607 => x"33",
          2608 => x"70",
          2609 => x"f2",
          2610 => x"33",
          2611 => x"70",
          2612 => x"e6",
          2613 => x"22",
          2614 => x"74",
          2615 => x"80",
          2616 => x"13",
          2617 => x"52",
          2618 => x"26",
          2619 => x"81",
          2620 => x"98",
          2621 => x"22",
          2622 => x"bc",
          2623 => x"33",
          2624 => x"b8",
          2625 => x"33",
          2626 => x"b4",
          2627 => x"33",
          2628 => x"b0",
          2629 => x"33",
          2630 => x"ac",
          2631 => x"33",
          2632 => x"a8",
          2633 => x"c0",
          2634 => x"73",
          2635 => x"a0",
          2636 => x"87",
          2637 => x"0c",
          2638 => x"82",
          2639 => x"86",
          2640 => x"f3",
          2641 => x"5b",
          2642 => x"9c",
          2643 => x"0c",
          2644 => x"bc",
          2645 => x"7b",
          2646 => x"98",
          2647 => x"79",
          2648 => x"87",
          2649 => x"08",
          2650 => x"1c",
          2651 => x"98",
          2652 => x"79",
          2653 => x"87",
          2654 => x"08",
          2655 => x"1c",
          2656 => x"98",
          2657 => x"79",
          2658 => x"87",
          2659 => x"08",
          2660 => x"1c",
          2661 => x"98",
          2662 => x"79",
          2663 => x"80",
          2664 => x"83",
          2665 => x"59",
          2666 => x"ff",
          2667 => x"1b",
          2668 => x"1b",
          2669 => x"1b",
          2670 => x"1b",
          2671 => x"1b",
          2672 => x"83",
          2673 => x"52",
          2674 => x"51",
          2675 => x"8f",
          2676 => x"ff",
          2677 => x"8f",
          2678 => x"30",
          2679 => x"51",
          2680 => x"0b",
          2681 => x"94",
          2682 => x"0d",
          2683 => x"0d",
          2684 => x"82",
          2685 => x"70",
          2686 => x"57",
          2687 => x"c0",
          2688 => x"74",
          2689 => x"38",
          2690 => x"94",
          2691 => x"70",
          2692 => x"81",
          2693 => x"52",
          2694 => x"8c",
          2695 => x"2a",
          2696 => x"51",
          2697 => x"38",
          2698 => x"70",
          2699 => x"51",
          2700 => x"8d",
          2701 => x"2a",
          2702 => x"51",
          2703 => x"be",
          2704 => x"ff",
          2705 => x"c0",
          2706 => x"70",
          2707 => x"38",
          2708 => x"90",
          2709 => x"0c",
          2710 => x"ec",
          2711 => x"0d",
          2712 => x"0d",
          2713 => x"33",
          2714 => x"89",
          2715 => x"81",
          2716 => x"55",
          2717 => x"94",
          2718 => x"80",
          2719 => x"87",
          2720 => x"51",
          2721 => x"96",
          2722 => x"06",
          2723 => x"70",
          2724 => x"38",
          2725 => x"70",
          2726 => x"51",
          2727 => x"72",
          2728 => x"81",
          2729 => x"70",
          2730 => x"38",
          2731 => x"70",
          2732 => x"51",
          2733 => x"38",
          2734 => x"06",
          2735 => x"94",
          2736 => x"80",
          2737 => x"87",
          2738 => x"52",
          2739 => x"87",
          2740 => x"f9",
          2741 => x"54",
          2742 => x"70",
          2743 => x"53",
          2744 => x"77",
          2745 => x"38",
          2746 => x"06",
          2747 => x"0b",
          2748 => x"33",
          2749 => x"06",
          2750 => x"58",
          2751 => x"84",
          2752 => x"2e",
          2753 => x"c0",
          2754 => x"70",
          2755 => x"2a",
          2756 => x"53",
          2757 => x"80",
          2758 => x"71",
          2759 => x"81",
          2760 => x"70",
          2761 => x"81",
          2762 => x"06",
          2763 => x"80",
          2764 => x"71",
          2765 => x"81",
          2766 => x"70",
          2767 => x"74",
          2768 => x"51",
          2769 => x"80",
          2770 => x"2e",
          2771 => x"c0",
          2772 => x"77",
          2773 => x"17",
          2774 => x"81",
          2775 => x"53",
          2776 => x"84",
          2777 => x"8c",
          2778 => x"3d",
          2779 => x"3d",
          2780 => x"82",
          2781 => x"70",
          2782 => x"54",
          2783 => x"94",
          2784 => x"80",
          2785 => x"87",
          2786 => x"51",
          2787 => x"82",
          2788 => x"06",
          2789 => x"70",
          2790 => x"38",
          2791 => x"06",
          2792 => x"94",
          2793 => x"80",
          2794 => x"87",
          2795 => x"52",
          2796 => x"81",
          2797 => x"8c",
          2798 => x"84",
          2799 => x"fe",
          2800 => x"0b",
          2801 => x"33",
          2802 => x"06",
          2803 => x"c0",
          2804 => x"70",
          2805 => x"38",
          2806 => x"94",
          2807 => x"70",
          2808 => x"81",
          2809 => x"51",
          2810 => x"80",
          2811 => x"72",
          2812 => x"51",
          2813 => x"80",
          2814 => x"2e",
          2815 => x"c0",
          2816 => x"71",
          2817 => x"2b",
          2818 => x"51",
          2819 => x"82",
          2820 => x"84",
          2821 => x"ff",
          2822 => x"c0",
          2823 => x"70",
          2824 => x"06",
          2825 => x"80",
          2826 => x"38",
          2827 => x"a4",
          2828 => x"98",
          2829 => x"9e",
          2830 => x"89",
          2831 => x"c0",
          2832 => x"82",
          2833 => x"87",
          2834 => x"08",
          2835 => x"0c",
          2836 => x"9c",
          2837 => x"a8",
          2838 => x"9e",
          2839 => x"89",
          2840 => x"c0",
          2841 => x"82",
          2842 => x"87",
          2843 => x"08",
          2844 => x"0c",
          2845 => x"b4",
          2846 => x"b8",
          2847 => x"9e",
          2848 => x"89",
          2849 => x"c0",
          2850 => x"82",
          2851 => x"87",
          2852 => x"08",
          2853 => x"0c",
          2854 => x"c4",
          2855 => x"c8",
          2856 => x"9e",
          2857 => x"70",
          2858 => x"23",
          2859 => x"84",
          2860 => x"d0",
          2861 => x"9e",
          2862 => x"89",
          2863 => x"c0",
          2864 => x"82",
          2865 => x"81",
          2866 => x"dc",
          2867 => x"87",
          2868 => x"08",
          2869 => x"0a",
          2870 => x"52",
          2871 => x"83",
          2872 => x"71",
          2873 => x"34",
          2874 => x"c0",
          2875 => x"70",
          2876 => x"06",
          2877 => x"70",
          2878 => x"38",
          2879 => x"82",
          2880 => x"80",
          2881 => x"9e",
          2882 => x"90",
          2883 => x"51",
          2884 => x"80",
          2885 => x"81",
          2886 => x"89",
          2887 => x"0b",
          2888 => x"90",
          2889 => x"80",
          2890 => x"52",
          2891 => x"2e",
          2892 => x"52",
          2893 => x"e0",
          2894 => x"87",
          2895 => x"08",
          2896 => x"80",
          2897 => x"52",
          2898 => x"83",
          2899 => x"71",
          2900 => x"34",
          2901 => x"c0",
          2902 => x"70",
          2903 => x"06",
          2904 => x"70",
          2905 => x"38",
          2906 => x"82",
          2907 => x"80",
          2908 => x"9e",
          2909 => x"84",
          2910 => x"51",
          2911 => x"80",
          2912 => x"81",
          2913 => x"89",
          2914 => x"0b",
          2915 => x"90",
          2916 => x"80",
          2917 => x"52",
          2918 => x"2e",
          2919 => x"52",
          2920 => x"e4",
          2921 => x"87",
          2922 => x"08",
          2923 => x"80",
          2924 => x"52",
          2925 => x"83",
          2926 => x"71",
          2927 => x"34",
          2928 => x"c0",
          2929 => x"70",
          2930 => x"06",
          2931 => x"70",
          2932 => x"38",
          2933 => x"82",
          2934 => x"80",
          2935 => x"9e",
          2936 => x"a0",
          2937 => x"52",
          2938 => x"2e",
          2939 => x"52",
          2940 => x"e7",
          2941 => x"9e",
          2942 => x"98",
          2943 => x"8a",
          2944 => x"51",
          2945 => x"e8",
          2946 => x"87",
          2947 => x"08",
          2948 => x"06",
          2949 => x"70",
          2950 => x"38",
          2951 => x"82",
          2952 => x"87",
          2953 => x"08",
          2954 => x"06",
          2955 => x"51",
          2956 => x"82",
          2957 => x"80",
          2958 => x"9e",
          2959 => x"88",
          2960 => x"52",
          2961 => x"83",
          2962 => x"71",
          2963 => x"34",
          2964 => x"90",
          2965 => x"06",
          2966 => x"82",
          2967 => x"83",
          2968 => x"fb",
          2969 => x"f6",
          2970 => x"c7",
          2971 => x"dc",
          2972 => x"80",
          2973 => x"81",
          2974 => x"85",
          2975 => x"f6",
          2976 => x"af",
          2977 => x"de",
          2978 => x"80",
          2979 => x"82",
          2980 => x"82",
          2981 => x"11",
          2982 => x"f6",
          2983 => x"f7",
          2984 => x"e3",
          2985 => x"80",
          2986 => x"82",
          2987 => x"82",
          2988 => x"11",
          2989 => x"f6",
          2990 => x"db",
          2991 => x"e0",
          2992 => x"80",
          2993 => x"82",
          2994 => x"82",
          2995 => x"11",
          2996 => x"f6",
          2997 => x"bf",
          2998 => x"e1",
          2999 => x"80",
          3000 => x"82",
          3001 => x"82",
          3002 => x"11",
          3003 => x"f7",
          3004 => x"a3",
          3005 => x"e2",
          3006 => x"80",
          3007 => x"82",
          3008 => x"82",
          3009 => x"11",
          3010 => x"f7",
          3011 => x"87",
          3012 => x"e7",
          3013 => x"80",
          3014 => x"82",
          3015 => x"52",
          3016 => x"51",
          3017 => x"82",
          3018 => x"54",
          3019 => x"8d",
          3020 => x"ec",
          3021 => x"f7",
          3022 => x"db",
          3023 => x"e9",
          3024 => x"80",
          3025 => x"82",
          3026 => x"52",
          3027 => x"51",
          3028 => x"82",
          3029 => x"54",
          3030 => x"88",
          3031 => x"b0",
          3032 => x"3f",
          3033 => x"33",
          3034 => x"2e",
          3035 => x"f8",
          3036 => x"bf",
          3037 => x"e4",
          3038 => x"80",
          3039 => x"81",
          3040 => x"83",
          3041 => x"89",
          3042 => x"73",
          3043 => x"38",
          3044 => x"51",
          3045 => x"82",
          3046 => x"54",
          3047 => x"88",
          3048 => x"e8",
          3049 => x"3f",
          3050 => x"51",
          3051 => x"82",
          3052 => x"52",
          3053 => x"51",
          3054 => x"82",
          3055 => x"52",
          3056 => x"51",
          3057 => x"82",
          3058 => x"52",
          3059 => x"51",
          3060 => x"81",
          3061 => x"82",
          3062 => x"89",
          3063 => x"81",
          3064 => x"88",
          3065 => x"89",
          3066 => x"bd",
          3067 => x"75",
          3068 => x"3f",
          3069 => x"08",
          3070 => x"29",
          3071 => x"54",
          3072 => x"ec",
          3073 => x"fa",
          3074 => x"8b",
          3075 => x"e3",
          3076 => x"80",
          3077 => x"82",
          3078 => x"56",
          3079 => x"52",
          3080 => x"95",
          3081 => x"ec",
          3082 => x"c0",
          3083 => x"31",
          3084 => x"8c",
          3085 => x"81",
          3086 => x"87",
          3087 => x"89",
          3088 => x"73",
          3089 => x"38",
          3090 => x"08",
          3091 => x"c0",
          3092 => x"e9",
          3093 => x"8c",
          3094 => x"84",
          3095 => x"71",
          3096 => x"82",
          3097 => x"52",
          3098 => x"51",
          3099 => x"82",
          3100 => x"81",
          3101 => x"3d",
          3102 => x"3d",
          3103 => x"05",
          3104 => x"52",
          3105 => x"ac",
          3106 => x"29",
          3107 => x"f5",
          3108 => x"71",
          3109 => x"fb",
          3110 => x"39",
          3111 => x"51",
          3112 => x"fb",
          3113 => x"39",
          3114 => x"51",
          3115 => x"fb",
          3116 => x"39",
          3117 => x"51",
          3118 => x"84",
          3119 => x"71",
          3120 => x"04",
          3121 => x"c0",
          3122 => x"04",
          3123 => x"08",
          3124 => x"84",
          3125 => x"3d",
          3126 => x"05",
          3127 => x"8a",
          3128 => x"06",
          3129 => x"51",
          3130 => x"8d",
          3131 => x"71",
          3132 => x"38",
          3133 => x"82",
          3134 => x"81",
          3135 => x"84",
          3136 => x"82",
          3137 => x"52",
          3138 => x"85",
          3139 => x"71",
          3140 => x"0d",
          3141 => x"0d",
          3142 => x"33",
          3143 => x"08",
          3144 => x"fc",
          3145 => x"ff",
          3146 => x"82",
          3147 => x"84",
          3148 => x"fd",
          3149 => x"54",
          3150 => x"81",
          3151 => x"53",
          3152 => x"8e",
          3153 => x"ff",
          3154 => x"14",
          3155 => x"3f",
          3156 => x"3d",
          3157 => x"3d",
          3158 => x"8c",
          3159 => x"82",
          3160 => x"56",
          3161 => x"70",
          3162 => x"53",
          3163 => x"2e",
          3164 => x"81",
          3165 => x"81",
          3166 => x"da",
          3167 => x"74",
          3168 => x"0c",
          3169 => x"04",
          3170 => x"66",
          3171 => x"78",
          3172 => x"5a",
          3173 => x"80",
          3174 => x"38",
          3175 => x"09",
          3176 => x"de",
          3177 => x"7a",
          3178 => x"5c",
          3179 => x"5b",
          3180 => x"09",
          3181 => x"38",
          3182 => x"39",
          3183 => x"09",
          3184 => x"38",
          3185 => x"70",
          3186 => x"33",
          3187 => x"2e",
          3188 => x"92",
          3189 => x"19",
          3190 => x"70",
          3191 => x"33",
          3192 => x"53",
          3193 => x"16",
          3194 => x"26",
          3195 => x"88",
          3196 => x"05",
          3197 => x"05",
          3198 => x"05",
          3199 => x"5b",
          3200 => x"80",
          3201 => x"30",
          3202 => x"80",
          3203 => x"cc",
          3204 => x"70",
          3205 => x"25",
          3206 => x"54",
          3207 => x"53",
          3208 => x"8c",
          3209 => x"07",
          3210 => x"05",
          3211 => x"5a",
          3212 => x"83",
          3213 => x"54",
          3214 => x"27",
          3215 => x"16",
          3216 => x"06",
          3217 => x"80",
          3218 => x"aa",
          3219 => x"cf",
          3220 => x"73",
          3221 => x"81",
          3222 => x"80",
          3223 => x"38",
          3224 => x"2e",
          3225 => x"81",
          3226 => x"80",
          3227 => x"8a",
          3228 => x"39",
          3229 => x"2e",
          3230 => x"73",
          3231 => x"8a",
          3232 => x"d3",
          3233 => x"80",
          3234 => x"80",
          3235 => x"ee",
          3236 => x"39",
          3237 => x"71",
          3238 => x"53",
          3239 => x"54",
          3240 => x"2e",
          3241 => x"15",
          3242 => x"33",
          3243 => x"72",
          3244 => x"81",
          3245 => x"39",
          3246 => x"56",
          3247 => x"27",
          3248 => x"51",
          3249 => x"75",
          3250 => x"72",
          3251 => x"38",
          3252 => x"df",
          3253 => x"16",
          3254 => x"7b",
          3255 => x"38",
          3256 => x"f2",
          3257 => x"77",
          3258 => x"12",
          3259 => x"53",
          3260 => x"5c",
          3261 => x"5c",
          3262 => x"5c",
          3263 => x"5c",
          3264 => x"51",
          3265 => x"fd",
          3266 => x"82",
          3267 => x"06",
          3268 => x"80",
          3269 => x"77",
          3270 => x"53",
          3271 => x"18",
          3272 => x"72",
          3273 => x"c4",
          3274 => x"70",
          3275 => x"25",
          3276 => x"55",
          3277 => x"8d",
          3278 => x"2e",
          3279 => x"30",
          3280 => x"5b",
          3281 => x"8f",
          3282 => x"7b",
          3283 => x"e4",
          3284 => x"8c",
          3285 => x"ff",
          3286 => x"75",
          3287 => x"d9",
          3288 => x"ec",
          3289 => x"74",
          3290 => x"a7",
          3291 => x"80",
          3292 => x"38",
          3293 => x"72",
          3294 => x"54",
          3295 => x"72",
          3296 => x"05",
          3297 => x"17",
          3298 => x"77",
          3299 => x"51",
          3300 => x"9f",
          3301 => x"72",
          3302 => x"79",
          3303 => x"81",
          3304 => x"72",
          3305 => x"38",
          3306 => x"05",
          3307 => x"ad",
          3308 => x"17",
          3309 => x"81",
          3310 => x"b0",
          3311 => x"38",
          3312 => x"81",
          3313 => x"06",
          3314 => x"9f",
          3315 => x"55",
          3316 => x"97",
          3317 => x"f9",
          3318 => x"81",
          3319 => x"8b",
          3320 => x"16",
          3321 => x"73",
          3322 => x"96",
          3323 => x"e0",
          3324 => x"17",
          3325 => x"33",
          3326 => x"f9",
          3327 => x"f2",
          3328 => x"16",
          3329 => x"7b",
          3330 => x"38",
          3331 => x"c6",
          3332 => x"96",
          3333 => x"fd",
          3334 => x"3d",
          3335 => x"05",
          3336 => x"52",
          3337 => x"e0",
          3338 => x"0d",
          3339 => x"0d",
          3340 => x"84",
          3341 => x"88",
          3342 => x"51",
          3343 => x"82",
          3344 => x"53",
          3345 => x"80",
          3346 => x"84",
          3347 => x"0d",
          3348 => x"0d",
          3349 => x"08",
          3350 => x"fc",
          3351 => x"88",
          3352 => x"52",
          3353 => x"3f",
          3354 => x"fc",
          3355 => x"0d",
          3356 => x"0d",
          3357 => x"8d",
          3358 => x"56",
          3359 => x"80",
          3360 => x"2e",
          3361 => x"82",
          3362 => x"52",
          3363 => x"8c",
          3364 => x"ff",
          3365 => x"80",
          3366 => x"38",
          3367 => x"b9",
          3368 => x"32",
          3369 => x"80",
          3370 => x"52",
          3371 => x"8b",
          3372 => x"2e",
          3373 => x"14",
          3374 => x"9f",
          3375 => x"38",
          3376 => x"73",
          3377 => x"38",
          3378 => x"72",
          3379 => x"14",
          3380 => x"f8",
          3381 => x"af",
          3382 => x"52",
          3383 => x"8a",
          3384 => x"3f",
          3385 => x"82",
          3386 => x"87",
          3387 => x"fe",
          3388 => x"8d",
          3389 => x"82",
          3390 => x"77",
          3391 => x"53",
          3392 => x"72",
          3393 => x"0c",
          3394 => x"04",
          3395 => x"7a",
          3396 => x"80",
          3397 => x"58",
          3398 => x"33",
          3399 => x"a0",
          3400 => x"06",
          3401 => x"13",
          3402 => x"39",
          3403 => x"09",
          3404 => x"38",
          3405 => x"11",
          3406 => x"08",
          3407 => x"54",
          3408 => x"2e",
          3409 => x"80",
          3410 => x"08",
          3411 => x"0c",
          3412 => x"33",
          3413 => x"80",
          3414 => x"38",
          3415 => x"80",
          3416 => x"38",
          3417 => x"57",
          3418 => x"0c",
          3419 => x"33",
          3420 => x"39",
          3421 => x"74",
          3422 => x"38",
          3423 => x"80",
          3424 => x"89",
          3425 => x"38",
          3426 => x"d0",
          3427 => x"55",
          3428 => x"80",
          3429 => x"39",
          3430 => x"d9",
          3431 => x"80",
          3432 => x"27",
          3433 => x"80",
          3434 => x"89",
          3435 => x"70",
          3436 => x"55",
          3437 => x"70",
          3438 => x"55",
          3439 => x"27",
          3440 => x"14",
          3441 => x"06",
          3442 => x"74",
          3443 => x"73",
          3444 => x"38",
          3445 => x"14",
          3446 => x"05",
          3447 => x"08",
          3448 => x"54",
          3449 => x"39",
          3450 => x"84",
          3451 => x"55",
          3452 => x"81",
          3453 => x"8c",
          3454 => x"3d",
          3455 => x"3d",
          3456 => x"5a",
          3457 => x"7a",
          3458 => x"08",
          3459 => x"53",
          3460 => x"09",
          3461 => x"38",
          3462 => x"0c",
          3463 => x"ad",
          3464 => x"06",
          3465 => x"76",
          3466 => x"0c",
          3467 => x"33",
          3468 => x"73",
          3469 => x"81",
          3470 => x"38",
          3471 => x"05",
          3472 => x"08",
          3473 => x"53",
          3474 => x"2e",
          3475 => x"57",
          3476 => x"2e",
          3477 => x"39",
          3478 => x"13",
          3479 => x"08",
          3480 => x"53",
          3481 => x"55",
          3482 => x"80",
          3483 => x"14",
          3484 => x"88",
          3485 => x"27",
          3486 => x"eb",
          3487 => x"53",
          3488 => x"89",
          3489 => x"38",
          3490 => x"55",
          3491 => x"8a",
          3492 => x"a0",
          3493 => x"c2",
          3494 => x"74",
          3495 => x"e0",
          3496 => x"ff",
          3497 => x"d0",
          3498 => x"ff",
          3499 => x"90",
          3500 => x"38",
          3501 => x"81",
          3502 => x"53",
          3503 => x"ca",
          3504 => x"27",
          3505 => x"77",
          3506 => x"08",
          3507 => x"0c",
          3508 => x"33",
          3509 => x"ff",
          3510 => x"80",
          3511 => x"74",
          3512 => x"79",
          3513 => x"74",
          3514 => x"0c",
          3515 => x"04",
          3516 => x"02",
          3517 => x"51",
          3518 => x"72",
          3519 => x"82",
          3520 => x"33",
          3521 => x"8c",
          3522 => x"3d",
          3523 => x"3d",
          3524 => x"05",
          3525 => x"05",
          3526 => x"56",
          3527 => x"72",
          3528 => x"e0",
          3529 => x"2b",
          3530 => x"8c",
          3531 => x"88",
          3532 => x"2e",
          3533 => x"88",
          3534 => x"0c",
          3535 => x"8c",
          3536 => x"71",
          3537 => x"87",
          3538 => x"0c",
          3539 => x"08",
          3540 => x"51",
          3541 => x"2e",
          3542 => x"c0",
          3543 => x"51",
          3544 => x"71",
          3545 => x"80",
          3546 => x"92",
          3547 => x"98",
          3548 => x"70",
          3549 => x"38",
          3550 => x"f4",
          3551 => x"89",
          3552 => x"51",
          3553 => x"ec",
          3554 => x"0d",
          3555 => x"0d",
          3556 => x"02",
          3557 => x"05",
          3558 => x"58",
          3559 => x"52",
          3560 => x"3f",
          3561 => x"08",
          3562 => x"54",
          3563 => x"be",
          3564 => x"75",
          3565 => x"c0",
          3566 => x"87",
          3567 => x"12",
          3568 => x"84",
          3569 => x"40",
          3570 => x"85",
          3571 => x"98",
          3572 => x"7d",
          3573 => x"0c",
          3574 => x"85",
          3575 => x"06",
          3576 => x"71",
          3577 => x"38",
          3578 => x"71",
          3579 => x"05",
          3580 => x"19",
          3581 => x"a2",
          3582 => x"71",
          3583 => x"38",
          3584 => x"83",
          3585 => x"38",
          3586 => x"8a",
          3587 => x"98",
          3588 => x"71",
          3589 => x"c0",
          3590 => x"52",
          3591 => x"87",
          3592 => x"80",
          3593 => x"81",
          3594 => x"c0",
          3595 => x"53",
          3596 => x"82",
          3597 => x"71",
          3598 => x"1a",
          3599 => x"84",
          3600 => x"19",
          3601 => x"06",
          3602 => x"79",
          3603 => x"38",
          3604 => x"80",
          3605 => x"87",
          3606 => x"26",
          3607 => x"73",
          3608 => x"06",
          3609 => x"2e",
          3610 => x"52",
          3611 => x"82",
          3612 => x"8f",
          3613 => x"f3",
          3614 => x"62",
          3615 => x"05",
          3616 => x"57",
          3617 => x"83",
          3618 => x"52",
          3619 => x"3f",
          3620 => x"08",
          3621 => x"54",
          3622 => x"2e",
          3623 => x"81",
          3624 => x"74",
          3625 => x"c0",
          3626 => x"87",
          3627 => x"12",
          3628 => x"84",
          3629 => x"5f",
          3630 => x"0b",
          3631 => x"8c",
          3632 => x"0c",
          3633 => x"80",
          3634 => x"70",
          3635 => x"81",
          3636 => x"54",
          3637 => x"8c",
          3638 => x"81",
          3639 => x"7c",
          3640 => x"58",
          3641 => x"70",
          3642 => x"52",
          3643 => x"8a",
          3644 => x"98",
          3645 => x"71",
          3646 => x"c0",
          3647 => x"52",
          3648 => x"87",
          3649 => x"80",
          3650 => x"81",
          3651 => x"c0",
          3652 => x"53",
          3653 => x"82",
          3654 => x"71",
          3655 => x"19",
          3656 => x"81",
          3657 => x"ff",
          3658 => x"19",
          3659 => x"78",
          3660 => x"38",
          3661 => x"80",
          3662 => x"87",
          3663 => x"26",
          3664 => x"73",
          3665 => x"06",
          3666 => x"2e",
          3667 => x"52",
          3668 => x"82",
          3669 => x"8f",
          3670 => x"fa",
          3671 => x"02",
          3672 => x"05",
          3673 => x"05",
          3674 => x"71",
          3675 => x"57",
          3676 => x"82",
          3677 => x"81",
          3678 => x"54",
          3679 => x"38",
          3680 => x"c0",
          3681 => x"81",
          3682 => x"2e",
          3683 => x"71",
          3684 => x"38",
          3685 => x"87",
          3686 => x"11",
          3687 => x"80",
          3688 => x"80",
          3689 => x"83",
          3690 => x"38",
          3691 => x"72",
          3692 => x"2a",
          3693 => x"51",
          3694 => x"80",
          3695 => x"87",
          3696 => x"08",
          3697 => x"38",
          3698 => x"8c",
          3699 => x"96",
          3700 => x"0c",
          3701 => x"8c",
          3702 => x"08",
          3703 => x"51",
          3704 => x"38",
          3705 => x"56",
          3706 => x"80",
          3707 => x"85",
          3708 => x"77",
          3709 => x"83",
          3710 => x"75",
          3711 => x"8c",
          3712 => x"3d",
          3713 => x"3d",
          3714 => x"11",
          3715 => x"71",
          3716 => x"82",
          3717 => x"53",
          3718 => x"0d",
          3719 => x"0d",
          3720 => x"33",
          3721 => x"71",
          3722 => x"88",
          3723 => x"14",
          3724 => x"07",
          3725 => x"33",
          3726 => x"8c",
          3727 => x"53",
          3728 => x"52",
          3729 => x"04",
          3730 => x"73",
          3731 => x"92",
          3732 => x"52",
          3733 => x"81",
          3734 => x"70",
          3735 => x"70",
          3736 => x"3d",
          3737 => x"3d",
          3738 => x"52",
          3739 => x"70",
          3740 => x"34",
          3741 => x"51",
          3742 => x"81",
          3743 => x"70",
          3744 => x"70",
          3745 => x"05",
          3746 => x"88",
          3747 => x"72",
          3748 => x"0d",
          3749 => x"0d",
          3750 => x"54",
          3751 => x"80",
          3752 => x"71",
          3753 => x"53",
          3754 => x"81",
          3755 => x"ff",
          3756 => x"39",
          3757 => x"04",
          3758 => x"75",
          3759 => x"52",
          3760 => x"70",
          3761 => x"34",
          3762 => x"70",
          3763 => x"3d",
          3764 => x"3d",
          3765 => x"79",
          3766 => x"74",
          3767 => x"56",
          3768 => x"81",
          3769 => x"71",
          3770 => x"16",
          3771 => x"52",
          3772 => x"86",
          3773 => x"2e",
          3774 => x"82",
          3775 => x"86",
          3776 => x"fe",
          3777 => x"76",
          3778 => x"39",
          3779 => x"8a",
          3780 => x"51",
          3781 => x"71",
          3782 => x"33",
          3783 => x"0c",
          3784 => x"04",
          3785 => x"8c",
          3786 => x"80",
          3787 => x"ec",
          3788 => x"3d",
          3789 => x"80",
          3790 => x"33",
          3791 => x"7a",
          3792 => x"38",
          3793 => x"16",
          3794 => x"16",
          3795 => x"17",
          3796 => x"fa",
          3797 => x"8c",
          3798 => x"2e",
          3799 => x"b7",
          3800 => x"ec",
          3801 => x"34",
          3802 => x"70",
          3803 => x"31",
          3804 => x"59",
          3805 => x"77",
          3806 => x"82",
          3807 => x"74",
          3808 => x"81",
          3809 => x"81",
          3810 => x"53",
          3811 => x"16",
          3812 => x"e3",
          3813 => x"81",
          3814 => x"8c",
          3815 => x"3d",
          3816 => x"3d",
          3817 => x"56",
          3818 => x"74",
          3819 => x"2e",
          3820 => x"51",
          3821 => x"82",
          3822 => x"57",
          3823 => x"08",
          3824 => x"54",
          3825 => x"16",
          3826 => x"33",
          3827 => x"3f",
          3828 => x"08",
          3829 => x"38",
          3830 => x"57",
          3831 => x"0c",
          3832 => x"ec",
          3833 => x"0d",
          3834 => x"0d",
          3835 => x"57",
          3836 => x"82",
          3837 => x"58",
          3838 => x"08",
          3839 => x"76",
          3840 => x"83",
          3841 => x"06",
          3842 => x"84",
          3843 => x"78",
          3844 => x"81",
          3845 => x"38",
          3846 => x"82",
          3847 => x"52",
          3848 => x"52",
          3849 => x"3f",
          3850 => x"52",
          3851 => x"51",
          3852 => x"84",
          3853 => x"d2",
          3854 => x"fc",
          3855 => x"8a",
          3856 => x"52",
          3857 => x"51",
          3858 => x"90",
          3859 => x"84",
          3860 => x"fc",
          3861 => x"17",
          3862 => x"a0",
          3863 => x"86",
          3864 => x"08",
          3865 => x"b0",
          3866 => x"55",
          3867 => x"81",
          3868 => x"f8",
          3869 => x"84",
          3870 => x"53",
          3871 => x"17",
          3872 => x"d7",
          3873 => x"ec",
          3874 => x"83",
          3875 => x"77",
          3876 => x"0c",
          3877 => x"04",
          3878 => x"77",
          3879 => x"12",
          3880 => x"55",
          3881 => x"56",
          3882 => x"8d",
          3883 => x"22",
          3884 => x"ac",
          3885 => x"57",
          3886 => x"8c",
          3887 => x"3d",
          3888 => x"3d",
          3889 => x"70",
          3890 => x"57",
          3891 => x"81",
          3892 => x"98",
          3893 => x"81",
          3894 => x"74",
          3895 => x"72",
          3896 => x"f5",
          3897 => x"24",
          3898 => x"81",
          3899 => x"81",
          3900 => x"83",
          3901 => x"38",
          3902 => x"76",
          3903 => x"70",
          3904 => x"16",
          3905 => x"74",
          3906 => x"96",
          3907 => x"ec",
          3908 => x"38",
          3909 => x"06",
          3910 => x"33",
          3911 => x"89",
          3912 => x"08",
          3913 => x"54",
          3914 => x"fc",
          3915 => x"8c",
          3916 => x"fe",
          3917 => x"ff",
          3918 => x"11",
          3919 => x"2b",
          3920 => x"81",
          3921 => x"2a",
          3922 => x"51",
          3923 => x"e2",
          3924 => x"ff",
          3925 => x"da",
          3926 => x"2a",
          3927 => x"05",
          3928 => x"fc",
          3929 => x"8c",
          3930 => x"c6",
          3931 => x"83",
          3932 => x"05",
          3933 => x"f9",
          3934 => x"8c",
          3935 => x"ff",
          3936 => x"ae",
          3937 => x"2a",
          3938 => x"05",
          3939 => x"fc",
          3940 => x"8c",
          3941 => x"38",
          3942 => x"83",
          3943 => x"05",
          3944 => x"f8",
          3945 => x"8c",
          3946 => x"0a",
          3947 => x"39",
          3948 => x"82",
          3949 => x"89",
          3950 => x"f8",
          3951 => x"7c",
          3952 => x"56",
          3953 => x"77",
          3954 => x"38",
          3955 => x"08",
          3956 => x"38",
          3957 => x"72",
          3958 => x"9d",
          3959 => x"24",
          3960 => x"81",
          3961 => x"82",
          3962 => x"83",
          3963 => x"38",
          3964 => x"76",
          3965 => x"70",
          3966 => x"18",
          3967 => x"76",
          3968 => x"9e",
          3969 => x"ec",
          3970 => x"8c",
          3971 => x"d9",
          3972 => x"ff",
          3973 => x"05",
          3974 => x"81",
          3975 => x"54",
          3976 => x"80",
          3977 => x"77",
          3978 => x"f0",
          3979 => x"8f",
          3980 => x"51",
          3981 => x"34",
          3982 => x"17",
          3983 => x"2a",
          3984 => x"05",
          3985 => x"fa",
          3986 => x"8c",
          3987 => x"82",
          3988 => x"81",
          3989 => x"83",
          3990 => x"b4",
          3991 => x"2a",
          3992 => x"8f",
          3993 => x"2a",
          3994 => x"f0",
          3995 => x"06",
          3996 => x"72",
          3997 => x"ec",
          3998 => x"2a",
          3999 => x"05",
          4000 => x"fa",
          4001 => x"8c",
          4002 => x"82",
          4003 => x"80",
          4004 => x"83",
          4005 => x"52",
          4006 => x"fe",
          4007 => x"b4",
          4008 => x"a4",
          4009 => x"76",
          4010 => x"17",
          4011 => x"75",
          4012 => x"3f",
          4013 => x"08",
          4014 => x"ec",
          4015 => x"77",
          4016 => x"77",
          4017 => x"fc",
          4018 => x"b4",
          4019 => x"51",
          4020 => x"c9",
          4021 => x"ec",
          4022 => x"06",
          4023 => x"72",
          4024 => x"3f",
          4025 => x"17",
          4026 => x"8c",
          4027 => x"3d",
          4028 => x"3d",
          4029 => x"7e",
          4030 => x"56",
          4031 => x"75",
          4032 => x"74",
          4033 => x"27",
          4034 => x"80",
          4035 => x"ff",
          4036 => x"75",
          4037 => x"3f",
          4038 => x"08",
          4039 => x"ec",
          4040 => x"38",
          4041 => x"54",
          4042 => x"81",
          4043 => x"39",
          4044 => x"08",
          4045 => x"39",
          4046 => x"51",
          4047 => x"82",
          4048 => x"58",
          4049 => x"08",
          4050 => x"c7",
          4051 => x"ec",
          4052 => x"d2",
          4053 => x"ec",
          4054 => x"cf",
          4055 => x"74",
          4056 => x"fc",
          4057 => x"8c",
          4058 => x"38",
          4059 => x"fe",
          4060 => x"08",
          4061 => x"74",
          4062 => x"38",
          4063 => x"17",
          4064 => x"33",
          4065 => x"73",
          4066 => x"77",
          4067 => x"26",
          4068 => x"80",
          4069 => x"8c",
          4070 => x"3d",
          4071 => x"3d",
          4072 => x"71",
          4073 => x"5b",
          4074 => x"8c",
          4075 => x"77",
          4076 => x"38",
          4077 => x"78",
          4078 => x"81",
          4079 => x"79",
          4080 => x"f9",
          4081 => x"55",
          4082 => x"ec",
          4083 => x"e0",
          4084 => x"ec",
          4085 => x"8c",
          4086 => x"2e",
          4087 => x"98",
          4088 => x"8c",
          4089 => x"82",
          4090 => x"58",
          4091 => x"70",
          4092 => x"80",
          4093 => x"38",
          4094 => x"09",
          4095 => x"e2",
          4096 => x"56",
          4097 => x"76",
          4098 => x"82",
          4099 => x"7a",
          4100 => x"3f",
          4101 => x"8c",
          4102 => x"2e",
          4103 => x"86",
          4104 => x"ec",
          4105 => x"8c",
          4106 => x"70",
          4107 => x"07",
          4108 => x"7c",
          4109 => x"ec",
          4110 => x"51",
          4111 => x"81",
          4112 => x"8c",
          4113 => x"2e",
          4114 => x"17",
          4115 => x"74",
          4116 => x"73",
          4117 => x"27",
          4118 => x"58",
          4119 => x"80",
          4120 => x"56",
          4121 => x"98",
          4122 => x"26",
          4123 => x"56",
          4124 => x"81",
          4125 => x"52",
          4126 => x"c6",
          4127 => x"ec",
          4128 => x"b8",
          4129 => x"82",
          4130 => x"81",
          4131 => x"06",
          4132 => x"8c",
          4133 => x"82",
          4134 => x"09",
          4135 => x"72",
          4136 => x"70",
          4137 => x"51",
          4138 => x"80",
          4139 => x"78",
          4140 => x"06",
          4141 => x"73",
          4142 => x"39",
          4143 => x"52",
          4144 => x"f7",
          4145 => x"ec",
          4146 => x"ec",
          4147 => x"82",
          4148 => x"07",
          4149 => x"55",
          4150 => x"2e",
          4151 => x"80",
          4152 => x"75",
          4153 => x"76",
          4154 => x"3f",
          4155 => x"08",
          4156 => x"38",
          4157 => x"0c",
          4158 => x"fe",
          4159 => x"08",
          4160 => x"74",
          4161 => x"ff",
          4162 => x"0c",
          4163 => x"81",
          4164 => x"84",
          4165 => x"39",
          4166 => x"81",
          4167 => x"8c",
          4168 => x"8c",
          4169 => x"ec",
          4170 => x"39",
          4171 => x"55",
          4172 => x"ec",
          4173 => x"0d",
          4174 => x"0d",
          4175 => x"55",
          4176 => x"82",
          4177 => x"58",
          4178 => x"8c",
          4179 => x"d8",
          4180 => x"74",
          4181 => x"3f",
          4182 => x"08",
          4183 => x"08",
          4184 => x"59",
          4185 => x"77",
          4186 => x"70",
          4187 => x"c8",
          4188 => x"84",
          4189 => x"56",
          4190 => x"58",
          4191 => x"97",
          4192 => x"75",
          4193 => x"52",
          4194 => x"51",
          4195 => x"82",
          4196 => x"80",
          4197 => x"8a",
          4198 => x"32",
          4199 => x"72",
          4200 => x"2a",
          4201 => x"56",
          4202 => x"ec",
          4203 => x"0d",
          4204 => x"0d",
          4205 => x"08",
          4206 => x"74",
          4207 => x"26",
          4208 => x"74",
          4209 => x"72",
          4210 => x"74",
          4211 => x"88",
          4212 => x"73",
          4213 => x"33",
          4214 => x"27",
          4215 => x"16",
          4216 => x"9b",
          4217 => x"2a",
          4218 => x"88",
          4219 => x"58",
          4220 => x"80",
          4221 => x"16",
          4222 => x"0c",
          4223 => x"8a",
          4224 => x"89",
          4225 => x"72",
          4226 => x"38",
          4227 => x"51",
          4228 => x"82",
          4229 => x"54",
          4230 => x"08",
          4231 => x"38",
          4232 => x"8c",
          4233 => x"8b",
          4234 => x"08",
          4235 => x"08",
          4236 => x"82",
          4237 => x"74",
          4238 => x"cb",
          4239 => x"75",
          4240 => x"3f",
          4241 => x"08",
          4242 => x"73",
          4243 => x"98",
          4244 => x"82",
          4245 => x"2e",
          4246 => x"39",
          4247 => x"39",
          4248 => x"13",
          4249 => x"74",
          4250 => x"16",
          4251 => x"18",
          4252 => x"77",
          4253 => x"0c",
          4254 => x"04",
          4255 => x"7a",
          4256 => x"12",
          4257 => x"59",
          4258 => x"80",
          4259 => x"86",
          4260 => x"98",
          4261 => x"14",
          4262 => x"55",
          4263 => x"81",
          4264 => x"83",
          4265 => x"77",
          4266 => x"81",
          4267 => x"0c",
          4268 => x"55",
          4269 => x"76",
          4270 => x"17",
          4271 => x"74",
          4272 => x"9b",
          4273 => x"39",
          4274 => x"ff",
          4275 => x"2a",
          4276 => x"81",
          4277 => x"52",
          4278 => x"e6",
          4279 => x"ec",
          4280 => x"55",
          4281 => x"8c",
          4282 => x"80",
          4283 => x"55",
          4284 => x"08",
          4285 => x"f4",
          4286 => x"08",
          4287 => x"08",
          4288 => x"38",
          4289 => x"77",
          4290 => x"84",
          4291 => x"39",
          4292 => x"52",
          4293 => x"86",
          4294 => x"ec",
          4295 => x"55",
          4296 => x"08",
          4297 => x"c4",
          4298 => x"82",
          4299 => x"81",
          4300 => x"81",
          4301 => x"ec",
          4302 => x"b0",
          4303 => x"ec",
          4304 => x"51",
          4305 => x"82",
          4306 => x"a0",
          4307 => x"15",
          4308 => x"75",
          4309 => x"3f",
          4310 => x"08",
          4311 => x"76",
          4312 => x"77",
          4313 => x"9c",
          4314 => x"55",
          4315 => x"ec",
          4316 => x"0d",
          4317 => x"0d",
          4318 => x"08",
          4319 => x"80",
          4320 => x"fc",
          4321 => x"8c",
          4322 => x"82",
          4323 => x"80",
          4324 => x"8c",
          4325 => x"98",
          4326 => x"78",
          4327 => x"3f",
          4328 => x"08",
          4329 => x"ec",
          4330 => x"38",
          4331 => x"08",
          4332 => x"70",
          4333 => x"58",
          4334 => x"2e",
          4335 => x"83",
          4336 => x"82",
          4337 => x"55",
          4338 => x"81",
          4339 => x"07",
          4340 => x"2e",
          4341 => x"16",
          4342 => x"2e",
          4343 => x"88",
          4344 => x"82",
          4345 => x"56",
          4346 => x"51",
          4347 => x"82",
          4348 => x"54",
          4349 => x"08",
          4350 => x"9b",
          4351 => x"2e",
          4352 => x"83",
          4353 => x"73",
          4354 => x"0c",
          4355 => x"04",
          4356 => x"76",
          4357 => x"54",
          4358 => x"82",
          4359 => x"83",
          4360 => x"76",
          4361 => x"53",
          4362 => x"2e",
          4363 => x"90",
          4364 => x"51",
          4365 => x"82",
          4366 => x"90",
          4367 => x"53",
          4368 => x"ec",
          4369 => x"0d",
          4370 => x"0d",
          4371 => x"83",
          4372 => x"54",
          4373 => x"55",
          4374 => x"3f",
          4375 => x"51",
          4376 => x"2e",
          4377 => x"8b",
          4378 => x"2a",
          4379 => x"51",
          4380 => x"86",
          4381 => x"f7",
          4382 => x"7d",
          4383 => x"75",
          4384 => x"98",
          4385 => x"2e",
          4386 => x"98",
          4387 => x"78",
          4388 => x"3f",
          4389 => x"08",
          4390 => x"ec",
          4391 => x"38",
          4392 => x"70",
          4393 => x"73",
          4394 => x"58",
          4395 => x"8b",
          4396 => x"bf",
          4397 => x"ff",
          4398 => x"53",
          4399 => x"34",
          4400 => x"08",
          4401 => x"e5",
          4402 => x"81",
          4403 => x"2e",
          4404 => x"70",
          4405 => x"57",
          4406 => x"9e",
          4407 => x"2e",
          4408 => x"8c",
          4409 => x"df",
          4410 => x"72",
          4411 => x"81",
          4412 => x"76",
          4413 => x"2e",
          4414 => x"52",
          4415 => x"fc",
          4416 => x"ec",
          4417 => x"8c",
          4418 => x"38",
          4419 => x"fe",
          4420 => x"39",
          4421 => x"16",
          4422 => x"8c",
          4423 => x"3d",
          4424 => x"3d",
          4425 => x"08",
          4426 => x"52",
          4427 => x"c5",
          4428 => x"ec",
          4429 => x"8c",
          4430 => x"38",
          4431 => x"52",
          4432 => x"de",
          4433 => x"ec",
          4434 => x"8c",
          4435 => x"38",
          4436 => x"8c",
          4437 => x"9c",
          4438 => x"ea",
          4439 => x"53",
          4440 => x"9c",
          4441 => x"ea",
          4442 => x"0b",
          4443 => x"74",
          4444 => x"0c",
          4445 => x"04",
          4446 => x"75",
          4447 => x"12",
          4448 => x"53",
          4449 => x"9a",
          4450 => x"ec",
          4451 => x"9c",
          4452 => x"e5",
          4453 => x"0b",
          4454 => x"85",
          4455 => x"fa",
          4456 => x"7a",
          4457 => x"0b",
          4458 => x"98",
          4459 => x"2e",
          4460 => x"80",
          4461 => x"55",
          4462 => x"17",
          4463 => x"33",
          4464 => x"51",
          4465 => x"2e",
          4466 => x"85",
          4467 => x"06",
          4468 => x"e5",
          4469 => x"2e",
          4470 => x"8b",
          4471 => x"70",
          4472 => x"34",
          4473 => x"71",
          4474 => x"05",
          4475 => x"15",
          4476 => x"27",
          4477 => x"15",
          4478 => x"80",
          4479 => x"34",
          4480 => x"52",
          4481 => x"88",
          4482 => x"17",
          4483 => x"52",
          4484 => x"3f",
          4485 => x"08",
          4486 => x"12",
          4487 => x"3f",
          4488 => x"08",
          4489 => x"98",
          4490 => x"da",
          4491 => x"ec",
          4492 => x"23",
          4493 => x"04",
          4494 => x"7f",
          4495 => x"5b",
          4496 => x"33",
          4497 => x"73",
          4498 => x"38",
          4499 => x"80",
          4500 => x"38",
          4501 => x"8c",
          4502 => x"08",
          4503 => x"aa",
          4504 => x"41",
          4505 => x"33",
          4506 => x"73",
          4507 => x"81",
          4508 => x"81",
          4509 => x"dc",
          4510 => x"70",
          4511 => x"07",
          4512 => x"73",
          4513 => x"88",
          4514 => x"70",
          4515 => x"73",
          4516 => x"38",
          4517 => x"ab",
          4518 => x"52",
          4519 => x"91",
          4520 => x"ec",
          4521 => x"98",
          4522 => x"61",
          4523 => x"5a",
          4524 => x"a0",
          4525 => x"e7",
          4526 => x"70",
          4527 => x"79",
          4528 => x"73",
          4529 => x"81",
          4530 => x"38",
          4531 => x"33",
          4532 => x"ae",
          4533 => x"70",
          4534 => x"82",
          4535 => x"51",
          4536 => x"54",
          4537 => x"79",
          4538 => x"74",
          4539 => x"57",
          4540 => x"af",
          4541 => x"70",
          4542 => x"51",
          4543 => x"dc",
          4544 => x"73",
          4545 => x"38",
          4546 => x"82",
          4547 => x"19",
          4548 => x"54",
          4549 => x"82",
          4550 => x"54",
          4551 => x"78",
          4552 => x"81",
          4553 => x"54",
          4554 => x"81",
          4555 => x"af",
          4556 => x"77",
          4557 => x"70",
          4558 => x"25",
          4559 => x"07",
          4560 => x"51",
          4561 => x"2e",
          4562 => x"39",
          4563 => x"80",
          4564 => x"33",
          4565 => x"73",
          4566 => x"81",
          4567 => x"81",
          4568 => x"dc",
          4569 => x"70",
          4570 => x"07",
          4571 => x"73",
          4572 => x"b5",
          4573 => x"2e",
          4574 => x"83",
          4575 => x"76",
          4576 => x"07",
          4577 => x"2e",
          4578 => x"8b",
          4579 => x"77",
          4580 => x"30",
          4581 => x"71",
          4582 => x"53",
          4583 => x"55",
          4584 => x"38",
          4585 => x"5c",
          4586 => x"75",
          4587 => x"73",
          4588 => x"38",
          4589 => x"06",
          4590 => x"11",
          4591 => x"75",
          4592 => x"3f",
          4593 => x"08",
          4594 => x"38",
          4595 => x"33",
          4596 => x"54",
          4597 => x"e6",
          4598 => x"8c",
          4599 => x"2e",
          4600 => x"ff",
          4601 => x"74",
          4602 => x"38",
          4603 => x"75",
          4604 => x"17",
          4605 => x"57",
          4606 => x"a7",
          4607 => x"81",
          4608 => x"e5",
          4609 => x"8c",
          4610 => x"38",
          4611 => x"54",
          4612 => x"89",
          4613 => x"70",
          4614 => x"57",
          4615 => x"54",
          4616 => x"81",
          4617 => x"f7",
          4618 => x"7e",
          4619 => x"2e",
          4620 => x"33",
          4621 => x"e5",
          4622 => x"06",
          4623 => x"7a",
          4624 => x"a0",
          4625 => x"38",
          4626 => x"55",
          4627 => x"84",
          4628 => x"39",
          4629 => x"8b",
          4630 => x"7b",
          4631 => x"7a",
          4632 => x"3f",
          4633 => x"08",
          4634 => x"ec",
          4635 => x"38",
          4636 => x"52",
          4637 => x"aa",
          4638 => x"ec",
          4639 => x"8c",
          4640 => x"c2",
          4641 => x"08",
          4642 => x"55",
          4643 => x"ff",
          4644 => x"15",
          4645 => x"54",
          4646 => x"34",
          4647 => x"70",
          4648 => x"81",
          4649 => x"58",
          4650 => x"8b",
          4651 => x"74",
          4652 => x"3f",
          4653 => x"08",
          4654 => x"38",
          4655 => x"51",
          4656 => x"ff",
          4657 => x"ab",
          4658 => x"55",
          4659 => x"bb",
          4660 => x"2e",
          4661 => x"80",
          4662 => x"85",
          4663 => x"06",
          4664 => x"58",
          4665 => x"80",
          4666 => x"75",
          4667 => x"73",
          4668 => x"b5",
          4669 => x"0b",
          4670 => x"80",
          4671 => x"39",
          4672 => x"54",
          4673 => x"85",
          4674 => x"75",
          4675 => x"81",
          4676 => x"73",
          4677 => x"1b",
          4678 => x"2a",
          4679 => x"51",
          4680 => x"80",
          4681 => x"90",
          4682 => x"ff",
          4683 => x"05",
          4684 => x"f5",
          4685 => x"8c",
          4686 => x"1c",
          4687 => x"39",
          4688 => x"ec",
          4689 => x"0d",
          4690 => x"0d",
          4691 => x"7b",
          4692 => x"73",
          4693 => x"55",
          4694 => x"2e",
          4695 => x"75",
          4696 => x"57",
          4697 => x"26",
          4698 => x"ba",
          4699 => x"70",
          4700 => x"ba",
          4701 => x"06",
          4702 => x"73",
          4703 => x"70",
          4704 => x"51",
          4705 => x"89",
          4706 => x"82",
          4707 => x"ff",
          4708 => x"56",
          4709 => x"2e",
          4710 => x"80",
          4711 => x"ac",
          4712 => x"08",
          4713 => x"76",
          4714 => x"58",
          4715 => x"81",
          4716 => x"ff",
          4717 => x"53",
          4718 => x"26",
          4719 => x"13",
          4720 => x"06",
          4721 => x"9f",
          4722 => x"99",
          4723 => x"e0",
          4724 => x"ff",
          4725 => x"72",
          4726 => x"2a",
          4727 => x"72",
          4728 => x"06",
          4729 => x"ff",
          4730 => x"30",
          4731 => x"70",
          4732 => x"07",
          4733 => x"9f",
          4734 => x"54",
          4735 => x"80",
          4736 => x"81",
          4737 => x"59",
          4738 => x"25",
          4739 => x"8b",
          4740 => x"24",
          4741 => x"76",
          4742 => x"78",
          4743 => x"82",
          4744 => x"51",
          4745 => x"ec",
          4746 => x"0d",
          4747 => x"0d",
          4748 => x"0b",
          4749 => x"ff",
          4750 => x"0c",
          4751 => x"51",
          4752 => x"84",
          4753 => x"ec",
          4754 => x"38",
          4755 => x"51",
          4756 => x"82",
          4757 => x"83",
          4758 => x"54",
          4759 => x"82",
          4760 => x"09",
          4761 => x"e3",
          4762 => x"b4",
          4763 => x"57",
          4764 => x"2e",
          4765 => x"83",
          4766 => x"74",
          4767 => x"70",
          4768 => x"25",
          4769 => x"51",
          4770 => x"38",
          4771 => x"2e",
          4772 => x"b5",
          4773 => x"81",
          4774 => x"80",
          4775 => x"e0",
          4776 => x"8c",
          4777 => x"82",
          4778 => x"80",
          4779 => x"85",
          4780 => x"f0",
          4781 => x"16",
          4782 => x"3f",
          4783 => x"08",
          4784 => x"ec",
          4785 => x"83",
          4786 => x"74",
          4787 => x"0c",
          4788 => x"04",
          4789 => x"61",
          4790 => x"80",
          4791 => x"58",
          4792 => x"0c",
          4793 => x"e1",
          4794 => x"ec",
          4795 => x"56",
          4796 => x"8c",
          4797 => x"86",
          4798 => x"8c",
          4799 => x"29",
          4800 => x"05",
          4801 => x"53",
          4802 => x"80",
          4803 => x"38",
          4804 => x"76",
          4805 => x"74",
          4806 => x"72",
          4807 => x"38",
          4808 => x"51",
          4809 => x"82",
          4810 => x"81",
          4811 => x"81",
          4812 => x"72",
          4813 => x"80",
          4814 => x"38",
          4815 => x"70",
          4816 => x"53",
          4817 => x"86",
          4818 => x"a7",
          4819 => x"34",
          4820 => x"34",
          4821 => x"14",
          4822 => x"b2",
          4823 => x"ec",
          4824 => x"06",
          4825 => x"54",
          4826 => x"72",
          4827 => x"76",
          4828 => x"38",
          4829 => x"70",
          4830 => x"53",
          4831 => x"85",
          4832 => x"70",
          4833 => x"5b",
          4834 => x"82",
          4835 => x"81",
          4836 => x"76",
          4837 => x"81",
          4838 => x"38",
          4839 => x"56",
          4840 => x"83",
          4841 => x"70",
          4842 => x"80",
          4843 => x"83",
          4844 => x"dc",
          4845 => x"8c",
          4846 => x"76",
          4847 => x"05",
          4848 => x"16",
          4849 => x"56",
          4850 => x"d7",
          4851 => x"8d",
          4852 => x"72",
          4853 => x"54",
          4854 => x"57",
          4855 => x"95",
          4856 => x"73",
          4857 => x"3f",
          4858 => x"08",
          4859 => x"57",
          4860 => x"89",
          4861 => x"56",
          4862 => x"d7",
          4863 => x"76",
          4864 => x"f1",
          4865 => x"76",
          4866 => x"e9",
          4867 => x"51",
          4868 => x"82",
          4869 => x"83",
          4870 => x"53",
          4871 => x"2e",
          4872 => x"84",
          4873 => x"ca",
          4874 => x"da",
          4875 => x"ec",
          4876 => x"ff",
          4877 => x"8d",
          4878 => x"14",
          4879 => x"3f",
          4880 => x"08",
          4881 => x"15",
          4882 => x"14",
          4883 => x"34",
          4884 => x"33",
          4885 => x"81",
          4886 => x"54",
          4887 => x"72",
          4888 => x"91",
          4889 => x"ff",
          4890 => x"29",
          4891 => x"33",
          4892 => x"72",
          4893 => x"72",
          4894 => x"38",
          4895 => x"06",
          4896 => x"2e",
          4897 => x"56",
          4898 => x"80",
          4899 => x"da",
          4900 => x"8c",
          4901 => x"82",
          4902 => x"88",
          4903 => x"8f",
          4904 => x"56",
          4905 => x"38",
          4906 => x"51",
          4907 => x"82",
          4908 => x"83",
          4909 => x"55",
          4910 => x"80",
          4911 => x"da",
          4912 => x"8c",
          4913 => x"80",
          4914 => x"da",
          4915 => x"8c",
          4916 => x"ff",
          4917 => x"8d",
          4918 => x"2e",
          4919 => x"88",
          4920 => x"14",
          4921 => x"05",
          4922 => x"75",
          4923 => x"38",
          4924 => x"52",
          4925 => x"51",
          4926 => x"3f",
          4927 => x"08",
          4928 => x"ec",
          4929 => x"82",
          4930 => x"8c",
          4931 => x"ff",
          4932 => x"26",
          4933 => x"57",
          4934 => x"f5",
          4935 => x"82",
          4936 => x"f5",
          4937 => x"81",
          4938 => x"8d",
          4939 => x"2e",
          4940 => x"82",
          4941 => x"16",
          4942 => x"16",
          4943 => x"70",
          4944 => x"7a",
          4945 => x"0c",
          4946 => x"83",
          4947 => x"06",
          4948 => x"de",
          4949 => x"ae",
          4950 => x"ec",
          4951 => x"ff",
          4952 => x"56",
          4953 => x"38",
          4954 => x"38",
          4955 => x"51",
          4956 => x"82",
          4957 => x"a8",
          4958 => x"82",
          4959 => x"39",
          4960 => x"80",
          4961 => x"38",
          4962 => x"15",
          4963 => x"53",
          4964 => x"8d",
          4965 => x"15",
          4966 => x"76",
          4967 => x"51",
          4968 => x"13",
          4969 => x"8d",
          4970 => x"15",
          4971 => x"c5",
          4972 => x"90",
          4973 => x"0b",
          4974 => x"ff",
          4975 => x"15",
          4976 => x"2e",
          4977 => x"81",
          4978 => x"e4",
          4979 => x"b6",
          4980 => x"ec",
          4981 => x"ff",
          4982 => x"81",
          4983 => x"06",
          4984 => x"81",
          4985 => x"51",
          4986 => x"82",
          4987 => x"80",
          4988 => x"8c",
          4989 => x"15",
          4990 => x"14",
          4991 => x"3f",
          4992 => x"08",
          4993 => x"06",
          4994 => x"d4",
          4995 => x"81",
          4996 => x"38",
          4997 => x"d8",
          4998 => x"8c",
          4999 => x"8b",
          5000 => x"2e",
          5001 => x"b3",
          5002 => x"14",
          5003 => x"3f",
          5004 => x"08",
          5005 => x"e4",
          5006 => x"81",
          5007 => x"84",
          5008 => x"d7",
          5009 => x"8c",
          5010 => x"15",
          5011 => x"14",
          5012 => x"3f",
          5013 => x"08",
          5014 => x"76",
          5015 => x"8d",
          5016 => x"05",
          5017 => x"8d",
          5018 => x"86",
          5019 => x"0b",
          5020 => x"80",
          5021 => x"8c",
          5022 => x"3d",
          5023 => x"3d",
          5024 => x"89",
          5025 => x"2e",
          5026 => x"08",
          5027 => x"2e",
          5028 => x"33",
          5029 => x"2e",
          5030 => x"13",
          5031 => x"22",
          5032 => x"76",
          5033 => x"06",
          5034 => x"13",
          5035 => x"c0",
          5036 => x"ec",
          5037 => x"52",
          5038 => x"71",
          5039 => x"55",
          5040 => x"53",
          5041 => x"0c",
          5042 => x"8c",
          5043 => x"3d",
          5044 => x"3d",
          5045 => x"05",
          5046 => x"89",
          5047 => x"52",
          5048 => x"3f",
          5049 => x"0b",
          5050 => x"08",
          5051 => x"82",
          5052 => x"84",
          5053 => x"88",
          5054 => x"55",
          5055 => x"2e",
          5056 => x"74",
          5057 => x"73",
          5058 => x"38",
          5059 => x"78",
          5060 => x"54",
          5061 => x"92",
          5062 => x"89",
          5063 => x"84",
          5064 => x"b0",
          5065 => x"ec",
          5066 => x"82",
          5067 => x"88",
          5068 => x"eb",
          5069 => x"02",
          5070 => x"e7",
          5071 => x"59",
          5072 => x"80",
          5073 => x"38",
          5074 => x"70",
          5075 => x"d0",
          5076 => x"3d",
          5077 => x"58",
          5078 => x"82",
          5079 => x"55",
          5080 => x"08",
          5081 => x"7a",
          5082 => x"8c",
          5083 => x"56",
          5084 => x"82",
          5085 => x"55",
          5086 => x"08",
          5087 => x"80",
          5088 => x"70",
          5089 => x"57",
          5090 => x"83",
          5091 => x"77",
          5092 => x"73",
          5093 => x"ab",
          5094 => x"2e",
          5095 => x"84",
          5096 => x"06",
          5097 => x"51",
          5098 => x"82",
          5099 => x"55",
          5100 => x"b2",
          5101 => x"06",
          5102 => x"b8",
          5103 => x"2a",
          5104 => x"51",
          5105 => x"2e",
          5106 => x"55",
          5107 => x"77",
          5108 => x"74",
          5109 => x"77",
          5110 => x"81",
          5111 => x"73",
          5112 => x"af",
          5113 => x"7a",
          5114 => x"3f",
          5115 => x"08",
          5116 => x"b2",
          5117 => x"8e",
          5118 => x"ea",
          5119 => x"a0",
          5120 => x"34",
          5121 => x"52",
          5122 => x"bd",
          5123 => x"62",
          5124 => x"d4",
          5125 => x"54",
          5126 => x"15",
          5127 => x"2e",
          5128 => x"7a",
          5129 => x"51",
          5130 => x"75",
          5131 => x"d4",
          5132 => x"be",
          5133 => x"ec",
          5134 => x"8c",
          5135 => x"ca",
          5136 => x"74",
          5137 => x"02",
          5138 => x"70",
          5139 => x"81",
          5140 => x"56",
          5141 => x"86",
          5142 => x"82",
          5143 => x"81",
          5144 => x"06",
          5145 => x"80",
          5146 => x"75",
          5147 => x"73",
          5148 => x"38",
          5149 => x"92",
          5150 => x"7a",
          5151 => x"3f",
          5152 => x"08",
          5153 => x"8c",
          5154 => x"55",
          5155 => x"08",
          5156 => x"77",
          5157 => x"81",
          5158 => x"73",
          5159 => x"38",
          5160 => x"07",
          5161 => x"11",
          5162 => x"0c",
          5163 => x"0c",
          5164 => x"52",
          5165 => x"3f",
          5166 => x"08",
          5167 => x"08",
          5168 => x"63",
          5169 => x"5a",
          5170 => x"82",
          5171 => x"82",
          5172 => x"8c",
          5173 => x"7a",
          5174 => x"17",
          5175 => x"23",
          5176 => x"34",
          5177 => x"1a",
          5178 => x"9c",
          5179 => x"0b",
          5180 => x"77",
          5181 => x"81",
          5182 => x"73",
          5183 => x"8d",
          5184 => x"ec",
          5185 => x"81",
          5186 => x"8c",
          5187 => x"1a",
          5188 => x"22",
          5189 => x"7b",
          5190 => x"a8",
          5191 => x"78",
          5192 => x"3f",
          5193 => x"08",
          5194 => x"ec",
          5195 => x"83",
          5196 => x"82",
          5197 => x"ff",
          5198 => x"06",
          5199 => x"55",
          5200 => x"56",
          5201 => x"76",
          5202 => x"51",
          5203 => x"27",
          5204 => x"70",
          5205 => x"5a",
          5206 => x"76",
          5207 => x"74",
          5208 => x"83",
          5209 => x"73",
          5210 => x"38",
          5211 => x"51",
          5212 => x"82",
          5213 => x"85",
          5214 => x"8e",
          5215 => x"2a",
          5216 => x"08",
          5217 => x"0c",
          5218 => x"79",
          5219 => x"73",
          5220 => x"0c",
          5221 => x"04",
          5222 => x"60",
          5223 => x"40",
          5224 => x"80",
          5225 => x"3d",
          5226 => x"78",
          5227 => x"3f",
          5228 => x"08",
          5229 => x"ec",
          5230 => x"91",
          5231 => x"74",
          5232 => x"38",
          5233 => x"c4",
          5234 => x"33",
          5235 => x"87",
          5236 => x"2e",
          5237 => x"95",
          5238 => x"91",
          5239 => x"56",
          5240 => x"81",
          5241 => x"34",
          5242 => x"a0",
          5243 => x"08",
          5244 => x"31",
          5245 => x"27",
          5246 => x"5c",
          5247 => x"82",
          5248 => x"19",
          5249 => x"ff",
          5250 => x"74",
          5251 => x"7e",
          5252 => x"ff",
          5253 => x"2a",
          5254 => x"79",
          5255 => x"87",
          5256 => x"08",
          5257 => x"98",
          5258 => x"78",
          5259 => x"3f",
          5260 => x"08",
          5261 => x"27",
          5262 => x"74",
          5263 => x"a3",
          5264 => x"1a",
          5265 => x"08",
          5266 => x"d4",
          5267 => x"8c",
          5268 => x"2e",
          5269 => x"82",
          5270 => x"1a",
          5271 => x"59",
          5272 => x"2e",
          5273 => x"77",
          5274 => x"11",
          5275 => x"55",
          5276 => x"85",
          5277 => x"31",
          5278 => x"76",
          5279 => x"81",
          5280 => x"ca",
          5281 => x"8c",
          5282 => x"d7",
          5283 => x"11",
          5284 => x"74",
          5285 => x"38",
          5286 => x"77",
          5287 => x"78",
          5288 => x"84",
          5289 => x"16",
          5290 => x"08",
          5291 => x"2b",
          5292 => x"cf",
          5293 => x"89",
          5294 => x"39",
          5295 => x"0c",
          5296 => x"83",
          5297 => x"80",
          5298 => x"55",
          5299 => x"83",
          5300 => x"9c",
          5301 => x"7e",
          5302 => x"3f",
          5303 => x"08",
          5304 => x"75",
          5305 => x"08",
          5306 => x"1f",
          5307 => x"7c",
          5308 => x"3f",
          5309 => x"7e",
          5310 => x"0c",
          5311 => x"1b",
          5312 => x"1c",
          5313 => x"fd",
          5314 => x"56",
          5315 => x"ec",
          5316 => x"0d",
          5317 => x"0d",
          5318 => x"64",
          5319 => x"58",
          5320 => x"90",
          5321 => x"52",
          5322 => x"d2",
          5323 => x"ec",
          5324 => x"8c",
          5325 => x"38",
          5326 => x"55",
          5327 => x"86",
          5328 => x"83",
          5329 => x"18",
          5330 => x"2a",
          5331 => x"51",
          5332 => x"56",
          5333 => x"83",
          5334 => x"39",
          5335 => x"19",
          5336 => x"83",
          5337 => x"0b",
          5338 => x"81",
          5339 => x"39",
          5340 => x"7c",
          5341 => x"74",
          5342 => x"38",
          5343 => x"7b",
          5344 => x"ec",
          5345 => x"08",
          5346 => x"06",
          5347 => x"81",
          5348 => x"8a",
          5349 => x"05",
          5350 => x"06",
          5351 => x"bf",
          5352 => x"38",
          5353 => x"55",
          5354 => x"7a",
          5355 => x"98",
          5356 => x"77",
          5357 => x"3f",
          5358 => x"08",
          5359 => x"ec",
          5360 => x"82",
          5361 => x"81",
          5362 => x"38",
          5363 => x"ff",
          5364 => x"98",
          5365 => x"18",
          5366 => x"74",
          5367 => x"7e",
          5368 => x"08",
          5369 => x"2e",
          5370 => x"8d",
          5371 => x"ce",
          5372 => x"8c",
          5373 => x"ee",
          5374 => x"08",
          5375 => x"d1",
          5376 => x"8c",
          5377 => x"2e",
          5378 => x"82",
          5379 => x"1b",
          5380 => x"5a",
          5381 => x"2e",
          5382 => x"78",
          5383 => x"11",
          5384 => x"55",
          5385 => x"85",
          5386 => x"31",
          5387 => x"76",
          5388 => x"81",
          5389 => x"c8",
          5390 => x"8c",
          5391 => x"a6",
          5392 => x"11",
          5393 => x"56",
          5394 => x"27",
          5395 => x"80",
          5396 => x"08",
          5397 => x"2b",
          5398 => x"b4",
          5399 => x"b5",
          5400 => x"80",
          5401 => x"34",
          5402 => x"56",
          5403 => x"8c",
          5404 => x"19",
          5405 => x"38",
          5406 => x"b6",
          5407 => x"ec",
          5408 => x"38",
          5409 => x"12",
          5410 => x"9c",
          5411 => x"18",
          5412 => x"06",
          5413 => x"31",
          5414 => x"76",
          5415 => x"7b",
          5416 => x"08",
          5417 => x"cd",
          5418 => x"8c",
          5419 => x"b6",
          5420 => x"7c",
          5421 => x"08",
          5422 => x"1f",
          5423 => x"cb",
          5424 => x"55",
          5425 => x"16",
          5426 => x"31",
          5427 => x"7f",
          5428 => x"94",
          5429 => x"70",
          5430 => x"8c",
          5431 => x"58",
          5432 => x"76",
          5433 => x"75",
          5434 => x"19",
          5435 => x"39",
          5436 => x"80",
          5437 => x"74",
          5438 => x"80",
          5439 => x"8c",
          5440 => x"3d",
          5441 => x"3d",
          5442 => x"3d",
          5443 => x"70",
          5444 => x"ea",
          5445 => x"ec",
          5446 => x"8c",
          5447 => x"fb",
          5448 => x"33",
          5449 => x"70",
          5450 => x"55",
          5451 => x"2e",
          5452 => x"a0",
          5453 => x"78",
          5454 => x"3f",
          5455 => x"08",
          5456 => x"ec",
          5457 => x"38",
          5458 => x"8b",
          5459 => x"07",
          5460 => x"8b",
          5461 => x"16",
          5462 => x"52",
          5463 => x"dd",
          5464 => x"16",
          5465 => x"15",
          5466 => x"3f",
          5467 => x"0a",
          5468 => x"51",
          5469 => x"76",
          5470 => x"51",
          5471 => x"78",
          5472 => x"83",
          5473 => x"51",
          5474 => x"82",
          5475 => x"90",
          5476 => x"bf",
          5477 => x"73",
          5478 => x"76",
          5479 => x"0c",
          5480 => x"04",
          5481 => x"76",
          5482 => x"fe",
          5483 => x"8c",
          5484 => x"82",
          5485 => x"9c",
          5486 => x"fc",
          5487 => x"51",
          5488 => x"82",
          5489 => x"53",
          5490 => x"08",
          5491 => x"8c",
          5492 => x"0c",
          5493 => x"ec",
          5494 => x"0d",
          5495 => x"0d",
          5496 => x"e6",
          5497 => x"52",
          5498 => x"8c",
          5499 => x"8b",
          5500 => x"ec",
          5501 => x"9c",
          5502 => x"71",
          5503 => x"0c",
          5504 => x"04",
          5505 => x"80",
          5506 => x"d0",
          5507 => x"3d",
          5508 => x"3f",
          5509 => x"08",
          5510 => x"ec",
          5511 => x"38",
          5512 => x"52",
          5513 => x"05",
          5514 => x"3f",
          5515 => x"08",
          5516 => x"ec",
          5517 => x"02",
          5518 => x"33",
          5519 => x"55",
          5520 => x"25",
          5521 => x"7a",
          5522 => x"54",
          5523 => x"a2",
          5524 => x"84",
          5525 => x"06",
          5526 => x"73",
          5527 => x"38",
          5528 => x"70",
          5529 => x"a8",
          5530 => x"ec",
          5531 => x"0c",
          5532 => x"8c",
          5533 => x"2e",
          5534 => x"83",
          5535 => x"74",
          5536 => x"0c",
          5537 => x"04",
          5538 => x"6f",
          5539 => x"80",
          5540 => x"53",
          5541 => x"b8",
          5542 => x"3d",
          5543 => x"3f",
          5544 => x"08",
          5545 => x"ec",
          5546 => x"38",
          5547 => x"7c",
          5548 => x"47",
          5549 => x"54",
          5550 => x"81",
          5551 => x"52",
          5552 => x"52",
          5553 => x"3f",
          5554 => x"08",
          5555 => x"ec",
          5556 => x"38",
          5557 => x"51",
          5558 => x"82",
          5559 => x"57",
          5560 => x"08",
          5561 => x"69",
          5562 => x"da",
          5563 => x"8c",
          5564 => x"76",
          5565 => x"d5",
          5566 => x"8c",
          5567 => x"82",
          5568 => x"82",
          5569 => x"52",
          5570 => x"eb",
          5571 => x"ec",
          5572 => x"8c",
          5573 => x"38",
          5574 => x"51",
          5575 => x"73",
          5576 => x"08",
          5577 => x"76",
          5578 => x"d6",
          5579 => x"8c",
          5580 => x"82",
          5581 => x"80",
          5582 => x"76",
          5583 => x"81",
          5584 => x"82",
          5585 => x"39",
          5586 => x"38",
          5587 => x"bc",
          5588 => x"51",
          5589 => x"76",
          5590 => x"11",
          5591 => x"51",
          5592 => x"73",
          5593 => x"38",
          5594 => x"55",
          5595 => x"16",
          5596 => x"56",
          5597 => x"38",
          5598 => x"73",
          5599 => x"90",
          5600 => x"2e",
          5601 => x"16",
          5602 => x"ff",
          5603 => x"ff",
          5604 => x"58",
          5605 => x"74",
          5606 => x"75",
          5607 => x"18",
          5608 => x"58",
          5609 => x"fe",
          5610 => x"7b",
          5611 => x"06",
          5612 => x"18",
          5613 => x"58",
          5614 => x"80",
          5615 => x"9c",
          5616 => x"29",
          5617 => x"05",
          5618 => x"33",
          5619 => x"56",
          5620 => x"2e",
          5621 => x"16",
          5622 => x"33",
          5623 => x"73",
          5624 => x"16",
          5625 => x"26",
          5626 => x"55",
          5627 => x"91",
          5628 => x"54",
          5629 => x"70",
          5630 => x"34",
          5631 => x"ec",
          5632 => x"70",
          5633 => x"34",
          5634 => x"09",
          5635 => x"38",
          5636 => x"39",
          5637 => x"19",
          5638 => x"33",
          5639 => x"05",
          5640 => x"78",
          5641 => x"80",
          5642 => x"82",
          5643 => x"9e",
          5644 => x"f7",
          5645 => x"7d",
          5646 => x"05",
          5647 => x"57",
          5648 => x"3f",
          5649 => x"08",
          5650 => x"ec",
          5651 => x"38",
          5652 => x"53",
          5653 => x"38",
          5654 => x"54",
          5655 => x"92",
          5656 => x"33",
          5657 => x"70",
          5658 => x"54",
          5659 => x"38",
          5660 => x"15",
          5661 => x"70",
          5662 => x"58",
          5663 => x"82",
          5664 => x"8a",
          5665 => x"89",
          5666 => x"53",
          5667 => x"b7",
          5668 => x"ff",
          5669 => x"99",
          5670 => x"8c",
          5671 => x"15",
          5672 => x"53",
          5673 => x"99",
          5674 => x"8c",
          5675 => x"26",
          5676 => x"30",
          5677 => x"70",
          5678 => x"77",
          5679 => x"18",
          5680 => x"51",
          5681 => x"88",
          5682 => x"73",
          5683 => x"52",
          5684 => x"ca",
          5685 => x"ec",
          5686 => x"8c",
          5687 => x"2e",
          5688 => x"82",
          5689 => x"ff",
          5690 => x"38",
          5691 => x"08",
          5692 => x"73",
          5693 => x"73",
          5694 => x"9c",
          5695 => x"27",
          5696 => x"75",
          5697 => x"16",
          5698 => x"17",
          5699 => x"33",
          5700 => x"70",
          5701 => x"55",
          5702 => x"80",
          5703 => x"73",
          5704 => x"cc",
          5705 => x"8c",
          5706 => x"82",
          5707 => x"94",
          5708 => x"ec",
          5709 => x"39",
          5710 => x"51",
          5711 => x"82",
          5712 => x"54",
          5713 => x"be",
          5714 => x"27",
          5715 => x"53",
          5716 => x"08",
          5717 => x"73",
          5718 => x"ff",
          5719 => x"15",
          5720 => x"16",
          5721 => x"ff",
          5722 => x"80",
          5723 => x"73",
          5724 => x"c6",
          5725 => x"8c",
          5726 => x"38",
          5727 => x"16",
          5728 => x"80",
          5729 => x"0b",
          5730 => x"81",
          5731 => x"75",
          5732 => x"8c",
          5733 => x"58",
          5734 => x"54",
          5735 => x"74",
          5736 => x"73",
          5737 => x"90",
          5738 => x"c0",
          5739 => x"90",
          5740 => x"83",
          5741 => x"72",
          5742 => x"38",
          5743 => x"08",
          5744 => x"77",
          5745 => x"80",
          5746 => x"8c",
          5747 => x"3d",
          5748 => x"3d",
          5749 => x"89",
          5750 => x"2e",
          5751 => x"80",
          5752 => x"fc",
          5753 => x"3d",
          5754 => x"e1",
          5755 => x"8c",
          5756 => x"82",
          5757 => x"80",
          5758 => x"76",
          5759 => x"75",
          5760 => x"3f",
          5761 => x"08",
          5762 => x"ec",
          5763 => x"38",
          5764 => x"70",
          5765 => x"57",
          5766 => x"a2",
          5767 => x"33",
          5768 => x"70",
          5769 => x"55",
          5770 => x"2e",
          5771 => x"16",
          5772 => x"51",
          5773 => x"82",
          5774 => x"88",
          5775 => x"54",
          5776 => x"84",
          5777 => x"52",
          5778 => x"e5",
          5779 => x"ec",
          5780 => x"84",
          5781 => x"06",
          5782 => x"55",
          5783 => x"80",
          5784 => x"80",
          5785 => x"54",
          5786 => x"ec",
          5787 => x"0d",
          5788 => x"0d",
          5789 => x"fc",
          5790 => x"52",
          5791 => x"3f",
          5792 => x"08",
          5793 => x"8c",
          5794 => x"0c",
          5795 => x"04",
          5796 => x"77",
          5797 => x"fc",
          5798 => x"53",
          5799 => x"de",
          5800 => x"ec",
          5801 => x"8c",
          5802 => x"df",
          5803 => x"38",
          5804 => x"08",
          5805 => x"cd",
          5806 => x"8c",
          5807 => x"80",
          5808 => x"8c",
          5809 => x"73",
          5810 => x"3f",
          5811 => x"08",
          5812 => x"ec",
          5813 => x"09",
          5814 => x"38",
          5815 => x"39",
          5816 => x"08",
          5817 => x"52",
          5818 => x"b3",
          5819 => x"73",
          5820 => x"3f",
          5821 => x"08",
          5822 => x"30",
          5823 => x"9f",
          5824 => x"8c",
          5825 => x"51",
          5826 => x"72",
          5827 => x"0c",
          5828 => x"04",
          5829 => x"65",
          5830 => x"89",
          5831 => x"96",
          5832 => x"df",
          5833 => x"8c",
          5834 => x"82",
          5835 => x"b2",
          5836 => x"75",
          5837 => x"3f",
          5838 => x"08",
          5839 => x"ec",
          5840 => x"02",
          5841 => x"33",
          5842 => x"55",
          5843 => x"25",
          5844 => x"55",
          5845 => x"80",
          5846 => x"76",
          5847 => x"d4",
          5848 => x"82",
          5849 => x"94",
          5850 => x"f0",
          5851 => x"65",
          5852 => x"53",
          5853 => x"05",
          5854 => x"51",
          5855 => x"82",
          5856 => x"5b",
          5857 => x"08",
          5858 => x"7c",
          5859 => x"08",
          5860 => x"fe",
          5861 => x"08",
          5862 => x"55",
          5863 => x"91",
          5864 => x"0c",
          5865 => x"81",
          5866 => x"39",
          5867 => x"c7",
          5868 => x"ec",
          5869 => x"55",
          5870 => x"2e",
          5871 => x"bf",
          5872 => x"5f",
          5873 => x"92",
          5874 => x"51",
          5875 => x"82",
          5876 => x"ff",
          5877 => x"82",
          5878 => x"81",
          5879 => x"82",
          5880 => x"30",
          5881 => x"ec",
          5882 => x"25",
          5883 => x"19",
          5884 => x"5a",
          5885 => x"08",
          5886 => x"38",
          5887 => x"a4",
          5888 => x"8c",
          5889 => x"58",
          5890 => x"77",
          5891 => x"7d",
          5892 => x"bf",
          5893 => x"8c",
          5894 => x"82",
          5895 => x"80",
          5896 => x"70",
          5897 => x"ff",
          5898 => x"56",
          5899 => x"2e",
          5900 => x"9e",
          5901 => x"51",
          5902 => x"3f",
          5903 => x"08",
          5904 => x"06",
          5905 => x"80",
          5906 => x"19",
          5907 => x"54",
          5908 => x"14",
          5909 => x"c5",
          5910 => x"ec",
          5911 => x"06",
          5912 => x"80",
          5913 => x"19",
          5914 => x"54",
          5915 => x"06",
          5916 => x"79",
          5917 => x"78",
          5918 => x"79",
          5919 => x"84",
          5920 => x"07",
          5921 => x"84",
          5922 => x"82",
          5923 => x"92",
          5924 => x"f9",
          5925 => x"8a",
          5926 => x"53",
          5927 => x"e3",
          5928 => x"8c",
          5929 => x"82",
          5930 => x"81",
          5931 => x"17",
          5932 => x"81",
          5933 => x"17",
          5934 => x"2a",
          5935 => x"51",
          5936 => x"55",
          5937 => x"81",
          5938 => x"17",
          5939 => x"8c",
          5940 => x"81",
          5941 => x"9b",
          5942 => x"ec",
          5943 => x"17",
          5944 => x"51",
          5945 => x"82",
          5946 => x"74",
          5947 => x"56",
          5948 => x"98",
          5949 => x"76",
          5950 => x"c6",
          5951 => x"ec",
          5952 => x"09",
          5953 => x"38",
          5954 => x"8c",
          5955 => x"2e",
          5956 => x"85",
          5957 => x"a3",
          5958 => x"38",
          5959 => x"8c",
          5960 => x"15",
          5961 => x"38",
          5962 => x"53",
          5963 => x"08",
          5964 => x"c3",
          5965 => x"8c",
          5966 => x"94",
          5967 => x"18",
          5968 => x"33",
          5969 => x"54",
          5970 => x"34",
          5971 => x"85",
          5972 => x"18",
          5973 => x"74",
          5974 => x"0c",
          5975 => x"04",
          5976 => x"82",
          5977 => x"ff",
          5978 => x"a1",
          5979 => x"e4",
          5980 => x"ec",
          5981 => x"8c",
          5982 => x"f5",
          5983 => x"a1",
          5984 => x"95",
          5985 => x"58",
          5986 => x"82",
          5987 => x"55",
          5988 => x"08",
          5989 => x"02",
          5990 => x"33",
          5991 => x"70",
          5992 => x"55",
          5993 => x"73",
          5994 => x"75",
          5995 => x"80",
          5996 => x"bd",
          5997 => x"d6",
          5998 => x"81",
          5999 => x"87",
          6000 => x"ad",
          6001 => x"78",
          6002 => x"3f",
          6003 => x"08",
          6004 => x"70",
          6005 => x"55",
          6006 => x"2e",
          6007 => x"78",
          6008 => x"ec",
          6009 => x"08",
          6010 => x"38",
          6011 => x"8c",
          6012 => x"76",
          6013 => x"70",
          6014 => x"b5",
          6015 => x"ec",
          6016 => x"8c",
          6017 => x"e9",
          6018 => x"ec",
          6019 => x"51",
          6020 => x"82",
          6021 => x"55",
          6022 => x"08",
          6023 => x"55",
          6024 => x"82",
          6025 => x"84",
          6026 => x"82",
          6027 => x"80",
          6028 => x"51",
          6029 => x"82",
          6030 => x"82",
          6031 => x"30",
          6032 => x"ec",
          6033 => x"25",
          6034 => x"75",
          6035 => x"38",
          6036 => x"8f",
          6037 => x"75",
          6038 => x"c1",
          6039 => x"8c",
          6040 => x"74",
          6041 => x"51",
          6042 => x"3f",
          6043 => x"08",
          6044 => x"8c",
          6045 => x"3d",
          6046 => x"3d",
          6047 => x"99",
          6048 => x"52",
          6049 => x"d8",
          6050 => x"8c",
          6051 => x"82",
          6052 => x"82",
          6053 => x"5e",
          6054 => x"3d",
          6055 => x"cf",
          6056 => x"8c",
          6057 => x"82",
          6058 => x"86",
          6059 => x"82",
          6060 => x"8c",
          6061 => x"2e",
          6062 => x"82",
          6063 => x"80",
          6064 => x"70",
          6065 => x"06",
          6066 => x"54",
          6067 => x"38",
          6068 => x"52",
          6069 => x"52",
          6070 => x"3f",
          6071 => x"08",
          6072 => x"82",
          6073 => x"83",
          6074 => x"82",
          6075 => x"81",
          6076 => x"06",
          6077 => x"54",
          6078 => x"08",
          6079 => x"81",
          6080 => x"81",
          6081 => x"39",
          6082 => x"38",
          6083 => x"08",
          6084 => x"c4",
          6085 => x"8c",
          6086 => x"82",
          6087 => x"81",
          6088 => x"53",
          6089 => x"19",
          6090 => x"8c",
          6091 => x"ae",
          6092 => x"34",
          6093 => x"0b",
          6094 => x"82",
          6095 => x"52",
          6096 => x"51",
          6097 => x"3f",
          6098 => x"b4",
          6099 => x"c9",
          6100 => x"53",
          6101 => x"53",
          6102 => x"51",
          6103 => x"3f",
          6104 => x"0b",
          6105 => x"34",
          6106 => x"80",
          6107 => x"51",
          6108 => x"78",
          6109 => x"83",
          6110 => x"51",
          6111 => x"82",
          6112 => x"54",
          6113 => x"08",
          6114 => x"88",
          6115 => x"64",
          6116 => x"ff",
          6117 => x"75",
          6118 => x"78",
          6119 => x"3f",
          6120 => x"0b",
          6121 => x"78",
          6122 => x"83",
          6123 => x"51",
          6124 => x"3f",
          6125 => x"08",
          6126 => x"80",
          6127 => x"76",
          6128 => x"ae",
          6129 => x"8c",
          6130 => x"3d",
          6131 => x"3d",
          6132 => x"84",
          6133 => x"f1",
          6134 => x"a8",
          6135 => x"05",
          6136 => x"51",
          6137 => x"82",
          6138 => x"55",
          6139 => x"08",
          6140 => x"78",
          6141 => x"08",
          6142 => x"70",
          6143 => x"b8",
          6144 => x"ec",
          6145 => x"8c",
          6146 => x"b9",
          6147 => x"9b",
          6148 => x"a0",
          6149 => x"55",
          6150 => x"38",
          6151 => x"3d",
          6152 => x"3d",
          6153 => x"51",
          6154 => x"3f",
          6155 => x"52",
          6156 => x"52",
          6157 => x"dd",
          6158 => x"08",
          6159 => x"cb",
          6160 => x"8c",
          6161 => x"82",
          6162 => x"95",
          6163 => x"2e",
          6164 => x"88",
          6165 => x"3d",
          6166 => x"38",
          6167 => x"e5",
          6168 => x"ec",
          6169 => x"09",
          6170 => x"b8",
          6171 => x"c9",
          6172 => x"8c",
          6173 => x"82",
          6174 => x"81",
          6175 => x"56",
          6176 => x"3d",
          6177 => x"52",
          6178 => x"ff",
          6179 => x"02",
          6180 => x"8b",
          6181 => x"16",
          6182 => x"2a",
          6183 => x"51",
          6184 => x"89",
          6185 => x"07",
          6186 => x"17",
          6187 => x"81",
          6188 => x"34",
          6189 => x"70",
          6190 => x"81",
          6191 => x"55",
          6192 => x"80",
          6193 => x"64",
          6194 => x"38",
          6195 => x"51",
          6196 => x"82",
          6197 => x"52",
          6198 => x"b7",
          6199 => x"55",
          6200 => x"08",
          6201 => x"dd",
          6202 => x"ec",
          6203 => x"51",
          6204 => x"3f",
          6205 => x"08",
          6206 => x"11",
          6207 => x"82",
          6208 => x"80",
          6209 => x"16",
          6210 => x"ae",
          6211 => x"06",
          6212 => x"53",
          6213 => x"51",
          6214 => x"78",
          6215 => x"83",
          6216 => x"39",
          6217 => x"08",
          6218 => x"51",
          6219 => x"82",
          6220 => x"55",
          6221 => x"08",
          6222 => x"51",
          6223 => x"3f",
          6224 => x"08",
          6225 => x"8c",
          6226 => x"3d",
          6227 => x"3d",
          6228 => x"db",
          6229 => x"84",
          6230 => x"05",
          6231 => x"82",
          6232 => x"d0",
          6233 => x"3d",
          6234 => x"3f",
          6235 => x"08",
          6236 => x"ec",
          6237 => x"38",
          6238 => x"52",
          6239 => x"05",
          6240 => x"3f",
          6241 => x"08",
          6242 => x"ec",
          6243 => x"02",
          6244 => x"33",
          6245 => x"54",
          6246 => x"aa",
          6247 => x"06",
          6248 => x"8b",
          6249 => x"06",
          6250 => x"07",
          6251 => x"56",
          6252 => x"34",
          6253 => x"0b",
          6254 => x"78",
          6255 => x"a9",
          6256 => x"ec",
          6257 => x"82",
          6258 => x"95",
          6259 => x"ef",
          6260 => x"56",
          6261 => x"3d",
          6262 => x"94",
          6263 => x"f4",
          6264 => x"ec",
          6265 => x"8c",
          6266 => x"cb",
          6267 => x"63",
          6268 => x"d4",
          6269 => x"c0",
          6270 => x"ec",
          6271 => x"8c",
          6272 => x"38",
          6273 => x"05",
          6274 => x"06",
          6275 => x"73",
          6276 => x"16",
          6277 => x"22",
          6278 => x"07",
          6279 => x"1f",
          6280 => x"c2",
          6281 => x"81",
          6282 => x"34",
          6283 => x"b3",
          6284 => x"8c",
          6285 => x"74",
          6286 => x"0c",
          6287 => x"04",
          6288 => x"69",
          6289 => x"80",
          6290 => x"d0",
          6291 => x"3d",
          6292 => x"3f",
          6293 => x"08",
          6294 => x"08",
          6295 => x"8c",
          6296 => x"80",
          6297 => x"57",
          6298 => x"81",
          6299 => x"70",
          6300 => x"55",
          6301 => x"80",
          6302 => x"5d",
          6303 => x"52",
          6304 => x"52",
          6305 => x"a9",
          6306 => x"ec",
          6307 => x"8c",
          6308 => x"d1",
          6309 => x"73",
          6310 => x"3f",
          6311 => x"08",
          6312 => x"ec",
          6313 => x"82",
          6314 => x"82",
          6315 => x"65",
          6316 => x"78",
          6317 => x"7b",
          6318 => x"55",
          6319 => x"34",
          6320 => x"8a",
          6321 => x"38",
          6322 => x"1a",
          6323 => x"34",
          6324 => x"9e",
          6325 => x"70",
          6326 => x"51",
          6327 => x"a0",
          6328 => x"8e",
          6329 => x"2e",
          6330 => x"86",
          6331 => x"34",
          6332 => x"30",
          6333 => x"80",
          6334 => x"7a",
          6335 => x"c1",
          6336 => x"2e",
          6337 => x"a0",
          6338 => x"51",
          6339 => x"3f",
          6340 => x"08",
          6341 => x"ec",
          6342 => x"7b",
          6343 => x"55",
          6344 => x"73",
          6345 => x"38",
          6346 => x"73",
          6347 => x"38",
          6348 => x"15",
          6349 => x"ff",
          6350 => x"82",
          6351 => x"7b",
          6352 => x"8c",
          6353 => x"3d",
          6354 => x"3d",
          6355 => x"9c",
          6356 => x"05",
          6357 => x"51",
          6358 => x"82",
          6359 => x"82",
          6360 => x"56",
          6361 => x"ec",
          6362 => x"38",
          6363 => x"52",
          6364 => x"52",
          6365 => x"c0",
          6366 => x"70",
          6367 => x"ff",
          6368 => x"55",
          6369 => x"27",
          6370 => x"78",
          6371 => x"ff",
          6372 => x"05",
          6373 => x"55",
          6374 => x"3f",
          6375 => x"08",
          6376 => x"38",
          6377 => x"70",
          6378 => x"ff",
          6379 => x"82",
          6380 => x"80",
          6381 => x"74",
          6382 => x"07",
          6383 => x"4e",
          6384 => x"82",
          6385 => x"55",
          6386 => x"70",
          6387 => x"06",
          6388 => x"99",
          6389 => x"e0",
          6390 => x"ff",
          6391 => x"54",
          6392 => x"27",
          6393 => x"fb",
          6394 => x"55",
          6395 => x"a3",
          6396 => x"81",
          6397 => x"ff",
          6398 => x"82",
          6399 => x"93",
          6400 => x"75",
          6401 => x"76",
          6402 => x"38",
          6403 => x"77",
          6404 => x"86",
          6405 => x"39",
          6406 => x"27",
          6407 => x"88",
          6408 => x"78",
          6409 => x"5a",
          6410 => x"57",
          6411 => x"81",
          6412 => x"81",
          6413 => x"33",
          6414 => x"06",
          6415 => x"57",
          6416 => x"fe",
          6417 => x"3d",
          6418 => x"55",
          6419 => x"2e",
          6420 => x"76",
          6421 => x"38",
          6422 => x"55",
          6423 => x"33",
          6424 => x"a0",
          6425 => x"06",
          6426 => x"17",
          6427 => x"38",
          6428 => x"43",
          6429 => x"3d",
          6430 => x"ff",
          6431 => x"82",
          6432 => x"54",
          6433 => x"08",
          6434 => x"81",
          6435 => x"ff",
          6436 => x"82",
          6437 => x"54",
          6438 => x"08",
          6439 => x"80",
          6440 => x"54",
          6441 => x"80",
          6442 => x"8c",
          6443 => x"2e",
          6444 => x"80",
          6445 => x"54",
          6446 => x"80",
          6447 => x"52",
          6448 => x"bd",
          6449 => x"8c",
          6450 => x"82",
          6451 => x"b1",
          6452 => x"82",
          6453 => x"52",
          6454 => x"ab",
          6455 => x"54",
          6456 => x"15",
          6457 => x"78",
          6458 => x"ff",
          6459 => x"79",
          6460 => x"83",
          6461 => x"51",
          6462 => x"3f",
          6463 => x"08",
          6464 => x"74",
          6465 => x"0c",
          6466 => x"04",
          6467 => x"60",
          6468 => x"05",
          6469 => x"33",
          6470 => x"05",
          6471 => x"40",
          6472 => x"da",
          6473 => x"ec",
          6474 => x"8c",
          6475 => x"bd",
          6476 => x"33",
          6477 => x"b5",
          6478 => x"2e",
          6479 => x"1a",
          6480 => x"90",
          6481 => x"33",
          6482 => x"70",
          6483 => x"55",
          6484 => x"38",
          6485 => x"97",
          6486 => x"82",
          6487 => x"58",
          6488 => x"7e",
          6489 => x"70",
          6490 => x"55",
          6491 => x"56",
          6492 => x"c5",
          6493 => x"7d",
          6494 => x"70",
          6495 => x"2a",
          6496 => x"08",
          6497 => x"08",
          6498 => x"5d",
          6499 => x"77",
          6500 => x"98",
          6501 => x"26",
          6502 => x"57",
          6503 => x"59",
          6504 => x"52",
          6505 => x"ae",
          6506 => x"15",
          6507 => x"98",
          6508 => x"26",
          6509 => x"55",
          6510 => x"08",
          6511 => x"99",
          6512 => x"ec",
          6513 => x"ff",
          6514 => x"8c",
          6515 => x"38",
          6516 => x"75",
          6517 => x"81",
          6518 => x"93",
          6519 => x"80",
          6520 => x"2e",
          6521 => x"ff",
          6522 => x"58",
          6523 => x"7d",
          6524 => x"38",
          6525 => x"55",
          6526 => x"b4",
          6527 => x"56",
          6528 => x"09",
          6529 => x"38",
          6530 => x"53",
          6531 => x"51",
          6532 => x"3f",
          6533 => x"08",
          6534 => x"ec",
          6535 => x"38",
          6536 => x"ff",
          6537 => x"5c",
          6538 => x"84",
          6539 => x"5c",
          6540 => x"12",
          6541 => x"80",
          6542 => x"78",
          6543 => x"7c",
          6544 => x"90",
          6545 => x"c0",
          6546 => x"90",
          6547 => x"15",
          6548 => x"90",
          6549 => x"54",
          6550 => x"91",
          6551 => x"31",
          6552 => x"84",
          6553 => x"07",
          6554 => x"16",
          6555 => x"73",
          6556 => x"0c",
          6557 => x"04",
          6558 => x"6b",
          6559 => x"05",
          6560 => x"33",
          6561 => x"5a",
          6562 => x"bd",
          6563 => x"80",
          6564 => x"ec",
          6565 => x"f8",
          6566 => x"ec",
          6567 => x"82",
          6568 => x"70",
          6569 => x"74",
          6570 => x"38",
          6571 => x"82",
          6572 => x"81",
          6573 => x"81",
          6574 => x"ff",
          6575 => x"82",
          6576 => x"81",
          6577 => x"81",
          6578 => x"83",
          6579 => x"c0",
          6580 => x"2a",
          6581 => x"51",
          6582 => x"74",
          6583 => x"99",
          6584 => x"53",
          6585 => x"51",
          6586 => x"3f",
          6587 => x"08",
          6588 => x"55",
          6589 => x"92",
          6590 => x"80",
          6591 => x"38",
          6592 => x"06",
          6593 => x"2e",
          6594 => x"48",
          6595 => x"87",
          6596 => x"79",
          6597 => x"78",
          6598 => x"26",
          6599 => x"19",
          6600 => x"74",
          6601 => x"38",
          6602 => x"e4",
          6603 => x"2a",
          6604 => x"70",
          6605 => x"59",
          6606 => x"7a",
          6607 => x"56",
          6608 => x"80",
          6609 => x"51",
          6610 => x"74",
          6611 => x"99",
          6612 => x"53",
          6613 => x"51",
          6614 => x"3f",
          6615 => x"8c",
          6616 => x"ac",
          6617 => x"2a",
          6618 => x"82",
          6619 => x"43",
          6620 => x"83",
          6621 => x"66",
          6622 => x"60",
          6623 => x"90",
          6624 => x"31",
          6625 => x"80",
          6626 => x"8a",
          6627 => x"56",
          6628 => x"26",
          6629 => x"77",
          6630 => x"81",
          6631 => x"74",
          6632 => x"38",
          6633 => x"55",
          6634 => x"83",
          6635 => x"81",
          6636 => x"80",
          6637 => x"38",
          6638 => x"55",
          6639 => x"5e",
          6640 => x"89",
          6641 => x"5a",
          6642 => x"09",
          6643 => x"e1",
          6644 => x"38",
          6645 => x"57",
          6646 => x"fd",
          6647 => x"5a",
          6648 => x"9d",
          6649 => x"26",
          6650 => x"fd",
          6651 => x"10",
          6652 => x"22",
          6653 => x"74",
          6654 => x"38",
          6655 => x"ee",
          6656 => x"66",
          6657 => x"b1",
          6658 => x"ec",
          6659 => x"84",
          6660 => x"89",
          6661 => x"a0",
          6662 => x"82",
          6663 => x"fc",
          6664 => x"56",
          6665 => x"f0",
          6666 => x"80",
          6667 => x"d3",
          6668 => x"38",
          6669 => x"57",
          6670 => x"fd",
          6671 => x"5a",
          6672 => x"9d",
          6673 => x"26",
          6674 => x"fd",
          6675 => x"10",
          6676 => x"22",
          6677 => x"74",
          6678 => x"38",
          6679 => x"ee",
          6680 => x"66",
          6681 => x"d1",
          6682 => x"ec",
          6683 => x"05",
          6684 => x"ec",
          6685 => x"26",
          6686 => x"0b",
          6687 => x"08",
          6688 => x"ec",
          6689 => x"11",
          6690 => x"05",
          6691 => x"83",
          6692 => x"2a",
          6693 => x"a0",
          6694 => x"7d",
          6695 => x"69",
          6696 => x"05",
          6697 => x"72",
          6698 => x"5c",
          6699 => x"59",
          6700 => x"2e",
          6701 => x"89",
          6702 => x"60",
          6703 => x"84",
          6704 => x"5d",
          6705 => x"18",
          6706 => x"68",
          6707 => x"74",
          6708 => x"af",
          6709 => x"31",
          6710 => x"53",
          6711 => x"52",
          6712 => x"d5",
          6713 => x"ec",
          6714 => x"83",
          6715 => x"06",
          6716 => x"8c",
          6717 => x"ff",
          6718 => x"dd",
          6719 => x"83",
          6720 => x"2a",
          6721 => x"be",
          6722 => x"39",
          6723 => x"09",
          6724 => x"c5",
          6725 => x"f5",
          6726 => x"ec",
          6727 => x"38",
          6728 => x"79",
          6729 => x"80",
          6730 => x"38",
          6731 => x"96",
          6732 => x"06",
          6733 => x"2e",
          6734 => x"5e",
          6735 => x"82",
          6736 => x"9f",
          6737 => x"38",
          6738 => x"38",
          6739 => x"81",
          6740 => x"fc",
          6741 => x"ab",
          6742 => x"7d",
          6743 => x"81",
          6744 => x"7d",
          6745 => x"78",
          6746 => x"74",
          6747 => x"8e",
          6748 => x"9c",
          6749 => x"53",
          6750 => x"51",
          6751 => x"3f",
          6752 => x"fb",
          6753 => x"51",
          6754 => x"3f",
          6755 => x"8b",
          6756 => x"a1",
          6757 => x"8d",
          6758 => x"83",
          6759 => x"52",
          6760 => x"ff",
          6761 => x"81",
          6762 => x"34",
          6763 => x"70",
          6764 => x"2a",
          6765 => x"54",
          6766 => x"1b",
          6767 => x"88",
          6768 => x"74",
          6769 => x"26",
          6770 => x"83",
          6771 => x"52",
          6772 => x"ff",
          6773 => x"8a",
          6774 => x"a0",
          6775 => x"a1",
          6776 => x"0b",
          6777 => x"bf",
          6778 => x"51",
          6779 => x"3f",
          6780 => x"9a",
          6781 => x"a0",
          6782 => x"52",
          6783 => x"ff",
          6784 => x"7d",
          6785 => x"81",
          6786 => x"38",
          6787 => x"0a",
          6788 => x"1b",
          6789 => x"ce",
          6790 => x"a4",
          6791 => x"a0",
          6792 => x"52",
          6793 => x"ff",
          6794 => x"81",
          6795 => x"51",
          6796 => x"3f",
          6797 => x"1b",
          6798 => x"8c",
          6799 => x"0b",
          6800 => x"34",
          6801 => x"c2",
          6802 => x"53",
          6803 => x"52",
          6804 => x"51",
          6805 => x"88",
          6806 => x"a7",
          6807 => x"a0",
          6808 => x"83",
          6809 => x"52",
          6810 => x"ff",
          6811 => x"ff",
          6812 => x"1c",
          6813 => x"a6",
          6814 => x"53",
          6815 => x"52",
          6816 => x"ff",
          6817 => x"82",
          6818 => x"83",
          6819 => x"52",
          6820 => x"b4",
          6821 => x"60",
          6822 => x"7e",
          6823 => x"d7",
          6824 => x"82",
          6825 => x"83",
          6826 => x"83",
          6827 => x"06",
          6828 => x"75",
          6829 => x"05",
          6830 => x"7e",
          6831 => x"b7",
          6832 => x"53",
          6833 => x"51",
          6834 => x"3f",
          6835 => x"a4",
          6836 => x"51",
          6837 => x"3f",
          6838 => x"e4",
          6839 => x"e4",
          6840 => x"9f",
          6841 => x"18",
          6842 => x"1b",
          6843 => x"f6",
          6844 => x"83",
          6845 => x"ff",
          6846 => x"82",
          6847 => x"78",
          6848 => x"c4",
          6849 => x"60",
          6850 => x"7a",
          6851 => x"ff",
          6852 => x"75",
          6853 => x"53",
          6854 => x"51",
          6855 => x"3f",
          6856 => x"52",
          6857 => x"9f",
          6858 => x"56",
          6859 => x"83",
          6860 => x"06",
          6861 => x"52",
          6862 => x"9e",
          6863 => x"52",
          6864 => x"ff",
          6865 => x"f0",
          6866 => x"1b",
          6867 => x"87",
          6868 => x"55",
          6869 => x"83",
          6870 => x"74",
          6871 => x"ff",
          6872 => x"7c",
          6873 => x"74",
          6874 => x"38",
          6875 => x"54",
          6876 => x"52",
          6877 => x"99",
          6878 => x"8c",
          6879 => x"87",
          6880 => x"53",
          6881 => x"08",
          6882 => x"ff",
          6883 => x"76",
          6884 => x"31",
          6885 => x"cd",
          6886 => x"58",
          6887 => x"ff",
          6888 => x"55",
          6889 => x"83",
          6890 => x"61",
          6891 => x"26",
          6892 => x"57",
          6893 => x"53",
          6894 => x"51",
          6895 => x"3f",
          6896 => x"08",
          6897 => x"76",
          6898 => x"31",
          6899 => x"db",
          6900 => x"7d",
          6901 => x"38",
          6902 => x"83",
          6903 => x"8a",
          6904 => x"7d",
          6905 => x"38",
          6906 => x"81",
          6907 => x"80",
          6908 => x"80",
          6909 => x"7a",
          6910 => x"bc",
          6911 => x"d5",
          6912 => x"ff",
          6913 => x"83",
          6914 => x"77",
          6915 => x"0b",
          6916 => x"81",
          6917 => x"34",
          6918 => x"34",
          6919 => x"34",
          6920 => x"56",
          6921 => x"52",
          6922 => x"f2",
          6923 => x"0b",
          6924 => x"82",
          6925 => x"82",
          6926 => x"56",
          6927 => x"34",
          6928 => x"08",
          6929 => x"60",
          6930 => x"1b",
          6931 => x"96",
          6932 => x"83",
          6933 => x"ff",
          6934 => x"81",
          6935 => x"7a",
          6936 => x"ff",
          6937 => x"81",
          6938 => x"ec",
          6939 => x"80",
          6940 => x"7e",
          6941 => x"e3",
          6942 => x"82",
          6943 => x"90",
          6944 => x"8e",
          6945 => x"81",
          6946 => x"82",
          6947 => x"56",
          6948 => x"ec",
          6949 => x"0d",
          6950 => x"0d",
          6951 => x"59",
          6952 => x"ff",
          6953 => x"57",
          6954 => x"b4",
          6955 => x"f8",
          6956 => x"81",
          6957 => x"52",
          6958 => x"dc",
          6959 => x"2e",
          6960 => x"9c",
          6961 => x"33",
          6962 => x"2e",
          6963 => x"76",
          6964 => x"58",
          6965 => x"57",
          6966 => x"09",
          6967 => x"38",
          6968 => x"78",
          6969 => x"38",
          6970 => x"82",
          6971 => x"8d",
          6972 => x"fa",
          6973 => x"70",
          6974 => x"56",
          6975 => x"2e",
          6976 => x"8e",
          6977 => x"0c",
          6978 => x"53",
          6979 => x"81",
          6980 => x"75",
          6981 => x"73",
          6982 => x"38",
          6983 => x"30",
          6984 => x"77",
          6985 => x"72",
          6986 => x"a0",
          6987 => x"06",
          6988 => x"75",
          6989 => x"57",
          6990 => x"75",
          6991 => x"89",
          6992 => x"08",
          6993 => x"52",
          6994 => x"f6",
          6995 => x"ec",
          6996 => x"84",
          6997 => x"72",
          6998 => x"a9",
          6999 => x"70",
          7000 => x"57",
          7001 => x"27",
          7002 => x"53",
          7003 => x"ec",
          7004 => x"0d",
          7005 => x"0d",
          7006 => x"93",
          7007 => x"38",
          7008 => x"81",
          7009 => x"52",
          7010 => x"81",
          7011 => x"81",
          7012 => x"ff",
          7013 => x"f9",
          7014 => x"a8",
          7015 => x"39",
          7016 => x"51",
          7017 => x"81",
          7018 => x"80",
          7019 => x"ff",
          7020 => x"dd",
          7021 => x"f0",
          7022 => x"39",
          7023 => x"51",
          7024 => x"82",
          7025 => x"80",
          7026 => x"80",
          7027 => x"c1",
          7028 => x"c8",
          7029 => x"82",
          7030 => x"b5",
          7031 => x"f8",
          7032 => x"82",
          7033 => x"a9",
          7034 => x"b8",
          7035 => x"82",
          7036 => x"9d",
          7037 => x"ec",
          7038 => x"82",
          7039 => x"91",
          7040 => x"9c",
          7041 => x"82",
          7042 => x"85",
          7043 => x"c0",
          7044 => x"9f",
          7045 => x"0d",
          7046 => x"0d",
          7047 => x"56",
          7048 => x"26",
          7049 => x"52",
          7050 => x"29",
          7051 => x"87",
          7052 => x"51",
          7053 => x"3f",
          7054 => x"08",
          7055 => x"fe",
          7056 => x"82",
          7057 => x"54",
          7058 => x"52",
          7059 => x"51",
          7060 => x"3f",
          7061 => x"04",
          7062 => x"66",
          7063 => x"80",
          7064 => x"5b",
          7065 => x"78",
          7066 => x"07",
          7067 => x"57",
          7068 => x"56",
          7069 => x"26",
          7070 => x"56",
          7071 => x"70",
          7072 => x"51",
          7073 => x"74",
          7074 => x"81",
          7075 => x"8c",
          7076 => x"56",
          7077 => x"82",
          7078 => x"57",
          7079 => x"08",
          7080 => x"8c",
          7081 => x"c0",
          7082 => x"82",
          7083 => x"59",
          7084 => x"05",
          7085 => x"53",
          7086 => x"51",
          7087 => x"82",
          7088 => x"57",
          7089 => x"08",
          7090 => x"55",
          7091 => x"89",
          7092 => x"75",
          7093 => x"d8",
          7094 => x"d8",
          7095 => x"c4",
          7096 => x"70",
          7097 => x"25",
          7098 => x"9f",
          7099 => x"51",
          7100 => x"74",
          7101 => x"38",
          7102 => x"53",
          7103 => x"88",
          7104 => x"51",
          7105 => x"76",
          7106 => x"8c",
          7107 => x"3d",
          7108 => x"3d",
          7109 => x"84",
          7110 => x"33",
          7111 => x"57",
          7112 => x"52",
          7113 => x"b0",
          7114 => x"ec",
          7115 => x"75",
          7116 => x"38",
          7117 => x"98",
          7118 => x"60",
          7119 => x"82",
          7120 => x"7e",
          7121 => x"77",
          7122 => x"ec",
          7123 => x"39",
          7124 => x"82",
          7125 => x"89",
          7126 => x"f3",
          7127 => x"61",
          7128 => x"05",
          7129 => x"33",
          7130 => x"68",
          7131 => x"5c",
          7132 => x"7a",
          7133 => x"fc",
          7134 => x"9b",
          7135 => x"84",
          7136 => x"af",
          7137 => x"74",
          7138 => x"fc",
          7139 => x"2e",
          7140 => x"a0",
          7141 => x"80",
          7142 => x"18",
          7143 => x"27",
          7144 => x"22",
          7145 => x"88",
          7146 => x"eb",
          7147 => x"82",
          7148 => x"ff",
          7149 => x"82",
          7150 => x"c3",
          7151 => x"53",
          7152 => x"8e",
          7153 => x"52",
          7154 => x"51",
          7155 => x"3f",
          7156 => x"83",
          7157 => x"82",
          7158 => x"15",
          7159 => x"74",
          7160 => x"7a",
          7161 => x"72",
          7162 => x"83",
          7163 => x"88",
          7164 => x"39",
          7165 => x"51",
          7166 => x"3f",
          7167 => x"a0",
          7168 => x"d2",
          7169 => x"39",
          7170 => x"51",
          7171 => x"3f",
          7172 => x"79",
          7173 => x"74",
          7174 => x"55",
          7175 => x"72",
          7176 => x"38",
          7177 => x"53",
          7178 => x"83",
          7179 => x"75",
          7180 => x"81",
          7181 => x"53",
          7182 => x"8b",
          7183 => x"fe",
          7184 => x"73",
          7185 => x"a0",
          7186 => x"8a",
          7187 => x"55",
          7188 => x"83",
          7189 => x"81",
          7190 => x"18",
          7191 => x"58",
          7192 => x"3f",
          7193 => x"08",
          7194 => x"98",
          7195 => x"76",
          7196 => x"81",
          7197 => x"fe",
          7198 => x"82",
          7199 => x"98",
          7200 => x"2c",
          7201 => x"70",
          7202 => x"32",
          7203 => x"72",
          7204 => x"07",
          7205 => x"58",
          7206 => x"57",
          7207 => x"d7",
          7208 => x"2e",
          7209 => x"85",
          7210 => x"8c",
          7211 => x"53",
          7212 => x"fd",
          7213 => x"53",
          7214 => x"ec",
          7215 => x"0d",
          7216 => x"0d",
          7217 => x"33",
          7218 => x"53",
          7219 => x"52",
          7220 => x"c3",
          7221 => x"cc",
          7222 => x"ff",
          7223 => x"83",
          7224 => x"83",
          7225 => x"89",
          7226 => x"82",
          7227 => x"ff",
          7228 => x"74",
          7229 => x"38",
          7230 => x"3f",
          7231 => x"04",
          7232 => x"87",
          7233 => x"08",
          7234 => x"b8",
          7235 => x"fe",
          7236 => x"82",
          7237 => x"fe",
          7238 => x"80",
          7239 => x"b3",
          7240 => x"2a",
          7241 => x"51",
          7242 => x"2e",
          7243 => x"51",
          7244 => x"3f",
          7245 => x"51",
          7246 => x"3f",
          7247 => x"f1",
          7248 => x"82",
          7249 => x"06",
          7250 => x"80",
          7251 => x"81",
          7252 => x"ff",
          7253 => x"9c",
          7254 => x"f7",
          7255 => x"fe",
          7256 => x"72",
          7257 => x"81",
          7258 => x"71",
          7259 => x"38",
          7260 => x"f0",
          7261 => x"84",
          7262 => x"f2",
          7263 => x"51",
          7264 => x"3f",
          7265 => x"70",
          7266 => x"52",
          7267 => x"95",
          7268 => x"fe",
          7269 => x"82",
          7270 => x"fe",
          7271 => x"80",
          7272 => x"af",
          7273 => x"2a",
          7274 => x"51",
          7275 => x"2e",
          7276 => x"51",
          7277 => x"3f",
          7278 => x"51",
          7279 => x"3f",
          7280 => x"f0",
          7281 => x"86",
          7282 => x"06",
          7283 => x"80",
          7284 => x"81",
          7285 => x"fb",
          7286 => x"e8",
          7287 => x"f3",
          7288 => x"fe",
          7289 => x"72",
          7290 => x"81",
          7291 => x"71",
          7292 => x"38",
          7293 => x"ef",
          7294 => x"84",
          7295 => x"f1",
          7296 => x"51",
          7297 => x"3f",
          7298 => x"70",
          7299 => x"52",
          7300 => x"95",
          7301 => x"fe",
          7302 => x"82",
          7303 => x"fe",
          7304 => x"80",
          7305 => x"ab",
          7306 => x"a0",
          7307 => x"0d",
          7308 => x"0d",
          7309 => x"55",
          7310 => x"52",
          7311 => x"e8",
          7312 => x"89",
          7313 => x"73",
          7314 => x"53",
          7315 => x"52",
          7316 => x"51",
          7317 => x"3f",
          7318 => x"08",
          7319 => x"8c",
          7320 => x"80",
          7321 => x"31",
          7322 => x"73",
          7323 => x"34",
          7324 => x"33",
          7325 => x"2e",
          7326 => x"ac",
          7327 => x"f0",
          7328 => x"75",
          7329 => x"3f",
          7330 => x"08",
          7331 => x"38",
          7332 => x"08",
          7333 => x"9b",
          7334 => x"82",
          7335 => x"c6",
          7336 => x"0b",
          7337 => x"34",
          7338 => x"33",
          7339 => x"2e",
          7340 => x"89",
          7341 => x"75",
          7342 => x"b5",
          7343 => x"82",
          7344 => x"87",
          7345 => x"ce",
          7346 => x"70",
          7347 => x"ec",
          7348 => x"81",
          7349 => x"ff",
          7350 => x"82",
          7351 => x"81",
          7352 => x"78",
          7353 => x"81",
          7354 => x"82",
          7355 => x"96",
          7356 => x"59",
          7357 => x"3f",
          7358 => x"52",
          7359 => x"51",
          7360 => x"3f",
          7361 => x"08",
          7362 => x"38",
          7363 => x"51",
          7364 => x"81",
          7365 => x"82",
          7366 => x"fe",
          7367 => x"96",
          7368 => x"5a",
          7369 => x"79",
          7370 => x"3f",
          7371 => x"84",
          7372 => x"bf",
          7373 => x"ec",
          7374 => x"70",
          7375 => x"59",
          7376 => x"2e",
          7377 => x"78",
          7378 => x"b2",
          7379 => x"2e",
          7380 => x"78",
          7381 => x"38",
          7382 => x"ff",
          7383 => x"bc",
          7384 => x"38",
          7385 => x"78",
          7386 => x"83",
          7387 => x"80",
          7388 => x"dd",
          7389 => x"2e",
          7390 => x"8a",
          7391 => x"80",
          7392 => x"ea",
          7393 => x"f9",
          7394 => x"78",
          7395 => x"88",
          7396 => x"80",
          7397 => x"b1",
          7398 => x"39",
          7399 => x"2e",
          7400 => x"78",
          7401 => x"8b",
          7402 => x"82",
          7403 => x"38",
          7404 => x"78",
          7405 => x"8a",
          7406 => x"93",
          7407 => x"ff",
          7408 => x"ff",
          7409 => x"ff",
          7410 => x"82",
          7411 => x"80",
          7412 => x"38",
          7413 => x"fc",
          7414 => x"84",
          7415 => x"82",
          7416 => x"8c",
          7417 => x"2e",
          7418 => x"b4",
          7419 => x"11",
          7420 => x"05",
          7421 => x"94",
          7422 => x"ec",
          7423 => x"82",
          7424 => x"42",
          7425 => x"51",
          7426 => x"3f",
          7427 => x"5a",
          7428 => x"81",
          7429 => x"59",
          7430 => x"84",
          7431 => x"7a",
          7432 => x"38",
          7433 => x"b4",
          7434 => x"11",
          7435 => x"05",
          7436 => x"d8",
          7437 => x"ec",
          7438 => x"fd",
          7439 => x"3d",
          7440 => x"53",
          7441 => x"51",
          7442 => x"3f",
          7443 => x"08",
          7444 => x"c3",
          7445 => x"fe",
          7446 => x"ff",
          7447 => x"ff",
          7448 => x"82",
          7449 => x"80",
          7450 => x"38",
          7451 => x"51",
          7452 => x"3f",
          7453 => x"63",
          7454 => x"38",
          7455 => x"70",
          7456 => x"33",
          7457 => x"81",
          7458 => x"39",
          7459 => x"80",
          7460 => x"84",
          7461 => x"80",
          7462 => x"8c",
          7463 => x"2e",
          7464 => x"b4",
          7465 => x"11",
          7466 => x"05",
          7467 => x"dc",
          7468 => x"ec",
          7469 => x"fc",
          7470 => x"3d",
          7471 => x"53",
          7472 => x"51",
          7473 => x"3f",
          7474 => x"08",
          7475 => x"c7",
          7476 => x"bc",
          7477 => x"db",
          7478 => x"79",
          7479 => x"38",
          7480 => x"7b",
          7481 => x"5b",
          7482 => x"92",
          7483 => x"7a",
          7484 => x"53",
          7485 => x"86",
          7486 => x"fe",
          7487 => x"1a",
          7488 => x"43",
          7489 => x"82",
          7490 => x"82",
          7491 => x"3d",
          7492 => x"53",
          7493 => x"51",
          7494 => x"3f",
          7495 => x"08",
          7496 => x"82",
          7497 => x"59",
          7498 => x"89",
          7499 => x"98",
          7500 => x"cd",
          7501 => x"e1",
          7502 => x"80",
          7503 => x"82",
          7504 => x"44",
          7505 => x"89",
          7506 => x"78",
          7507 => x"38",
          7508 => x"08",
          7509 => x"82",
          7510 => x"59",
          7511 => x"88",
          7512 => x"b0",
          7513 => x"39",
          7514 => x"33",
          7515 => x"2e",
          7516 => x"89",
          7517 => x"89",
          7518 => x"c8",
          7519 => x"05",
          7520 => x"fe",
          7521 => x"ff",
          7522 => x"fe",
          7523 => x"82",
          7524 => x"80",
          7525 => x"89",
          7526 => x"78",
          7527 => x"38",
          7528 => x"08",
          7529 => x"39",
          7530 => x"33",
          7531 => x"2e",
          7532 => x"89",
          7533 => x"bb",
          7534 => x"e2",
          7535 => x"80",
          7536 => x"82",
          7537 => x"43",
          7538 => x"89",
          7539 => x"78",
          7540 => x"38",
          7541 => x"08",
          7542 => x"82",
          7543 => x"59",
          7544 => x"88",
          7545 => x"bc",
          7546 => x"39",
          7547 => x"08",
          7548 => x"b4",
          7549 => x"11",
          7550 => x"05",
          7551 => x"8c",
          7552 => x"ec",
          7553 => x"a7",
          7554 => x"5c",
          7555 => x"2e",
          7556 => x"5c",
          7557 => x"70",
          7558 => x"07",
          7559 => x"7f",
          7560 => x"5a",
          7561 => x"2e",
          7562 => x"a0",
          7563 => x"88",
          7564 => x"e8",
          7565 => x"fb",
          7566 => x"63",
          7567 => x"62",
          7568 => x"f2",
          7569 => x"86",
          7570 => x"f5",
          7571 => x"c7",
          7572 => x"ff",
          7573 => x"ff",
          7574 => x"fe",
          7575 => x"82",
          7576 => x"80",
          7577 => x"38",
          7578 => x"fc",
          7579 => x"84",
          7580 => x"fd",
          7581 => x"8c",
          7582 => x"2e",
          7583 => x"59",
          7584 => x"05",
          7585 => x"63",
          7586 => x"b4",
          7587 => x"11",
          7588 => x"05",
          7589 => x"f4",
          7590 => x"ec",
          7591 => x"f8",
          7592 => x"70",
          7593 => x"82",
          7594 => x"fe",
          7595 => x"80",
          7596 => x"51",
          7597 => x"3f",
          7598 => x"33",
          7599 => x"2e",
          7600 => x"9f",
          7601 => x"38",
          7602 => x"fc",
          7603 => x"84",
          7604 => x"fc",
          7605 => x"8c",
          7606 => x"2e",
          7607 => x"59",
          7608 => x"05",
          7609 => x"63",
          7610 => x"ff",
          7611 => x"87",
          7612 => x"f4",
          7613 => x"aa",
          7614 => x"fe",
          7615 => x"ff",
          7616 => x"fe",
          7617 => x"82",
          7618 => x"80",
          7619 => x"38",
          7620 => x"f0",
          7621 => x"84",
          7622 => x"fd",
          7623 => x"8c",
          7624 => x"2e",
          7625 => x"59",
          7626 => x"22",
          7627 => x"05",
          7628 => x"41",
          7629 => x"f0",
          7630 => x"84",
          7631 => x"fd",
          7632 => x"8c",
          7633 => x"38",
          7634 => x"60",
          7635 => x"52",
          7636 => x"51",
          7637 => x"3f",
          7638 => x"79",
          7639 => x"91",
          7640 => x"79",
          7641 => x"ae",
          7642 => x"38",
          7643 => x"87",
          7644 => x"05",
          7645 => x"b4",
          7646 => x"11",
          7647 => x"05",
          7648 => x"fa",
          7649 => x"ec",
          7650 => x"92",
          7651 => x"02",
          7652 => x"79",
          7653 => x"5b",
          7654 => x"ff",
          7655 => x"87",
          7656 => x"f3",
          7657 => x"a3",
          7658 => x"fe",
          7659 => x"ff",
          7660 => x"fe",
          7661 => x"82",
          7662 => x"80",
          7663 => x"38",
          7664 => x"f0",
          7665 => x"84",
          7666 => x"fc",
          7667 => x"8c",
          7668 => x"2e",
          7669 => x"60",
          7670 => x"60",
          7671 => x"b4",
          7672 => x"11",
          7673 => x"05",
          7674 => x"92",
          7675 => x"ec",
          7676 => x"f6",
          7677 => x"70",
          7678 => x"82",
          7679 => x"fe",
          7680 => x"80",
          7681 => x"51",
          7682 => x"3f",
          7683 => x"33",
          7684 => x"2e",
          7685 => x"9f",
          7686 => x"38",
          7687 => x"f0",
          7688 => x"84",
          7689 => x"fb",
          7690 => x"8c",
          7691 => x"2e",
          7692 => x"60",
          7693 => x"60",
          7694 => x"ff",
          7695 => x"87",
          7696 => x"f1",
          7697 => x"ae",
          7698 => x"ff",
          7699 => x"ff",
          7700 => x"fe",
          7701 => x"82",
          7702 => x"80",
          7703 => x"38",
          7704 => x"87",
          7705 => x"f7",
          7706 => x"59",
          7707 => x"3d",
          7708 => x"53",
          7709 => x"51",
          7710 => x"3f",
          7711 => x"08",
          7712 => x"93",
          7713 => x"82",
          7714 => x"fe",
          7715 => x"63",
          7716 => x"82",
          7717 => x"80",
          7718 => x"38",
          7719 => x"08",
          7720 => x"e8",
          7721 => x"ef",
          7722 => x"39",
          7723 => x"51",
          7724 => x"3f",
          7725 => x"3f",
          7726 => x"82",
          7727 => x"fe",
          7728 => x"80",
          7729 => x"39",
          7730 => x"3f",
          7731 => x"64",
          7732 => x"59",
          7733 => x"f4",
          7734 => x"7d",
          7735 => x"80",
          7736 => x"38",
          7737 => x"84",
          7738 => x"de",
          7739 => x"8c",
          7740 => x"81",
          7741 => x"2e",
          7742 => x"82",
          7743 => x"7a",
          7744 => x"38",
          7745 => x"7a",
          7746 => x"38",
          7747 => x"82",
          7748 => x"7b",
          7749 => x"b8",
          7750 => x"82",
          7751 => x"b4",
          7752 => x"05",
          7753 => x"85",
          7754 => x"82",
          7755 => x"b4",
          7756 => x"05",
          7757 => x"f5",
          7758 => x"7b",
          7759 => x"b8",
          7760 => x"82",
          7761 => x"b4",
          7762 => x"05",
          7763 => x"dd",
          7764 => x"7b",
          7765 => x"82",
          7766 => x"b4",
          7767 => x"05",
          7768 => x"c9",
          7769 => x"98",
          7770 => x"a0",
          7771 => x"64",
          7772 => x"81",
          7773 => x"54",
          7774 => x"53",
          7775 => x"52",
          7776 => x"b0",
          7777 => x"8a",
          7778 => x"ec",
          7779 => x"ec",
          7780 => x"30",
          7781 => x"80",
          7782 => x"5b",
          7783 => x"7a",
          7784 => x"38",
          7785 => x"7a",
          7786 => x"80",
          7787 => x"81",
          7788 => x"ff",
          7789 => x"7a",
          7790 => x"7d",
          7791 => x"81",
          7792 => x"78",
          7793 => x"ff",
          7794 => x"06",
          7795 => x"82",
          7796 => x"fe",
          7797 => x"f2",
          7798 => x"3d",
          7799 => x"82",
          7800 => x"87",
          7801 => x"70",
          7802 => x"87",
          7803 => x"72",
          7804 => x"c5",
          7805 => x"ec",
          7806 => x"75",
          7807 => x"87",
          7808 => x"73",
          7809 => x"b1",
          7810 => x"8c",
          7811 => x"75",
          7812 => x"94",
          7813 => x"54",
          7814 => x"80",
          7815 => x"fe",
          7816 => x"82",
          7817 => x"90",
          7818 => x"55",
          7819 => x"80",
          7820 => x"fe",
          7821 => x"72",
          7822 => x"08",
          7823 => x"8c",
          7824 => x"87",
          7825 => x"0c",
          7826 => x"0b",
          7827 => x"94",
          7828 => x"ea",
          7829 => x"fc",
          7830 => x"eb",
          7831 => x"80",
          7832 => x"b3",
          7833 => x"dc",
          7834 => x"f0",
          7835 => x"c3",
          7836 => x"fc",
          7837 => x"bb",
          7838 => x"fd",
          7839 => x"bf",
          7840 => x"ec",
          7841 => x"bf",
          7842 => x"00",
          7843 => x"00",
          7844 => x"00",
          7845 => x"00",
          7846 => x"00",
          7847 => x"00",
          7848 => x"00",
          7849 => x"00",
          7850 => x"00",
          7851 => x"00",
          7852 => x"00",
          7853 => x"00",
          7854 => x"00",
          7855 => x"00",
          7856 => x"00",
          7857 => x"00",
          7858 => x"00",
          7859 => x"00",
          7860 => x"00",
          7861 => x"00",
          7862 => x"00",
          7863 => x"00",
          7864 => x"00",
          7865 => x"00",
          7866 => x"00",
          7867 => x"25",
          7868 => x"64",
          7869 => x"20",
          7870 => x"25",
          7871 => x"64",
          7872 => x"25",
          7873 => x"53",
          7874 => x"43",
          7875 => x"69",
          7876 => x"61",
          7877 => x"6e",
          7878 => x"20",
          7879 => x"6f",
          7880 => x"6f",
          7881 => x"6f",
          7882 => x"67",
          7883 => x"3a",
          7884 => x"76",
          7885 => x"73",
          7886 => x"70",
          7887 => x"65",
          7888 => x"64",
          7889 => x"20",
          7890 => x"57",
          7891 => x"44",
          7892 => x"20",
          7893 => x"30",
          7894 => x"25",
          7895 => x"29",
          7896 => x"20",
          7897 => x"53",
          7898 => x"4d",
          7899 => x"20",
          7900 => x"30",
          7901 => x"25",
          7902 => x"29",
          7903 => x"20",
          7904 => x"49",
          7905 => x"20",
          7906 => x"4d",
          7907 => x"30",
          7908 => x"25",
          7909 => x"29",
          7910 => x"20",
          7911 => x"42",
          7912 => x"20",
          7913 => x"20",
          7914 => x"30",
          7915 => x"25",
          7916 => x"29",
          7917 => x"20",
          7918 => x"52",
          7919 => x"20",
          7920 => x"20",
          7921 => x"30",
          7922 => x"25",
          7923 => x"29",
          7924 => x"20",
          7925 => x"53",
          7926 => x"41",
          7927 => x"20",
          7928 => x"65",
          7929 => x"65",
          7930 => x"25",
          7931 => x"29",
          7932 => x"20",
          7933 => x"54",
          7934 => x"52",
          7935 => x"20",
          7936 => x"69",
          7937 => x"73",
          7938 => x"25",
          7939 => x"29",
          7940 => x"20",
          7941 => x"49",
          7942 => x"20",
          7943 => x"4c",
          7944 => x"68",
          7945 => x"65",
          7946 => x"25",
          7947 => x"29",
          7948 => x"20",
          7949 => x"57",
          7950 => x"42",
          7951 => x"20",
          7952 => x"0a",
          7953 => x"20",
          7954 => x"57",
          7955 => x"32",
          7956 => x"20",
          7957 => x"49",
          7958 => x"4c",
          7959 => x"20",
          7960 => x"50",
          7961 => x"00",
          7962 => x"20",
          7963 => x"53",
          7964 => x"00",
          7965 => x"41",
          7966 => x"65",
          7967 => x"73",
          7968 => x"20",
          7969 => x"43",
          7970 => x"52",
          7971 => x"74",
          7972 => x"63",
          7973 => x"20",
          7974 => x"72",
          7975 => x"20",
          7976 => x"30",
          7977 => x"00",
          7978 => x"20",
          7979 => x"43",
          7980 => x"4d",
          7981 => x"72",
          7982 => x"74",
          7983 => x"20",
          7984 => x"72",
          7985 => x"20",
          7986 => x"30",
          7987 => x"00",
          7988 => x"20",
          7989 => x"53",
          7990 => x"6b",
          7991 => x"61",
          7992 => x"41",
          7993 => x"65",
          7994 => x"20",
          7995 => x"20",
          7996 => x"30",
          7997 => x"00",
          7998 => x"4d",
          7999 => x"3a",
          8000 => x"20",
          8001 => x"5a",
          8002 => x"49",
          8003 => x"20",
          8004 => x"20",
          8005 => x"20",
          8006 => x"20",
          8007 => x"20",
          8008 => x"30",
          8009 => x"00",
          8010 => x"20",
          8011 => x"53",
          8012 => x"65",
          8013 => x"6c",
          8014 => x"20",
          8015 => x"71",
          8016 => x"20",
          8017 => x"20",
          8018 => x"64",
          8019 => x"34",
          8020 => x"7a",
          8021 => x"20",
          8022 => x"53",
          8023 => x"4d",
          8024 => x"6f",
          8025 => x"46",
          8026 => x"20",
          8027 => x"20",
          8028 => x"20",
          8029 => x"64",
          8030 => x"34",
          8031 => x"7a",
          8032 => x"20",
          8033 => x"57",
          8034 => x"62",
          8035 => x"20",
          8036 => x"41",
          8037 => x"6c",
          8038 => x"20",
          8039 => x"71",
          8040 => x"64",
          8041 => x"34",
          8042 => x"7a",
          8043 => x"53",
          8044 => x"6c",
          8045 => x"4d",
          8046 => x"75",
          8047 => x"46",
          8048 => x"00",
          8049 => x"45",
          8050 => x"45",
          8051 => x"69",
          8052 => x"55",
          8053 => x"6f",
          8054 => x"53",
          8055 => x"22",
          8056 => x"3a",
          8057 => x"3e",
          8058 => x"7c",
          8059 => x"46",
          8060 => x"46",
          8061 => x"32",
          8062 => x"eb",
          8063 => x"53",
          8064 => x"35",
          8065 => x"4e",
          8066 => x"41",
          8067 => x"20",
          8068 => x"41",
          8069 => x"20",
          8070 => x"4e",
          8071 => x"41",
          8072 => x"20",
          8073 => x"41",
          8074 => x"20",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"80",
          8080 => x"8e",
          8081 => x"45",
          8082 => x"49",
          8083 => x"90",
          8084 => x"99",
          8085 => x"59",
          8086 => x"9c",
          8087 => x"41",
          8088 => x"a5",
          8089 => x"a8",
          8090 => x"ac",
          8091 => x"b0",
          8092 => x"b4",
          8093 => x"b8",
          8094 => x"bc",
          8095 => x"c0",
          8096 => x"c4",
          8097 => x"c8",
          8098 => x"cc",
          8099 => x"d0",
          8100 => x"d4",
          8101 => x"d8",
          8102 => x"dc",
          8103 => x"e0",
          8104 => x"e4",
          8105 => x"e8",
          8106 => x"ec",
          8107 => x"f0",
          8108 => x"f4",
          8109 => x"f8",
          8110 => x"fc",
          8111 => x"2b",
          8112 => x"3d",
          8113 => x"5c",
          8114 => x"3c",
          8115 => x"7f",
          8116 => x"00",
          8117 => x"00",
          8118 => x"01",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"64",
          8125 => x"74",
          8126 => x"64",
          8127 => x"74",
          8128 => x"66",
          8129 => x"74",
          8130 => x"66",
          8131 => x"64",
          8132 => x"66",
          8133 => x"63",
          8134 => x"6d",
          8135 => x"61",
          8136 => x"6d",
          8137 => x"79",
          8138 => x"6d",
          8139 => x"66",
          8140 => x"6d",
          8141 => x"70",
          8142 => x"6d",
          8143 => x"6d",
          8144 => x"6d",
          8145 => x"68",
          8146 => x"68",
          8147 => x"68",
          8148 => x"68",
          8149 => x"63",
          8150 => x"00",
          8151 => x"6a",
          8152 => x"72",
          8153 => x"61",
          8154 => x"72",
          8155 => x"74",
          8156 => x"69",
          8157 => x"00",
          8158 => x"74",
          8159 => x"00",
          8160 => x"74",
          8161 => x"69",
          8162 => x"44",
          8163 => x"20",
          8164 => x"6f",
          8165 => x"49",
          8166 => x"72",
          8167 => x"20",
          8168 => x"6f",
          8169 => x"00",
          8170 => x"44",
          8171 => x"20",
          8172 => x"20",
          8173 => x"64",
          8174 => x"00",
          8175 => x"4e",
          8176 => x"69",
          8177 => x"66",
          8178 => x"64",
          8179 => x"4e",
          8180 => x"61",
          8181 => x"66",
          8182 => x"64",
          8183 => x"49",
          8184 => x"6c",
          8185 => x"66",
          8186 => x"6e",
          8187 => x"2e",
          8188 => x"41",
          8189 => x"73",
          8190 => x"65",
          8191 => x"64",
          8192 => x"46",
          8193 => x"20",
          8194 => x"65",
          8195 => x"20",
          8196 => x"73",
          8197 => x"0a",
          8198 => x"46",
          8199 => x"20",
          8200 => x"64",
          8201 => x"69",
          8202 => x"6c",
          8203 => x"0a",
          8204 => x"53",
          8205 => x"73",
          8206 => x"69",
          8207 => x"70",
          8208 => x"65",
          8209 => x"64",
          8210 => x"44",
          8211 => x"65",
          8212 => x"6d",
          8213 => x"20",
          8214 => x"69",
          8215 => x"6c",
          8216 => x"0a",
          8217 => x"44",
          8218 => x"20",
          8219 => x"20",
          8220 => x"62",
          8221 => x"2e",
          8222 => x"4e",
          8223 => x"6f",
          8224 => x"74",
          8225 => x"65",
          8226 => x"6c",
          8227 => x"73",
          8228 => x"20",
          8229 => x"6e",
          8230 => x"6e",
          8231 => x"73",
          8232 => x"00",
          8233 => x"46",
          8234 => x"61",
          8235 => x"62",
          8236 => x"65",
          8237 => x"00",
          8238 => x"54",
          8239 => x"6f",
          8240 => x"20",
          8241 => x"72",
          8242 => x"6f",
          8243 => x"61",
          8244 => x"6c",
          8245 => x"2e",
          8246 => x"46",
          8247 => x"20",
          8248 => x"6c",
          8249 => x"65",
          8250 => x"00",
          8251 => x"49",
          8252 => x"66",
          8253 => x"69",
          8254 => x"20",
          8255 => x"6f",
          8256 => x"0a",
          8257 => x"54",
          8258 => x"6d",
          8259 => x"20",
          8260 => x"6e",
          8261 => x"6c",
          8262 => x"0a",
          8263 => x"50",
          8264 => x"6d",
          8265 => x"72",
          8266 => x"6e",
          8267 => x"72",
          8268 => x"2e",
          8269 => x"53",
          8270 => x"65",
          8271 => x"0a",
          8272 => x"55",
          8273 => x"6f",
          8274 => x"65",
          8275 => x"72",
          8276 => x"0a",
          8277 => x"20",
          8278 => x"65",
          8279 => x"73",
          8280 => x"20",
          8281 => x"20",
          8282 => x"65",
          8283 => x"65",
          8284 => x"00",
          8285 => x"72",
          8286 => x"00",
          8287 => x"25",
          8288 => x"00",
          8289 => x"3a",
          8290 => x"25",
          8291 => x"00",
          8292 => x"20",
          8293 => x"20",
          8294 => x"00",
          8295 => x"25",
          8296 => x"00",
          8297 => x"20",
          8298 => x"20",
          8299 => x"7c",
          8300 => x"7a",
          8301 => x"0a",
          8302 => x"25",
          8303 => x"00",
          8304 => x"31",
          8305 => x"34",
          8306 => x"32",
          8307 => x"76",
          8308 => x"00",
          8309 => x"20",
          8310 => x"2c",
          8311 => x"76",
          8312 => x"32",
          8313 => x"25",
          8314 => x"73",
          8315 => x"0a",
          8316 => x"5a",
          8317 => x"49",
          8318 => x"72",
          8319 => x"74",
          8320 => x"6e",
          8321 => x"72",
          8322 => x"54",
          8323 => x"72",
          8324 => x"74",
          8325 => x"75",
          8326 => x"00",
          8327 => x"50",
          8328 => x"69",
          8329 => x"72",
          8330 => x"74",
          8331 => x"49",
          8332 => x"4c",
          8333 => x"20",
          8334 => x"65",
          8335 => x"70",
          8336 => x"49",
          8337 => x"4c",
          8338 => x"20",
          8339 => x"65",
          8340 => x"70",
          8341 => x"55",
          8342 => x"30",
          8343 => x"20",
          8344 => x"65",
          8345 => x"70",
          8346 => x"55",
          8347 => x"30",
          8348 => x"20",
          8349 => x"65",
          8350 => x"70",
          8351 => x"55",
          8352 => x"31",
          8353 => x"20",
          8354 => x"65",
          8355 => x"70",
          8356 => x"55",
          8357 => x"31",
          8358 => x"20",
          8359 => x"65",
          8360 => x"70",
          8361 => x"53",
          8362 => x"69",
          8363 => x"75",
          8364 => x"69",
          8365 => x"2e",
          8366 => x"00",
          8367 => x"45",
          8368 => x"6c",
          8369 => x"20",
          8370 => x"65",
          8371 => x"2e",
          8372 => x"61",
          8373 => x"65",
          8374 => x"2e",
          8375 => x"00",
          8376 => x"30",
          8377 => x"46",
          8378 => x"65",
          8379 => x"6f",
          8380 => x"69",
          8381 => x"6c",
          8382 => x"20",
          8383 => x"63",
          8384 => x"20",
          8385 => x"70",
          8386 => x"73",
          8387 => x"6e",
          8388 => x"6d",
          8389 => x"61",
          8390 => x"2e",
          8391 => x"2a",
          8392 => x"43",
          8393 => x"72",
          8394 => x"2e",
          8395 => x"00",
          8396 => x"43",
          8397 => x"69",
          8398 => x"2e",
          8399 => x"43",
          8400 => x"61",
          8401 => x"67",
          8402 => x"00",
          8403 => x"25",
          8404 => x"78",
          8405 => x"38",
          8406 => x"3e",
          8407 => x"6c",
          8408 => x"30",
          8409 => x"0a",
          8410 => x"44",
          8411 => x"20",
          8412 => x"6f",
          8413 => x"00",
          8414 => x"0a",
          8415 => x"70",
          8416 => x"65",
          8417 => x"25",
          8418 => x"20",
          8419 => x"58",
          8420 => x"3f",
          8421 => x"00",
          8422 => x"25",
          8423 => x"20",
          8424 => x"58",
          8425 => x"25",
          8426 => x"20",
          8427 => x"58",
          8428 => x"45",
          8429 => x"75",
          8430 => x"67",
          8431 => x"64",
          8432 => x"20",
          8433 => x"78",
          8434 => x"2e",
          8435 => x"43",
          8436 => x"69",
          8437 => x"63",
          8438 => x"20",
          8439 => x"30",
          8440 => x"2e",
          8441 => x"00",
          8442 => x"43",
          8443 => x"20",
          8444 => x"75",
          8445 => x"64",
          8446 => x"64",
          8447 => x"25",
          8448 => x"0a",
          8449 => x"52",
          8450 => x"61",
          8451 => x"6e",
          8452 => x"70",
          8453 => x"63",
          8454 => x"6f",
          8455 => x"2e",
          8456 => x"43",
          8457 => x"20",
          8458 => x"6f",
          8459 => x"6e",
          8460 => x"2e",
          8461 => x"5a",
          8462 => x"62",
          8463 => x"25",
          8464 => x"25",
          8465 => x"73",
          8466 => x"00",
          8467 => x"25",
          8468 => x"25",
          8469 => x"73",
          8470 => x"25",
          8471 => x"25",
          8472 => x"42",
          8473 => x"63",
          8474 => x"61",
          8475 => x"0a",
          8476 => x"52",
          8477 => x"69",
          8478 => x"2e",
          8479 => x"45",
          8480 => x"6c",
          8481 => x"20",
          8482 => x"65",
          8483 => x"70",
          8484 => x"2e",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"01",
          8495 => x"01",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"05",
          8501 => x"05",
          8502 => x"05",
          8503 => x"00",
          8504 => x"01",
          8505 => x"01",
          8506 => x"01",
          8507 => x"01",
          8508 => x"00",
          8509 => x"01",
          8510 => x"00",
          8511 => x"00",
          8512 => x"01",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"01",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"01",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"01",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"01",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"01",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"01",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"01",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"01",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"01",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"01",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"01",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"01",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"01",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"01",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"01",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"01",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"01",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"01",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"01",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"01",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"01",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"01",
          8601 => x"00",
          8602 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
