-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e9040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"cc738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cb2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8a",
           179 => x"fd2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"80040088",
           281 => x"e2040000",
           282 => x"009ff070",
           283 => x"a0a0278b",
           284 => x"38807170",
           285 => x"8405530c",
           286 => x"88eb0488",
           287 => x"e2519e99",
           288 => x"04940802",
           289 => x"940cfd3d",
           290 => x"0d805394",
           291 => x"088c0508",
           292 => x"52940888",
           293 => x"05085182",
           294 => x"de3f8808",
           295 => x"70880c54",
           296 => x"853d0d94",
           297 => x"0c049408",
           298 => x"02940cfd",
           299 => x"3d0d8153",
           300 => x"94088c05",
           301 => x"08529408",
           302 => x"88050851",
           303 => x"82b93f88",
           304 => x"0870880c",
           305 => x"54853d0d",
           306 => x"940c0494",
           307 => x"0802940c",
           308 => x"f93d0d80",
           309 => x"0b9408fc",
           310 => x"050c9408",
           311 => x"88050880",
           312 => x"25ab3894",
           313 => x"08880508",
           314 => x"30940888",
           315 => x"050c800b",
           316 => x"9408f405",
           317 => x"0c9408fc",
           318 => x"05088838",
           319 => x"810b9408",
           320 => x"f4050c94",
           321 => x"08f40508",
           322 => x"9408fc05",
           323 => x"0c94088c",
           324 => x"05088025",
           325 => x"ab389408",
           326 => x"8c050830",
           327 => x"94088c05",
           328 => x"0c800b94",
           329 => x"08f0050c",
           330 => x"9408fc05",
           331 => x"08883881",
           332 => x"0b9408f0",
           333 => x"050c9408",
           334 => x"f0050894",
           335 => x"08fc050c",
           336 => x"80539408",
           337 => x"8c050852",
           338 => x"94088805",
           339 => x"085181a7",
           340 => x"3f880870",
           341 => x"9408f805",
           342 => x"0c549408",
           343 => x"fc050880",
           344 => x"2e8c3894",
           345 => x"08f80508",
           346 => x"309408f8",
           347 => x"050c9408",
           348 => x"f8050870",
           349 => x"880c5489",
           350 => x"3d0d940c",
           351 => x"04940802",
           352 => x"940cfb3d",
           353 => x"0d800b94",
           354 => x"08fc050c",
           355 => x"94088805",
           356 => x"08802593",
           357 => x"38940888",
           358 => x"05083094",
           359 => x"0888050c",
           360 => x"810b9408",
           361 => x"fc050c94",
           362 => x"088c0508",
           363 => x"80258c38",
           364 => x"94088c05",
           365 => x"08309408",
           366 => x"8c050c81",
           367 => x"5394088c",
           368 => x"05085294",
           369 => x"08880508",
           370 => x"51ad3f88",
           371 => x"08709408",
           372 => x"f8050c54",
           373 => x"9408fc05",
           374 => x"08802e8c",
           375 => x"389408f8",
           376 => x"05083094",
           377 => x"08f8050c",
           378 => x"9408f805",
           379 => x"0870880c",
           380 => x"54873d0d",
           381 => x"940c0494",
           382 => x"0802940c",
           383 => x"fd3d0d81",
           384 => x"0b9408fc",
           385 => x"050c800b",
           386 => x"9408f805",
           387 => x"0c94088c",
           388 => x"05089408",
           389 => x"88050827",
           390 => x"ac389408",
           391 => x"fc050880",
           392 => x"2ea33880",
           393 => x"0b94088c",
           394 => x"05082499",
           395 => x"3894088c",
           396 => x"05081094",
           397 => x"088c050c",
           398 => x"9408fc05",
           399 => x"08109408",
           400 => x"fc050cc9",
           401 => x"399408fc",
           402 => x"0508802e",
           403 => x"80c93894",
           404 => x"088c0508",
           405 => x"94088805",
           406 => x"0826a138",
           407 => x"94088805",
           408 => x"0894088c",
           409 => x"05083194",
           410 => x"0888050c",
           411 => x"9408f805",
           412 => x"089408fc",
           413 => x"05080794",
           414 => x"08f8050c",
           415 => x"9408fc05",
           416 => x"08812a94",
           417 => x"08fc050c",
           418 => x"94088c05",
           419 => x"08812a94",
           420 => x"088c050c",
           421 => x"ffaf3994",
           422 => x"08900508",
           423 => x"802e8f38",
           424 => x"94088805",
           425 => x"08709408",
           426 => x"f4050c51",
           427 => x"8d399408",
           428 => x"f8050870",
           429 => x"9408f405",
           430 => x"0c519408",
           431 => x"f4050888",
           432 => x"0c853d0d",
           433 => x"940c04ff",
           434 => x"3d0d8188",
           435 => x"0b87c092",
           436 => x"8c0c810b",
           437 => x"87c0928c",
           438 => x"0c850b87",
           439 => x"c0988c0c",
           440 => x"87c0928c",
           441 => x"08708206",
           442 => x"51517080",
           443 => x"2e8a3887",
           444 => x"c0988c08",
           445 => x"5170e938",
           446 => x"87c0928c",
           447 => x"08fc8080",
           448 => x"06527193",
           449 => x"3887c098",
           450 => x"8c085170",
           451 => x"802e8838",
           452 => x"710b0b0b",
           453 => x"9fec340b",
           454 => x"0b0b9fec",
           455 => x"33880c83",
           456 => x"3d0d04fa",
           457 => x"3d0d787b",
           458 => x"7d565856",
           459 => x"800b0b0b",
           460 => x"0b9fec33",
           461 => x"81065255",
           462 => x"82527075",
           463 => x"2e098106",
           464 => x"819e3885",
           465 => x"0b87c098",
           466 => x"8c0c7987",
           467 => x"c092800c",
           468 => x"840b87c0",
           469 => x"928c0c87",
           470 => x"c0928c08",
           471 => x"70852a70",
           472 => x"81065152",
           473 => x"5370802e",
           474 => x"a73887c0",
           475 => x"92840870",
           476 => x"81ff0676",
           477 => x"79275253",
           478 => x"5173802e",
           479 => x"90387080",
           480 => x"2e8b3871",
           481 => x"76708105",
           482 => x"5834ff14",
           483 => x"54811555",
           484 => x"72a20651",
           485 => x"70802e8b",
           486 => x"3887c098",
           487 => x"8c085170",
           488 => x"ffb53887",
           489 => x"c0988c08",
           490 => x"51709538",
           491 => x"810b87c0",
           492 => x"928c0c87",
           493 => x"c0928c08",
           494 => x"70820651",
           495 => x"5170f438",
           496 => x"8073fc80",
           497 => x"80065252",
           498 => x"70722e09",
           499 => x"81068f38",
           500 => x"87c0988c",
           501 => x"08517072",
           502 => x"2e098106",
           503 => x"83388152",
           504 => x"71880c88",
           505 => x"3d0d04fe",
           506 => x"3d0d7481",
           507 => x"11337133",
           508 => x"71882b07",
           509 => x"880c5351",
           510 => x"843d0d04",
           511 => x"fd3d0d75",
           512 => x"83113382",
           513 => x"12337190",
           514 => x"2b71882b",
           515 => x"07811433",
           516 => x"70720788",
           517 => x"2b753371",
           518 => x"07880c52",
           519 => x"53545654",
           520 => x"52853d0d",
           521 => x"04f93d0d",
           522 => x"790b0b0b",
           523 => x"9ff00857",
           524 => x"57817727",
           525 => x"80ed3876",
           526 => x"88170827",
           527 => x"80e53875",
           528 => x"33557482",
           529 => x"2e893874",
           530 => x"832eae38",
           531 => x"80d53974",
           532 => x"54761083",
           533 => x"fe065376",
           534 => x"882a8c17",
           535 => x"08055288",
           536 => x"3d705255",
           537 => x"fdbd3f88",
           538 => x"08b93874",
           539 => x"51fef83f",
           540 => x"880883ff",
           541 => x"ff0655ad",
           542 => x"39845476",
           543 => x"822b83fc",
           544 => x"06537687",
           545 => x"2a8c1708",
           546 => x"0552883d",
           547 => x"705255fd",
           548 => x"923f8808",
           549 => x"8e387451",
           550 => x"fee23f88",
           551 => x"08f00a06",
           552 => x"55833981",
           553 => x"5574880c",
           554 => x"893d0d04",
           555 => x"fb3d0d0b",
           556 => x"0b0b9ff0",
           557 => x"08fe1988",
           558 => x"1208fe05",
           559 => x"55565480",
           560 => x"56747327",
           561 => x"8d388214",
           562 => x"33757129",
           563 => x"94160805",
           564 => x"57537588",
           565 => x"0c873d0d",
           566 => x"04fd3d0d",
           567 => x"7554800b",
           568 => x"0b0b0b9f",
           569 => x"f0087033",
           570 => x"51535371",
           571 => x"832e0981",
           572 => x"068c3894",
           573 => x"1451fdef",
           574 => x"3f880890",
           575 => x"2b539a14",
           576 => x"51fde43f",
           577 => x"880883ff",
           578 => x"ff067307",
           579 => x"880c853d",
           580 => x"0d04fc3d",
           581 => x"0d760b0b",
           582 => x"0b9ff008",
           583 => x"55558075",
           584 => x"23881508",
           585 => x"5372812e",
           586 => x"88388814",
           587 => x"08732685",
           588 => x"388152b0",
           589 => x"39729038",
           590 => x"73335271",
           591 => x"832e0981",
           592 => x"06853890",
           593 => x"14085372",
           594 => x"8c160c72",
           595 => x"802e8b38",
           596 => x"7251fed8",
           597 => x"3f880852",
           598 => x"85399014",
           599 => x"08527190",
           600 => x"160c8052",
           601 => x"71880c86",
           602 => x"3d0d04fa",
           603 => x"3d0d780b",
           604 => x"0b0b9ff0",
           605 => x"08712281",
           606 => x"057083ff",
           607 => x"ff065754",
           608 => x"57557380",
           609 => x"2e883890",
           610 => x"15085372",
           611 => x"86388352",
           612 => x"80dc3973",
           613 => x"8f065271",
           614 => x"80cf3881",
           615 => x"1390160c",
           616 => x"8c150853",
           617 => x"728f3883",
           618 => x"0b841722",
           619 => x"57527376",
           620 => x"27bc38b5",
           621 => x"39821633",
           622 => x"ff057484",
           623 => x"2a065271",
           624 => x"a8387251",
           625 => x"fcdf3f81",
           626 => x"52718808",
           627 => x"27a03883",
           628 => x"52880888",
           629 => x"17082796",
           630 => x"3888088c",
           631 => x"160c8808",
           632 => x"51fdc93f",
           633 => x"88089016",
           634 => x"0c737523",
           635 => x"80527188",
           636 => x"0c883d0d",
           637 => x"04f23d0d",
           638 => x"60626458",
           639 => x"5e5c7533",
           640 => x"5574a02e",
           641 => x"09810688",
           642 => x"38811670",
           643 => x"4456ef39",
           644 => x"62703356",
           645 => x"5674af2e",
           646 => x"09810684",
           647 => x"38811643",
           648 => x"800b881d",
           649 => x"0c627033",
           650 => x"5155749f",
           651 => x"268f387b",
           652 => x"51fddf3f",
           653 => x"88085680",
           654 => x"7d3482d3",
           655 => x"39933d84",
           656 => x"1d087058",
           657 => x"5a5f8a55",
           658 => x"a0767081",
           659 => x"055834ff",
           660 => x"155574ff",
           661 => x"2e098106",
           662 => x"ef388070",
           663 => x"595b887f",
           664 => x"085f5a7a",
           665 => x"811c7081",
           666 => x"ff066013",
           667 => x"703370af",
           668 => x"327030a0",
           669 => x"73277180",
           670 => x"25075151",
           671 => x"525b535d",
           672 => x"57557480",
           673 => x"c73876ae",
           674 => x"2e098106",
           675 => x"83388155",
           676 => x"777a2775",
           677 => x"07557480",
           678 => x"2e9f3879",
           679 => x"88327030",
           680 => x"78ae3270",
           681 => x"30707307",
           682 => x"9f2a5351",
           683 => x"57515675",
           684 => x"9b388858",
           685 => x"8b5affab",
           686 => x"39778119",
           687 => x"7081ff06",
           688 => x"721c535a",
           689 => x"57557675",
           690 => x"34ff9839",
           691 => x"7a1e7f0c",
           692 => x"805576a0",
           693 => x"26833881",
           694 => x"55748b1a",
           695 => x"347b51fc",
           696 => x"b13f8808",
           697 => x"80ef38a0",
           698 => x"547b2270",
           699 => x"852b83e0",
           700 => x"06545590",
           701 => x"1c08527c",
           702 => x"51f8a83f",
           703 => x"88085788",
           704 => x"0880fb38",
           705 => x"7c335574",
           706 => x"802e80ee",
           707 => x"388b1d33",
           708 => x"70832a70",
           709 => x"81065156",
           710 => x"5674b238",
           711 => x"8b7d841e",
           712 => x"08880859",
           713 => x"5b5b58ff",
           714 => x"185877ff",
           715 => x"2e9a3879",
           716 => x"7081055b",
           717 => x"33797081",
           718 => x"055b3371",
           719 => x"71315256",
           720 => x"5675802e",
           721 => x"e2388639",
           722 => x"75802e92",
           723 => x"387b51fc",
           724 => x"9a3fff8e",
           725 => x"39880856",
           726 => x"8808b438",
           727 => x"83397656",
           728 => x"841c088b",
           729 => x"11335155",
           730 => x"74a5388b",
           731 => x"1d337084",
           732 => x"2a708106",
           733 => x"51565674",
           734 => x"89388356",
           735 => x"92398156",
           736 => x"8e397c51",
           737 => x"fad33f88",
           738 => x"08881d0c",
           739 => x"fdaf3975",
           740 => x"880c903d",
           741 => x"0d04f93d",
           742 => x"0d797b59",
           743 => x"57825483",
           744 => x"fe537752",
           745 => x"7651f6fb",
           746 => x"3f835688",
           747 => x"0880e738",
           748 => x"7651f8b3",
           749 => x"3f880883",
           750 => x"ffff0655",
           751 => x"82567482",
           752 => x"d4d52e09",
           753 => x"810680ce",
           754 => x"387554b6",
           755 => x"53775276",
           756 => x"51f6d03f",
           757 => x"88085688",
           758 => x"08943876",
           759 => x"51f8883f",
           760 => x"880883ff",
           761 => x"ff065574",
           762 => x"8182c62e",
           763 => x"a9388254",
           764 => x"80d25377",
           765 => x"527651f6",
           766 => x"aa3f8808",
           767 => x"56880894",
           768 => x"387651f7",
           769 => x"e23f8808",
           770 => x"83ffff06",
           771 => x"55748182",
           772 => x"c62e8338",
           773 => x"81567588",
           774 => x"0c893d0d",
           775 => x"04ed3d0d",
           776 => x"6559800b",
           777 => x"0b0b0b9f",
           778 => x"f00cf59b",
           779 => x"3f880881",
           780 => x"06558256",
           781 => x"7482f238",
           782 => x"7475538d",
           783 => x"3d705357",
           784 => x"5afed33f",
           785 => x"880881ff",
           786 => x"06577681",
           787 => x"2e098106",
           788 => x"b3389054",
           789 => x"83be5374",
           790 => x"527551f5",
           791 => x"c63f8808",
           792 => x"ab388d3d",
           793 => x"33557480",
           794 => x"2eac3895",
           795 => x"3de40551",
           796 => x"f78a3f88",
           797 => x"08880853",
           798 => x"76525afe",
           799 => x"993f8808",
           800 => x"81ff0657",
           801 => x"76832e09",
           802 => x"81068638",
           803 => x"81568299",
           804 => x"3976802e",
           805 => x"86388656",
           806 => x"828f39a4",
           807 => x"548d5379",
           808 => x"527551f4",
           809 => x"fe3f8156",
           810 => x"880881fd",
           811 => x"38953de5",
           812 => x"0551f6b3",
           813 => x"3f880883",
           814 => x"ffff0658",
           815 => x"778c3895",
           816 => x"3df30551",
           817 => x"f6b63f88",
           818 => x"085802af",
           819 => x"05337871",
           820 => x"29028805",
           821 => x"ad057054",
           822 => x"52595bf6",
           823 => x"8a3f8808",
           824 => x"83ffff06",
           825 => x"7a058c1a",
           826 => x"0c8c3d33",
           827 => x"821a3495",
           828 => x"3de00551",
           829 => x"f5f13f88",
           830 => x"08841a23",
           831 => x"953de205",
           832 => x"51f5e43f",
           833 => x"880883ff",
           834 => x"ff065675",
           835 => x"8c38953d",
           836 => x"ef0551f5",
           837 => x"e73f8808",
           838 => x"567a51f5",
           839 => x"ca3f8808",
           840 => x"83ffff06",
           841 => x"76713179",
           842 => x"31841b22",
           843 => x"70842a82",
           844 => x"1d335672",
           845 => x"71315559",
           846 => x"5c5155ee",
           847 => x"c43f8808",
           848 => x"82057088",
           849 => x"1b0c8808",
           850 => x"e08a0556",
           851 => x"567483df",
           852 => x"fe268338",
           853 => x"825783ff",
           854 => x"f6762785",
           855 => x"38835789",
           856 => x"39865676",
           857 => x"802e80c1",
           858 => x"38767934",
           859 => x"76832e09",
           860 => x"81069038",
           861 => x"953dfb05",
           862 => x"51f5813f",
           863 => x"8808901a",
           864 => x"0c88398c",
           865 => x"19081890",
           866 => x"1a0c7983",
           867 => x"ffff068c",
           868 => x"1a081971",
           869 => x"842a0594",
           870 => x"1b0c5580",
           871 => x"0b811a34",
           872 => x"780b0b0b",
           873 => x"9ff00c80",
           874 => x"5675880c",
           875 => x"953d0d04",
           876 => x"ea3d0d0b",
           877 => x"0b0b9ff0",
           878 => x"08558554",
           879 => x"74802e80",
           880 => x"df38800b",
           881 => x"81163498",
           882 => x"3de01145",
           883 => x"6954893d",
           884 => x"705457ec",
           885 => x"0551f89d",
           886 => x"3f880854",
           887 => x"880880c0",
           888 => x"38883d33",
           889 => x"5473802e",
           890 => x"933802a7",
           891 => x"05337084",
           892 => x"2a708106",
           893 => x"51555773",
           894 => x"802e8538",
           895 => x"8354a139",
           896 => x"7551f5d5",
           897 => x"3f8808a0",
           898 => x"160c983d",
           899 => x"dc0551f3",
           900 => x"eb3f8808",
           901 => x"9c160c73",
           902 => x"98160c81",
           903 => x"0b811634",
           904 => x"73880c98",
           905 => x"3d0d04f6",
           906 => x"3d0d7d7f",
           907 => x"7e0b0b0b",
           908 => x"9ff00859",
           909 => x"5b5c5880",
           910 => x"7b0c8557",
           911 => x"75802e81",
           912 => x"d1388116",
           913 => x"33810655",
           914 => x"84577480",
           915 => x"2e81c338",
           916 => x"91397481",
           917 => x"17348639",
           918 => x"800b8117",
           919 => x"34815781",
           920 => x"b1399c16",
           921 => x"08981708",
           922 => x"31557478",
           923 => x"27833874",
           924 => x"5877802e",
           925 => x"819a3898",
           926 => x"16087083",
           927 => x"ff065657",
           928 => x"7480c738",
           929 => x"821633ff",
           930 => x"0577892a",
           931 => x"067081ff",
           932 => x"065b5579",
           933 => x"9e387687",
           934 => x"38a01608",
           935 => x"558b39a4",
           936 => x"160851f3",
           937 => x"803f8808",
           938 => x"55817527",
           939 => x"ffaa3874",
           940 => x"a4170ca4",
           941 => x"160851f3",
           942 => x"f33f8808",
           943 => x"55880880",
           944 => x"2eff8f38",
           945 => x"88081aa8",
           946 => x"170c9816",
           947 => x"0883ff06",
           948 => x"84807131",
           949 => x"51557775",
           950 => x"27833877",
           951 => x"55745498",
           952 => x"160883ff",
           953 => x"0653a816",
           954 => x"08527851",
           955 => x"f0b53f88",
           956 => x"08fee538",
           957 => x"98160815",
           958 => x"98170c77",
           959 => x"75317b08",
           960 => x"167c0c58",
           961 => x"78802efe",
           962 => x"e8387419",
           963 => x"59fee239",
           964 => x"80577688",
           965 => x"0c8c3d0d",
           966 => x"04fb3d0d",
           967 => x"87c0948c",
           968 => x"08548784",
           969 => x"80527351",
           970 => x"ead73f88",
           971 => x"08902b87",
           972 => x"c0948c08",
           973 => x"56548784",
           974 => x"80527451",
           975 => x"eac33f73",
           976 => x"88080787",
           977 => x"c0948c0c",
           978 => x"87c0949c",
           979 => x"08548784",
           980 => x"80527351",
           981 => x"eaab3f88",
           982 => x"08902b87",
           983 => x"c0949c08",
           984 => x"56548784",
           985 => x"80527451",
           986 => x"ea973f73",
           987 => x"88080787",
           988 => x"c0949c0c",
           989 => x"8c80830b",
           990 => x"87c09484",
           991 => x"0c8c8083",
           992 => x"0b87c094",
           993 => x"940c9ff4",
           994 => x"51f9923f",
           995 => x"8808b838",
           996 => x"9fdc51fc",
           997 => x"9b3f8808",
           998 => x"ae38a080",
           999 => x"0b880887",
          1000 => x"c098880c",
          1001 => x"55873dfc",
          1002 => x"05538480",
          1003 => x"527451fc",
          1004 => x"f63f8808",
          1005 => x"8d387554",
          1006 => x"73802e86",
          1007 => x"38731555",
          1008 => x"e439a080",
          1009 => x"54730480",
          1010 => x"54fb3900",
          1011 => x"00ffffff",
          1012 => x"ff00ffff",
          1013 => x"ffff00ff",
          1014 => x"ffffff00",
          1015 => x"424f4f54",
          1016 => x"54494e59",
          1017 => x"2e524f4d",
          1018 => x"00000000",
          1019 => x"01000000",
          2048 => x"0b0b0b92",
          2049 => x"d8040000",
          2050 => x"00000000",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b92",
          2121 => x"bc040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b929f",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b81c5",
          2210 => x"f0738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"92a40400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b0b93",
          2219 => x"dd2d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b0b95",
          2227 => x"c92d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"94040b0b",
          2317 => x"0b8ca304",
          2318 => x"0b0b0b8c",
          2319 => x"b2040b0b",
          2320 => x"0b8cc104",
          2321 => x"0b0b0b8c",
          2322 => x"d0040b0b",
          2323 => x"0b8cdf04",
          2324 => x"0b0b0b8c",
          2325 => x"ee040b0b",
          2326 => x"0b8cfd04",
          2327 => x"0b0b0b8d",
          2328 => x"8c040b0b",
          2329 => x"0b8d9b04",
          2330 => x"0b0b0b8d",
          2331 => x"aa040b0b",
          2332 => x"0b8db904",
          2333 => x"0b0b0b8d",
          2334 => x"c8040b0b",
          2335 => x"0b8dd704",
          2336 => x"0b0b0b8d",
          2337 => x"e6040b0b",
          2338 => x"0b8df504",
          2339 => x"0b0b0b8e",
          2340 => x"84040b0b",
          2341 => x"0b8e9404",
          2342 => x"0b0b0b8e",
          2343 => x"a4040b0b",
          2344 => x"0b8eb404",
          2345 => x"0b0b0b8e",
          2346 => x"c4040b0b",
          2347 => x"0b8ed404",
          2348 => x"0b0b0b8e",
          2349 => x"e4040b0b",
          2350 => x"0b8ef404",
          2351 => x"0b0b0b8f",
          2352 => x"84040b0b",
          2353 => x"0b8f9404",
          2354 => x"0b0b0b8f",
          2355 => x"a4040b0b",
          2356 => x"0b8fb404",
          2357 => x"0b0b0b8f",
          2358 => x"c4040b0b",
          2359 => x"0b8fd404",
          2360 => x"0b0b0b8f",
          2361 => x"e4040b0b",
          2362 => x"0b8ff404",
          2363 => x"0b0b0b90",
          2364 => x"84040b0b",
          2365 => x"0b909404",
          2366 => x"0b0b0b90",
          2367 => x"a4040b0b",
          2368 => x"0b90b404",
          2369 => x"0b0b0b90",
          2370 => x"c4040b0b",
          2371 => x"0b90d404",
          2372 => x"0b0b0b90",
          2373 => x"e4040b0b",
          2374 => x"0b90f404",
          2375 => x"0b0b0b91",
          2376 => x"84040b0b",
          2377 => x"0b919404",
          2378 => x"0b0b0b91",
          2379 => x"a3040b0b",
          2380 => x"0b91b204",
          2381 => x"0b0b0b91",
          2382 => x"c1040b0b",
          2383 => x"0b91d004",
          2384 => x"0b0b0b91",
          2385 => x"df040b0b",
          2386 => x"0b91ee04",
          2387 => x"ffffffff",
          2388 => x"ffffffff",
          2389 => x"ffffffff",
          2390 => x"ffffffff",
          2391 => x"ffffffff",
          2392 => x"ffffffff",
          2393 => x"ffffffff",
          2394 => x"ffffffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0481decc",
          2434 => x"0ca0ae2d",
          2435 => x"81decc08",
          2436 => x"82809004",
          2437 => x"81decc0c",
          2438 => x"ade22d81",
          2439 => x"decc0882",
          2440 => x"80900481",
          2441 => x"decc0cae",
          2442 => x"a12d81de",
          2443 => x"cc088280",
          2444 => x"900481de",
          2445 => x"cc0caebf",
          2446 => x"2d81decc",
          2447 => x"08828090",
          2448 => x"0481decc",
          2449 => x"0cb4fd2d",
          2450 => x"81decc08",
          2451 => x"82809004",
          2452 => x"81decc0c",
          2453 => x"b5fb2d81",
          2454 => x"decc0882",
          2455 => x"80900481",
          2456 => x"decc0cae",
          2457 => x"e22d81de",
          2458 => x"cc088280",
          2459 => x"900481de",
          2460 => x"cc0cb698",
          2461 => x"2d81decc",
          2462 => x"08828090",
          2463 => x"0481decc",
          2464 => x"0cb88a2d",
          2465 => x"81decc08",
          2466 => x"82809004",
          2467 => x"81decc0c",
          2468 => x"b4a32d81",
          2469 => x"decc0882",
          2470 => x"80900481",
          2471 => x"decc0cb4",
          2472 => x"b92d81de",
          2473 => x"cc088280",
          2474 => x"900481de",
          2475 => x"cc0cb4dd",
          2476 => x"2d81decc",
          2477 => x"08828090",
          2478 => x"0481decc",
          2479 => x"0ca2bb2d",
          2480 => x"81decc08",
          2481 => x"82809004",
          2482 => x"81decc0c",
          2483 => x"a38c2d81",
          2484 => x"decc0882",
          2485 => x"80900481",
          2486 => x"decc0c9b",
          2487 => x"a82d81de",
          2488 => x"cc088280",
          2489 => x"900481de",
          2490 => x"cc0c9cdd",
          2491 => x"2d81decc",
          2492 => x"08828090",
          2493 => x"0481decc",
          2494 => x"0c9e902d",
          2495 => x"81decc08",
          2496 => x"82809004",
          2497 => x"81decc0c",
          2498 => x"80eabf2d",
          2499 => x"81decc08",
          2500 => x"82809004",
          2501 => x"81decc0c",
          2502 => x"80f7b02d",
          2503 => x"81decc08",
          2504 => x"82809004",
          2505 => x"81decc0c",
          2506 => x"80efa42d",
          2507 => x"81decc08",
          2508 => x"82809004",
          2509 => x"81decc0c",
          2510 => x"80f2a12d",
          2511 => x"81decc08",
          2512 => x"82809004",
          2513 => x"81decc0c",
          2514 => x"80fcbf2d",
          2515 => x"81decc08",
          2516 => x"82809004",
          2517 => x"81decc0c",
          2518 => x"81859f2d",
          2519 => x"81decc08",
          2520 => x"82809004",
          2521 => x"81decc0c",
          2522 => x"80f6922d",
          2523 => x"81decc08",
          2524 => x"82809004",
          2525 => x"81decc0c",
          2526 => x"80ffde2d",
          2527 => x"81decc08",
          2528 => x"82809004",
          2529 => x"81decc0c",
          2530 => x"8180fd2d",
          2531 => x"81decc08",
          2532 => x"82809004",
          2533 => x"81decc0c",
          2534 => x"81819c2d",
          2535 => x"81decc08",
          2536 => x"82809004",
          2537 => x"81decc0c",
          2538 => x"8189862d",
          2539 => x"81decc08",
          2540 => x"82809004",
          2541 => x"81decc0c",
          2542 => x"8186ec2d",
          2543 => x"81decc08",
          2544 => x"82809004",
          2545 => x"81decc0c",
          2546 => x"818bda2d",
          2547 => x"81decc08",
          2548 => x"82809004",
          2549 => x"81decc0c",
          2550 => x"8182a02d",
          2551 => x"81decc08",
          2552 => x"82809004",
          2553 => x"81decc0c",
          2554 => x"818eda2d",
          2555 => x"81decc08",
          2556 => x"82809004",
          2557 => x"81decc0c",
          2558 => x"818fdb2d",
          2559 => x"81decc08",
          2560 => x"82809004",
          2561 => x"81decc0c",
          2562 => x"80f8902d",
          2563 => x"81decc08",
          2564 => x"82809004",
          2565 => x"81decc0c",
          2566 => x"80f7e92d",
          2567 => x"81decc08",
          2568 => x"82809004",
          2569 => x"81decc0c",
          2570 => x"80f9942d",
          2571 => x"81decc08",
          2572 => x"82809004",
          2573 => x"81decc0c",
          2574 => x"8182f72d",
          2575 => x"81decc08",
          2576 => x"82809004",
          2577 => x"81decc0c",
          2578 => x"8190cc2d",
          2579 => x"81decc08",
          2580 => x"82809004",
          2581 => x"81decc0c",
          2582 => x"8192d62d",
          2583 => x"81decc08",
          2584 => x"82809004",
          2585 => x"81decc0c",
          2586 => x"8196982d",
          2587 => x"81decc08",
          2588 => x"82809004",
          2589 => x"81decc0c",
          2590 => x"80e9de2d",
          2591 => x"81decc08",
          2592 => x"82809004",
          2593 => x"81decc0c",
          2594 => x"8199842d",
          2595 => x"81decc08",
          2596 => x"82809004",
          2597 => x"81decc0c",
          2598 => x"bb992d81",
          2599 => x"decc0882",
          2600 => x"80900481",
          2601 => x"decc0cbd",
          2602 => x"832d81de",
          2603 => x"cc088280",
          2604 => x"900481de",
          2605 => x"cc0cbee7",
          2606 => x"2d81decc",
          2607 => x"08828090",
          2608 => x"0481decc",
          2609 => x"0c9bd12d",
          2610 => x"81decc08",
          2611 => x"82809004",
          2612 => x"81decc0c",
          2613 => x"9cb32d81",
          2614 => x"decc0882",
          2615 => x"80900481",
          2616 => x"decc0c9f",
          2617 => x"a02d81de",
          2618 => x"cc088280",
          2619 => x"900481de",
          2620 => x"cc0c81a5",
          2621 => x"ff2d81de",
          2622 => x"cc088280",
          2623 => x"90043c04",
          2624 => x"10101010",
          2625 => x"10101010",
          2626 => x"10101010",
          2627 => x"10101010",
          2628 => x"10101010",
          2629 => x"10101010",
          2630 => x"10101010",
          2631 => x"10101053",
          2632 => x"51040000",
          2633 => x"7381ff06",
          2634 => x"73830609",
          2635 => x"81058305",
          2636 => x"1010102b",
          2637 => x"0772fc06",
          2638 => x"0c515104",
          2639 => x"72728072",
          2640 => x"8106ff05",
          2641 => x"09720605",
          2642 => x"71105272",
          2643 => x"0a100a53",
          2644 => x"72ed3851",
          2645 => x"51535104",
          2646 => x"81dec070",
          2647 => x"81f5ec27",
          2648 => x"8e388071",
          2649 => x"70840553",
          2650 => x"0c0b0b0b",
          2651 => x"92db048c",
          2652 => x"815181c4",
          2653 => x"be040081",
          2654 => x"decc0802",
          2655 => x"81decc0c",
          2656 => x"fd3d0d80",
          2657 => x"5381decc",
          2658 => x"088c0508",
          2659 => x"5281decc",
          2660 => x"08880508",
          2661 => x"5183d43f",
          2662 => x"81dec008",
          2663 => x"7081dec0",
          2664 => x"0c54853d",
          2665 => x"0d81decc",
          2666 => x"0c0481de",
          2667 => x"cc080281",
          2668 => x"decc0cfd",
          2669 => x"3d0d8153",
          2670 => x"81decc08",
          2671 => x"8c050852",
          2672 => x"81decc08",
          2673 => x"88050851",
          2674 => x"83a13f81",
          2675 => x"dec00870",
          2676 => x"81dec00c",
          2677 => x"54853d0d",
          2678 => x"81decc0c",
          2679 => x"0481decc",
          2680 => x"080281de",
          2681 => x"cc0cf93d",
          2682 => x"0d800b81",
          2683 => x"decc08fc",
          2684 => x"050c81de",
          2685 => x"cc088805",
          2686 => x"088025b9",
          2687 => x"3881decc",
          2688 => x"08880508",
          2689 => x"3081decc",
          2690 => x"0888050c",
          2691 => x"800b81de",
          2692 => x"cc08f405",
          2693 => x"0c81decc",
          2694 => x"08fc0508",
          2695 => x"8a38810b",
          2696 => x"81decc08",
          2697 => x"f4050c81",
          2698 => x"decc08f4",
          2699 => x"050881de",
          2700 => x"cc08fc05",
          2701 => x"0c81decc",
          2702 => x"088c0508",
          2703 => x"8025b938",
          2704 => x"81decc08",
          2705 => x"8c050830",
          2706 => x"81decc08",
          2707 => x"8c050c80",
          2708 => x"0b81decc",
          2709 => x"08f0050c",
          2710 => x"81decc08",
          2711 => x"fc05088a",
          2712 => x"38810b81",
          2713 => x"decc08f0",
          2714 => x"050c81de",
          2715 => x"cc08f005",
          2716 => x"0881decc",
          2717 => x"08fc050c",
          2718 => x"805381de",
          2719 => x"cc088c05",
          2720 => x"085281de",
          2721 => x"cc088805",
          2722 => x"085181df",
          2723 => x"3f81dec0",
          2724 => x"087081de",
          2725 => x"cc08f805",
          2726 => x"0c5481de",
          2727 => x"cc08fc05",
          2728 => x"08802e90",
          2729 => x"3881decc",
          2730 => x"08f80508",
          2731 => x"3081decc",
          2732 => x"08f8050c",
          2733 => x"81decc08",
          2734 => x"f8050870",
          2735 => x"81dec00c",
          2736 => x"54893d0d",
          2737 => x"81decc0c",
          2738 => x"0481decc",
          2739 => x"080281de",
          2740 => x"cc0cfb3d",
          2741 => x"0d800b81",
          2742 => x"decc08fc",
          2743 => x"050c81de",
          2744 => x"cc088805",
          2745 => x"08802599",
          2746 => x"3881decc",
          2747 => x"08880508",
          2748 => x"3081decc",
          2749 => x"0888050c",
          2750 => x"810b81de",
          2751 => x"cc08fc05",
          2752 => x"0c81decc",
          2753 => x"088c0508",
          2754 => x"80259038",
          2755 => x"81decc08",
          2756 => x"8c050830",
          2757 => x"81decc08",
          2758 => x"8c050c81",
          2759 => x"5381decc",
          2760 => x"088c0508",
          2761 => x"5281decc",
          2762 => x"08880508",
          2763 => x"51bd3f81",
          2764 => x"dec00870",
          2765 => x"81decc08",
          2766 => x"f8050c54",
          2767 => x"81decc08",
          2768 => x"fc050880",
          2769 => x"2e903881",
          2770 => x"decc08f8",
          2771 => x"05083081",
          2772 => x"decc08f8",
          2773 => x"050c81de",
          2774 => x"cc08f805",
          2775 => x"087081de",
          2776 => x"c00c5487",
          2777 => x"3d0d81de",
          2778 => x"cc0c0481",
          2779 => x"decc0802",
          2780 => x"81decc0c",
          2781 => x"fd3d0d81",
          2782 => x"0b81decc",
          2783 => x"08fc050c",
          2784 => x"800b81de",
          2785 => x"cc08f805",
          2786 => x"0c81decc",
          2787 => x"088c0508",
          2788 => x"81decc08",
          2789 => x"88050827",
          2790 => x"b93881de",
          2791 => x"cc08fc05",
          2792 => x"08802eae",
          2793 => x"38800b81",
          2794 => x"decc088c",
          2795 => x"050824a2",
          2796 => x"3881decc",
          2797 => x"088c0508",
          2798 => x"1081decc",
          2799 => x"088c050c",
          2800 => x"81decc08",
          2801 => x"fc050810",
          2802 => x"81decc08",
          2803 => x"fc050cff",
          2804 => x"b83981de",
          2805 => x"cc08fc05",
          2806 => x"08802e80",
          2807 => x"e13881de",
          2808 => x"cc088c05",
          2809 => x"0881decc",
          2810 => x"08880508",
          2811 => x"26ad3881",
          2812 => x"decc0888",
          2813 => x"050881de",
          2814 => x"cc088c05",
          2815 => x"083181de",
          2816 => x"cc088805",
          2817 => x"0c81decc",
          2818 => x"08f80508",
          2819 => x"81decc08",
          2820 => x"fc050807",
          2821 => x"81decc08",
          2822 => x"f8050c81",
          2823 => x"decc08fc",
          2824 => x"0508812a",
          2825 => x"81decc08",
          2826 => x"fc050c81",
          2827 => x"decc088c",
          2828 => x"0508812a",
          2829 => x"81decc08",
          2830 => x"8c050cff",
          2831 => x"953981de",
          2832 => x"cc089005",
          2833 => x"08802e93",
          2834 => x"3881decc",
          2835 => x"08880508",
          2836 => x"7081decc",
          2837 => x"08f4050c",
          2838 => x"51913981",
          2839 => x"decc08f8",
          2840 => x"05087081",
          2841 => x"decc08f4",
          2842 => x"050c5181",
          2843 => x"decc08f4",
          2844 => x"050881de",
          2845 => x"c00c853d",
          2846 => x"0d81decc",
          2847 => x"0c04fc3d",
          2848 => x"0d767971",
          2849 => x"028c059f",
          2850 => x"05335755",
          2851 => x"53558372",
          2852 => x"278a3874",
          2853 => x"83065170",
          2854 => x"802ea438",
          2855 => x"ff125271",
          2856 => x"ff2e9338",
          2857 => x"73737081",
          2858 => x"055534ff",
          2859 => x"125271ff",
          2860 => x"2e098106",
          2861 => x"ef387481",
          2862 => x"dec00c86",
          2863 => x"3d0d0474",
          2864 => x"74882b75",
          2865 => x"07707190",
          2866 => x"2b075154",
          2867 => x"518f7227",
          2868 => x"a5387271",
          2869 => x"70840553",
          2870 => x"0c727170",
          2871 => x"8405530c",
          2872 => x"72717084",
          2873 => x"05530c72",
          2874 => x"71708405",
          2875 => x"530cf012",
          2876 => x"52718f26",
          2877 => x"dd388372",
          2878 => x"27903872",
          2879 => x"71708405",
          2880 => x"530cfc12",
          2881 => x"52718326",
          2882 => x"f2387053",
          2883 => x"ff8e39fb",
          2884 => x"3d0d7779",
          2885 => x"70720783",
          2886 => x"06535452",
          2887 => x"70933871",
          2888 => x"73730854",
          2889 => x"56547173",
          2890 => x"082e80c6",
          2891 => x"38737554",
          2892 => x"52713370",
          2893 => x"81ff0652",
          2894 => x"5470802e",
          2895 => x"9d387233",
          2896 => x"5570752e",
          2897 => x"09810695",
          2898 => x"38811281",
          2899 => x"14713370",
          2900 => x"81ff0654",
          2901 => x"56545270",
          2902 => x"e5387233",
          2903 => x"557381ff",
          2904 => x"067581ff",
          2905 => x"06717131",
          2906 => x"81dec00c",
          2907 => x"5252873d",
          2908 => x"0d047109",
          2909 => x"70f7fbfd",
          2910 => x"ff140670",
          2911 => x"f8848281",
          2912 => x"80065151",
          2913 => x"51709738",
          2914 => x"84148416",
          2915 => x"71085456",
          2916 => x"54717508",
          2917 => x"2edc3873",
          2918 => x"755452ff",
          2919 => x"9439800b",
          2920 => x"81dec00c",
          2921 => x"873d0d04",
          2922 => x"fe3d0d80",
          2923 => x"52835371",
          2924 => x"882b5287",
          2925 => x"863f81de",
          2926 => x"c00881ff",
          2927 => x"067207ff",
          2928 => x"14545272",
          2929 => x"8025e838",
          2930 => x"7181dec0",
          2931 => x"0c843d0d",
          2932 => x"04fb3d0d",
          2933 => x"77700870",
          2934 => x"53535671",
          2935 => x"802e80ca",
          2936 => x"38713351",
          2937 => x"70a02e09",
          2938 => x"81068638",
          2939 => x"811252f1",
          2940 => x"39715384",
          2941 => x"39811353",
          2942 => x"80733370",
          2943 => x"81ff0653",
          2944 => x"555570a0",
          2945 => x"2e833881",
          2946 => x"5570802e",
          2947 => x"843874e5",
          2948 => x"387381ff",
          2949 => x"065170a0",
          2950 => x"2e098106",
          2951 => x"88388073",
          2952 => x"70810555",
          2953 => x"3472760c",
          2954 => x"71517081",
          2955 => x"dec00c87",
          2956 => x"3d0d04fc",
          2957 => x"3d0d7653",
          2958 => x"7208802e",
          2959 => x"9138863d",
          2960 => x"fc055272",
          2961 => x"519bc33f",
          2962 => x"81dec008",
          2963 => x"85388053",
          2964 => x"83397453",
          2965 => x"7281dec0",
          2966 => x"0c863d0d",
          2967 => x"04fc3d0d",
          2968 => x"76821133",
          2969 => x"ff055253",
          2970 => x"8152708b",
          2971 => x"26819838",
          2972 => x"831333ff",
          2973 => x"05518252",
          2974 => x"709e2681",
          2975 => x"8a388413",
          2976 => x"33518352",
          2977 => x"70972680",
          2978 => x"fe388513",
          2979 => x"33518452",
          2980 => x"70bb2680",
          2981 => x"f2388613",
          2982 => x"33518552",
          2983 => x"70bb2680",
          2984 => x"e6388813",
          2985 => x"22558652",
          2986 => x"7487e726",
          2987 => x"80d9388a",
          2988 => x"13225487",
          2989 => x"527387e7",
          2990 => x"2680cc38",
          2991 => x"810b87c0",
          2992 => x"989c0c72",
          2993 => x"2287c098",
          2994 => x"bc0c8213",
          2995 => x"3387c098",
          2996 => x"b80c8313",
          2997 => x"3387c098",
          2998 => x"b40c8413",
          2999 => x"3387c098",
          3000 => x"b00c8513",
          3001 => x"3387c098",
          3002 => x"ac0c8613",
          3003 => x"3387c098",
          3004 => x"a80c7487",
          3005 => x"c098a40c",
          3006 => x"7387c098",
          3007 => x"a00c800b",
          3008 => x"87c0989c",
          3009 => x"0c805271",
          3010 => x"81dec00c",
          3011 => x"863d0d04",
          3012 => x"f33d0d7f",
          3013 => x"5b87c098",
          3014 => x"9c5d817d",
          3015 => x"0c87c098",
          3016 => x"bc085e7d",
          3017 => x"7b2387c0",
          3018 => x"98b8085a",
          3019 => x"79821c34",
          3020 => x"87c098b4",
          3021 => x"085a7983",
          3022 => x"1c3487c0",
          3023 => x"98b0085a",
          3024 => x"79841c34",
          3025 => x"87c098ac",
          3026 => x"085a7985",
          3027 => x"1c3487c0",
          3028 => x"98a8085a",
          3029 => x"79861c34",
          3030 => x"87c098a4",
          3031 => x"085c7b88",
          3032 => x"1c2387c0",
          3033 => x"98a0085a",
          3034 => x"798a1c23",
          3035 => x"807d0c79",
          3036 => x"83ffff06",
          3037 => x"597b83ff",
          3038 => x"ff065886",
          3039 => x"1b335785",
          3040 => x"1b335684",
          3041 => x"1b335583",
          3042 => x"1b335482",
          3043 => x"1b33537d",
          3044 => x"83ffff06",
          3045 => x"5281c6e4",
          3046 => x"5195883f",
          3047 => x"8f3d0d04",
          3048 => x"ff3d0d02",
          3049 => x"8f053370",
          3050 => x"30709f2a",
          3051 => x"51525270",
          3052 => x"0b0b81db",
          3053 => x"8834833d",
          3054 => x"0d04fb3d",
          3055 => x"0d770b0b",
          3056 => x"81db8833",
          3057 => x"7081ff06",
          3058 => x"57555687",
          3059 => x"c0948451",
          3060 => x"74802e86",
          3061 => x"3887c094",
          3062 => x"94517008",
          3063 => x"70962a70",
          3064 => x"81065354",
          3065 => x"5270802e",
          3066 => x"8c387191",
          3067 => x"2a708106",
          3068 => x"515170d7",
          3069 => x"38728132",
          3070 => x"70810651",
          3071 => x"5170802e",
          3072 => x"8d387193",
          3073 => x"2a708106",
          3074 => x"515170ff",
          3075 => x"be387381",
          3076 => x"ff065187",
          3077 => x"c0948052",
          3078 => x"70802e86",
          3079 => x"3887c094",
          3080 => x"90527572",
          3081 => x"0c7581de",
          3082 => x"c00c873d",
          3083 => x"0d04fb3d",
          3084 => x"0d029f05",
          3085 => x"330b0b81",
          3086 => x"db883370",
          3087 => x"81ff0657",
          3088 => x"555687c0",
          3089 => x"94845174",
          3090 => x"802e8638",
          3091 => x"87c09494",
          3092 => x"51700870",
          3093 => x"962a7081",
          3094 => x"06535452",
          3095 => x"70802e8c",
          3096 => x"3871912a",
          3097 => x"70810651",
          3098 => x"5170d738",
          3099 => x"72813270",
          3100 => x"81065151",
          3101 => x"70802e8d",
          3102 => x"3871932a",
          3103 => x"70810651",
          3104 => x"5170ffbe",
          3105 => x"387381ff",
          3106 => x"065187c0",
          3107 => x"94805270",
          3108 => x"802e8638",
          3109 => x"87c09490",
          3110 => x"5275720c",
          3111 => x"873d0d04",
          3112 => x"f93d0d79",
          3113 => x"54807433",
          3114 => x"7081ff06",
          3115 => x"53535770",
          3116 => x"772e80fe",
          3117 => x"387181ff",
          3118 => x"0681150b",
          3119 => x"0b81db88",
          3120 => x"337081ff",
          3121 => x"06595755",
          3122 => x"5887c094",
          3123 => x"84517580",
          3124 => x"2e863887",
          3125 => x"c0949451",
          3126 => x"70087096",
          3127 => x"2a708106",
          3128 => x"53545270",
          3129 => x"802e8c38",
          3130 => x"71912a70",
          3131 => x"81065151",
          3132 => x"70d73872",
          3133 => x"81327081",
          3134 => x"06515170",
          3135 => x"802e8d38",
          3136 => x"71932a70",
          3137 => x"81065151",
          3138 => x"70ffbe38",
          3139 => x"7481ff06",
          3140 => x"5187c094",
          3141 => x"80527080",
          3142 => x"2e863887",
          3143 => x"c0949052",
          3144 => x"77720c81",
          3145 => x"17743370",
          3146 => x"81ff0653",
          3147 => x"535770ff",
          3148 => x"84387681",
          3149 => x"dec00c89",
          3150 => x"3d0d04fe",
          3151 => x"3d0d0b0b",
          3152 => x"81db8833",
          3153 => x"7081ff06",
          3154 => x"545287c0",
          3155 => x"94845172",
          3156 => x"802e8638",
          3157 => x"87c09494",
          3158 => x"51700870",
          3159 => x"822a7081",
          3160 => x"06515151",
          3161 => x"70802ee2",
          3162 => x"387181ff",
          3163 => x"065187c0",
          3164 => x"94805270",
          3165 => x"802e8638",
          3166 => x"87c09490",
          3167 => x"52710870",
          3168 => x"81ff0681",
          3169 => x"dec00c51",
          3170 => x"843d0d04",
          3171 => x"fe3d0d0b",
          3172 => x"0b81db88",
          3173 => x"337081ff",
          3174 => x"06525387",
          3175 => x"c0948452",
          3176 => x"70802e86",
          3177 => x"3887c094",
          3178 => x"94527108",
          3179 => x"70822a70",
          3180 => x"81065151",
          3181 => x"51ff5270",
          3182 => x"802ea038",
          3183 => x"7281ff06",
          3184 => x"5187c094",
          3185 => x"80527080",
          3186 => x"2e863887",
          3187 => x"c0949052",
          3188 => x"71087098",
          3189 => x"2b70982c",
          3190 => x"51535171",
          3191 => x"81dec00c",
          3192 => x"843d0d04",
          3193 => x"ff3d0d87",
          3194 => x"c09e8008",
          3195 => x"709c2a8a",
          3196 => x"06515170",
          3197 => x"802e84b4",
          3198 => x"3887c09e",
          3199 => x"a40881db",
          3200 => x"8c0c87c0",
          3201 => x"9ea80881",
          3202 => x"db900c87",
          3203 => x"c09e9408",
          3204 => x"81db940c",
          3205 => x"87c09e98",
          3206 => x"0881db98",
          3207 => x"0c87c09e",
          3208 => x"9c0881db",
          3209 => x"9c0c87c0",
          3210 => x"9ea00881",
          3211 => x"dba00c87",
          3212 => x"c09eac08",
          3213 => x"81dba40c",
          3214 => x"87c09eb0",
          3215 => x"0881dba8",
          3216 => x"0c87c09e",
          3217 => x"b40881db",
          3218 => x"ac0c87c0",
          3219 => x"9eb80881",
          3220 => x"dbb00c87",
          3221 => x"c09ebc08",
          3222 => x"81dbb40c",
          3223 => x"87c09ec0",
          3224 => x"0881dbb8",
          3225 => x"0c87c09e",
          3226 => x"c40881db",
          3227 => x"bc0c87c0",
          3228 => x"9e800851",
          3229 => x"7081dbc0",
          3230 => x"2387c09e",
          3231 => x"840881db",
          3232 => x"c40c87c0",
          3233 => x"9e880881",
          3234 => x"dbc80c87",
          3235 => x"c09e8c08",
          3236 => x"81dbcc0c",
          3237 => x"810b81db",
          3238 => x"d034800b",
          3239 => x"87c09e90",
          3240 => x"08708480",
          3241 => x"0a065152",
          3242 => x"5270802e",
          3243 => x"83388152",
          3244 => x"7181dbd1",
          3245 => x"34800b87",
          3246 => x"c09e9008",
          3247 => x"7088800a",
          3248 => x"06515252",
          3249 => x"70802e83",
          3250 => x"38815271",
          3251 => x"81dbd234",
          3252 => x"800b87c0",
          3253 => x"9e900870",
          3254 => x"90800a06",
          3255 => x"51525270",
          3256 => x"802e8338",
          3257 => x"81527181",
          3258 => x"dbd33480",
          3259 => x"0b87c09e",
          3260 => x"90087088",
          3261 => x"80800651",
          3262 => x"52527080",
          3263 => x"2e833881",
          3264 => x"527181db",
          3265 => x"d434800b",
          3266 => x"87c09e90",
          3267 => x"0870a080",
          3268 => x"80065152",
          3269 => x"5270802e",
          3270 => x"83388152",
          3271 => x"7181dbd5",
          3272 => x"34800b87",
          3273 => x"c09e9008",
          3274 => x"70908080",
          3275 => x"06515252",
          3276 => x"70802e83",
          3277 => x"38815271",
          3278 => x"81dbd634",
          3279 => x"800b87c0",
          3280 => x"9e900870",
          3281 => x"84808006",
          3282 => x"51525270",
          3283 => x"802e8338",
          3284 => x"81527181",
          3285 => x"dbd73480",
          3286 => x"0b87c09e",
          3287 => x"90087082",
          3288 => x"80800651",
          3289 => x"52527080",
          3290 => x"2e833881",
          3291 => x"527181db",
          3292 => x"d834800b",
          3293 => x"87c09e90",
          3294 => x"08708180",
          3295 => x"80065152",
          3296 => x"5270802e",
          3297 => x"83388152",
          3298 => x"7181dbd9",
          3299 => x"34800b87",
          3300 => x"c09e9008",
          3301 => x"7080c080",
          3302 => x"06515252",
          3303 => x"70802e83",
          3304 => x"38815271",
          3305 => x"81dbda34",
          3306 => x"800b87c0",
          3307 => x"9e900870",
          3308 => x"a0800651",
          3309 => x"52527080",
          3310 => x"2e833881",
          3311 => x"527181db",
          3312 => x"db3487c0",
          3313 => x"9e900870",
          3314 => x"98800670",
          3315 => x"8a2a5151",
          3316 => x"517081db",
          3317 => x"dc34800b",
          3318 => x"87c09e90",
          3319 => x"08708480",
          3320 => x"06515252",
          3321 => x"70802e83",
          3322 => x"38815271",
          3323 => x"81dbdd34",
          3324 => x"87c09e90",
          3325 => x"087083f0",
          3326 => x"0670842a",
          3327 => x"51515170",
          3328 => x"81dbde34",
          3329 => x"800b87c0",
          3330 => x"9e900870",
          3331 => x"88065152",
          3332 => x"5270802e",
          3333 => x"83388152",
          3334 => x"7181dbdf",
          3335 => x"3487c09e",
          3336 => x"90087087",
          3337 => x"06515170",
          3338 => x"81dbe034",
          3339 => x"833d0d04",
          3340 => x"fb3d0d81",
          3341 => x"c6fc5186",
          3342 => x"863f81db",
          3343 => x"d0335473",
          3344 => x"802e8838",
          3345 => x"81c79051",
          3346 => x"85f53f81",
          3347 => x"c7a45185",
          3348 => x"ee3f81db",
          3349 => x"d2335473",
          3350 => x"802e9338",
          3351 => x"81dbac08",
          3352 => x"81dbb008",
          3353 => x"11545281",
          3354 => x"c7bc518b",
          3355 => x"b63f81db",
          3356 => x"d7335473",
          3357 => x"802e9338",
          3358 => x"81dba408",
          3359 => x"81dba808",
          3360 => x"11545281",
          3361 => x"c7d8518b",
          3362 => x"9a3f81db",
          3363 => x"d4335473",
          3364 => x"802e9338",
          3365 => x"81db8c08",
          3366 => x"81db9008",
          3367 => x"11545281",
          3368 => x"c7f4518a",
          3369 => x"fe3f81db",
          3370 => x"d5335473",
          3371 => x"802e9338",
          3372 => x"81db9408",
          3373 => x"81db9808",
          3374 => x"11545281",
          3375 => x"c890518a",
          3376 => x"e23f81db",
          3377 => x"d6335473",
          3378 => x"802e9338",
          3379 => x"81db9c08",
          3380 => x"81dba008",
          3381 => x"11545281",
          3382 => x"c8ac518a",
          3383 => x"c63f81db",
          3384 => x"db335473",
          3385 => x"802e8d38",
          3386 => x"81dbdc33",
          3387 => x"5281c8c8",
          3388 => x"518ab03f",
          3389 => x"81dbdf33",
          3390 => x"5473802e",
          3391 => x"8d3881db",
          3392 => x"e0335281",
          3393 => x"c8e8518a",
          3394 => x"9a3f81db",
          3395 => x"dd335473",
          3396 => x"802e8d38",
          3397 => x"81dbde33",
          3398 => x"5281c988",
          3399 => x"518a843f",
          3400 => x"81dbd133",
          3401 => x"5473802e",
          3402 => x"883881c9",
          3403 => x"a851848f",
          3404 => x"3f81dbd3",
          3405 => x"33547380",
          3406 => x"2e883881",
          3407 => x"c9bc5183",
          3408 => x"fe3f81db",
          3409 => x"d8335473",
          3410 => x"802e8838",
          3411 => x"81c9c851",
          3412 => x"83ed3f81",
          3413 => x"dbd93354",
          3414 => x"73802e88",
          3415 => x"3881c9d4",
          3416 => x"5183dc3f",
          3417 => x"81dbda33",
          3418 => x"5473802e",
          3419 => x"883881c9",
          3420 => x"e05183cb",
          3421 => x"3f81c9ec",
          3422 => x"5183c43f",
          3423 => x"81dbb408",
          3424 => x"5281c9f8",
          3425 => x"51899c3f",
          3426 => x"81dbb808",
          3427 => x"5281caa0",
          3428 => x"5189903f",
          3429 => x"81dbbc08",
          3430 => x"5281cac8",
          3431 => x"5189843f",
          3432 => x"81caf051",
          3433 => x"f5fa3f81",
          3434 => x"dbc02252",
          3435 => x"81caf851",
          3436 => x"88f13f81",
          3437 => x"dbc40856",
          3438 => x"bd84c052",
          3439 => x"7551e7b7",
          3440 => x"3f81dec0",
          3441 => x"08bd84c0",
          3442 => x"29767131",
          3443 => x"545481de",
          3444 => x"c0085281",
          3445 => x"cba05188",
          3446 => x"ca3f81db",
          3447 => x"d7335473",
          3448 => x"802ea838",
          3449 => x"81dbc808",
          3450 => x"56bd84c0",
          3451 => x"527551e7",
          3452 => x"863f81de",
          3453 => x"c008bd84",
          3454 => x"c0297671",
          3455 => x"31545481",
          3456 => x"dec00852",
          3457 => x"81cbcc51",
          3458 => x"88993f81",
          3459 => x"dbd23354",
          3460 => x"73802ea8",
          3461 => x"3881dbcc",
          3462 => x"0856bd84",
          3463 => x"c0527551",
          3464 => x"e6d53f81",
          3465 => x"dec008bd",
          3466 => x"84c02976",
          3467 => x"71315454",
          3468 => x"81dec008",
          3469 => x"5281cbf8",
          3470 => x"5187e83f",
          3471 => x"81d79c51",
          3472 => x"81fd3f87",
          3473 => x"3d0d04fe",
          3474 => x"3d0d0292",
          3475 => x"0533ff05",
          3476 => x"52718426",
          3477 => x"aa387184",
          3478 => x"2981c680",
          3479 => x"05527108",
          3480 => x"0481cca4",
          3481 => x"519d3981",
          3482 => x"ccac5197",
          3483 => x"3981ccb4",
          3484 => x"51913981",
          3485 => x"ccbc518b",
          3486 => x"3981ccc0",
          3487 => x"51853981",
          3488 => x"ccc851f4",
          3489 => x"9b3f843d",
          3490 => x"0d047188",
          3491 => x"800c0480",
          3492 => x"0b87c096",
          3493 => x"840c04ff",
          3494 => x"3d0d87c0",
          3495 => x"96847008",
          3496 => x"52528072",
          3497 => x"0c707407",
          3498 => x"7081dbe4",
          3499 => x"0c720c83",
          3500 => x"3d0d04ff",
          3501 => x"3d0d87c0",
          3502 => x"96847008",
          3503 => x"81dbe40c",
          3504 => x"5280720c",
          3505 => x"73097081",
          3506 => x"dbe40806",
          3507 => x"7081dbe4",
          3508 => x"0c730c51",
          3509 => x"833d0d04",
          3510 => x"81dbe408",
          3511 => x"87c09684",
          3512 => x"0c04fe3d",
          3513 => x"0d029305",
          3514 => x"3353728a",
          3515 => x"2e098106",
          3516 => x"85388d51",
          3517 => x"ed3f81de",
          3518 => x"d8085271",
          3519 => x"802e9038",
          3520 => x"72723481",
          3521 => x"ded80881",
          3522 => x"0581ded8",
          3523 => x"0c8f3981",
          3524 => x"ded00852",
          3525 => x"71802e85",
          3526 => x"38725171",
          3527 => x"2d843d0d",
          3528 => x"04fe3d0d",
          3529 => x"02970533",
          3530 => x"81ded008",
          3531 => x"7681ded0",
          3532 => x"0c5451ff",
          3533 => x"ad3f7281",
          3534 => x"ded00c84",
          3535 => x"3d0d04fd",
          3536 => x"3d0d7554",
          3537 => x"73337081",
          3538 => x"ff065353",
          3539 => x"71802e8e",
          3540 => x"387281ff",
          3541 => x"06518114",
          3542 => x"54ff873f",
          3543 => x"e739853d",
          3544 => x"0d04fc3d",
          3545 => x"0d7781de",
          3546 => x"d0087881",
          3547 => x"ded00c56",
          3548 => x"54733370",
          3549 => x"81ff0653",
          3550 => x"5371802e",
          3551 => x"8e387281",
          3552 => x"ff065181",
          3553 => x"1454feda",
          3554 => x"3fe73974",
          3555 => x"81ded00c",
          3556 => x"863d0d04",
          3557 => x"ec3d0d66",
          3558 => x"68595978",
          3559 => x"7081055a",
          3560 => x"33567580",
          3561 => x"2e84f838",
          3562 => x"75a52e09",
          3563 => x"810682de",
          3564 => x"3880707a",
          3565 => x"7081055c",
          3566 => x"33585b5b",
          3567 => x"75b02e09",
          3568 => x"81068538",
          3569 => x"815a8b39",
          3570 => x"75ad2e09",
          3571 => x"81068a38",
          3572 => x"825a7870",
          3573 => x"81055a33",
          3574 => x"5675aa2e",
          3575 => x"09810692",
          3576 => x"38778419",
          3577 => x"71087b70",
          3578 => x"81055d33",
          3579 => x"595d5953",
          3580 => x"9d39d016",
          3581 => x"53728926",
          3582 => x"95387a88",
          3583 => x"297b1005",
          3584 => x"7605d005",
          3585 => x"79708105",
          3586 => x"5b33575b",
          3587 => x"e5397580",
          3588 => x"ec327030",
          3589 => x"70720780",
          3590 => x"257880cc",
          3591 => x"32703070",
          3592 => x"72078025",
          3593 => x"73075354",
          3594 => x"58515553",
          3595 => x"73802e8c",
          3596 => x"38798407",
          3597 => x"79708105",
          3598 => x"5b33575a",
          3599 => x"75802e83",
          3600 => x"de387554",
          3601 => x"80e07627",
          3602 => x"8938e016",
          3603 => x"7081ff06",
          3604 => x"55537380",
          3605 => x"cf2e81aa",
          3606 => x"387380cf",
          3607 => x"24a23873",
          3608 => x"80c32e81",
          3609 => x"8e387380",
          3610 => x"c3248b38",
          3611 => x"7380c22e",
          3612 => x"818c3881",
          3613 => x"99397380",
          3614 => x"c42e818a",
          3615 => x"38818f39",
          3616 => x"7380d52e",
          3617 => x"81803873",
          3618 => x"80d5248a",
          3619 => x"387380d3",
          3620 => x"2e8e3880",
          3621 => x"f9397380",
          3622 => x"d82e80ee",
          3623 => x"3880ef39",
          3624 => x"77841971",
          3625 => x"08565953",
          3626 => x"80743354",
          3627 => x"5572752e",
          3628 => x"8d388115",
          3629 => x"70157033",
          3630 => x"51545572",
          3631 => x"f5387981",
          3632 => x"2a569039",
          3633 => x"74811656",
          3634 => x"53727b27",
          3635 => x"8f38a051",
          3636 => x"fc903f75",
          3637 => x"81065372",
          3638 => x"802ee938",
          3639 => x"7351fcdf",
          3640 => x"3f748116",
          3641 => x"5653727b",
          3642 => x"27fdb038",
          3643 => x"a051fbf2",
          3644 => x"3fef3977",
          3645 => x"84198312",
          3646 => x"33535953",
          3647 => x"9339825c",
          3648 => x"9539885c",
          3649 => x"91398a5c",
          3650 => x"8d39905c",
          3651 => x"89397551",
          3652 => x"fbd03ffd",
          3653 => x"86397982",
          3654 => x"2a708106",
          3655 => x"51537280",
          3656 => x"2e883877",
          3657 => x"84195953",
          3658 => x"86398418",
          3659 => x"78545872",
          3660 => x"087480c4",
          3661 => x"32703070",
          3662 => x"72078025",
          3663 => x"51555555",
          3664 => x"7480258d",
          3665 => x"3872802e",
          3666 => x"88387430",
          3667 => x"7a90075b",
          3668 => x"55800b8f",
          3669 => x"3d5e577b",
          3670 => x"527451e0",
          3671 => x"cd3f81de",
          3672 => x"c00881ff",
          3673 => x"067c5375",
          3674 => x"5254e08b",
          3675 => x"3f81dec0",
          3676 => x"08558974",
          3677 => x"279238a7",
          3678 => x"14537580",
          3679 => x"f82e8438",
          3680 => x"87145372",
          3681 => x"81ff0654",
          3682 => x"b0145372",
          3683 => x"7d708105",
          3684 => x"5f348117",
          3685 => x"75307077",
          3686 => x"079f2a51",
          3687 => x"5457769f",
          3688 => x"26853872",
          3689 => x"ffb13879",
          3690 => x"842a7081",
          3691 => x"06515372",
          3692 => x"802e8e38",
          3693 => x"963d7705",
          3694 => x"e00553ad",
          3695 => x"73348117",
          3696 => x"57767a81",
          3697 => x"065455b0",
          3698 => x"54728338",
          3699 => x"a0547981",
          3700 => x"2a708106",
          3701 => x"5456729f",
          3702 => x"38811755",
          3703 => x"767b2797",
          3704 => x"387351f9",
          3705 => x"fd3f7581",
          3706 => x"0653728b",
          3707 => x"38748116",
          3708 => x"56537a73",
          3709 => x"26eb3896",
          3710 => x"3d7705e0",
          3711 => x"0553ff17",
          3712 => x"ff147033",
          3713 => x"535457f9",
          3714 => x"d93f76f2",
          3715 => x"38748116",
          3716 => x"5653727b",
          3717 => x"27fb8438",
          3718 => x"a051f9c6",
          3719 => x"3fef3996",
          3720 => x"3d0d04fd",
          3721 => x"3d0d863d",
          3722 => x"70708405",
          3723 => x"52085552",
          3724 => x"7351fae0",
          3725 => x"3f853d0d",
          3726 => x"04fe3d0d",
          3727 => x"7481ded8",
          3728 => x"0c853d88",
          3729 => x"05527551",
          3730 => x"faca3f81",
          3731 => x"ded80853",
          3732 => x"80733480",
          3733 => x"0b81ded8",
          3734 => x"0c843d0d",
          3735 => x"04fd3d0d",
          3736 => x"81ded008",
          3737 => x"7681ded0",
          3738 => x"0c873d88",
          3739 => x"05537752",
          3740 => x"53faa13f",
          3741 => x"7281ded0",
          3742 => x"0c853d0d",
          3743 => x"04fb3d0d",
          3744 => x"777981de",
          3745 => x"d4087056",
          3746 => x"54575580",
          3747 => x"5471802e",
          3748 => x"80e03881",
          3749 => x"ded40852",
          3750 => x"712d81de",
          3751 => x"c00881ff",
          3752 => x"06537280",
          3753 => x"2e80cb38",
          3754 => x"728d2eb9",
          3755 => x"38728832",
          3756 => x"70307080",
          3757 => x"25515152",
          3758 => x"73802e8b",
          3759 => x"3871802e",
          3760 => x"8638ff14",
          3761 => x"5497399f",
          3762 => x"7325c838",
          3763 => x"ff165273",
          3764 => x"7225c038",
          3765 => x"74145272",
          3766 => x"72348114",
          3767 => x"547251f8",
          3768 => x"813fffaf",
          3769 => x"39731552",
          3770 => x"8072348a",
          3771 => x"51f7f33f",
          3772 => x"81537281",
          3773 => x"dec00c87",
          3774 => x"3d0d04fe",
          3775 => x"3d0d81de",
          3776 => x"d4087581",
          3777 => x"ded40c77",
          3778 => x"53765253",
          3779 => x"feef3f72",
          3780 => x"81ded40c",
          3781 => x"843d0d04",
          3782 => x"f83d0d7a",
          3783 => x"7c5a5680",
          3784 => x"707a0c58",
          3785 => x"75087033",
          3786 => x"555373a0",
          3787 => x"2e098106",
          3788 => x"87388113",
          3789 => x"760ced39",
          3790 => x"73ad2e09",
          3791 => x"81068e38",
          3792 => x"81760811",
          3793 => x"770c7608",
          3794 => x"70335654",
          3795 => x"5873b02e",
          3796 => x"09810680",
          3797 => x"c2387508",
          3798 => x"8105760c",
          3799 => x"75087033",
          3800 => x"55537380",
          3801 => x"e22e8b38",
          3802 => x"90577380",
          3803 => x"f82e8538",
          3804 => x"8f398257",
          3805 => x"8113760c",
          3806 => x"75087033",
          3807 => x"5553ac39",
          3808 => x"8155a074",
          3809 => x"2780fa38",
          3810 => x"d0145380",
          3811 => x"55885789",
          3812 => x"73279838",
          3813 => x"80eb39d0",
          3814 => x"14538055",
          3815 => x"72892680",
          3816 => x"e0388639",
          3817 => x"805580d9",
          3818 => x"398a5780",
          3819 => x"55a07427",
          3820 => x"80c23880",
          3821 => x"e0742789",
          3822 => x"38e01470",
          3823 => x"81ff0655",
          3824 => x"53d01470",
          3825 => x"81ff0655",
          3826 => x"53907427",
          3827 => x"8e38f914",
          3828 => x"7081ff06",
          3829 => x"55538974",
          3830 => x"27ca3873",
          3831 => x"7727c538",
          3832 => x"74772914",
          3833 => x"76088105",
          3834 => x"770c7608",
          3835 => x"70335654",
          3836 => x"55ffba39",
          3837 => x"77802e84",
          3838 => x"38743055",
          3839 => x"74790c81",
          3840 => x"557481de",
          3841 => x"c00c8a3d",
          3842 => x"0d04f83d",
          3843 => x"0d7a7c5a",
          3844 => x"5680707a",
          3845 => x"0c587508",
          3846 => x"70335553",
          3847 => x"73a02e09",
          3848 => x"81068738",
          3849 => x"8113760c",
          3850 => x"ed3973ad",
          3851 => x"2e098106",
          3852 => x"8e388176",
          3853 => x"0811770c",
          3854 => x"76087033",
          3855 => x"56545873",
          3856 => x"b02e0981",
          3857 => x"0680c238",
          3858 => x"75088105",
          3859 => x"760c7508",
          3860 => x"70335553",
          3861 => x"7380e22e",
          3862 => x"8b389057",
          3863 => x"7380f82e",
          3864 => x"85388f39",
          3865 => x"82578113",
          3866 => x"760c7508",
          3867 => x"70335553",
          3868 => x"ac398155",
          3869 => x"a0742780",
          3870 => x"fa38d014",
          3871 => x"53805588",
          3872 => x"57897327",
          3873 => x"983880eb",
          3874 => x"39d01453",
          3875 => x"80557289",
          3876 => x"2680e038",
          3877 => x"86398055",
          3878 => x"80d9398a",
          3879 => x"578055a0",
          3880 => x"742780c2",
          3881 => x"3880e074",
          3882 => x"278938e0",
          3883 => x"147081ff",
          3884 => x"065553d0",
          3885 => x"147081ff",
          3886 => x"06555390",
          3887 => x"74278e38",
          3888 => x"f9147081",
          3889 => x"ff065553",
          3890 => x"897427ca",
          3891 => x"38737727",
          3892 => x"c5387477",
          3893 => x"29147608",
          3894 => x"8105770c",
          3895 => x"76087033",
          3896 => x"565455ff",
          3897 => x"ba397780",
          3898 => x"2e843874",
          3899 => x"30557479",
          3900 => x"0c815574",
          3901 => x"81dec00c",
          3902 => x"8a3d0d04",
          3903 => x"ff3d0d02",
          3904 => x"8f053351",
          3905 => x"81527072",
          3906 => x"26873881",
          3907 => x"dbe81133",
          3908 => x"527181de",
          3909 => x"c00c833d",
          3910 => x"0d04fc3d",
          3911 => x"0d029b05",
          3912 => x"33028405",
          3913 => x"9f053356",
          3914 => x"53835172",
          3915 => x"812680e0",
          3916 => x"3872842b",
          3917 => x"87c0928c",
          3918 => x"11535188",
          3919 => x"5474802e",
          3920 => x"84388188",
          3921 => x"5473720c",
          3922 => x"87c0928c",
          3923 => x"11518171",
          3924 => x"0c850b87",
          3925 => x"c0988c0c",
          3926 => x"70527108",
          3927 => x"70820651",
          3928 => x"5170802e",
          3929 => x"8a3887c0",
          3930 => x"988c0851",
          3931 => x"70ec3871",
          3932 => x"08fc8080",
          3933 => x"06527192",
          3934 => x"3887c098",
          3935 => x"8c085170",
          3936 => x"802e8738",
          3937 => x"7181dbe8",
          3938 => x"143481db",
          3939 => x"e8133351",
          3940 => x"7081dec0",
          3941 => x"0c863d0d",
          3942 => x"04f33d0d",
          3943 => x"60626402",
          3944 => x"8c05bf05",
          3945 => x"33574058",
          3946 => x"5b837452",
          3947 => x"5afecd3f",
          3948 => x"81dec008",
          3949 => x"81067a54",
          3950 => x"527181be",
          3951 => x"38717275",
          3952 => x"842b87c0",
          3953 => x"92801187",
          3954 => x"c0928c12",
          3955 => x"87c09284",
          3956 => x"13415a40",
          3957 => x"575a5885",
          3958 => x"0b87c098",
          3959 => x"8c0c767d",
          3960 => x"0c84760c",
          3961 => x"75087085",
          3962 => x"2a708106",
          3963 => x"51535471",
          3964 => x"802e8e38",
          3965 => x"7b085271",
          3966 => x"7b708105",
          3967 => x"5d348119",
          3968 => x"598074a2",
          3969 => x"06535371",
          3970 => x"732e8338",
          3971 => x"81537883",
          3972 => x"ff268f38",
          3973 => x"72802e8a",
          3974 => x"3887c098",
          3975 => x"8c085271",
          3976 => x"c33887c0",
          3977 => x"988c0852",
          3978 => x"71802e87",
          3979 => x"38788480",
          3980 => x"2e993881",
          3981 => x"760c87c0",
          3982 => x"928c1553",
          3983 => x"72087082",
          3984 => x"06515271",
          3985 => x"f738ff1a",
          3986 => x"5a8d3984",
          3987 => x"80178119",
          3988 => x"7081ff06",
          3989 => x"5a535779",
          3990 => x"802e9038",
          3991 => x"73fc8080",
          3992 => x"06527187",
          3993 => x"387d7826",
          3994 => x"feed3873",
          3995 => x"fc808006",
          3996 => x"5271802e",
          3997 => x"83388152",
          3998 => x"71537281",
          3999 => x"dec00c8f",
          4000 => x"3d0d04f3",
          4001 => x"3d0d6062",
          4002 => x"64028c05",
          4003 => x"bf053357",
          4004 => x"40585b83",
          4005 => x"59807452",
          4006 => x"58fce13f",
          4007 => x"81dec008",
          4008 => x"81067954",
          4009 => x"5271782e",
          4010 => x"09810681",
          4011 => x"b1387774",
          4012 => x"842b87c0",
          4013 => x"92801187",
          4014 => x"c0928c12",
          4015 => x"87c09284",
          4016 => x"1340595f",
          4017 => x"565a850b",
          4018 => x"87c0988c",
          4019 => x"0c767d0c",
          4020 => x"82760c80",
          4021 => x"58750870",
          4022 => x"842a7081",
          4023 => x"06515354",
          4024 => x"71802e8c",
          4025 => x"387a7081",
          4026 => x"055c337c",
          4027 => x"0c811858",
          4028 => x"73812a70",
          4029 => x"81065152",
          4030 => x"71802e8a",
          4031 => x"3887c098",
          4032 => x"8c085271",
          4033 => x"d03887c0",
          4034 => x"988c0852",
          4035 => x"71802e87",
          4036 => x"38778480",
          4037 => x"2e993881",
          4038 => x"760c87c0",
          4039 => x"928c1553",
          4040 => x"72087082",
          4041 => x"06515271",
          4042 => x"f738ff19",
          4043 => x"598d3981",
          4044 => x"1a7081ff",
          4045 => x"06848019",
          4046 => x"595b5278",
          4047 => x"802e9038",
          4048 => x"73fc8080",
          4049 => x"06527187",
          4050 => x"387d7a26",
          4051 => x"fef83873",
          4052 => x"fc808006",
          4053 => x"5271802e",
          4054 => x"83388152",
          4055 => x"71537281",
          4056 => x"dec00c8f",
          4057 => x"3d0d04f6",
          4058 => x"3d0d7e02",
          4059 => x"8405b305",
          4060 => x"33028805",
          4061 => x"b7053371",
          4062 => x"54545657",
          4063 => x"fafe3f81",
          4064 => x"dec00881",
          4065 => x"06538354",
          4066 => x"7280fe38",
          4067 => x"850b87c0",
          4068 => x"988c0c81",
          4069 => x"5671762e",
          4070 => x"80dc3871",
          4071 => x"76249338",
          4072 => x"74842b87",
          4073 => x"c0928c11",
          4074 => x"54547180",
          4075 => x"2e8d3880",
          4076 => x"d4397183",
          4077 => x"2e80c638",
          4078 => x"80cb3972",
          4079 => x"0870812a",
          4080 => x"70810651",
          4081 => x"51527180",
          4082 => x"2e8a3887",
          4083 => x"c0988c08",
          4084 => x"5271e838",
          4085 => x"87c0988c",
          4086 => x"08527196",
          4087 => x"3881730c",
          4088 => x"87c0928c",
          4089 => x"14537208",
          4090 => x"70820651",
          4091 => x"5271f738",
          4092 => x"96398056",
          4093 => x"92398880",
          4094 => x"0a770c85",
          4095 => x"39818077",
          4096 => x"0c725683",
          4097 => x"39845675",
          4098 => x"547381de",
          4099 => x"c00c8c3d",
          4100 => x"0d04fe3d",
          4101 => x"0d748111",
          4102 => x"33713371",
          4103 => x"882b0781",
          4104 => x"dec00c53",
          4105 => x"51843d0d",
          4106 => x"04fd3d0d",
          4107 => x"75831133",
          4108 => x"82123371",
          4109 => x"902b7188",
          4110 => x"2b078114",
          4111 => x"33707207",
          4112 => x"882b7533",
          4113 => x"710781de",
          4114 => x"c00c5253",
          4115 => x"54565452",
          4116 => x"853d0d04",
          4117 => x"ff3d0d73",
          4118 => x"02840592",
          4119 => x"05225252",
          4120 => x"70727081",
          4121 => x"05543470",
          4122 => x"882a5170",
          4123 => x"7234833d",
          4124 => x"0d04ff3d",
          4125 => x"0d737552",
          4126 => x"52707270",
          4127 => x"81055434",
          4128 => x"70882a51",
          4129 => x"70727081",
          4130 => x"05543470",
          4131 => x"882a5170",
          4132 => x"72708105",
          4133 => x"54347088",
          4134 => x"2a517072",
          4135 => x"34833d0d",
          4136 => x"04fe3d0d",
          4137 => x"76757754",
          4138 => x"54517080",
          4139 => x"2e923871",
          4140 => x"70810553",
          4141 => x"33737081",
          4142 => x"055534ff",
          4143 => x"1151eb39",
          4144 => x"843d0d04",
          4145 => x"fe3d0d75",
          4146 => x"77765452",
          4147 => x"53727270",
          4148 => x"81055434",
          4149 => x"ff115170",
          4150 => x"f438843d",
          4151 => x"0d04fc3d",
          4152 => x"0d787779",
          4153 => x"56565374",
          4154 => x"70810556",
          4155 => x"33747081",
          4156 => x"05563371",
          4157 => x"7131ff16",
          4158 => x"56525252",
          4159 => x"72802e86",
          4160 => x"3871802e",
          4161 => x"e2387181",
          4162 => x"dec00c86",
          4163 => x"3d0d04fe",
          4164 => x"3d0d7476",
          4165 => x"54518939",
          4166 => x"71732e8a",
          4167 => x"38811151",
          4168 => x"70335271",
          4169 => x"f3387033",
          4170 => x"81dec00c",
          4171 => x"843d0d04",
          4172 => x"800b81de",
          4173 => x"c00c0480",
          4174 => x"0b81dec0",
          4175 => x"0c04f73d",
          4176 => x"0d7b5680",
          4177 => x"0b831733",
          4178 => x"565a747a",
          4179 => x"2e80d638",
          4180 => x"8154b016",
          4181 => x"0853b416",
          4182 => x"70538117",
          4183 => x"335259fa",
          4184 => x"a23f81de",
          4185 => x"c0087a2e",
          4186 => x"098106b7",
          4187 => x"3881dec0",
          4188 => x"08831734",
          4189 => x"b0160870",
          4190 => x"a4180831",
          4191 => x"9c180859",
          4192 => x"56587477",
          4193 => x"279f3882",
          4194 => x"16335574",
          4195 => x"822e0981",
          4196 => x"06933881",
          4197 => x"54761853",
          4198 => x"78528116",
          4199 => x"3351f9e3",
          4200 => x"3f833981",
          4201 => x"5a7981de",
          4202 => x"c00c8b3d",
          4203 => x"0d04fa3d",
          4204 => x"0d787a56",
          4205 => x"56805774",
          4206 => x"b017082e",
          4207 => x"af387551",
          4208 => x"fefc3f81",
          4209 => x"dec00857",
          4210 => x"81dec008",
          4211 => x"9f388154",
          4212 => x"7453b416",
          4213 => x"52811633",
          4214 => x"51f7be3f",
          4215 => x"81dec008",
          4216 => x"802e8538",
          4217 => x"ff558157",
          4218 => x"74b0170c",
          4219 => x"7681dec0",
          4220 => x"0c883d0d",
          4221 => x"04f83d0d",
          4222 => x"7a705257",
          4223 => x"fec03f81",
          4224 => x"dec00858",
          4225 => x"81dec008",
          4226 => x"81913876",
          4227 => x"33557483",
          4228 => x"2e098106",
          4229 => x"80f03884",
          4230 => x"17335978",
          4231 => x"812e0981",
          4232 => x"0680e338",
          4233 => x"84805381",
          4234 => x"dec00852",
          4235 => x"b4177052",
          4236 => x"56fd913f",
          4237 => x"82d4d552",
          4238 => x"84b21751",
          4239 => x"fc963f84",
          4240 => x"8b85a4d2",
          4241 => x"527551fc",
          4242 => x"a93f868a",
          4243 => x"85e4f252",
          4244 => x"84981751",
          4245 => x"fc9c3f90",
          4246 => x"17085284",
          4247 => x"9c1751fc",
          4248 => x"913f8c17",
          4249 => x"085284a0",
          4250 => x"1751fc86",
          4251 => x"3fa01708",
          4252 => x"810570b0",
          4253 => x"190c7955",
          4254 => x"53755281",
          4255 => x"173351f8",
          4256 => x"823f7784",
          4257 => x"18348053",
          4258 => x"80528117",
          4259 => x"3351f9d7",
          4260 => x"3f81dec0",
          4261 => x"08802e83",
          4262 => x"38815877",
          4263 => x"81dec00c",
          4264 => x"8a3d0d04",
          4265 => x"fb3d0d77",
          4266 => x"fe1a9812",
          4267 => x"08fe0555",
          4268 => x"56548056",
          4269 => x"7473278d",
          4270 => x"388a1422",
          4271 => x"757129ac",
          4272 => x"16080557",
          4273 => x"537581de",
          4274 => x"c00c873d",
          4275 => x"0d04f93d",
          4276 => x"0d7a7a70",
          4277 => x"08565457",
          4278 => x"81772781",
          4279 => x"df387698",
          4280 => x"15082781",
          4281 => x"d738ff74",
          4282 => x"33545872",
          4283 => x"822e80f5",
          4284 => x"38728224",
          4285 => x"89387281",
          4286 => x"2e8d3881",
          4287 => x"bf397283",
          4288 => x"2e818e38",
          4289 => x"81b63976",
          4290 => x"812a1770",
          4291 => x"892aa416",
          4292 => x"08055374",
          4293 => x"5255fd96",
          4294 => x"3f81dec0",
          4295 => x"08819f38",
          4296 => x"7483ff06",
          4297 => x"14b41133",
          4298 => x"81177089",
          4299 => x"2aa41808",
          4300 => x"05557654",
          4301 => x"575753fc",
          4302 => x"f53f81de",
          4303 => x"c00880fe",
          4304 => x"387483ff",
          4305 => x"0614b411",
          4306 => x"3370882b",
          4307 => x"78077981",
          4308 => x"0671842a",
          4309 => x"5c525851",
          4310 => x"537280e2",
          4311 => x"38759fff",
          4312 => x"065880da",
          4313 => x"3976882a",
          4314 => x"a4150805",
          4315 => x"527351fc",
          4316 => x"bd3f81de",
          4317 => x"c00880c6",
          4318 => x"38761083",
          4319 => x"fe067405",
          4320 => x"b40551f9",
          4321 => x"8d3f81de",
          4322 => x"c00883ff",
          4323 => x"ff0658ae",
          4324 => x"3976872a",
          4325 => x"a4150805",
          4326 => x"527351fc",
          4327 => x"913f81de",
          4328 => x"c0089b38",
          4329 => x"76822b83",
          4330 => x"fc067405",
          4331 => x"b40551f8",
          4332 => x"f83f81de",
          4333 => x"c008f00a",
          4334 => x"06588339",
          4335 => x"81587781",
          4336 => x"dec00c89",
          4337 => x"3d0d04f8",
          4338 => x"3d0d7a7c",
          4339 => x"7e5a5856",
          4340 => x"82598177",
          4341 => x"27829e38",
          4342 => x"76981708",
          4343 => x"27829638",
          4344 => x"75335372",
          4345 => x"792e819d",
          4346 => x"38727924",
          4347 => x"89387281",
          4348 => x"2e8d3882",
          4349 => x"80397283",
          4350 => x"2e81b838",
          4351 => x"81f73976",
          4352 => x"812a1770",
          4353 => x"892aa418",
          4354 => x"08055376",
          4355 => x"5255fb9e",
          4356 => x"3f81dec0",
          4357 => x"085981de",
          4358 => x"c00881d9",
          4359 => x"387483ff",
          4360 => x"0616b405",
          4361 => x"81167881",
          4362 => x"06595654",
          4363 => x"77537680",
          4364 => x"2e8f3877",
          4365 => x"842b9ff0",
          4366 => x"0674338f",
          4367 => x"06710751",
          4368 => x"53727434",
          4369 => x"810b8317",
          4370 => x"3474892a",
          4371 => x"a4170805",
          4372 => x"527551fa",
          4373 => x"d93f81de",
          4374 => x"c0085981",
          4375 => x"dec00881",
          4376 => x"94387483",
          4377 => x"ff0616b4",
          4378 => x"0578842a",
          4379 => x"5454768f",
          4380 => x"3877882a",
          4381 => x"743381f0",
          4382 => x"06718f06",
          4383 => x"07515372",
          4384 => x"743480ec",
          4385 => x"3976882a",
          4386 => x"a4170805",
          4387 => x"527551fa",
          4388 => x"9d3f81de",
          4389 => x"c0085981",
          4390 => x"dec00880",
          4391 => x"d8387783",
          4392 => x"ffff0652",
          4393 => x"761083fe",
          4394 => x"067605b4",
          4395 => x"0551f7a4",
          4396 => x"3fbe3976",
          4397 => x"872aa417",
          4398 => x"08055275",
          4399 => x"51f9ef3f",
          4400 => x"81dec008",
          4401 => x"5981dec0",
          4402 => x"08ab3877",
          4403 => x"f00a0677",
          4404 => x"822b83fc",
          4405 => x"067018b4",
          4406 => x"05705451",
          4407 => x"5454f6c9",
          4408 => x"3f81dec0",
          4409 => x"088f0a06",
          4410 => x"74075272",
          4411 => x"51f7833f",
          4412 => x"810b8317",
          4413 => x"347881de",
          4414 => x"c00c8a3d",
          4415 => x"0d04f83d",
          4416 => x"0d7a7c7e",
          4417 => x"72085956",
          4418 => x"56598175",
          4419 => x"27a43874",
          4420 => x"98170827",
          4421 => x"9d387380",
          4422 => x"2eaa38ff",
          4423 => x"53735275",
          4424 => x"51fda43f",
          4425 => x"81dec008",
          4426 => x"5481dec0",
          4427 => x"0880f238",
          4428 => x"93398254",
          4429 => x"80eb3981",
          4430 => x"5480e639",
          4431 => x"81dec008",
          4432 => x"5480de39",
          4433 => x"74527851",
          4434 => x"fb843f81",
          4435 => x"dec00858",
          4436 => x"81dec008",
          4437 => x"802e80c7",
          4438 => x"3881dec0",
          4439 => x"08812ed2",
          4440 => x"3881dec0",
          4441 => x"08ff2ecf",
          4442 => x"38805374",
          4443 => x"527551fc",
          4444 => x"d63f81de",
          4445 => x"c008c538",
          4446 => x"981608fe",
          4447 => x"11901808",
          4448 => x"57555774",
          4449 => x"74279038",
          4450 => x"81159017",
          4451 => x"0c841633",
          4452 => x"81075473",
          4453 => x"84173477",
          4454 => x"55767826",
          4455 => x"ffa63880",
          4456 => x"547381de",
          4457 => x"c00c8a3d",
          4458 => x"0d04f63d",
          4459 => x"0d7c7e71",
          4460 => x"08595b5b",
          4461 => x"7995388c",
          4462 => x"17085877",
          4463 => x"802e8838",
          4464 => x"98170878",
          4465 => x"26b23881",
          4466 => x"58ae3979",
          4467 => x"527a51f9",
          4468 => x"fd3f8155",
          4469 => x"7481dec0",
          4470 => x"082782e0",
          4471 => x"3881dec0",
          4472 => x"085581de",
          4473 => x"c008ff2e",
          4474 => x"82d23898",
          4475 => x"170881de",
          4476 => x"c0082682",
          4477 => x"c7387958",
          4478 => x"90170870",
          4479 => x"56547380",
          4480 => x"2e82b938",
          4481 => x"777a2e09",
          4482 => x"810680e2",
          4483 => x"38811a56",
          4484 => x"98170876",
          4485 => x"26833882",
          4486 => x"5675527a",
          4487 => x"51f9af3f",
          4488 => x"805981de",
          4489 => x"c008812e",
          4490 => x"09810686",
          4491 => x"3881dec0",
          4492 => x"085981de",
          4493 => x"c0080970",
          4494 => x"30707207",
          4495 => x"8025707c",
          4496 => x"0781dec0",
          4497 => x"08545151",
          4498 => x"55557381",
          4499 => x"ef3881de",
          4500 => x"c008802e",
          4501 => x"95388c17",
          4502 => x"08548174",
          4503 => x"27903873",
          4504 => x"98180827",
          4505 => x"89387358",
          4506 => x"85397580",
          4507 => x"db387756",
          4508 => x"81165698",
          4509 => x"17087626",
          4510 => x"89388256",
          4511 => x"75782681",
          4512 => x"ac387552",
          4513 => x"7a51f8c6",
          4514 => x"3f81dec0",
          4515 => x"08802eb8",
          4516 => x"38805981",
          4517 => x"dec00881",
          4518 => x"2e098106",
          4519 => x"863881de",
          4520 => x"c0085981",
          4521 => x"dec00809",
          4522 => x"70307072",
          4523 => x"07802570",
          4524 => x"7c075151",
          4525 => x"55557380",
          4526 => x"f8387578",
          4527 => x"2e098106",
          4528 => x"ffae3873",
          4529 => x"5580f539",
          4530 => x"ff537552",
          4531 => x"7651f9f7",
          4532 => x"3f81dec0",
          4533 => x"0881dec0",
          4534 => x"08307081",
          4535 => x"dec00807",
          4536 => x"80255155",
          4537 => x"5579802e",
          4538 => x"94387380",
          4539 => x"2e8f3875",
          4540 => x"53795276",
          4541 => x"51f9d03f",
          4542 => x"81dec008",
          4543 => x"5574a538",
          4544 => x"758c180c",
          4545 => x"981708fe",
          4546 => x"05901808",
          4547 => x"56547474",
          4548 => x"268638ff",
          4549 => x"1590180c",
          4550 => x"84173381",
          4551 => x"07547384",
          4552 => x"18349739",
          4553 => x"ff567481",
          4554 => x"2e90388c",
          4555 => x"3980558c",
          4556 => x"3981dec0",
          4557 => x"08558539",
          4558 => x"81567555",
          4559 => x"7481dec0",
          4560 => x"0c8c3d0d",
          4561 => x"04f83d0d",
          4562 => x"7a705255",
          4563 => x"f3f03f81",
          4564 => x"dec00858",
          4565 => x"815681de",
          4566 => x"c00880d8",
          4567 => x"387b5274",
          4568 => x"51f6c13f",
          4569 => x"81dec008",
          4570 => x"81dec008",
          4571 => x"b0170c59",
          4572 => x"84805377",
          4573 => x"52b41570",
          4574 => x"5257f2c8",
          4575 => x"3f775684",
          4576 => x"39811656",
          4577 => x"8a152258",
          4578 => x"75782797",
          4579 => x"38815475",
          4580 => x"19537652",
          4581 => x"81153351",
          4582 => x"ede93f81",
          4583 => x"dec00880",
          4584 => x"2edf388a",
          4585 => x"15227632",
          4586 => x"70307072",
          4587 => x"07709f2a",
          4588 => x"53515656",
          4589 => x"7581dec0",
          4590 => x"0c8a3d0d",
          4591 => x"04f83d0d",
          4592 => x"7a7c7108",
          4593 => x"58565774",
          4594 => x"f0800a26",
          4595 => x"80f13874",
          4596 => x"9f065372",
          4597 => x"80e93874",
          4598 => x"90180c88",
          4599 => x"17085473",
          4600 => x"aa387533",
          4601 => x"53827327",
          4602 => x"8838a816",
          4603 => x"0854739b",
          4604 => x"3874852a",
          4605 => x"53820b88",
          4606 => x"17225a58",
          4607 => x"72792780",
          4608 => x"fe38a816",
          4609 => x"0898180c",
          4610 => x"80cd398a",
          4611 => x"16227089",
          4612 => x"2b545872",
          4613 => x"7526b238",
          4614 => x"73527651",
          4615 => x"f5b03f81",
          4616 => x"dec00854",
          4617 => x"81dec008",
          4618 => x"ff2ebd38",
          4619 => x"810b81de",
          4620 => x"c008278b",
          4621 => x"38981608",
          4622 => x"81dec008",
          4623 => x"26853882",
          4624 => x"58bd3974",
          4625 => x"733155cb",
          4626 => x"39735275",
          4627 => x"51f4d53f",
          4628 => x"81dec008",
          4629 => x"98180c73",
          4630 => x"94180c98",
          4631 => x"17085382",
          4632 => x"5872802e",
          4633 => x"9a388539",
          4634 => x"81589439",
          4635 => x"74892a13",
          4636 => x"98180c74",
          4637 => x"83ff0616",
          4638 => x"b4059c18",
          4639 => x"0c805877",
          4640 => x"81dec00c",
          4641 => x"8a3d0d04",
          4642 => x"f83d0d7a",
          4643 => x"70089012",
          4644 => x"08a00559",
          4645 => x"5754f080",
          4646 => x"0a772786",
          4647 => x"38800b98",
          4648 => x"150c9814",
          4649 => x"08538455",
          4650 => x"72802e81",
          4651 => x"cb387683",
          4652 => x"ff065877",
          4653 => x"81b53881",
          4654 => x"1398150c",
          4655 => x"94140855",
          4656 => x"74923876",
          4657 => x"852a8817",
          4658 => x"22565374",
          4659 => x"7326819b",
          4660 => x"3880c039",
          4661 => x"8a1622ff",
          4662 => x"0577892a",
          4663 => x"06537281",
          4664 => x"8a387452",
          4665 => x"7351f3e6",
          4666 => x"3f81dec0",
          4667 => x"08538255",
          4668 => x"810b81de",
          4669 => x"c0082780",
          4670 => x"ff388155",
          4671 => x"81dec008",
          4672 => x"ff2e80f4",
          4673 => x"38981608",
          4674 => x"81dec008",
          4675 => x"2680ca38",
          4676 => x"7b8a3877",
          4677 => x"98150c84",
          4678 => x"5580dd39",
          4679 => x"94140852",
          4680 => x"7351f986",
          4681 => x"3f81dec0",
          4682 => x"08538755",
          4683 => x"81dec008",
          4684 => x"802e80c4",
          4685 => x"38825581",
          4686 => x"dec00881",
          4687 => x"2eba3881",
          4688 => x"5581dec0",
          4689 => x"08ff2eb0",
          4690 => x"3881dec0",
          4691 => x"08527551",
          4692 => x"fbf33f81",
          4693 => x"dec008a0",
          4694 => x"38729415",
          4695 => x"0c725275",
          4696 => x"51f2c13f",
          4697 => x"81dec008",
          4698 => x"98150c76",
          4699 => x"90150c77",
          4700 => x"16b4059c",
          4701 => x"150c8055",
          4702 => x"7481dec0",
          4703 => x"0c8a3d0d",
          4704 => x"04f73d0d",
          4705 => x"7b7d7108",
          4706 => x"5b5b5780",
          4707 => x"527651fc",
          4708 => x"ac3f81de",
          4709 => x"c0085481",
          4710 => x"dec00880",
          4711 => x"ec3881de",
          4712 => x"c0085698",
          4713 => x"17085278",
          4714 => x"51f0833f",
          4715 => x"81dec008",
          4716 => x"5481dec0",
          4717 => x"0880d238",
          4718 => x"81dec008",
          4719 => x"9c180870",
          4720 => x"33515458",
          4721 => x"7281e52e",
          4722 => x"09810683",
          4723 => x"38815881",
          4724 => x"dec00855",
          4725 => x"72833881",
          4726 => x"55777507",
          4727 => x"5372802e",
          4728 => x"8e388116",
          4729 => x"56757a2e",
          4730 => x"09810688",
          4731 => x"38a53981",
          4732 => x"dec00856",
          4733 => x"81527651",
          4734 => x"fd8e3f81",
          4735 => x"dec00854",
          4736 => x"81dec008",
          4737 => x"802eff9b",
          4738 => x"3873842e",
          4739 => x"09810683",
          4740 => x"38875473",
          4741 => x"81dec00c",
          4742 => x"8b3d0d04",
          4743 => x"fd3d0d76",
          4744 => x"9a115254",
          4745 => x"ebec3f81",
          4746 => x"dec00883",
          4747 => x"ffff0676",
          4748 => x"70335153",
          4749 => x"5371832e",
          4750 => x"09810690",
          4751 => x"38941451",
          4752 => x"ebd03f81",
          4753 => x"dec00890",
          4754 => x"2b730753",
          4755 => x"7281dec0",
          4756 => x"0c853d0d",
          4757 => x"04fc3d0d",
          4758 => x"77797083",
          4759 => x"ffff0654",
          4760 => x"9a125355",
          4761 => x"55ebed3f",
          4762 => x"76703351",
          4763 => x"5372832e",
          4764 => x"0981068b",
          4765 => x"3873902a",
          4766 => x"52941551",
          4767 => x"ebd63f86",
          4768 => x"3d0d04f7",
          4769 => x"3d0d7b7d",
          4770 => x"5b558475",
          4771 => x"085a5898",
          4772 => x"1508802e",
          4773 => x"818a3898",
          4774 => x"15085278",
          4775 => x"51ee8f3f",
          4776 => x"81dec008",
          4777 => x"5881dec0",
          4778 => x"0880f538",
          4779 => x"9c150870",
          4780 => x"33555373",
          4781 => x"86388458",
          4782 => x"80e6398b",
          4783 => x"133370bf",
          4784 => x"067081ff",
          4785 => x"06585153",
          4786 => x"72861634",
          4787 => x"81dec008",
          4788 => x"537381e5",
          4789 => x"2e833881",
          4790 => x"5373ae2e",
          4791 => x"a9388170",
          4792 => x"74065457",
          4793 => x"72802e9e",
          4794 => x"38758f2e",
          4795 => x"993881de",
          4796 => x"c00876df",
          4797 => x"06545472",
          4798 => x"882e0981",
          4799 => x"06833876",
          4800 => x"54737a2e",
          4801 => x"a0388052",
          4802 => x"7451fafc",
          4803 => x"3f81dec0",
          4804 => x"085881de",
          4805 => x"c0088938",
          4806 => x"981508fe",
          4807 => x"fa388639",
          4808 => x"800b9816",
          4809 => x"0c7781de",
          4810 => x"c00c8b3d",
          4811 => x"0d04fb3d",
          4812 => x"0d777008",
          4813 => x"57548152",
          4814 => x"7351fcc5",
          4815 => x"3f81dec0",
          4816 => x"085581de",
          4817 => x"c008b438",
          4818 => x"98140852",
          4819 => x"7551ecde",
          4820 => x"3f81dec0",
          4821 => x"085581de",
          4822 => x"c008a038",
          4823 => x"a05381de",
          4824 => x"c008529c",
          4825 => x"140851ea",
          4826 => x"db3f8b53",
          4827 => x"a014529c",
          4828 => x"140851ea",
          4829 => x"ac3f810b",
          4830 => x"83173474",
          4831 => x"81dec00c",
          4832 => x"873d0d04",
          4833 => x"fd3d0d75",
          4834 => x"70089812",
          4835 => x"08547053",
          4836 => x"5553ec9a",
          4837 => x"3f81dec0",
          4838 => x"088d389c",
          4839 => x"130853e5",
          4840 => x"7334810b",
          4841 => x"83153485",
          4842 => x"3d0d04fa",
          4843 => x"3d0d787a",
          4844 => x"5757800b",
          4845 => x"89173498",
          4846 => x"1708802e",
          4847 => x"81823880",
          4848 => x"70891855",
          4849 => x"55559c17",
          4850 => x"08147033",
          4851 => x"81165651",
          4852 => x"5271a02e",
          4853 => x"a8387185",
          4854 => x"2e098106",
          4855 => x"843881e5",
          4856 => x"5273892e",
          4857 => x"0981068b",
          4858 => x"38ae7370",
          4859 => x"81055534",
          4860 => x"81155571",
          4861 => x"73708105",
          4862 => x"55348115",
          4863 => x"558a7427",
          4864 => x"c5387515",
          4865 => x"88055280",
          4866 => x"0b811334",
          4867 => x"9c170852",
          4868 => x"8b123388",
          4869 => x"17349c17",
          4870 => x"089c1152",
          4871 => x"52e88a3f",
          4872 => x"81dec008",
          4873 => x"760c9612",
          4874 => x"51e7e73f",
          4875 => x"81dec008",
          4876 => x"86172398",
          4877 => x"1251e7da",
          4878 => x"3f81dec0",
          4879 => x"08841723",
          4880 => x"883d0d04",
          4881 => x"f33d0d7f",
          4882 => x"70085e5b",
          4883 => x"80617033",
          4884 => x"51555573",
          4885 => x"af2e8338",
          4886 => x"81557380",
          4887 => x"dc2e9138",
          4888 => x"74802e8c",
          4889 => x"38941d08",
          4890 => x"881c0caa",
          4891 => x"39811541",
          4892 => x"80617033",
          4893 => x"56565673",
          4894 => x"af2e0981",
          4895 => x"06833881",
          4896 => x"567380dc",
          4897 => x"32703070",
          4898 => x"80257807",
          4899 => x"51515473",
          4900 => x"dc387388",
          4901 => x"1c0c6070",
          4902 => x"33515473",
          4903 => x"9f269638",
          4904 => x"ff800bab",
          4905 => x"1c348052",
          4906 => x"7a51f691",
          4907 => x"3f81dec0",
          4908 => x"08558598",
          4909 => x"39913d61",
          4910 => x"a01d5c5a",
          4911 => x"5e8b53a0",
          4912 => x"527951e7",
          4913 => x"ff3f8070",
          4914 => x"59578879",
          4915 => x"33555c73",
          4916 => x"ae2e0981",
          4917 => x"0680d438",
          4918 => x"78187033",
          4919 => x"811a71ae",
          4920 => x"32703070",
          4921 => x"9f2a7382",
          4922 => x"26075151",
          4923 => x"535a5754",
          4924 => x"738c3879",
          4925 => x"17547574",
          4926 => x"34811757",
          4927 => x"db3975af",
          4928 => x"32703070",
          4929 => x"9f2a5151",
          4930 => x"547580dc",
          4931 => x"2e8c3873",
          4932 => x"802e8738",
          4933 => x"75a02682",
          4934 => x"bd387719",
          4935 => x"7e0ca454",
          4936 => x"a0762782",
          4937 => x"bd38a054",
          4938 => x"82b83978",
          4939 => x"18703381",
          4940 => x"1a5a5754",
          4941 => x"a0762781",
          4942 => x"fc3875af",
          4943 => x"32703077",
          4944 => x"80dc3270",
          4945 => x"30728025",
          4946 => x"71802507",
          4947 => x"51515651",
          4948 => x"5573802e",
          4949 => x"ac388439",
          4950 => x"81185880",
          4951 => x"781a7033",
          4952 => x"51555573",
          4953 => x"af2e0981",
          4954 => x"06833881",
          4955 => x"557380dc",
          4956 => x"32703070",
          4957 => x"80257707",
          4958 => x"51515473",
          4959 => x"db3881b5",
          4960 => x"3975ae2e",
          4961 => x"09810683",
          4962 => x"38815476",
          4963 => x"7c277407",
          4964 => x"5473802e",
          4965 => x"a2387b8b",
          4966 => x"32703077",
          4967 => x"ae327030",
          4968 => x"72802571",
          4969 => x"9f2a0753",
          4970 => x"51565155",
          4971 => x"7481a738",
          4972 => x"88578b5c",
          4973 => x"fef53975",
          4974 => x"982b5473",
          4975 => x"80258c38",
          4976 => x"7580ff06",
          4977 => x"81cdb411",
          4978 => x"33575475",
          4979 => x"51e6e13f",
          4980 => x"81dec008",
          4981 => x"802eb238",
          4982 => x"78187033",
          4983 => x"811a7154",
          4984 => x"5a5654e6",
          4985 => x"d23f81de",
          4986 => x"c008802e",
          4987 => x"80e838ff",
          4988 => x"1c547674",
          4989 => x"2780df38",
          4990 => x"79175475",
          4991 => x"74348117",
          4992 => x"7a115557",
          4993 => x"747434a7",
          4994 => x"39755281",
          4995 => x"ccd451e5",
          4996 => x"fe3f81de",
          4997 => x"c008bf38",
          4998 => x"ff9f1654",
          4999 => x"73992689",
          5000 => x"38e01670",
          5001 => x"81ff0657",
          5002 => x"54791754",
          5003 => x"75743481",
          5004 => x"1757fdf7",
          5005 => x"3977197e",
          5006 => x"0c76802e",
          5007 => x"99387933",
          5008 => x"547381e5",
          5009 => x"2e098106",
          5010 => x"8438857a",
          5011 => x"348454a0",
          5012 => x"76278f38",
          5013 => x"8b398655",
          5014 => x"81f23984",
          5015 => x"5680f339",
          5016 => x"8054738b",
          5017 => x"1b34807b",
          5018 => x"0858527a",
          5019 => x"51f2ce3f",
          5020 => x"81dec008",
          5021 => x"5681dec0",
          5022 => x"0880d738",
          5023 => x"981b0852",
          5024 => x"7651e6aa",
          5025 => x"3f81dec0",
          5026 => x"085681de",
          5027 => x"c00880c2",
          5028 => x"389c1b08",
          5029 => x"70335555",
          5030 => x"73802eff",
          5031 => x"be388b15",
          5032 => x"33bf0654",
          5033 => x"73861c34",
          5034 => x"8b153370",
          5035 => x"832a7081",
          5036 => x"06515558",
          5037 => x"7392388b",
          5038 => x"53795274",
          5039 => x"51e49f3f",
          5040 => x"81dec008",
          5041 => x"802e8b38",
          5042 => x"75527a51",
          5043 => x"f3ba3fff",
          5044 => x"9f3975ab",
          5045 => x"1c335755",
          5046 => x"74802ebb",
          5047 => x"3874842e",
          5048 => x"09810680",
          5049 => x"e7387585",
          5050 => x"2a708106",
          5051 => x"77822a58",
          5052 => x"51547380",
          5053 => x"2e963875",
          5054 => x"81065473",
          5055 => x"802efbb5",
          5056 => x"38ff800b",
          5057 => x"ab1c3480",
          5058 => x"5580c139",
          5059 => x"75810654",
          5060 => x"73ba3885",
          5061 => x"55b63975",
          5062 => x"822a7081",
          5063 => x"06515473",
          5064 => x"ab38861b",
          5065 => x"3370842a",
          5066 => x"70810651",
          5067 => x"55557380",
          5068 => x"2ee13890",
          5069 => x"1b0883ff",
          5070 => x"061db405",
          5071 => x"527c51f5",
          5072 => x"db3f81de",
          5073 => x"c008881c",
          5074 => x"0cfaea39",
          5075 => x"7481dec0",
          5076 => x"0c8f3d0d",
          5077 => x"04f63d0d",
          5078 => x"7c5bff7b",
          5079 => x"08707173",
          5080 => x"55595c55",
          5081 => x"5973802e",
          5082 => x"81c63875",
          5083 => x"70810557",
          5084 => x"3370a026",
          5085 => x"525271ba",
          5086 => x"2e8d3870",
          5087 => x"ee3871ba",
          5088 => x"2e098106",
          5089 => x"81a53873",
          5090 => x"33d01170",
          5091 => x"81ff0651",
          5092 => x"52537089",
          5093 => x"26913882",
          5094 => x"147381ff",
          5095 => x"06d00556",
          5096 => x"5271762e",
          5097 => x"80f73880",
          5098 => x"0b81cda4",
          5099 => x"59557708",
          5100 => x"7a555776",
          5101 => x"70810558",
          5102 => x"33747081",
          5103 => x"055633ff",
          5104 => x"9f125353",
          5105 => x"53709926",
          5106 => x"8938e013",
          5107 => x"7081ff06",
          5108 => x"5451ff9f",
          5109 => x"12517099",
          5110 => x"268938e0",
          5111 => x"127081ff",
          5112 => x"06535172",
          5113 => x"30709f2a",
          5114 => x"51517272",
          5115 => x"2e098106",
          5116 => x"853870ff",
          5117 => x"be387230",
          5118 => x"74773270",
          5119 => x"30707207",
          5120 => x"9f2a739f",
          5121 => x"2a075354",
          5122 => x"54517080",
          5123 => x"2e8f3881",
          5124 => x"15841959",
          5125 => x"55837525",
          5126 => x"ff94388b",
          5127 => x"39748324",
          5128 => x"86387476",
          5129 => x"7c0c5978",
          5130 => x"51863981",
          5131 => x"def03351",
          5132 => x"7081dec0",
          5133 => x"0c8c3d0d",
          5134 => x"04fa3d0d",
          5135 => x"7856800b",
          5136 => x"831734ff",
          5137 => x"0bb0170c",
          5138 => x"79527551",
          5139 => x"e2e03f84",
          5140 => x"5581dec0",
          5141 => x"08818038",
          5142 => x"84b21651",
          5143 => x"dfb43f81",
          5144 => x"dec00883",
          5145 => x"ffff0654",
          5146 => x"83557382",
          5147 => x"d4d52e09",
          5148 => x"810680e3",
          5149 => x"38800bb4",
          5150 => x"17335657",
          5151 => x"7481e92e",
          5152 => x"09810683",
          5153 => x"38815774",
          5154 => x"81eb3270",
          5155 => x"30708025",
          5156 => x"79075151",
          5157 => x"54738a38",
          5158 => x"7481e82e",
          5159 => x"098106b5",
          5160 => x"38835381",
          5161 => x"cce45280",
          5162 => x"ea1651e0",
          5163 => x"b13f81de",
          5164 => x"c0085581",
          5165 => x"dec00880",
          5166 => x"2e9d3885",
          5167 => x"5381cce8",
          5168 => x"52818616",
          5169 => x"51e0973f",
          5170 => x"81dec008",
          5171 => x"5581dec0",
          5172 => x"08802e83",
          5173 => x"38825574",
          5174 => x"81dec00c",
          5175 => x"883d0d04",
          5176 => x"f23d0d61",
          5177 => x"02840580",
          5178 => x"cb053358",
          5179 => x"5580750c",
          5180 => x"6051fce1",
          5181 => x"3f81dec0",
          5182 => x"08588b56",
          5183 => x"800b81de",
          5184 => x"c0082486",
          5185 => x"fc3881de",
          5186 => x"c0088429",
          5187 => x"81dedc05",
          5188 => x"70085553",
          5189 => x"8c567380",
          5190 => x"2e86e638",
          5191 => x"73750c76",
          5192 => x"81fe0674",
          5193 => x"33545772",
          5194 => x"802eae38",
          5195 => x"81143351",
          5196 => x"d7ca3f81",
          5197 => x"dec00881",
          5198 => x"ff067081",
          5199 => x"06545572",
          5200 => x"98387680",
          5201 => x"2e86b838",
          5202 => x"74822a70",
          5203 => x"81065153",
          5204 => x"8a567286",
          5205 => x"ac3886a7",
          5206 => x"39807434",
          5207 => x"77811534",
          5208 => x"81528114",
          5209 => x"3351d7b2",
          5210 => x"3f81dec0",
          5211 => x"0881ff06",
          5212 => x"70810654",
          5213 => x"55835672",
          5214 => x"86873876",
          5215 => x"802e8f38",
          5216 => x"74822a70",
          5217 => x"81065153",
          5218 => x"8a567285",
          5219 => x"f4388070",
          5220 => x"5374525b",
          5221 => x"fda33f81",
          5222 => x"dec00881",
          5223 => x"ff065776",
          5224 => x"822e0981",
          5225 => x"0680e238",
          5226 => x"8c3d7456",
          5227 => x"58835683",
          5228 => x"f6153370",
          5229 => x"58537280",
          5230 => x"2e8d3883",
          5231 => x"fa1551dc",
          5232 => x"e83f81de",
          5233 => x"c0085776",
          5234 => x"78708405",
          5235 => x"5a0cff16",
          5236 => x"90165656",
          5237 => x"758025d7",
          5238 => x"38800b8d",
          5239 => x"3d545672",
          5240 => x"70840554",
          5241 => x"085b8357",
          5242 => x"7a802e95",
          5243 => x"387a5273",
          5244 => x"51fcc63f",
          5245 => x"81dec008",
          5246 => x"81ff0657",
          5247 => x"81772789",
          5248 => x"38811656",
          5249 => x"837627d7",
          5250 => x"38815676",
          5251 => x"842e84f1",
          5252 => x"388d5676",
          5253 => x"812684e9",
          5254 => x"38bf1451",
          5255 => x"dbf43f81",
          5256 => x"dec00883",
          5257 => x"ffff0653",
          5258 => x"7284802e",
          5259 => x"09810684",
          5260 => x"d03880ca",
          5261 => x"1451dbda",
          5262 => x"3f81dec0",
          5263 => x"0883ffff",
          5264 => x"0658778d",
          5265 => x"3880d814",
          5266 => x"51dbde3f",
          5267 => x"81dec008",
          5268 => x"58779c15",
          5269 => x"0c80c414",
          5270 => x"33821534",
          5271 => x"80c41433",
          5272 => x"ff117081",
          5273 => x"ff065154",
          5274 => x"558d5672",
          5275 => x"81268491",
          5276 => x"387481ff",
          5277 => x"06787129",
          5278 => x"80c11633",
          5279 => x"52595372",
          5280 => x"8a152372",
          5281 => x"802e8b38",
          5282 => x"ff137306",
          5283 => x"5372802e",
          5284 => x"86388d56",
          5285 => x"83eb3980",
          5286 => x"c51451da",
          5287 => x"f53f81de",
          5288 => x"c0085381",
          5289 => x"dec00888",
          5290 => x"1523728f",
          5291 => x"06578d56",
          5292 => x"7683ce38",
          5293 => x"80c71451",
          5294 => x"dad83f81",
          5295 => x"dec00883",
          5296 => x"ffff0655",
          5297 => x"748d3880",
          5298 => x"d41451da",
          5299 => x"dc3f81de",
          5300 => x"c0085580",
          5301 => x"c21451da",
          5302 => x"b93f81de",
          5303 => x"c00883ff",
          5304 => x"ff06538d",
          5305 => x"5672802e",
          5306 => x"83973888",
          5307 => x"14227814",
          5308 => x"71842a05",
          5309 => x"5a5a7875",
          5310 => x"26838638",
          5311 => x"8a142252",
          5312 => x"74793151",
          5313 => x"ffacf03f",
          5314 => x"81dec008",
          5315 => x"5581dec0",
          5316 => x"08802e82",
          5317 => x"ec3881de",
          5318 => x"c00880ff",
          5319 => x"fffff526",
          5320 => x"83388357",
          5321 => x"7483fff5",
          5322 => x"26833882",
          5323 => x"57749ff5",
          5324 => x"26853881",
          5325 => x"5789398d",
          5326 => x"5676802e",
          5327 => x"82c33882",
          5328 => x"15709816",
          5329 => x"0c7ba016",
          5330 => x"0c731c70",
          5331 => x"a4170c7a",
          5332 => x"1dac170c",
          5333 => x"54557683",
          5334 => x"2e098106",
          5335 => x"af3880de",
          5336 => x"1451d9ae",
          5337 => x"3f81dec0",
          5338 => x"0883ffff",
          5339 => x"06538d56",
          5340 => x"72828e38",
          5341 => x"79828a38",
          5342 => x"80e01451",
          5343 => x"d9ab3f81",
          5344 => x"dec008a8",
          5345 => x"150c7482",
          5346 => x"2b53a239",
          5347 => x"8d567980",
          5348 => x"2e81ee38",
          5349 => x"7713a815",
          5350 => x"0c741553",
          5351 => x"76822e8d",
          5352 => x"38741015",
          5353 => x"70812a76",
          5354 => x"81060551",
          5355 => x"5383ff13",
          5356 => x"892a538d",
          5357 => x"56729c15",
          5358 => x"082681c5",
          5359 => x"38ff0b90",
          5360 => x"150cff0b",
          5361 => x"8c150cff",
          5362 => x"800b8415",
          5363 => x"3476832e",
          5364 => x"09810681",
          5365 => x"923880e4",
          5366 => x"1451d8b6",
          5367 => x"3f81dec0",
          5368 => x"0883ffff",
          5369 => x"06537281",
          5370 => x"2e098106",
          5371 => x"80f93881",
          5372 => x"1b527351",
          5373 => x"dbb83f81",
          5374 => x"dec00880",
          5375 => x"ea3881de",
          5376 => x"c0088415",
          5377 => x"3484b214",
          5378 => x"51d8873f",
          5379 => x"81dec008",
          5380 => x"83ffff06",
          5381 => x"537282d4",
          5382 => x"d52e0981",
          5383 => x"0680c838",
          5384 => x"b41451d8",
          5385 => x"843f81de",
          5386 => x"c008848b",
          5387 => x"85a4d22e",
          5388 => x"098106b3",
          5389 => x"38849814",
          5390 => x"51d7ee3f",
          5391 => x"81dec008",
          5392 => x"868a85e4",
          5393 => x"f22e0981",
          5394 => x"069d3884",
          5395 => x"9c1451d7",
          5396 => x"d83f81de",
          5397 => x"c0089015",
          5398 => x"0c84a014",
          5399 => x"51d7ca3f",
          5400 => x"81dec008",
          5401 => x"8c150c76",
          5402 => x"743481de",
          5403 => x"ec228105",
          5404 => x"537281de",
          5405 => x"ec237286",
          5406 => x"1523800b",
          5407 => x"94150c80",
          5408 => x"567581de",
          5409 => x"c00c903d",
          5410 => x"0d04fb3d",
          5411 => x"0d775489",
          5412 => x"5573802e",
          5413 => x"b9387308",
          5414 => x"5372802e",
          5415 => x"b1387233",
          5416 => x"5271802e",
          5417 => x"a9388613",
          5418 => x"22841522",
          5419 => x"57527176",
          5420 => x"2e098106",
          5421 => x"99388113",
          5422 => x"3351d0c0",
          5423 => x"3f81dec0",
          5424 => x"08810652",
          5425 => x"71883871",
          5426 => x"74085455",
          5427 => x"83398053",
          5428 => x"7873710c",
          5429 => x"527481de",
          5430 => x"c00c873d",
          5431 => x"0d04fa3d",
          5432 => x"0d02ab05",
          5433 => x"337a5889",
          5434 => x"3dfc0552",
          5435 => x"56f4e63f",
          5436 => x"8b54800b",
          5437 => x"81dec008",
          5438 => x"24bc3881",
          5439 => x"dec00884",
          5440 => x"2981dedc",
          5441 => x"05700855",
          5442 => x"5573802e",
          5443 => x"84388074",
          5444 => x"34785473",
          5445 => x"802e8438",
          5446 => x"80743478",
          5447 => x"750c7554",
          5448 => x"75802e92",
          5449 => x"38805389",
          5450 => x"3d705384",
          5451 => x"0551f7b0",
          5452 => x"3f81dec0",
          5453 => x"08547381",
          5454 => x"dec00c88",
          5455 => x"3d0d04eb",
          5456 => x"3d0d6702",
          5457 => x"840580e7",
          5458 => x"05335959",
          5459 => x"89547880",
          5460 => x"2e84c838",
          5461 => x"77bf0670",
          5462 => x"54983dd0",
          5463 => x"0553993d",
          5464 => x"84055258",
          5465 => x"f6fa3f81",
          5466 => x"dec00855",
          5467 => x"81dec008",
          5468 => x"84a4387a",
          5469 => x"5c68528c",
          5470 => x"3d705256",
          5471 => x"edc63f81",
          5472 => x"dec00855",
          5473 => x"81dec008",
          5474 => x"92380280",
          5475 => x"d7053370",
          5476 => x"982b5557",
          5477 => x"73802583",
          5478 => x"38865577",
          5479 => x"9c065473",
          5480 => x"802e81ab",
          5481 => x"3874802e",
          5482 => x"95387484",
          5483 => x"2e098106",
          5484 => x"aa387551",
          5485 => x"eaf83f81",
          5486 => x"dec00855",
          5487 => x"9e3902b2",
          5488 => x"05339106",
          5489 => x"547381b8",
          5490 => x"3877822a",
          5491 => x"70810651",
          5492 => x"5473802e",
          5493 => x"8e388855",
          5494 => x"83bc3977",
          5495 => x"88075874",
          5496 => x"83b43877",
          5497 => x"832a7081",
          5498 => x"06515473",
          5499 => x"802e81af",
          5500 => x"3862527a",
          5501 => x"51e8a53f",
          5502 => x"81dec008",
          5503 => x"568288b2",
          5504 => x"0a52628e",
          5505 => x"0551d4ea",
          5506 => x"3f6254a0",
          5507 => x"0b8b1534",
          5508 => x"80536252",
          5509 => x"7a51e8bd",
          5510 => x"3f805262",
          5511 => x"9c0551d4",
          5512 => x"d13f7a54",
          5513 => x"810b8315",
          5514 => x"3475802e",
          5515 => x"80f1387a",
          5516 => x"b0110851",
          5517 => x"54805375",
          5518 => x"52973dd4",
          5519 => x"0551ddbe",
          5520 => x"3f81dec0",
          5521 => x"085581de",
          5522 => x"c00882ca",
          5523 => x"38b73974",
          5524 => x"82c43802",
          5525 => x"b2053370",
          5526 => x"842a7081",
          5527 => x"06515556",
          5528 => x"73802e86",
          5529 => x"38845582",
          5530 => x"ad397781",
          5531 => x"2a708106",
          5532 => x"51547380",
          5533 => x"2ea93875",
          5534 => x"81065473",
          5535 => x"802ea038",
          5536 => x"87558292",
          5537 => x"3973527a",
          5538 => x"51d6a33f",
          5539 => x"81dec008",
          5540 => x"7bff188c",
          5541 => x"120c5555",
          5542 => x"81dec008",
          5543 => x"81f83877",
          5544 => x"832a7081",
          5545 => x"06515473",
          5546 => x"802e8638",
          5547 => x"7780c007",
          5548 => x"587ab011",
          5549 => x"08a01b0c",
          5550 => x"63a41b0c",
          5551 => x"63537052",
          5552 => x"57e6d93f",
          5553 => x"81dec008",
          5554 => x"81dec008",
          5555 => x"881b0c63",
          5556 => x"9c05525a",
          5557 => x"d2d33f81",
          5558 => x"dec00881",
          5559 => x"dec0088c",
          5560 => x"1b0c777a",
          5561 => x"0c568617",
          5562 => x"22841a23",
          5563 => x"77901a34",
          5564 => x"800b911a",
          5565 => x"34800b9c",
          5566 => x"1a0c800b",
          5567 => x"941a0c77",
          5568 => x"852a7081",
          5569 => x"06515473",
          5570 => x"802e818d",
          5571 => x"3881dec0",
          5572 => x"08802e81",
          5573 => x"843881de",
          5574 => x"c008941a",
          5575 => x"0c8a1722",
          5576 => x"70892b7b",
          5577 => x"525957a8",
          5578 => x"39765278",
          5579 => x"51d79f3f",
          5580 => x"81dec008",
          5581 => x"5781dec0",
          5582 => x"08812683",
          5583 => x"38825581",
          5584 => x"dec008ff",
          5585 => x"2e098106",
          5586 => x"83387955",
          5587 => x"75783156",
          5588 => x"74307076",
          5589 => x"07802551",
          5590 => x"54777627",
          5591 => x"8a388170",
          5592 => x"7506555a",
          5593 => x"73c33876",
          5594 => x"981a0c74",
          5595 => x"a9387583",
          5596 => x"ff065473",
          5597 => x"802ea238",
          5598 => x"76527a51",
          5599 => x"d6a63f81",
          5600 => x"dec00885",
          5601 => x"3882558e",
          5602 => x"3975892a",
          5603 => x"81dec008",
          5604 => x"059c1a0c",
          5605 => x"84398079",
          5606 => x"0c745473",
          5607 => x"81dec00c",
          5608 => x"973d0d04",
          5609 => x"f23d0d60",
          5610 => x"63656440",
          5611 => x"405d5980",
          5612 => x"7e0c903d",
          5613 => x"fc055278",
          5614 => x"51f9cf3f",
          5615 => x"81dec008",
          5616 => x"5581dec0",
          5617 => x"088a3891",
          5618 => x"19335574",
          5619 => x"802e8638",
          5620 => x"745682c4",
          5621 => x"39901933",
          5622 => x"81065587",
          5623 => x"5674802e",
          5624 => x"82b63895",
          5625 => x"39820b91",
          5626 => x"1a348256",
          5627 => x"82aa3981",
          5628 => x"0b911a34",
          5629 => x"815682a0",
          5630 => x"398c1908",
          5631 => x"941a0831",
          5632 => x"55747c27",
          5633 => x"8338745c",
          5634 => x"7b802e82",
          5635 => x"89389419",
          5636 => x"087083ff",
          5637 => x"06565674",
          5638 => x"81b2387e",
          5639 => x"8a1122ff",
          5640 => x"0577892a",
          5641 => x"065b5579",
          5642 => x"a8387587",
          5643 => x"38881908",
          5644 => x"558f3998",
          5645 => x"19085278",
          5646 => x"51d5933f",
          5647 => x"81dec008",
          5648 => x"55817527",
          5649 => x"ff9f3874",
          5650 => x"ff2effa3",
          5651 => x"3874981a",
          5652 => x"0c981908",
          5653 => x"527e51d4",
          5654 => x"cb3f81de",
          5655 => x"c008802e",
          5656 => x"ff833881",
          5657 => x"dec0081a",
          5658 => x"7c892a59",
          5659 => x"5777802e",
          5660 => x"80d63877",
          5661 => x"1a7f8a11",
          5662 => x"22585c55",
          5663 => x"75752785",
          5664 => x"38757a31",
          5665 => x"58775476",
          5666 => x"537c5281",
          5667 => x"1b3351ca",
          5668 => x"883f81de",
          5669 => x"c008fed7",
          5670 => x"387e8311",
          5671 => x"33565674",
          5672 => x"802e9f38",
          5673 => x"b0160877",
          5674 => x"31557478",
          5675 => x"27943884",
          5676 => x"8053b416",
          5677 => x"52b01608",
          5678 => x"7731892b",
          5679 => x"7d0551cf",
          5680 => x"e03f7789",
          5681 => x"2b56b939",
          5682 => x"769c1a0c",
          5683 => x"94190883",
          5684 => x"ff068480",
          5685 => x"71315755",
          5686 => x"7b762783",
          5687 => x"387b569c",
          5688 => x"1908527e",
          5689 => x"51d1c73f",
          5690 => x"81dec008",
          5691 => x"fe813875",
          5692 => x"53941908",
          5693 => x"83ff061f",
          5694 => x"b405527c",
          5695 => x"51cfa23f",
          5696 => x"7b76317e",
          5697 => x"08177f0c",
          5698 => x"761e941b",
          5699 => x"0818941c",
          5700 => x"0c5e5cfd",
          5701 => x"f3398056",
          5702 => x"7581dec0",
          5703 => x"0c903d0d",
          5704 => x"04f23d0d",
          5705 => x"60636564",
          5706 => x"40405d58",
          5707 => x"807e0c90",
          5708 => x"3dfc0552",
          5709 => x"7751f6d2",
          5710 => x"3f81dec0",
          5711 => x"085581de",
          5712 => x"c0088a38",
          5713 => x"91183355",
          5714 => x"74802e86",
          5715 => x"38745683",
          5716 => x"b8399018",
          5717 => x"3370812a",
          5718 => x"70810651",
          5719 => x"56568756",
          5720 => x"74802e83",
          5721 => x"a4389539",
          5722 => x"820b9119",
          5723 => x"34825683",
          5724 => x"9839810b",
          5725 => x"91193481",
          5726 => x"56838e39",
          5727 => x"9418087c",
          5728 => x"11565674",
          5729 => x"76278438",
          5730 => x"75095c7b",
          5731 => x"802e82ec",
          5732 => x"38941808",
          5733 => x"7083ff06",
          5734 => x"56567481",
          5735 => x"fd387e8a",
          5736 => x"1122ff05",
          5737 => x"77892a06",
          5738 => x"5c557abf",
          5739 => x"38758c38",
          5740 => x"88180855",
          5741 => x"749c387a",
          5742 => x"52853998",
          5743 => x"18085277",
          5744 => x"51d7e73f",
          5745 => x"81dec008",
          5746 => x"5581dec0",
          5747 => x"08802e82",
          5748 => x"ab387481",
          5749 => x"2eff9138",
          5750 => x"74ff2eff",
          5751 => x"95387498",
          5752 => x"190c8818",
          5753 => x"08853874",
          5754 => x"88190c7e",
          5755 => x"55b01508",
          5756 => x"9c19082e",
          5757 => x"0981068d",
          5758 => x"387451ce",
          5759 => x"c13f81de",
          5760 => x"c008feee",
          5761 => x"38981808",
          5762 => x"527e51d1",
          5763 => x"973f81de",
          5764 => x"c008802e",
          5765 => x"fed23881",
          5766 => x"dec0081b",
          5767 => x"7c892a5a",
          5768 => x"5778802e",
          5769 => x"80d53878",
          5770 => x"1b7f8a11",
          5771 => x"22585b55",
          5772 => x"75752785",
          5773 => x"38757b31",
          5774 => x"59785476",
          5775 => x"537c5281",
          5776 => x"1a3351c8",
          5777 => x"be3f81de",
          5778 => x"c008fea6",
          5779 => x"387eb011",
          5780 => x"08783156",
          5781 => x"56747927",
          5782 => x"9b388480",
          5783 => x"53b01608",
          5784 => x"7731892b",
          5785 => x"7d0552b4",
          5786 => x"1651ccb5",
          5787 => x"3f7e5580",
          5788 => x"0b831634",
          5789 => x"78892b56",
          5790 => x"80db398c",
          5791 => x"18089419",
          5792 => x"08269338",
          5793 => x"7e51cdb6",
          5794 => x"3f81dec0",
          5795 => x"08fde338",
          5796 => x"7e77b012",
          5797 => x"0c55769c",
          5798 => x"190c9418",
          5799 => x"0883ff06",
          5800 => x"84807131",
          5801 => x"57557b76",
          5802 => x"2783387b",
          5803 => x"569c1808",
          5804 => x"527e51cd",
          5805 => x"f93f81de",
          5806 => x"c008fdb6",
          5807 => x"3875537c",
          5808 => x"52941808",
          5809 => x"83ff061f",
          5810 => x"b40551cb",
          5811 => x"d43f7e55",
          5812 => x"810b8316",
          5813 => x"347b7631",
          5814 => x"7e08177f",
          5815 => x"0c761e94",
          5816 => x"1a081870",
          5817 => x"941c0c8c",
          5818 => x"1b085858",
          5819 => x"5e5c7476",
          5820 => x"27833875",
          5821 => x"55748c19",
          5822 => x"0cfd9039",
          5823 => x"90183380",
          5824 => x"c0075574",
          5825 => x"90193480",
          5826 => x"567581de",
          5827 => x"c00c903d",
          5828 => x"0d04f83d",
          5829 => x"0d7a8b3d",
          5830 => x"fc055370",
          5831 => x"5256f2ea",
          5832 => x"3f81dec0",
          5833 => x"085781de",
          5834 => x"c00880fb",
          5835 => x"38901633",
          5836 => x"70862a70",
          5837 => x"81065155",
          5838 => x"5573802e",
          5839 => x"80e938a0",
          5840 => x"16085278",
          5841 => x"51cce73f",
          5842 => x"81dec008",
          5843 => x"5781dec0",
          5844 => x"0880d438",
          5845 => x"a416088b",
          5846 => x"1133a007",
          5847 => x"5555738b",
          5848 => x"16348816",
          5849 => x"08537452",
          5850 => x"750851dd",
          5851 => x"e83f8c16",
          5852 => x"08529c15",
          5853 => x"51c9fb3f",
          5854 => x"8288b20a",
          5855 => x"52961551",
          5856 => x"c9f03f76",
          5857 => x"52921551",
          5858 => x"c9ca3f78",
          5859 => x"54810b83",
          5860 => x"15347851",
          5861 => x"ccdf3f81",
          5862 => x"dec00890",
          5863 => x"173381bf",
          5864 => x"06555773",
          5865 => x"90173476",
          5866 => x"81dec00c",
          5867 => x"8a3d0d04",
          5868 => x"fc3d0d76",
          5869 => x"705254fe",
          5870 => x"d93f81de",
          5871 => x"c0085381",
          5872 => x"dec0089c",
          5873 => x"38863dfc",
          5874 => x"05527351",
          5875 => x"f1bc3f81",
          5876 => x"dec00853",
          5877 => x"81dec008",
          5878 => x"873881de",
          5879 => x"c008740c",
          5880 => x"7281dec0",
          5881 => x"0c863d0d",
          5882 => x"04ff3d0d",
          5883 => x"843d51e6",
          5884 => x"e43f8b52",
          5885 => x"800b81de",
          5886 => x"c008248b",
          5887 => x"3881dec0",
          5888 => x"0881def0",
          5889 => x"34805271",
          5890 => x"81dec00c",
          5891 => x"833d0d04",
          5892 => x"ef3d0d80",
          5893 => x"53933dd0",
          5894 => x"0552943d",
          5895 => x"51e9c13f",
          5896 => x"81dec008",
          5897 => x"5581dec0",
          5898 => x"0880e038",
          5899 => x"76586352",
          5900 => x"933dd405",
          5901 => x"51e08d3f",
          5902 => x"81dec008",
          5903 => x"5581dec0",
          5904 => x"08bc3802",
          5905 => x"80c70533",
          5906 => x"70982b55",
          5907 => x"56738025",
          5908 => x"8938767a",
          5909 => x"94120c54",
          5910 => x"b23902a2",
          5911 => x"05337084",
          5912 => x"2a708106",
          5913 => x"51555673",
          5914 => x"802e9e38",
          5915 => x"767f5370",
          5916 => x"5254dba8",
          5917 => x"3f81dec0",
          5918 => x"0894150c",
          5919 => x"8e3981de",
          5920 => x"c008842e",
          5921 => x"09810683",
          5922 => x"38855574",
          5923 => x"81dec00c",
          5924 => x"933d0d04",
          5925 => x"e43d0d6f",
          5926 => x"6f5b5b80",
          5927 => x"7a348053",
          5928 => x"9e3dffb8",
          5929 => x"05529f3d",
          5930 => x"51e8b53f",
          5931 => x"81dec008",
          5932 => x"5781dec0",
          5933 => x"0882fc38",
          5934 => x"7b437a7c",
          5935 => x"94110847",
          5936 => x"55586454",
          5937 => x"73802e81",
          5938 => x"ed38a052",
          5939 => x"933d7052",
          5940 => x"55d5ea3f",
          5941 => x"81dec008",
          5942 => x"5781dec0",
          5943 => x"0882d438",
          5944 => x"68527b51",
          5945 => x"c9c83f81",
          5946 => x"dec00857",
          5947 => x"81dec008",
          5948 => x"82c13869",
          5949 => x"527b51da",
          5950 => x"a33f81de",
          5951 => x"c0084576",
          5952 => x"527451d5",
          5953 => x"b83f81de",
          5954 => x"c0085781",
          5955 => x"dec00882",
          5956 => x"a2388052",
          5957 => x"7451daeb",
          5958 => x"3f81dec0",
          5959 => x"085781de",
          5960 => x"c008a438",
          5961 => x"69527b51",
          5962 => x"d9f23f73",
          5963 => x"81dec008",
          5964 => x"2ea63876",
          5965 => x"527451d6",
          5966 => x"cf3f81de",
          5967 => x"c0085781",
          5968 => x"dec00880",
          5969 => x"2ecc3876",
          5970 => x"842e0981",
          5971 => x"06863882",
          5972 => x"5781e039",
          5973 => x"7681dc38",
          5974 => x"9e3dffbc",
          5975 => x"05527451",
          5976 => x"dcc93f76",
          5977 => x"903d7811",
          5978 => x"81113351",
          5979 => x"565a5673",
          5980 => x"802e9138",
          5981 => x"02b90555",
          5982 => x"81168116",
          5983 => x"70335656",
          5984 => x"5673f538",
          5985 => x"81165473",
          5986 => x"78268190",
          5987 => x"3875802e",
          5988 => x"99387816",
          5989 => x"810555ff",
          5990 => x"186f11ff",
          5991 => x"18ff1858",
          5992 => x"58555874",
          5993 => x"33743475",
          5994 => x"ee38ff18",
          5995 => x"6f115558",
          5996 => x"af7434fe",
          5997 => x"8d39777b",
          5998 => x"2e098106",
          5999 => x"8a38ff18",
          6000 => x"6f115558",
          6001 => x"af743480",
          6002 => x"0b81def0",
          6003 => x"33708429",
          6004 => x"81cda405",
          6005 => x"70087033",
          6006 => x"525c5656",
          6007 => x"5673762e",
          6008 => x"8d388116",
          6009 => x"701a7033",
          6010 => x"51555673",
          6011 => x"f5388216",
          6012 => x"54737826",
          6013 => x"a7388055",
          6014 => x"74762791",
          6015 => x"38741954",
          6016 => x"73337a70",
          6017 => x"81055c34",
          6018 => x"811555ec",
          6019 => x"39ba7a70",
          6020 => x"81055c34",
          6021 => x"74ff2e09",
          6022 => x"81068538",
          6023 => x"91579439",
          6024 => x"6e188119",
          6025 => x"59547333",
          6026 => x"7a708105",
          6027 => x"5c347a78",
          6028 => x"26ee3880",
          6029 => x"7a347681",
          6030 => x"dec00c9e",
          6031 => x"3d0d04f7",
          6032 => x"3d0d7b7d",
          6033 => x"8d3dfc05",
          6034 => x"54715357",
          6035 => x"55ecbb3f",
          6036 => x"81dec008",
          6037 => x"5381dec0",
          6038 => x"0882fa38",
          6039 => x"91153353",
          6040 => x"7282f238",
          6041 => x"8c150854",
          6042 => x"73762792",
          6043 => x"38901533",
          6044 => x"70812a70",
          6045 => x"81065154",
          6046 => x"57728338",
          6047 => x"73569415",
          6048 => x"08548070",
          6049 => x"94170c58",
          6050 => x"75782e82",
          6051 => x"9738798a",
          6052 => x"11227089",
          6053 => x"2b595153",
          6054 => x"73782eb7",
          6055 => x"387652ff",
          6056 => x"1651ff95",
          6057 => x"d23f81de",
          6058 => x"c008ff15",
          6059 => x"78547053",
          6060 => x"5553ff95",
          6061 => x"c23f81de",
          6062 => x"c0087326",
          6063 => x"96387630",
          6064 => x"70750670",
          6065 => x"94180c77",
          6066 => x"71319818",
          6067 => x"08575851",
          6068 => x"53b13988",
          6069 => x"15085473",
          6070 => x"a6387352",
          6071 => x"7451cdca",
          6072 => x"3f81dec0",
          6073 => x"085481de",
          6074 => x"c008812e",
          6075 => x"819a3881",
          6076 => x"dec008ff",
          6077 => x"2e819b38",
          6078 => x"81dec008",
          6079 => x"88160c73",
          6080 => x"98160c73",
          6081 => x"802e819c",
          6082 => x"38767627",
          6083 => x"80dc3875",
          6084 => x"77319416",
          6085 => x"08189417",
          6086 => x"0c901633",
          6087 => x"70812a70",
          6088 => x"81065155",
          6089 => x"5a567280",
          6090 => x"2e9a3873",
          6091 => x"527451cc",
          6092 => x"f93f81de",
          6093 => x"c0085481",
          6094 => x"dec00894",
          6095 => x"3881dec0",
          6096 => x"0856a739",
          6097 => x"73527451",
          6098 => x"c7843f81",
          6099 => x"dec00854",
          6100 => x"73ff2ebe",
          6101 => x"38817427",
          6102 => x"af387953",
          6103 => x"73981408",
          6104 => x"27a63873",
          6105 => x"98160cff",
          6106 => x"a0399415",
          6107 => x"08169416",
          6108 => x"0c7583ff",
          6109 => x"06537280",
          6110 => x"2eaa3873",
          6111 => x"527951c6",
          6112 => x"a33f81de",
          6113 => x"c0089438",
          6114 => x"820b9116",
          6115 => x"34825380",
          6116 => x"c439810b",
          6117 => x"91163481",
          6118 => x"53bb3975",
          6119 => x"892a81de",
          6120 => x"c0080558",
          6121 => x"94150854",
          6122 => x"8c150874",
          6123 => x"27903873",
          6124 => x"8c160c90",
          6125 => x"153380c0",
          6126 => x"07537290",
          6127 => x"16347383",
          6128 => x"ff065372",
          6129 => x"802e8c38",
          6130 => x"779c1608",
          6131 => x"2e853877",
          6132 => x"9c160c80",
          6133 => x"537281de",
          6134 => x"c00c8b3d",
          6135 => x"0d04f93d",
          6136 => x"0d795689",
          6137 => x"5475802e",
          6138 => x"818a3880",
          6139 => x"53893dfc",
          6140 => x"05528a3d",
          6141 => x"840551e1",
          6142 => x"e73f81de",
          6143 => x"c0085581",
          6144 => x"dec00880",
          6145 => x"ea387776",
          6146 => x"0c7a5275",
          6147 => x"51d8b53f",
          6148 => x"81dec008",
          6149 => x"5581dec0",
          6150 => x"0880c338",
          6151 => x"ab163370",
          6152 => x"982b5557",
          6153 => x"807424a2",
          6154 => x"38861633",
          6155 => x"70842a70",
          6156 => x"81065155",
          6157 => x"5773802e",
          6158 => x"ad389c16",
          6159 => x"08527751",
          6160 => x"d3da3f81",
          6161 => x"dec00888",
          6162 => x"170c7754",
          6163 => x"86142284",
          6164 => x"17237452",
          6165 => x"7551cee5",
          6166 => x"3f81dec0",
          6167 => x"08557484",
          6168 => x"2e098106",
          6169 => x"85388555",
          6170 => x"86397480",
          6171 => x"2e843880",
          6172 => x"760c7454",
          6173 => x"7381dec0",
          6174 => x"0c893d0d",
          6175 => x"04fc3d0d",
          6176 => x"76873dfc",
          6177 => x"05537052",
          6178 => x"53e7ff3f",
          6179 => x"81dec008",
          6180 => x"873881de",
          6181 => x"c008730c",
          6182 => x"863d0d04",
          6183 => x"fb3d0d77",
          6184 => x"79893dfc",
          6185 => x"05547153",
          6186 => x"5654e7de",
          6187 => x"3f81dec0",
          6188 => x"085381de",
          6189 => x"c00880df",
          6190 => x"38749338",
          6191 => x"81dec008",
          6192 => x"527351cd",
          6193 => x"f83f81de",
          6194 => x"c0085380",
          6195 => x"ca3981de",
          6196 => x"c0085273",
          6197 => x"51d3ac3f",
          6198 => x"81dec008",
          6199 => x"5381dec0",
          6200 => x"08842e09",
          6201 => x"81068538",
          6202 => x"80538739",
          6203 => x"81dec008",
          6204 => x"a6387452",
          6205 => x"7351d5b3",
          6206 => x"3f725273",
          6207 => x"51cf893f",
          6208 => x"81dec008",
          6209 => x"84327030",
          6210 => x"7072079f",
          6211 => x"2c7081de",
          6212 => x"c0080651",
          6213 => x"51545472",
          6214 => x"81dec00c",
          6215 => x"873d0d04",
          6216 => x"ee3d0d65",
          6217 => x"57805389",
          6218 => x"3d705396",
          6219 => x"3d5256df",
          6220 => x"af3f81de",
          6221 => x"c0085581",
          6222 => x"dec008b2",
          6223 => x"38645275",
          6224 => x"51d6813f",
          6225 => x"81dec008",
          6226 => x"5581dec0",
          6227 => x"08a03802",
          6228 => x"80cb0533",
          6229 => x"70982b55",
          6230 => x"58738025",
          6231 => x"85388655",
          6232 => x"8d397680",
          6233 => x"2e883876",
          6234 => x"527551d4",
          6235 => x"be3f7481",
          6236 => x"dec00c94",
          6237 => x"3d0d04f0",
          6238 => x"3d0d6365",
          6239 => x"555c8053",
          6240 => x"923dec05",
          6241 => x"52933d51",
          6242 => x"ded63f81",
          6243 => x"dec0085b",
          6244 => x"81dec008",
          6245 => x"8280387c",
          6246 => x"740c7308",
          6247 => x"981108fe",
          6248 => x"11901308",
          6249 => x"59565855",
          6250 => x"75742691",
          6251 => x"38757c0c",
          6252 => x"81e43981",
          6253 => x"5b81cc39",
          6254 => x"825b81c7",
          6255 => x"3981dec0",
          6256 => x"08753355",
          6257 => x"5973812e",
          6258 => x"098106bf",
          6259 => x"3882755f",
          6260 => x"57765292",
          6261 => x"3df00551",
          6262 => x"c1f43f81",
          6263 => x"dec008ff",
          6264 => x"2ed13881",
          6265 => x"dec00881",
          6266 => x"2ece3881",
          6267 => x"dec00830",
          6268 => x"7081dec0",
          6269 => x"08078025",
          6270 => x"7a058119",
          6271 => x"7f53595a",
          6272 => x"54981408",
          6273 => x"7726ca38",
          6274 => x"80f939a4",
          6275 => x"150881de",
          6276 => x"c0085758",
          6277 => x"75983877",
          6278 => x"5281187d",
          6279 => x"5258ffbf",
          6280 => x"8d3f81de",
          6281 => x"c0085b81",
          6282 => x"dec00880",
          6283 => x"d6387c70",
          6284 => x"337712ff",
          6285 => x"1a5d5256",
          6286 => x"5474822e",
          6287 => x"0981069e",
          6288 => x"38b41451",
          6289 => x"ffbbcb3f",
          6290 => x"81dec008",
          6291 => x"83ffff06",
          6292 => x"70307080",
          6293 => x"251b8219",
          6294 => x"595b5154",
          6295 => x"9b39b414",
          6296 => x"51ffbbc5",
          6297 => x"3f81dec0",
          6298 => x"08f00a06",
          6299 => x"70307080",
          6300 => x"251b8419",
          6301 => x"595b5154",
          6302 => x"7583ff06",
          6303 => x"7a585679",
          6304 => x"ff923878",
          6305 => x"7c0c7c79",
          6306 => x"90120c84",
          6307 => x"11338107",
          6308 => x"56547484",
          6309 => x"15347a81",
          6310 => x"dec00c92",
          6311 => x"3d0d04f9",
          6312 => x"3d0d798a",
          6313 => x"3dfc0553",
          6314 => x"705257e3",
          6315 => x"dd3f81de",
          6316 => x"c0085681",
          6317 => x"dec00881",
          6318 => x"a8389117",
          6319 => x"33567581",
          6320 => x"a0389017",
          6321 => x"3370812a",
          6322 => x"70810651",
          6323 => x"55558755",
          6324 => x"73802e81",
          6325 => x"8e389417",
          6326 => x"0854738c",
          6327 => x"18082781",
          6328 => x"8038739b",
          6329 => x"3881dec0",
          6330 => x"08538817",
          6331 => x"08527651",
          6332 => x"c48c3f81",
          6333 => x"dec00874",
          6334 => x"88190c56",
          6335 => x"80c93998",
          6336 => x"17085276",
          6337 => x"51ffbfc6",
          6338 => x"3f81dec0",
          6339 => x"08ff2e09",
          6340 => x"81068338",
          6341 => x"815681de",
          6342 => x"c008812e",
          6343 => x"09810685",
          6344 => x"388256a3",
          6345 => x"3975a038",
          6346 => x"775481de",
          6347 => x"c0089815",
          6348 => x"08279438",
          6349 => x"98170853",
          6350 => x"81dec008",
          6351 => x"527651c3",
          6352 => x"bd3f81de",
          6353 => x"c0085694",
          6354 => x"17088c18",
          6355 => x"0c901733",
          6356 => x"80c00754",
          6357 => x"73901834",
          6358 => x"75802e85",
          6359 => x"38759118",
          6360 => x"34755574",
          6361 => x"81dec00c",
          6362 => x"893d0d04",
          6363 => x"e23d0d82",
          6364 => x"53a03dff",
          6365 => x"a40552a1",
          6366 => x"3d51dae4",
          6367 => x"3f81dec0",
          6368 => x"085581de",
          6369 => x"c00881f5",
          6370 => x"387845a1",
          6371 => x"3d085295",
          6372 => x"3d705258",
          6373 => x"d1ae3f81",
          6374 => x"dec00855",
          6375 => x"81dec008",
          6376 => x"81db3802",
          6377 => x"80fb0533",
          6378 => x"70852a70",
          6379 => x"81065155",
          6380 => x"56865573",
          6381 => x"81c73875",
          6382 => x"982b5480",
          6383 => x"742481bd",
          6384 => x"380280d6",
          6385 => x"05337081",
          6386 => x"06585487",
          6387 => x"557681ad",
          6388 => x"386b5278",
          6389 => x"51ccc53f",
          6390 => x"81dec008",
          6391 => x"74842a70",
          6392 => x"81065155",
          6393 => x"5673802e",
          6394 => x"80d43878",
          6395 => x"5481dec0",
          6396 => x"08941508",
          6397 => x"2e818638",
          6398 => x"735a81de",
          6399 => x"c0085c76",
          6400 => x"528a3d70",
          6401 => x"5254c7b5",
          6402 => x"3f81dec0",
          6403 => x"085581de",
          6404 => x"c00880e9",
          6405 => x"3881dec0",
          6406 => x"08527351",
          6407 => x"cce53f81",
          6408 => x"dec00855",
          6409 => x"81dec008",
          6410 => x"86388755",
          6411 => x"80cf3981",
          6412 => x"dec00884",
          6413 => x"2e883881",
          6414 => x"dec00880",
          6415 => x"c0387751",
          6416 => x"cec23f81",
          6417 => x"dec00881",
          6418 => x"dec00830",
          6419 => x"7081dec0",
          6420 => x"08078025",
          6421 => x"51555575",
          6422 => x"802e9438",
          6423 => x"73802e8f",
          6424 => x"38805375",
          6425 => x"527751c1",
          6426 => x"953f81de",
          6427 => x"c0085574",
          6428 => x"8c387851",
          6429 => x"ffbafe3f",
          6430 => x"81dec008",
          6431 => x"557481de",
          6432 => x"c00ca03d",
          6433 => x"0d04e93d",
          6434 => x"0d825399",
          6435 => x"3dc00552",
          6436 => x"9a3d51d8",
          6437 => x"cb3f81de",
          6438 => x"c0085481",
          6439 => x"dec00882",
          6440 => x"b038785e",
          6441 => x"69528e3d",
          6442 => x"705258cf",
          6443 => x"973f81de",
          6444 => x"c0085481",
          6445 => x"dec00886",
          6446 => x"38885482",
          6447 => x"943981de",
          6448 => x"c008842e",
          6449 => x"09810682",
          6450 => x"88380280",
          6451 => x"df053370",
          6452 => x"852a8106",
          6453 => x"51558654",
          6454 => x"7481f638",
          6455 => x"785a7452",
          6456 => x"8a3d7052",
          6457 => x"57c1c33f",
          6458 => x"81dec008",
          6459 => x"75555681",
          6460 => x"dec00883",
          6461 => x"38875481",
          6462 => x"dec00881",
          6463 => x"2e098106",
          6464 => x"83388254",
          6465 => x"81dec008",
          6466 => x"ff2e0981",
          6467 => x"06863881",
          6468 => x"5481b439",
          6469 => x"7381b038",
          6470 => x"81dec008",
          6471 => x"527851c4",
          6472 => x"a43f81de",
          6473 => x"c0085481",
          6474 => x"dec00881",
          6475 => x"9a388b53",
          6476 => x"a052b419",
          6477 => x"51ffb78c",
          6478 => x"3f7854ae",
          6479 => x"0bb41534",
          6480 => x"7854900b",
          6481 => x"bf153482",
          6482 => x"88b20a52",
          6483 => x"80ca1951",
          6484 => x"ffb69f3f",
          6485 => x"755378b4",
          6486 => x"115351c9",
          6487 => x"f83fa053",
          6488 => x"78b41153",
          6489 => x"80d40551",
          6490 => x"ffb6b63f",
          6491 => x"7854ae0b",
          6492 => x"80d51534",
          6493 => x"7f537880",
          6494 => x"d4115351",
          6495 => x"c9d73f78",
          6496 => x"54810b83",
          6497 => x"15347751",
          6498 => x"cba43f81",
          6499 => x"dec00854",
          6500 => x"81dec008",
          6501 => x"b2388288",
          6502 => x"b20a5264",
          6503 => x"960551ff",
          6504 => x"b5d03f75",
          6505 => x"53645278",
          6506 => x"51c9aa3f",
          6507 => x"6454900b",
          6508 => x"8b153478",
          6509 => x"54810b83",
          6510 => x"15347851",
          6511 => x"ffb8b63f",
          6512 => x"81dec008",
          6513 => x"548b3980",
          6514 => x"53755276",
          6515 => x"51ffbeae",
          6516 => x"3f7381de",
          6517 => x"c00c993d",
          6518 => x"0d04da3d",
          6519 => x"0da93d84",
          6520 => x"0551d2f1",
          6521 => x"3f8253a8",
          6522 => x"3dff8405",
          6523 => x"52a93d51",
          6524 => x"d5ee3f81",
          6525 => x"dec00855",
          6526 => x"81dec008",
          6527 => x"82d33878",
          6528 => x"4da93d08",
          6529 => x"529d3d70",
          6530 => x"5258ccb8",
          6531 => x"3f81dec0",
          6532 => x"085581de",
          6533 => x"c00882b9",
          6534 => x"3802819b",
          6535 => x"053381a0",
          6536 => x"06548655",
          6537 => x"7382aa38",
          6538 => x"a053a43d",
          6539 => x"0852a83d",
          6540 => x"ff880551",
          6541 => x"ffb4ea3f",
          6542 => x"ac537752",
          6543 => x"923d7052",
          6544 => x"54ffb4dd",
          6545 => x"3faa3d08",
          6546 => x"527351cb",
          6547 => x"f73f81de",
          6548 => x"c0085581",
          6549 => x"dec00895",
          6550 => x"38636f2e",
          6551 => x"09810688",
          6552 => x"3865a23d",
          6553 => x"082e9238",
          6554 => x"885581e5",
          6555 => x"3981dec0",
          6556 => x"08842e09",
          6557 => x"810681b8",
          6558 => x"387351c9",
          6559 => x"b13f81de",
          6560 => x"c0085581",
          6561 => x"dec00881",
          6562 => x"c8386856",
          6563 => x"9353a83d",
          6564 => x"ff950552",
          6565 => x"8d1651ff",
          6566 => x"b4873f02",
          6567 => x"af05338b",
          6568 => x"17348b16",
          6569 => x"3370842a",
          6570 => x"70810651",
          6571 => x"55557389",
          6572 => x"3874a007",
          6573 => x"54738b17",
          6574 => x"34785481",
          6575 => x"0b831534",
          6576 => x"8b163370",
          6577 => x"842a7081",
          6578 => x"06515555",
          6579 => x"73802e80",
          6580 => x"e5386e64",
          6581 => x"2e80df38",
          6582 => x"75527851",
          6583 => x"c6be3f81",
          6584 => x"dec00852",
          6585 => x"7851ffb7",
          6586 => x"bb3f8255",
          6587 => x"81dec008",
          6588 => x"802e80dd",
          6589 => x"3881dec0",
          6590 => x"08527851",
          6591 => x"ffb5af3f",
          6592 => x"81dec008",
          6593 => x"7980d411",
          6594 => x"58585581",
          6595 => x"dec00880",
          6596 => x"c0388116",
          6597 => x"335473ae",
          6598 => x"2e098106",
          6599 => x"99386353",
          6600 => x"75527651",
          6601 => x"c6af3f78",
          6602 => x"54810b83",
          6603 => x"15348739",
          6604 => x"81dec008",
          6605 => x"9c387751",
          6606 => x"c8ca3f81",
          6607 => x"dec00855",
          6608 => x"81dec008",
          6609 => x"8c387851",
          6610 => x"ffb5aa3f",
          6611 => x"81dec008",
          6612 => x"557481de",
          6613 => x"c00ca83d",
          6614 => x"0d04ed3d",
          6615 => x"0d0280db",
          6616 => x"05330284",
          6617 => x"0580df05",
          6618 => x"33575782",
          6619 => x"53953dd0",
          6620 => x"0552963d",
          6621 => x"51d2e93f",
          6622 => x"81dec008",
          6623 => x"5581dec0",
          6624 => x"0880cf38",
          6625 => x"785a6552",
          6626 => x"953dd405",
          6627 => x"51c9b53f",
          6628 => x"81dec008",
          6629 => x"5581dec0",
          6630 => x"08b83802",
          6631 => x"80cf0533",
          6632 => x"81a00654",
          6633 => x"865573aa",
          6634 => x"3875a706",
          6635 => x"6171098b",
          6636 => x"12337106",
          6637 => x"7a740607",
          6638 => x"51575556",
          6639 => x"748b1534",
          6640 => x"7854810b",
          6641 => x"83153478",
          6642 => x"51ffb4a9",
          6643 => x"3f81dec0",
          6644 => x"08557481",
          6645 => x"dec00c95",
          6646 => x"3d0d04ef",
          6647 => x"3d0d6456",
          6648 => x"8253933d",
          6649 => x"d0055294",
          6650 => x"3d51d1f4",
          6651 => x"3f81dec0",
          6652 => x"085581de",
          6653 => x"c00880cb",
          6654 => x"38765863",
          6655 => x"52933dd4",
          6656 => x"0551c8c0",
          6657 => x"3f81dec0",
          6658 => x"085581de",
          6659 => x"c008b438",
          6660 => x"0280c705",
          6661 => x"3381a006",
          6662 => x"54865573",
          6663 => x"a6388416",
          6664 => x"22861722",
          6665 => x"71902b07",
          6666 => x"5354961f",
          6667 => x"51ffb0c2",
          6668 => x"3f765481",
          6669 => x"0b831534",
          6670 => x"7651ffb3",
          6671 => x"b83f81de",
          6672 => x"c0085574",
          6673 => x"81dec00c",
          6674 => x"933d0d04",
          6675 => x"ea3d0d69",
          6676 => x"6b5c5a80",
          6677 => x"53983dd0",
          6678 => x"0552993d",
          6679 => x"51d1813f",
          6680 => x"81dec008",
          6681 => x"81dec008",
          6682 => x"307081de",
          6683 => x"c0080780",
          6684 => x"25515557",
          6685 => x"79802e81",
          6686 => x"85388170",
          6687 => x"75065555",
          6688 => x"73802e80",
          6689 => x"f9387b5d",
          6690 => x"805f8052",
          6691 => x"8d3d7052",
          6692 => x"54ffbea9",
          6693 => x"3f81dec0",
          6694 => x"085781de",
          6695 => x"c00880d1",
          6696 => x"38745273",
          6697 => x"51c3dc3f",
          6698 => x"81dec008",
          6699 => x"5781dec0",
          6700 => x"08bf3881",
          6701 => x"dec00881",
          6702 => x"dec00865",
          6703 => x"5b595678",
          6704 => x"1881197b",
          6705 => x"18565955",
          6706 => x"74337434",
          6707 => x"8116568a",
          6708 => x"7827ec38",
          6709 => x"8b56751a",
          6710 => x"54807434",
          6711 => x"75802e9e",
          6712 => x"38ff1670",
          6713 => x"1b703351",
          6714 => x"555673a0",
          6715 => x"2ee8388e",
          6716 => x"3976842e",
          6717 => x"09810686",
          6718 => x"38807a34",
          6719 => x"80577630",
          6720 => x"70780780",
          6721 => x"2551547a",
          6722 => x"802e80c1",
          6723 => x"3873802e",
          6724 => x"bc387ba0",
          6725 => x"11085351",
          6726 => x"ffb1933f",
          6727 => x"81dec008",
          6728 => x"5781dec0",
          6729 => x"08a7387b",
          6730 => x"70335555",
          6731 => x"80c35673",
          6732 => x"832e8b38",
          6733 => x"80e45673",
          6734 => x"842e8338",
          6735 => x"a7567515",
          6736 => x"b40551ff",
          6737 => x"ade33f81",
          6738 => x"dec0087b",
          6739 => x"0c7681de",
          6740 => x"c00c983d",
          6741 => x"0d04e63d",
          6742 => x"0d82539c",
          6743 => x"3dffb805",
          6744 => x"529d3d51",
          6745 => x"cefa3f81",
          6746 => x"dec00881",
          6747 => x"dec00856",
          6748 => x"5481dec0",
          6749 => x"08839838",
          6750 => x"8b53a052",
          6751 => x"8b3d7052",
          6752 => x"59ffaec0",
          6753 => x"3f736d70",
          6754 => x"337081ff",
          6755 => x"06525755",
          6756 => x"579f7427",
          6757 => x"81bc3878",
          6758 => x"587481ff",
          6759 => x"066d8105",
          6760 => x"4e705255",
          6761 => x"ffaf893f",
          6762 => x"81dec008",
          6763 => x"802ea538",
          6764 => x"6c703370",
          6765 => x"535754ff",
          6766 => x"aefd3f81",
          6767 => x"dec00880",
          6768 => x"2e8d3874",
          6769 => x"882b7607",
          6770 => x"6d81054e",
          6771 => x"55863981",
          6772 => x"dec00855",
          6773 => x"ff9f1570",
          6774 => x"83ffff06",
          6775 => x"51547399",
          6776 => x"268a38e0",
          6777 => x"157083ff",
          6778 => x"ff065654",
          6779 => x"80ff7527",
          6780 => x"873881cc",
          6781 => x"b4153355",
          6782 => x"74802ea3",
          6783 => x"38745281",
          6784 => x"ceb451ff",
          6785 => x"ae893f81",
          6786 => x"dec00893",
          6787 => x"3881ff75",
          6788 => x"27883876",
          6789 => x"89268838",
          6790 => x"8b398a77",
          6791 => x"27863886",
          6792 => x"5581ec39",
          6793 => x"81ff7527",
          6794 => x"8f387488",
          6795 => x"2a547378",
          6796 => x"7081055a",
          6797 => x"34811757",
          6798 => x"74787081",
          6799 => x"055a3481",
          6800 => x"176d7033",
          6801 => x"7081ff06",
          6802 => x"52575557",
          6803 => x"739f26fe",
          6804 => x"c8388b3d",
          6805 => x"33548655",
          6806 => x"7381e52e",
          6807 => x"81b13876",
          6808 => x"802e9938",
          6809 => x"02a70555",
          6810 => x"76157033",
          6811 => x"515473a0",
          6812 => x"2e098106",
          6813 => x"8738ff17",
          6814 => x"5776ed38",
          6815 => x"79418043",
          6816 => x"8052913d",
          6817 => x"705255ff",
          6818 => x"bab33f81",
          6819 => x"dec00854",
          6820 => x"81dec008",
          6821 => x"80f73881",
          6822 => x"527451ff",
          6823 => x"bfe53f81",
          6824 => x"dec00854",
          6825 => x"81dec008",
          6826 => x"8d387680",
          6827 => x"c4386754",
          6828 => x"e5743480",
          6829 => x"c63981de",
          6830 => x"c008842e",
          6831 => x"09810680",
          6832 => x"cc388054",
          6833 => x"76742e80",
          6834 => x"c4388152",
          6835 => x"7451ffbd",
          6836 => x"b03f81de",
          6837 => x"c0085481",
          6838 => x"dec008b1",
          6839 => x"38a05381",
          6840 => x"dec00852",
          6841 => x"6751ffab",
          6842 => x"db3f6754",
          6843 => x"880b8b15",
          6844 => x"348b5378",
          6845 => x"526751ff",
          6846 => x"aba73f79",
          6847 => x"54810b83",
          6848 => x"15347951",
          6849 => x"ffadee3f",
          6850 => x"81dec008",
          6851 => x"54735574",
          6852 => x"81dec00c",
          6853 => x"9c3d0d04",
          6854 => x"f23d0d60",
          6855 => x"62028805",
          6856 => x"80cb0533",
          6857 => x"933dfc05",
          6858 => x"55725440",
          6859 => x"5e5ad2da",
          6860 => x"3f81dec0",
          6861 => x"085881de",
          6862 => x"c00882bd",
          6863 => x"38911a33",
          6864 => x"587782b5",
          6865 => x"387c802e",
          6866 => x"97388c1a",
          6867 => x"08597890",
          6868 => x"38901a33",
          6869 => x"70812a70",
          6870 => x"81065155",
          6871 => x"55739038",
          6872 => x"87548297",
          6873 => x"39825882",
          6874 => x"90398158",
          6875 => x"828b397e",
          6876 => x"8a112270",
          6877 => x"892b7055",
          6878 => x"7f545656",
          6879 => x"56fefbf7",
          6880 => x"3fff147d",
          6881 => x"06703070",
          6882 => x"72079f2a",
          6883 => x"81dec008",
          6884 => x"058c1908",
          6885 => x"7c405a5d",
          6886 => x"55558177",
          6887 => x"27883898",
          6888 => x"16087726",
          6889 => x"83388257",
          6890 => x"76775659",
          6891 => x"80567452",
          6892 => x"7951ffae",
          6893 => x"993f8115",
          6894 => x"7f555598",
          6895 => x"14087526",
          6896 => x"83388255",
          6897 => x"81dec008",
          6898 => x"812eff99",
          6899 => x"3881dec0",
          6900 => x"08ff2eff",
          6901 => x"953881de",
          6902 => x"c0088e38",
          6903 => x"81165675",
          6904 => x"7b2e0981",
          6905 => x"06873893",
          6906 => x"39745980",
          6907 => x"5674772e",
          6908 => x"098106ff",
          6909 => x"b9388758",
          6910 => x"80ff397d",
          6911 => x"802eba38",
          6912 => x"787b5555",
          6913 => x"7a802eb4",
          6914 => x"38811556",
          6915 => x"73812e09",
          6916 => x"81068338",
          6917 => x"ff567553",
          6918 => x"74527e51",
          6919 => x"ffafa83f",
          6920 => x"81dec008",
          6921 => x"5881dec0",
          6922 => x"0880ce38",
          6923 => x"748116ff",
          6924 => x"1656565c",
          6925 => x"73d33884",
          6926 => x"39ff195c",
          6927 => x"7e7c8c12",
          6928 => x"0c557d80",
          6929 => x"2eb33878",
          6930 => x"881b0c7c",
          6931 => x"8c1b0c90",
          6932 => x"1a3380c0",
          6933 => x"07547390",
          6934 => x"1b349815",
          6935 => x"08fe0590",
          6936 => x"16085754",
          6937 => x"75742691",
          6938 => x"38757b31",
          6939 => x"90160c84",
          6940 => x"15338107",
          6941 => x"54738416",
          6942 => x"34775473",
          6943 => x"81dec00c",
          6944 => x"903d0d04",
          6945 => x"e93d0d6b",
          6946 => x"6d028805",
          6947 => x"80eb0533",
          6948 => x"9d3d545a",
          6949 => x"5c59c5bd",
          6950 => x"3f8b5680",
          6951 => x"0b81dec0",
          6952 => x"08248bf8",
          6953 => x"3881dec0",
          6954 => x"08842981",
          6955 => x"dedc0570",
          6956 => x"08515574",
          6957 => x"802e8438",
          6958 => x"80753481",
          6959 => x"dec00881",
          6960 => x"ff065f81",
          6961 => x"527e51ff",
          6962 => x"a0d03f81",
          6963 => x"dec00881",
          6964 => x"ff067081",
          6965 => x"06565783",
          6966 => x"56748bc0",
          6967 => x"3876822a",
          6968 => x"70810651",
          6969 => x"558a5674",
          6970 => x"8bb23899",
          6971 => x"3dfc0553",
          6972 => x"83527e51",
          6973 => x"ffa4f03f",
          6974 => x"81dec008",
          6975 => x"99386755",
          6976 => x"74802e92",
          6977 => x"38748280",
          6978 => x"80268b38",
          6979 => x"ff157506",
          6980 => x"5574802e",
          6981 => x"83388148",
          6982 => x"78802e87",
          6983 => x"38848079",
          6984 => x"26923878",
          6985 => x"81800a26",
          6986 => x"8b38ff19",
          6987 => x"79065574",
          6988 => x"802e8638",
          6989 => x"93568ae4",
          6990 => x"3978892a",
          6991 => x"6e892a70",
          6992 => x"892b7759",
          6993 => x"4843597a",
          6994 => x"83388156",
          6995 => x"61307080",
          6996 => x"25770751",
          6997 => x"55915674",
          6998 => x"8ac23899",
          6999 => x"3df80553",
          7000 => x"81527e51",
          7001 => x"ffa4803f",
          7002 => x"815681de",
          7003 => x"c0088aac",
          7004 => x"3877832a",
          7005 => x"70770681",
          7006 => x"dec00843",
          7007 => x"56457483",
          7008 => x"38bf4166",
          7009 => x"558e5660",
          7010 => x"75268a90",
          7011 => x"38746131",
          7012 => x"70485580",
          7013 => x"ff75278a",
          7014 => x"83389356",
          7015 => x"78818026",
          7016 => x"89fa3877",
          7017 => x"812a7081",
          7018 => x"06564374",
          7019 => x"802e9538",
          7020 => x"77870655",
          7021 => x"74822e83",
          7022 => x"8d387781",
          7023 => x"06557480",
          7024 => x"2e838338",
          7025 => x"77810655",
          7026 => x"9356825e",
          7027 => x"74802e89",
          7028 => x"cb38785a",
          7029 => x"7d832e09",
          7030 => x"810680e1",
          7031 => x"3878ae38",
          7032 => x"66912a57",
          7033 => x"810b81ce",
          7034 => x"d822565a",
          7035 => x"74802e9d",
          7036 => x"38747726",
          7037 => x"983881ce",
          7038 => x"d8567910",
          7039 => x"82177022",
          7040 => x"57575a74",
          7041 => x"802e8638",
          7042 => x"767527ee",
          7043 => x"38795266",
          7044 => x"51fef6e3",
          7045 => x"3f81dec0",
          7046 => x"08842984",
          7047 => x"87057089",
          7048 => x"2a5e55a0",
          7049 => x"5c800b81",
          7050 => x"dec008fc",
          7051 => x"808a0556",
          7052 => x"44fdfff0",
          7053 => x"0a752780",
          7054 => x"ec3888d3",
          7055 => x"3978ae38",
          7056 => x"668c2a57",
          7057 => x"810b81ce",
          7058 => x"c822565a",
          7059 => x"74802e9d",
          7060 => x"38747726",
          7061 => x"983881ce",
          7062 => x"c8567910",
          7063 => x"82177022",
          7064 => x"57575a74",
          7065 => x"802e8638",
          7066 => x"767527ee",
          7067 => x"38795266",
          7068 => x"51fef683",
          7069 => x"3f81dec0",
          7070 => x"08108405",
          7071 => x"5781dec0",
          7072 => x"089ff526",
          7073 => x"9638810b",
          7074 => x"81dec008",
          7075 => x"1081dec0",
          7076 => x"08057111",
          7077 => x"722a8305",
          7078 => x"59565e83",
          7079 => x"ff17892a",
          7080 => x"5d815ca0",
          7081 => x"44601c7d",
          7082 => x"11650569",
          7083 => x"7012ff05",
          7084 => x"71307072",
          7085 => x"0674315c",
          7086 => x"52595759",
          7087 => x"407d832e",
          7088 => x"09810689",
          7089 => x"38761c60",
          7090 => x"18415c84",
          7091 => x"39761d5d",
          7092 => x"79902918",
          7093 => x"70623168",
          7094 => x"58515574",
          7095 => x"762687af",
          7096 => x"38757c31",
          7097 => x"7d317a53",
          7098 => x"70653152",
          7099 => x"55fef587",
          7100 => x"3f81dec0",
          7101 => x"08587d83",
          7102 => x"2e098106",
          7103 => x"9b3881de",
          7104 => x"c00883ff",
          7105 => x"f52680dd",
          7106 => x"38788783",
          7107 => x"3879812a",
          7108 => x"5978fdbe",
          7109 => x"3886f839",
          7110 => x"7d822e09",
          7111 => x"810680c5",
          7112 => x"3883fff5",
          7113 => x"0b81dec0",
          7114 => x"0827a038",
          7115 => x"788f3879",
          7116 => x"1a557480",
          7117 => x"c0268638",
          7118 => x"7459fd96",
          7119 => x"39628106",
          7120 => x"5574802e",
          7121 => x"8f38835e",
          7122 => x"fd883981",
          7123 => x"dec0089f",
          7124 => x"f5269238",
          7125 => x"7886b838",
          7126 => x"791a5981",
          7127 => x"807927fc",
          7128 => x"f13886ab",
          7129 => x"3980557d",
          7130 => x"812e0981",
          7131 => x"0683387d",
          7132 => x"559ff578",
          7133 => x"278b3874",
          7134 => x"8106558e",
          7135 => x"5674869c",
          7136 => x"38848053",
          7137 => x"80527a51",
          7138 => x"ffa2b93f",
          7139 => x"8b5381cc",
          7140 => x"f0527a51",
          7141 => x"ffa28a3f",
          7142 => x"8480528b",
          7143 => x"1b51ffa1",
          7144 => x"b33f798d",
          7145 => x"1c347b83",
          7146 => x"ffff0652",
          7147 => x"8e1b51ff",
          7148 => x"a1a23f81",
          7149 => x"0b901c34",
          7150 => x"7d833270",
          7151 => x"3070962a",
          7152 => x"84800654",
          7153 => x"5155911b",
          7154 => x"51ffa188",
          7155 => x"3f665574",
          7156 => x"83ffff26",
          7157 => x"90387483",
          7158 => x"ffff0652",
          7159 => x"931b51ff",
          7160 => x"a0f23f8a",
          7161 => x"397452a0",
          7162 => x"1b51ffa1",
          7163 => x"853ff80b",
          7164 => x"951c34bf",
          7165 => x"52981b51",
          7166 => x"ffa0d93f",
          7167 => x"81ff529a",
          7168 => x"1b51ffa0",
          7169 => x"cf3f6052",
          7170 => x"9c1b51ff",
          7171 => x"a0e43f7d",
          7172 => x"832e0981",
          7173 => x"0680cb38",
          7174 => x"8288b20a",
          7175 => x"5280c31b",
          7176 => x"51ffa0ce",
          7177 => x"3f7c52a4",
          7178 => x"1b51ffa0",
          7179 => x"c53f8252",
          7180 => x"ac1b51ff",
          7181 => x"a0bc3f81",
          7182 => x"52b01b51",
          7183 => x"ffa0953f",
          7184 => x"8652b21b",
          7185 => x"51ffa08c",
          7186 => x"3fff800b",
          7187 => x"80c01c34",
          7188 => x"a90b80c2",
          7189 => x"1c349353",
          7190 => x"81ccfc52",
          7191 => x"80c71b51",
          7192 => x"ae398288",
          7193 => x"b20a52a7",
          7194 => x"1b51ffa0",
          7195 => x"853f7c83",
          7196 => x"ffff0652",
          7197 => x"961b51ff",
          7198 => x"9fda3fff",
          7199 => x"800ba41c",
          7200 => x"34a90ba6",
          7201 => x"1c349353",
          7202 => x"81cd9052",
          7203 => x"ab1b51ff",
          7204 => x"a08f3f82",
          7205 => x"d4d55283",
          7206 => x"fe1b7052",
          7207 => x"59ff9fb4",
          7208 => x"3f815460",
          7209 => x"537a527e",
          7210 => x"51ff9bd7",
          7211 => x"3f815681",
          7212 => x"dec00883",
          7213 => x"e7387d83",
          7214 => x"2e098106",
          7215 => x"80ee3875",
          7216 => x"54608605",
          7217 => x"537a527e",
          7218 => x"51ff9bb7",
          7219 => x"3f848053",
          7220 => x"80527a51",
          7221 => x"ff9fed3f",
          7222 => x"848b85a4",
          7223 => x"d2527a51",
          7224 => x"ff9f8f3f",
          7225 => x"868a85e4",
          7226 => x"f25283e4",
          7227 => x"1b51ff9f",
          7228 => x"813fff18",
          7229 => x"5283e81b",
          7230 => x"51ff9ef6",
          7231 => x"3f825283",
          7232 => x"ec1b51ff",
          7233 => x"9eec3f82",
          7234 => x"d4d55278",
          7235 => x"51ff9ec4",
          7236 => x"3f755460",
          7237 => x"8705537a",
          7238 => x"527e51ff",
          7239 => x"9ae53f75",
          7240 => x"54601653",
          7241 => x"7a527e51",
          7242 => x"ff9ad83f",
          7243 => x"65538052",
          7244 => x"7a51ff9f",
          7245 => x"8f3f7f56",
          7246 => x"80587d83",
          7247 => x"2e098106",
          7248 => x"9a38f852",
          7249 => x"7a51ff9e",
          7250 => x"a93fff52",
          7251 => x"841b51ff",
          7252 => x"9ea03ff0",
          7253 => x"0a52881b",
          7254 => x"51913987",
          7255 => x"fffff855",
          7256 => x"7d812e83",
          7257 => x"38f85574",
          7258 => x"527a51ff",
          7259 => x"9e843f7c",
          7260 => x"55615774",
          7261 => x"62268338",
          7262 => x"74577654",
          7263 => x"75537a52",
          7264 => x"7e51ff99",
          7265 => x"fe3f81de",
          7266 => x"c0088287",
          7267 => x"38848053",
          7268 => x"81dec008",
          7269 => x"527a51ff",
          7270 => x"9eaa3f76",
          7271 => x"16757831",
          7272 => x"565674cd",
          7273 => x"38811858",
          7274 => x"77802eff",
          7275 => x"8d387955",
          7276 => x"7d832e83",
          7277 => x"38635561",
          7278 => x"57746226",
          7279 => x"83387457",
          7280 => x"76547553",
          7281 => x"7a527e51",
          7282 => x"ff99b83f",
          7283 => x"81dec008",
          7284 => x"81c13876",
          7285 => x"16757831",
          7286 => x"565674db",
          7287 => x"388c567d",
          7288 => x"832e9338",
          7289 => x"86566683",
          7290 => x"ffff268a",
          7291 => x"3884567d",
          7292 => x"822e8338",
          7293 => x"81566481",
          7294 => x"06587780",
          7295 => x"fe388480",
          7296 => x"5377527a",
          7297 => x"51ff9dbc",
          7298 => x"3f82d4d5",
          7299 => x"527851ff",
          7300 => x"9cc23f83",
          7301 => x"be1b5577",
          7302 => x"7534810b",
          7303 => x"81163481",
          7304 => x"0b821634",
          7305 => x"77831634",
          7306 => x"75841634",
          7307 => x"60670556",
          7308 => x"80fdc152",
          7309 => x"7551feee",
          7310 => x"be3ffe0b",
          7311 => x"85163481",
          7312 => x"dec00882",
          7313 => x"2abf0756",
          7314 => x"75861634",
          7315 => x"81dec008",
          7316 => x"87163460",
          7317 => x"5283c61b",
          7318 => x"51ff9c96",
          7319 => x"3f665283",
          7320 => x"ca1b51ff",
          7321 => x"9c8c3f81",
          7322 => x"5477537a",
          7323 => x"527e51ff",
          7324 => x"98913f81",
          7325 => x"5681dec0",
          7326 => x"08a23880",
          7327 => x"5380527e",
          7328 => x"51ff99e3",
          7329 => x"3f815681",
          7330 => x"dec00890",
          7331 => x"3889398e",
          7332 => x"568a3981",
          7333 => x"56863981",
          7334 => x"dec00856",
          7335 => x"7581dec0",
          7336 => x"0c993d0d",
          7337 => x"04f53d0d",
          7338 => x"7d605b59",
          7339 => x"807960ff",
          7340 => x"055a5757",
          7341 => x"767825b4",
          7342 => x"388d3df8",
          7343 => x"11555581",
          7344 => x"53fc1552",
          7345 => x"7951c9dc",
          7346 => x"3f7a812e",
          7347 => x"0981069c",
          7348 => x"388c3d33",
          7349 => x"55748d2e",
          7350 => x"db387476",
          7351 => x"70810558",
          7352 => x"34811757",
          7353 => x"748a2e09",
          7354 => x"8106c938",
          7355 => x"80763478",
          7356 => x"55768338",
          7357 => x"76557481",
          7358 => x"dec00c8d",
          7359 => x"3d0d04ff",
          7360 => x"3d0d7352",
          7361 => x"71932681",
          7362 => x"8e387184",
          7363 => x"2981c694",
          7364 => x"05527108",
          7365 => x"0481cff0",
          7366 => x"51818039",
          7367 => x"81cffc51",
          7368 => x"80f93981",
          7369 => x"d0905180",
          7370 => x"f23981d0",
          7371 => x"a45180eb",
          7372 => x"3981d0b4",
          7373 => x"5180e439",
          7374 => x"81d0c451",
          7375 => x"80dd3981",
          7376 => x"d0d85180",
          7377 => x"d63981d0",
          7378 => x"e85180cf",
          7379 => x"3981d180",
          7380 => x"5180c839",
          7381 => x"81d19851",
          7382 => x"80c13981",
          7383 => x"d1b051bb",
          7384 => x"3981d1cc",
          7385 => x"51b53981",
          7386 => x"d1e051af",
          7387 => x"3981d28c",
          7388 => x"51a93981",
          7389 => x"d2a051a3",
          7390 => x"3981d2c0",
          7391 => x"519d3981",
          7392 => x"d2d45197",
          7393 => x"3981d2ec",
          7394 => x"51913981",
          7395 => x"d384518b",
          7396 => x"3981d39c",
          7397 => x"51853981",
          7398 => x"d3a851ff",
          7399 => x"87a13f83",
          7400 => x"3d0d04fb",
          7401 => x"3d0d7779",
          7402 => x"56567487",
          7403 => x"e7268a38",
          7404 => x"74527587",
          7405 => x"e8295191",
          7406 => x"3987e852",
          7407 => x"7451feeb",
          7408 => x"b63f81de",
          7409 => x"c0085275",
          7410 => x"51feebab",
          7411 => x"3f81dec0",
          7412 => x"08547953",
          7413 => x"755281d3",
          7414 => x"b851ff8c",
          7415 => x"c63f873d",
          7416 => x"0d04f53d",
          7417 => x"0d7d7f61",
          7418 => x"028c0580",
          7419 => x"c7053373",
          7420 => x"7315665f",
          7421 => x"5d5a5a5c",
          7422 => x"5c5c7852",
          7423 => x"81d3dc51",
          7424 => x"ff8ca03f",
          7425 => x"81d3e451",
          7426 => x"ff86b43f",
          7427 => x"80557477",
          7428 => x"2780fc38",
          7429 => x"79902e89",
          7430 => x"3879a02e",
          7431 => x"a73880c6",
          7432 => x"39741653",
          7433 => x"7278278e",
          7434 => x"38722252",
          7435 => x"81d3e851",
          7436 => x"ff8bf03f",
          7437 => x"893981d3",
          7438 => x"f451ff86",
          7439 => x"823f8215",
          7440 => x"5580c339",
          7441 => x"74165372",
          7442 => x"78278e38",
          7443 => x"72085281",
          7444 => x"d3dc51ff",
          7445 => x"8bcd3f89",
          7446 => x"3981d3f0",
          7447 => x"51ff85df",
          7448 => x"3f841555",
          7449 => x"a1397416",
          7450 => x"53727827",
          7451 => x"8e387233",
          7452 => x"5281d3fc",
          7453 => x"51ff8bab",
          7454 => x"3f893981",
          7455 => x"d48451ff",
          7456 => x"85bd3f81",
          7457 => x"1555a051",
          7458 => x"fef6af3f",
          7459 => x"ff803981",
          7460 => x"d48851ff",
          7461 => x"85a93f80",
          7462 => x"55747727",
          7463 => x"aa387416",
          7464 => x"70337972",
          7465 => x"26525553",
          7466 => x"9f742790",
          7467 => x"3872802e",
          7468 => x"8b387380",
          7469 => x"fe268538",
          7470 => x"73518339",
          7471 => x"a051fef5",
          7472 => x"f93f8115",
          7473 => x"55d33981",
          7474 => x"d48c51ff",
          7475 => x"84f13f76",
          7476 => x"16771a5a",
          7477 => x"56fef9b4",
          7478 => x"3f81dec0",
          7479 => x"08982b70",
          7480 => x"982c5155",
          7481 => x"74a02e09",
          7482 => x"8106a538",
          7483 => x"fef99d3f",
          7484 => x"81dec008",
          7485 => x"982b7098",
          7486 => x"2c70a032",
          7487 => x"70307072",
          7488 => x"079f2a51",
          7489 => x"56565155",
          7490 => x"749b2e8c",
          7491 => x"3872dd38",
          7492 => x"749b2e09",
          7493 => x"81068538",
          7494 => x"80538c39",
          7495 => x"7a1c5372",
          7496 => x"7626fdd6",
          7497 => x"38ff5372",
          7498 => x"81dec00c",
          7499 => x"8d3d0d04",
          7500 => x"ec3d0d66",
          7501 => x"02840580",
          7502 => x"e3053369",
          7503 => x"72307074",
          7504 => x"07802570",
          7505 => x"87ff7427",
          7506 => x"07515158",
          7507 => x"5a5b5693",
          7508 => x"577480fc",
          7509 => x"38815375",
          7510 => x"528c3d70",
          7511 => x"5257ffbf",
          7512 => x"de3f81de",
          7513 => x"c0085681",
          7514 => x"dec008b8",
          7515 => x"3881dec0",
          7516 => x"0887c098",
          7517 => x"880c81de",
          7518 => x"c0085996",
          7519 => x"3dd40554",
          7520 => x"84805377",
          7521 => x"527651c4",
          7522 => x"9b3f81de",
          7523 => x"c0085681",
          7524 => x"dec00890",
          7525 => x"387a5574",
          7526 => x"802e8938",
          7527 => x"74197519",
          7528 => x"5959d839",
          7529 => x"963dd805",
          7530 => x"51cc853f",
          7531 => x"75307077",
          7532 => x"07802551",
          7533 => x"5579802e",
          7534 => x"95387480",
          7535 => x"2e903881",
          7536 => x"d4905387",
          7537 => x"c0988808",
          7538 => x"527851fb",
          7539 => x"d63f7557",
          7540 => x"7681dec0",
          7541 => x"0c963d0d",
          7542 => x"04f93d0d",
          7543 => x"7b028405",
          7544 => x"b3053357",
          7545 => x"58ff5780",
          7546 => x"537a5279",
          7547 => x"51fec13f",
          7548 => x"81dec008",
          7549 => x"a4387580",
          7550 => x"2e883875",
          7551 => x"812e9838",
          7552 => x"98396055",
          7553 => x"7f5481de",
          7554 => x"c0537e52",
          7555 => x"7d51772d",
          7556 => x"81dec008",
          7557 => x"57833977",
          7558 => x"047681de",
          7559 => x"c00c893d",
          7560 => x"0d04fc3d",
          7561 => x"0d029b05",
          7562 => x"3381d498",
          7563 => x"5381d4a0",
          7564 => x"5255ff87",
          7565 => x"ee3f81db",
          7566 => x"c02251ff",
          7567 => x"80893f81",
          7568 => x"d4ac5481",
          7569 => x"d4b85381",
          7570 => x"dbc13352",
          7571 => x"81d4c051",
          7572 => x"ff87d03f",
          7573 => x"74802e85",
          7574 => x"38fefbd4",
          7575 => x"3f863d0d",
          7576 => x"04fe3d0d",
          7577 => x"87c09680",
          7578 => x"0853ff80",
          7579 => x"a23f8151",
          7580 => x"fef2ad3f",
          7581 => x"81d4dc51",
          7582 => x"fef4a53f",
          7583 => x"8051fef2",
          7584 => x"9f3f7281",
          7585 => x"2a708106",
          7586 => x"51527180",
          7587 => x"2e953881",
          7588 => x"51fef28c",
          7589 => x"3f81d4f8",
          7590 => x"51fef484",
          7591 => x"3f8051fe",
          7592 => x"f1fe3f72",
          7593 => x"822a7081",
          7594 => x"06515271",
          7595 => x"802e9538",
          7596 => x"8151fef1",
          7597 => x"eb3f81d5",
          7598 => x"8c51fef3",
          7599 => x"e33f8051",
          7600 => x"fef1dd3f",
          7601 => x"72832a70",
          7602 => x"81065152",
          7603 => x"71802e95",
          7604 => x"388151fe",
          7605 => x"f1ca3f81",
          7606 => x"d59c51fe",
          7607 => x"f3c23f80",
          7608 => x"51fef1bc",
          7609 => x"3f72842a",
          7610 => x"70810651",
          7611 => x"5271802e",
          7612 => x"95388151",
          7613 => x"fef1a93f",
          7614 => x"81d5b051",
          7615 => x"fef3a13f",
          7616 => x"8051fef1",
          7617 => x"9b3f7285",
          7618 => x"2a708106",
          7619 => x"51527180",
          7620 => x"2e953881",
          7621 => x"51fef188",
          7622 => x"3f81d5c4",
          7623 => x"51fef380",
          7624 => x"3f8051fe",
          7625 => x"f0fa3f72",
          7626 => x"862a7081",
          7627 => x"06515271",
          7628 => x"802e9538",
          7629 => x"8151fef0",
          7630 => x"e73f81d5",
          7631 => x"d851fef2",
          7632 => x"df3f8051",
          7633 => x"fef0d93f",
          7634 => x"72872a70",
          7635 => x"81065152",
          7636 => x"71802e95",
          7637 => x"388151fe",
          7638 => x"f0c63f81",
          7639 => x"d5ec51fe",
          7640 => x"f2be3f80",
          7641 => x"51fef0b8",
          7642 => x"3f72882a",
          7643 => x"70810651",
          7644 => x"5271802e",
          7645 => x"95388151",
          7646 => x"fef0a53f",
          7647 => x"81d68051",
          7648 => x"fef29d3f",
          7649 => x"8051fef0",
          7650 => x"973ffefe",
          7651 => x"cb3f843d",
          7652 => x"0d04fa3d",
          7653 => x"0d787008",
          7654 => x"70555557",
          7655 => x"73802e80",
          7656 => x"f0388e39",
          7657 => x"73770c85",
          7658 => x"15335380",
          7659 => x"e4398114",
          7660 => x"54807433",
          7661 => x"7081ff06",
          7662 => x"57575374",
          7663 => x"a02e8338",
          7664 => x"81537480",
          7665 => x"2e843872",
          7666 => x"e5387581",
          7667 => x"ff065372",
          7668 => x"a02e0981",
          7669 => x"06883880",
          7670 => x"74708105",
          7671 => x"56348056",
          7672 => x"75902981",
          7673 => x"dbf00577",
          7674 => x"08537008",
          7675 => x"5255feea",
          7676 => x"9e3f81de",
          7677 => x"c0088b38",
          7678 => x"84153353",
          7679 => x"72812eff",
          7680 => x"a3388116",
          7681 => x"7081ff06",
          7682 => x"57539476",
          7683 => x"27d238ff",
          7684 => x"537281de",
          7685 => x"c00c883d",
          7686 => x"0d04fb3d",
          7687 => x"0d777970",
          7688 => x"55565680",
          7689 => x"527551fe",
          7690 => x"e8d43f81",
          7691 => x"dbec3354",
          7692 => x"73a73881",
          7693 => x"5381d6c0",
          7694 => x"5281f5c4",
          7695 => x"51ffb9ff",
          7696 => x"3f81dec0",
          7697 => x"08307081",
          7698 => x"dec00807",
          7699 => x"80258271",
          7700 => x"31515154",
          7701 => x"7381dbec",
          7702 => x"3481dbec",
          7703 => x"33547381",
          7704 => x"2e098106",
          7705 => x"ac3881f5",
          7706 => x"c4537452",
          7707 => x"7551f4b5",
          7708 => x"3f81dec0",
          7709 => x"08802e8c",
          7710 => x"3881dec0",
          7711 => x"0851fefd",
          7712 => x"be3f8e39",
          7713 => x"81f5c451",
          7714 => x"c6a63f82",
          7715 => x"0b81dbec",
          7716 => x"3481dbec",
          7717 => x"33547382",
          7718 => x"2e098106",
          7719 => x"89387452",
          7720 => x"7551ff83",
          7721 => x"d83f800b",
          7722 => x"81dec00c",
          7723 => x"873d0d04",
          7724 => x"cb3d0d80",
          7725 => x"707181f5",
          7726 => x"c00c405d",
          7727 => x"81527c51",
          7728 => x"ff88d73f",
          7729 => x"81dec008",
          7730 => x"81ff0659",
          7731 => x"787d2e09",
          7732 => x"8106a238",
          7733 => x"81d6d052",
          7734 => x"993d7052",
          7735 => x"59ff82d9",
          7736 => x"3f7c5378",
          7737 => x"5281dff0",
          7738 => x"51ffb7f2",
          7739 => x"3f81dec0",
          7740 => x"087d2e88",
          7741 => x"3881d6d4",
          7742 => x"5192bc39",
          7743 => x"8170405d",
          7744 => x"81d78c51",
          7745 => x"fefcb83f",
          7746 => x"993d7046",
          7747 => x"5a80f852",
          7748 => x"7951fe86",
          7749 => x"3fb73dfe",
          7750 => x"f80551fc",
          7751 => x"f53f81de",
          7752 => x"c008902b",
          7753 => x"70902c51",
          7754 => x"597880c3",
          7755 => x"2e8ace38",
          7756 => x"7880c324",
          7757 => x"80dc3878",
          7758 => x"ab2e83bc",
          7759 => x"3878ab24",
          7760 => x"a4387882",
          7761 => x"2e81af38",
          7762 => x"7882248a",
          7763 => x"3878802e",
          7764 => x"ffae388f",
          7765 => x"de397884",
          7766 => x"2e828238",
          7767 => x"78942e82",
          7768 => x"ad388fcf",
          7769 => x"397880c0",
          7770 => x"2e858738",
          7771 => x"7880c024",
          7772 => x"903878b0",
          7773 => x"2e83a938",
          7774 => x"78bc2e84",
          7775 => x"8b388fb3",
          7776 => x"397880c1",
          7777 => x"2e879e38",
          7778 => x"7880c22e",
          7779 => x"88bf388f",
          7780 => x"a2397880",
          7781 => x"d52e8df3",
          7782 => x"387880d5",
          7783 => x"24a93878",
          7784 => x"80d02e8d",
          7785 => x"a7387880",
          7786 => x"d0248b38",
          7787 => x"7880c52e",
          7788 => x"8aeb388e",
          7789 => x"fe397880",
          7790 => x"d12e8da1",
          7791 => x"387880d4",
          7792 => x"2e8dab38",
          7793 => x"8eed3978",
          7794 => x"81822e8e",
          7795 => x"c3387881",
          7796 => x"82249238",
          7797 => x"7880f82e",
          7798 => x"8dce3878",
          7799 => x"80f92e8d",
          7800 => x"ec388ecf",
          7801 => x"39788183",
          7802 => x"2e8eb438",
          7803 => x"7881852e",
          7804 => x"8eba388e",
          7805 => x"be39b73d",
          7806 => x"fef41153",
          7807 => x"fef80551",
          7808 => x"ff82953f",
          7809 => x"81dec008",
          7810 => x"883881d7",
          7811 => x"905190a7",
          7812 => x"39b73dfe",
          7813 => x"f01153fe",
          7814 => x"f80551ff",
          7815 => x"81fa3f81",
          7816 => x"dec00880",
          7817 => x"2e883881",
          7818 => x"63258338",
          7819 => x"80430280",
          7820 => x"cb053352",
          7821 => x"0280cf05",
          7822 => x"3351ff85",
          7823 => x"dd3f81de",
          7824 => x"c00881ff",
          7825 => x"0659788e",
          7826 => x"3881d7a0",
          7827 => x"51fef9ef",
          7828 => x"3f815ffd",
          7829 => x"ab3981d7",
          7830 => x"b0518ca8",
          7831 => x"39b73dfe",
          7832 => x"f41153fe",
          7833 => x"f80551ff",
          7834 => x"81ae3f81",
          7835 => x"dec00880",
          7836 => x"2efd8d38",
          7837 => x"80538052",
          7838 => x"0280cf05",
          7839 => x"3351ff89",
          7840 => x"e63f81de",
          7841 => x"c0085281",
          7842 => x"d7c8518c",
          7843 => x"fc39b73d",
          7844 => x"fef41153",
          7845 => x"fef80551",
          7846 => x"ff80fd3f",
          7847 => x"81dec008",
          7848 => x"802e8738",
          7849 => x"638926fc",
          7850 => x"d738b73d",
          7851 => x"fef01153",
          7852 => x"fef80551",
          7853 => x"ff80e13f",
          7854 => x"81dec008",
          7855 => x"863881de",
          7856 => x"c0084363",
          7857 => x"5381d7d0",
          7858 => x"527951fe",
          7859 => x"feeb3f02",
          7860 => x"80cb0533",
          7861 => x"53795263",
          7862 => x"84b42981",
          7863 => x"dff00551",
          7864 => x"ffb3fb3f",
          7865 => x"81dec008",
          7866 => x"81933881",
          7867 => x"d7a051fe",
          7868 => x"f8cd3f81",
          7869 => x"5dfc8939",
          7870 => x"b73dfef8",
          7871 => x"0551fee5",
          7872 => x"d03f81de",
          7873 => x"c008b83d",
          7874 => x"fef80552",
          7875 => x"5bfee6a3",
          7876 => x"3f815381",
          7877 => x"dec00852",
          7878 => x"7a51f494",
          7879 => x"3f80d539",
          7880 => x"b73dfef8",
          7881 => x"0551fee5",
          7882 => x"a83f81de",
          7883 => x"c008b83d",
          7884 => x"fef80552",
          7885 => x"5bfee5fb",
          7886 => x"3f81dec0",
          7887 => x"08b83dfe",
          7888 => x"f805525a",
          7889 => x"fee5ec3f",
          7890 => x"81dec008",
          7891 => x"b83dfef8",
          7892 => x"055259fe",
          7893 => x"e5dd3f81",
          7894 => x"db8c5881",
          7895 => x"def45780",
          7896 => x"56805581",
          7897 => x"dec00881",
          7898 => x"ff065478",
          7899 => x"5379527a",
          7900 => x"51f4e63f",
          7901 => x"81dec008",
          7902 => x"802efb84",
          7903 => x"3881dec0",
          7904 => x"0851eefb",
          7905 => x"3ffaf939",
          7906 => x"b73dfef4",
          7907 => x"1153fef8",
          7908 => x"0551feff",
          7909 => x"833f81de",
          7910 => x"c008802e",
          7911 => x"fae238b7",
          7912 => x"3dfef011",
          7913 => x"53fef805",
          7914 => x"51fefeec",
          7915 => x"3f81dec0",
          7916 => x"08802efa",
          7917 => x"cb38b73d",
          7918 => x"feec1153",
          7919 => x"fef80551",
          7920 => x"fefed53f",
          7921 => x"81dec008",
          7922 => x"863881de",
          7923 => x"c0084281",
          7924 => x"d7d451fe",
          7925 => x"f6e93f63",
          7926 => x"635c5a79",
          7927 => x"7b2788e6",
          7928 => x"38615978",
          7929 => x"7a708405",
          7930 => x"5c0c7a7a",
          7931 => x"26f53888",
          7932 => x"d539b73d",
          7933 => x"fef41153",
          7934 => x"fef80551",
          7935 => x"fefe993f",
          7936 => x"81dec008",
          7937 => x"80df3881",
          7938 => x"dbd43359",
          7939 => x"78802e89",
          7940 => x"3881db8c",
          7941 => x"084480cd",
          7942 => x"3981dbd5",
          7943 => x"33597880",
          7944 => x"2e883881",
          7945 => x"db940844",
          7946 => x"bc3981db",
          7947 => x"d6335978",
          7948 => x"802e8838",
          7949 => x"81db9c08",
          7950 => x"44ab3981",
          7951 => x"dbd73359",
          7952 => x"78802e88",
          7953 => x"3881dba4",
          7954 => x"08449a39",
          7955 => x"81dbd233",
          7956 => x"5978802e",
          7957 => x"883881db",
          7958 => x"ac084489",
          7959 => x"3981dbbc",
          7960 => x"08fc8005",
          7961 => x"44b73dfe",
          7962 => x"f01153fe",
          7963 => x"f80551fe",
          7964 => x"fda63f81",
          7965 => x"dec00880",
          7966 => x"de3881db",
          7967 => x"d4335978",
          7968 => x"802e8938",
          7969 => x"81db9008",
          7970 => x"4380cc39",
          7971 => x"81dbd533",
          7972 => x"5978802e",
          7973 => x"883881db",
          7974 => x"980843bb",
          7975 => x"3981dbd6",
          7976 => x"33597880",
          7977 => x"2e883881",
          7978 => x"dba00843",
          7979 => x"aa3981db",
          7980 => x"d7335978",
          7981 => x"802e8838",
          7982 => x"81dba808",
          7983 => x"43993981",
          7984 => x"dbd23359",
          7985 => x"78802e88",
          7986 => x"3881dbb0",
          7987 => x"08438839",
          7988 => x"81dbbc08",
          7989 => x"880543b7",
          7990 => x"3dfeec11",
          7991 => x"53fef805",
          7992 => x"51fefcb4",
          7993 => x"3f81dec0",
          7994 => x"08802e9b",
          7995 => x"3880625b",
          7996 => x"5979882e",
          7997 => x"83388159",
          7998 => x"79902e8d",
          7999 => x"3878802e",
          8000 => x"883879a0",
          8001 => x"2e833888",
          8002 => x"4281d7e4",
          8003 => x"51fef4af",
          8004 => x"3fa05563",
          8005 => x"54615362",
          8006 => x"526351ed",
          8007 => x"c53f81d7",
          8008 => x"f45186e0",
          8009 => x"39b73dfe",
          8010 => x"f41153fe",
          8011 => x"f80551fe",
          8012 => x"fbe63f81",
          8013 => x"dec00880",
          8014 => x"2ef7c538",
          8015 => x"b73dfef0",
          8016 => x"1153fef8",
          8017 => x"0551fefb",
          8018 => x"cf3f81de",
          8019 => x"c008802e",
          8020 => x"a5386359",
          8021 => x"0280cb05",
          8022 => x"33793463",
          8023 => x"810544b7",
          8024 => x"3dfef011",
          8025 => x"53fef805",
          8026 => x"51fefbac",
          8027 => x"3f81dec0",
          8028 => x"08e038f7",
          8029 => x"8b396370",
          8030 => x"33545281",
          8031 => x"d88051fe",
          8032 => x"f9a13f80",
          8033 => x"f8527951",
          8034 => x"fef9f23f",
          8035 => x"79457933",
          8036 => x"5978ae2e",
          8037 => x"f6ea389f",
          8038 => x"7927a038",
          8039 => x"b73dfef0",
          8040 => x"1153fef8",
          8041 => x"0551fefa",
          8042 => x"ef3f81de",
          8043 => x"c008802e",
          8044 => x"91386359",
          8045 => x"0280cb05",
          8046 => x"33793463",
          8047 => x"810544ff",
          8048 => x"b53981d8",
          8049 => x"8c51fef2",
          8050 => x"f63fffaa",
          8051 => x"39b73dfe",
          8052 => x"e81153fe",
          8053 => x"f80551fe",
          8054 => x"fcb03f81",
          8055 => x"dec00880",
          8056 => x"2ef69d38",
          8057 => x"b73dfee4",
          8058 => x"1153fef8",
          8059 => x"0551fefc",
          8060 => x"993f81de",
          8061 => x"c008802e",
          8062 => x"a6386059",
          8063 => x"02be0522",
          8064 => x"79708205",
          8065 => x"5b237841",
          8066 => x"b73dfee4",
          8067 => x"1153fef8",
          8068 => x"0551fefb",
          8069 => x"f53f81de",
          8070 => x"c008df38",
          8071 => x"f5e23960",
          8072 => x"70225452",
          8073 => x"81d89451",
          8074 => x"fef7f83f",
          8075 => x"80f85279",
          8076 => x"51fef8c9",
          8077 => x"3f794579",
          8078 => x"335978ae",
          8079 => x"2ef5c138",
          8080 => x"789f2687",
          8081 => x"38608205",
          8082 => x"41d539b7",
          8083 => x"3dfee411",
          8084 => x"53fef805",
          8085 => x"51fefbb2",
          8086 => x"3f81dec0",
          8087 => x"08802e92",
          8088 => x"38605902",
          8089 => x"be052279",
          8090 => x"7082055b",
          8091 => x"237841ff",
          8092 => x"ae3981d8",
          8093 => x"8c51fef1",
          8094 => x"c63fffa3",
          8095 => x"39b73dfe",
          8096 => x"e81153fe",
          8097 => x"f80551fe",
          8098 => x"fb803f81",
          8099 => x"dec00880",
          8100 => x"2ef4ed38",
          8101 => x"b73dfee4",
          8102 => x"1153fef8",
          8103 => x"0551fefa",
          8104 => x"e93f81de",
          8105 => x"c008802e",
          8106 => x"a1386060",
          8107 => x"710c5960",
          8108 => x"840541b7",
          8109 => x"3dfee411",
          8110 => x"53fef805",
          8111 => x"51fefaca",
          8112 => x"3f81dec0",
          8113 => x"08e438f4",
          8114 => x"b7396070",
          8115 => x"08545281",
          8116 => x"d8a051fe",
          8117 => x"f6cd3f80",
          8118 => x"f8527951",
          8119 => x"fef79e3f",
          8120 => x"79457933",
          8121 => x"5978ae2e",
          8122 => x"f496389f",
          8123 => x"79279c38",
          8124 => x"b73dfee4",
          8125 => x"1153fef8",
          8126 => x"0551fefa",
          8127 => x"8d3f81de",
          8128 => x"c008802e",
          8129 => x"8d386060",
          8130 => x"710c5960",
          8131 => x"840541ff",
          8132 => x"b93981d8",
          8133 => x"8c51fef0",
          8134 => x"a63fffae",
          8135 => x"39b73dfe",
          8136 => x"f41153fe",
          8137 => x"f80551fe",
          8138 => x"f7ee3f81",
          8139 => x"dec00880",
          8140 => x"df3881db",
          8141 => x"d4335978",
          8142 => x"802e8938",
          8143 => x"81db8c08",
          8144 => x"4480cd39",
          8145 => x"81dbd533",
          8146 => x"5978802e",
          8147 => x"883881db",
          8148 => x"940844bc",
          8149 => x"3981dbd6",
          8150 => x"33597880",
          8151 => x"2e883881",
          8152 => x"db9c0844",
          8153 => x"ab3981db",
          8154 => x"d7335978",
          8155 => x"802e8838",
          8156 => x"81dba408",
          8157 => x"449a3981",
          8158 => x"dbd23359",
          8159 => x"78802e88",
          8160 => x"3881dbac",
          8161 => x"08448939",
          8162 => x"81dbbc08",
          8163 => x"fc800544",
          8164 => x"b73dfef0",
          8165 => x"1153fef8",
          8166 => x"0551fef6",
          8167 => x"fb3f81de",
          8168 => x"c00880de",
          8169 => x"3881dbd4",
          8170 => x"33597880",
          8171 => x"2e893881",
          8172 => x"db900843",
          8173 => x"80cc3981",
          8174 => x"dbd53359",
          8175 => x"78802e88",
          8176 => x"3881db98",
          8177 => x"0843bb39",
          8178 => x"81dbd633",
          8179 => x"5978802e",
          8180 => x"883881db",
          8181 => x"a00843aa",
          8182 => x"3981dbd7",
          8183 => x"33597880",
          8184 => x"2e883881",
          8185 => x"dba80843",
          8186 => x"993981db",
          8187 => x"d2335978",
          8188 => x"802e8838",
          8189 => x"81dbb008",
          8190 => x"43883981",
          8191 => x"dbbc0888",
          8192 => x"0543b73d",
          8193 => x"feec1153",
          8194 => x"fef80551",
          8195 => x"fef6893f",
          8196 => x"81dec008",
          8197 => x"863881de",
          8198 => x"c0084281",
          8199 => x"d8ac51fe",
          8200 => x"ee9d3f63",
          8201 => x"5a796327",
          8202 => x"9d387908",
          8203 => x"5978622e",
          8204 => x"0981068d",
          8205 => x"38785379",
          8206 => x"5281d8bc",
          8207 => x"51fef3e3",
          8208 => x"3f841a5a",
          8209 => x"e03981d7",
          8210 => x"9c51b939",
          8211 => x"81d8cc51",
          8212 => x"feedec3f",
          8213 => x"8251feec",
          8214 => x"da3ff1a4",
          8215 => x"3981d8e4",
          8216 => x"51feeddb",
          8217 => x"3fa251fe",
          8218 => x"ecad3ff1",
          8219 => x"93398480",
          8220 => x"810b87c0",
          8221 => x"94840c84",
          8222 => x"80810b87",
          8223 => x"c094940c",
          8224 => x"81d8fc51",
          8225 => x"feedb83f",
          8226 => x"f0f63981",
          8227 => x"d99051fe",
          8228 => x"edad3f8c",
          8229 => x"80830b87",
          8230 => x"c094840c",
          8231 => x"8c80830b",
          8232 => x"87c09494",
          8233 => x"0cf0d939",
          8234 => x"b73dfef4",
          8235 => x"1153fef8",
          8236 => x"0551fef4",
          8237 => x"e33f81de",
          8238 => x"c008802e",
          8239 => x"f0c23863",
          8240 => x"5281d9a4",
          8241 => x"51fef2db",
          8242 => x"3f635978",
          8243 => x"04b73dfe",
          8244 => x"f41153fe",
          8245 => x"f80551fe",
          8246 => x"f4be3f81",
          8247 => x"dec00880",
          8248 => x"2ef09d38",
          8249 => x"635281d9",
          8250 => x"c051fef2",
          8251 => x"b63f6359",
          8252 => x"782d81de",
          8253 => x"c0085e81",
          8254 => x"dec00880",
          8255 => x"2ef08138",
          8256 => x"81dec008",
          8257 => x"5281d9dc",
          8258 => x"51fef297",
          8259 => x"3feff139",
          8260 => x"81d9f851",
          8261 => x"feeca83f",
          8262 => x"febde53f",
          8263 => x"efe23981",
          8264 => x"da9451fe",
          8265 => x"ec993f80",
          8266 => x"59ffa039",
          8267 => x"fee6813f",
          8268 => x"efce3964",
          8269 => x"70335159",
          8270 => x"78802eef",
          8271 => x"c3387c80",
          8272 => x"2e81dc38",
          8273 => x"81706006",
          8274 => x"5a5a7880",
          8275 => x"2e81d038",
          8276 => x"b73dfef8",
          8277 => x"0551fed8",
          8278 => x"f83f81de",
          8279 => x"c0087a5d",
          8280 => x"5b7b822e",
          8281 => x"b2387b82",
          8282 => x"2489387b",
          8283 => x"812e8c38",
          8284 => x"80cd397b",
          8285 => x"832eb038",
          8286 => x"80c53981",
          8287 => x"daa8567a",
          8288 => x"5581daac",
          8289 => x"54805381",
          8290 => x"dab052b7",
          8291 => x"3dffb005",
          8292 => x"51fef1a5",
          8293 => x"3fbb3981",
          8294 => x"dad052b7",
          8295 => x"3dffb005",
          8296 => x"51fef195",
          8297 => x"3fab397a",
          8298 => x"5581daac",
          8299 => x"54805381",
          8300 => x"dac052b7",
          8301 => x"3dffb005",
          8302 => x"51fef0fd",
          8303 => x"3f93397a",
          8304 => x"54805381",
          8305 => x"dacc52b7",
          8306 => x"3dffb005",
          8307 => x"51fef0e9",
          8308 => x"3f81db8c",
          8309 => x"5881def4",
          8310 => x"57805664",
          8311 => x"81114681",
          8312 => x"05558054",
          8313 => x"82808053",
          8314 => x"82808052",
          8315 => x"b73dffb0",
          8316 => x"0551e7e5",
          8317 => x"3f81dec0",
          8318 => x"0881dec0",
          8319 => x"08097030",
          8320 => x"70720780",
          8321 => x"25515b5b",
          8322 => x"5e7b8326",
          8323 => x"92387880",
          8324 => x"2e8d3881",
          8325 => x"1c7081ff",
          8326 => x"065d597b",
          8327 => x"fec3387e",
          8328 => x"81327d81",
          8329 => x"32075978",
          8330 => x"8a387dff",
          8331 => x"2e098106",
          8332 => x"edce3881",
          8333 => x"dad451fe",
          8334 => x"efe93fed",
          8335 => x"c339fc3d",
          8336 => x"0d800b81",
          8337 => x"def43487",
          8338 => x"c0948c70",
          8339 => x"08545587",
          8340 => x"84805272",
          8341 => x"51fece9f",
          8342 => x"3f81dec0",
          8343 => x"08902b75",
          8344 => x"08555387",
          8345 => x"84805273",
          8346 => x"51fece8b",
          8347 => x"3f7281de",
          8348 => x"c0080775",
          8349 => x"0c87c094",
          8350 => x"9c700854",
          8351 => x"55878480",
          8352 => x"527251fe",
          8353 => x"cdf13f81",
          8354 => x"dec00890",
          8355 => x"2b750855",
          8356 => x"53878480",
          8357 => x"527351fe",
          8358 => x"cddd3f72",
          8359 => x"81dec008",
          8360 => x"07750c8c",
          8361 => x"80830b87",
          8362 => x"c094840c",
          8363 => x"8c80830b",
          8364 => x"87c09494",
          8365 => x"0c9fba0b",
          8366 => x"81ded00c",
          8367 => x"a2bb0b81",
          8368 => x"ded40cfe",
          8369 => x"de9e3ffe",
          8370 => x"e7c53f81",
          8371 => x"dae451fe",
          8372 => x"dbce3f81",
          8373 => x"daf051fe",
          8374 => x"e8e53f81",
          8375 => x"ace151fe",
          8376 => x"e7a83f81",
          8377 => x"51e6bb3f",
          8378 => x"ebc63f80",
          8379 => x"04000000",
          8380 => x"00ffffff",
          8381 => x"ff00ffff",
          8382 => x"ffff00ff",
          8383 => x"ffffff00",
          8384 => x"00001661",
          8385 => x"00001667",
          8386 => x"0000166d",
          8387 => x"00001673",
          8388 => x"00001679",
          8389 => x"00005391",
          8390 => x"00005315",
          8391 => x"0000531c",
          8392 => x"00005323",
          8393 => x"0000532a",
          8394 => x"00005331",
          8395 => x"00005338",
          8396 => x"0000533f",
          8397 => x"00005346",
          8398 => x"0000534d",
          8399 => x"00005354",
          8400 => x"0000535b",
          8401 => x"00005361",
          8402 => x"00005367",
          8403 => x"0000536d",
          8404 => x"00005373",
          8405 => x"00005379",
          8406 => x"0000537f",
          8407 => x"00005385",
          8408 => x"0000538b",
          8409 => x"25642f25",
          8410 => x"642f2564",
          8411 => x"2025643a",
          8412 => x"25643a25",
          8413 => x"642e2564",
          8414 => x"25640a00",
          8415 => x"536f4320",
          8416 => x"436f6e66",
          8417 => x"69677572",
          8418 => x"6174696f",
          8419 => x"6e000000",
          8420 => x"20286672",
          8421 => x"6f6d2053",
          8422 => x"6f432063",
          8423 => x"6f6e6669",
          8424 => x"67290000",
          8425 => x"3a0a4465",
          8426 => x"76696365",
          8427 => x"7320696d",
          8428 => x"706c656d",
          8429 => x"656e7465",
          8430 => x"643a0a00",
          8431 => x"20202020",
          8432 => x"57422053",
          8433 => x"4452414d",
          8434 => x"20202825",
          8435 => x"3038583a",
          8436 => x"25303858",
          8437 => x"292e0a00",
          8438 => x"20202020",
          8439 => x"53445241",
          8440 => x"4d202020",
          8441 => x"20202825",
          8442 => x"3038583a",
          8443 => x"25303858",
          8444 => x"292e0a00",
          8445 => x"20202020",
          8446 => x"494e534e",
          8447 => x"20425241",
          8448 => x"4d202825",
          8449 => x"3038583a",
          8450 => x"25303858",
          8451 => x"292e0a00",
          8452 => x"20202020",
          8453 => x"4252414d",
          8454 => x"20202020",
          8455 => x"20202825",
          8456 => x"3038583a",
          8457 => x"25303858",
          8458 => x"292e0a00",
          8459 => x"20202020",
          8460 => x"52414d20",
          8461 => x"20202020",
          8462 => x"20202825",
          8463 => x"3038583a",
          8464 => x"25303858",
          8465 => x"292e0a00",
          8466 => x"20202020",
          8467 => x"53442043",
          8468 => x"41524420",
          8469 => x"20202844",
          8470 => x"65766963",
          8471 => x"6573203d",
          8472 => x"25303264",
          8473 => x"292e0a00",
          8474 => x"20202020",
          8475 => x"54494d45",
          8476 => x"52312020",
          8477 => x"20202854",
          8478 => x"696d6572",
          8479 => x"7320203d",
          8480 => x"25303264",
          8481 => x"292e0a00",
          8482 => x"20202020",
          8483 => x"494e5452",
          8484 => x"20435452",
          8485 => x"4c202843",
          8486 => x"68616e6e",
          8487 => x"656c733d",
          8488 => x"25303264",
          8489 => x"292e0a00",
          8490 => x"20202020",
          8491 => x"57495348",
          8492 => x"424f4e45",
          8493 => x"20425553",
          8494 => x"0a000000",
          8495 => x"20202020",
          8496 => x"57422049",
          8497 => x"32430a00",
          8498 => x"20202020",
          8499 => x"494f4354",
          8500 => x"4c0a0000",
          8501 => x"20202020",
          8502 => x"5053320a",
          8503 => x"00000000",
          8504 => x"20202020",
          8505 => x"5350490a",
          8506 => x"00000000",
          8507 => x"41646472",
          8508 => x"65737365",
          8509 => x"733a0a00",
          8510 => x"20202020",
          8511 => x"43505520",
          8512 => x"52657365",
          8513 => x"74205665",
          8514 => x"63746f72",
          8515 => x"20416464",
          8516 => x"72657373",
          8517 => x"203d2025",
          8518 => x"3038580a",
          8519 => x"00000000",
          8520 => x"20202020",
          8521 => x"43505520",
          8522 => x"4d656d6f",
          8523 => x"72792053",
          8524 => x"74617274",
          8525 => x"20416464",
          8526 => x"72657373",
          8527 => x"203d2025",
          8528 => x"3038580a",
          8529 => x"00000000",
          8530 => x"20202020",
          8531 => x"53746163",
          8532 => x"6b205374",
          8533 => x"61727420",
          8534 => x"41646472",
          8535 => x"65737320",
          8536 => x"20202020",
          8537 => x"203d2025",
          8538 => x"3038580a",
          8539 => x"00000000",
          8540 => x"4d697363",
          8541 => x"3a0a0000",
          8542 => x"20202020",
          8543 => x"5a505520",
          8544 => x"49642020",
          8545 => x"20202020",
          8546 => x"20202020",
          8547 => x"20202020",
          8548 => x"20202020",
          8549 => x"203d2025",
          8550 => x"3034580a",
          8551 => x"00000000",
          8552 => x"20202020",
          8553 => x"53797374",
          8554 => x"656d2043",
          8555 => x"6c6f636b",
          8556 => x"20467265",
          8557 => x"71202020",
          8558 => x"20202020",
          8559 => x"203d2025",
          8560 => x"642e2530",
          8561 => x"34644d48",
          8562 => x"7a0a0000",
          8563 => x"20202020",
          8564 => x"53445241",
          8565 => x"4d20436c",
          8566 => x"6f636b20",
          8567 => x"46726571",
          8568 => x"20202020",
          8569 => x"20202020",
          8570 => x"203d2025",
          8571 => x"642e2530",
          8572 => x"34644d48",
          8573 => x"7a0a0000",
          8574 => x"20202020",
          8575 => x"57697368",
          8576 => x"626f6e65",
          8577 => x"20534452",
          8578 => x"414d2043",
          8579 => x"6c6f636b",
          8580 => x"20467265",
          8581 => x"713d2025",
          8582 => x"642e2530",
          8583 => x"34644d48",
          8584 => x"7a0a0000",
          8585 => x"536d616c",
          8586 => x"6c000000",
          8587 => x"4d656469",
          8588 => x"756d0000",
          8589 => x"466c6578",
          8590 => x"00000000",
          8591 => x"45564f00",
          8592 => x"45564f6d",
          8593 => x"696e0000",
          8594 => x"556e6b6e",
          8595 => x"6f776e00",
          8596 => x"53440000",
          8597 => x"222a2b2c",
          8598 => x"3a3b3c3d",
          8599 => x"3e3f5b5d",
          8600 => x"7c7f0000",
          8601 => x"46415400",
          8602 => x"46415433",
          8603 => x"32000000",
          8604 => x"ebfe904d",
          8605 => x"53444f53",
          8606 => x"352e3000",
          8607 => x"4e4f204e",
          8608 => x"414d4520",
          8609 => x"20202046",
          8610 => x"41543332",
          8611 => x"20202000",
          8612 => x"4e4f204e",
          8613 => x"414d4520",
          8614 => x"20202046",
          8615 => x"41542020",
          8616 => x"20202000",
          8617 => x"00006650",
          8618 => x"00000000",
          8619 => x"00000000",
          8620 => x"00000000",
          8621 => x"809a4541",
          8622 => x"8e418f80",
          8623 => x"45454549",
          8624 => x"49498e8f",
          8625 => x"9092924f",
          8626 => x"994f5555",
          8627 => x"59999a9b",
          8628 => x"9c9d9e9f",
          8629 => x"41494f55",
          8630 => x"a5a5a6a7",
          8631 => x"a8a9aaab",
          8632 => x"acadaeaf",
          8633 => x"b0b1b2b3",
          8634 => x"b4b5b6b7",
          8635 => x"b8b9babb",
          8636 => x"bcbdbebf",
          8637 => x"c0c1c2c3",
          8638 => x"c4c5c6c7",
          8639 => x"c8c9cacb",
          8640 => x"cccdcecf",
          8641 => x"d0d1d2d3",
          8642 => x"d4d5d6d7",
          8643 => x"d8d9dadb",
          8644 => x"dcdddedf",
          8645 => x"e0e1e2e3",
          8646 => x"e4e5e6e7",
          8647 => x"e8e9eaeb",
          8648 => x"ecedeeef",
          8649 => x"f0f1f2f3",
          8650 => x"f4f5f6f7",
          8651 => x"f8f9fafb",
          8652 => x"fcfdfeff",
          8653 => x"2b2e2c3b",
          8654 => x"3d5b5d2f",
          8655 => x"5c222a3a",
          8656 => x"3c3e3f7c",
          8657 => x"7f000000",
          8658 => x"00010004",
          8659 => x"00100040",
          8660 => x"01000200",
          8661 => x"00000000",
          8662 => x"00010002",
          8663 => x"00040008",
          8664 => x"00100020",
          8665 => x"00000000",
          8666 => x"64696e69",
          8667 => x"74000000",
          8668 => x"64696f63",
          8669 => x"746c0000",
          8670 => x"66696e69",
          8671 => x"74000000",
          8672 => x"666c6f61",
          8673 => x"64000000",
          8674 => x"66657865",
          8675 => x"63000000",
          8676 => x"6d636c65",
          8677 => x"61720000",
          8678 => x"6d64756d",
          8679 => x"70000000",
          8680 => x"6d737263",
          8681 => x"68000000",
          8682 => x"6d656200",
          8683 => x"6d656800",
          8684 => x"6d657700",
          8685 => x"68696400",
          8686 => x"68696500",
          8687 => x"68666400",
          8688 => x"68666500",
          8689 => x"63616c6c",
          8690 => x"00000000",
          8691 => x"6a6d7000",
          8692 => x"72657374",
          8693 => x"61727400",
          8694 => x"72657365",
          8695 => x"74000000",
          8696 => x"696e666f",
          8697 => x"00000000",
          8698 => x"74657374",
          8699 => x"00000000",
          8700 => x"4469736b",
          8701 => x"20457272",
          8702 => x"6f720a00",
          8703 => x"496e7465",
          8704 => x"726e616c",
          8705 => x"20657272",
          8706 => x"6f722e0a",
          8707 => x"00000000",
          8708 => x"4469736b",
          8709 => x"206e6f74",
          8710 => x"20726561",
          8711 => x"64792e0a",
          8712 => x"00000000",
          8713 => x"4e6f2066",
          8714 => x"696c6520",
          8715 => x"666f756e",
          8716 => x"642e0a00",
          8717 => x"4e6f2070",
          8718 => x"61746820",
          8719 => x"666f756e",
          8720 => x"642e0a00",
          8721 => x"496e7661",
          8722 => x"6c696420",
          8723 => x"66696c65",
          8724 => x"6e616d65",
          8725 => x"2e0a0000",
          8726 => x"41636365",
          8727 => x"73732064",
          8728 => x"656e6965",
          8729 => x"642e0a00",
          8730 => x"46696c65",
          8731 => x"20616c72",
          8732 => x"65616479",
          8733 => x"20657869",
          8734 => x"7374732e",
          8735 => x"0a000000",
          8736 => x"46696c65",
          8737 => x"2068616e",
          8738 => x"646c6520",
          8739 => x"696e7661",
          8740 => x"6c69642e",
          8741 => x"0a000000",
          8742 => x"53442069",
          8743 => x"73207772",
          8744 => x"69746520",
          8745 => x"70726f74",
          8746 => x"65637465",
          8747 => x"642e0a00",
          8748 => x"44726976",
          8749 => x"65206e75",
          8750 => x"6d626572",
          8751 => x"20697320",
          8752 => x"696e7661",
          8753 => x"6c69642e",
          8754 => x"0a000000",
          8755 => x"4469736b",
          8756 => x"206e6f74",
          8757 => x"20656e61",
          8758 => x"626c6564",
          8759 => x"2e0a0000",
          8760 => x"4e6f2063",
          8761 => x"6f6d7061",
          8762 => x"7469626c",
          8763 => x"65206669",
          8764 => x"6c657379",
          8765 => x"7374656d",
          8766 => x"20666f75",
          8767 => x"6e64206f",
          8768 => x"6e206469",
          8769 => x"736b2e0a",
          8770 => x"00000000",
          8771 => x"466f726d",
          8772 => x"61742061",
          8773 => x"626f7274",
          8774 => x"65642e0a",
          8775 => x"00000000",
          8776 => x"54696d65",
          8777 => x"6f75742c",
          8778 => x"206f7065",
          8779 => x"72617469",
          8780 => x"6f6e2063",
          8781 => x"616e6365",
          8782 => x"6c6c6564",
          8783 => x"2e0a0000",
          8784 => x"46696c65",
          8785 => x"20697320",
          8786 => x"6c6f636b",
          8787 => x"65642e0a",
          8788 => x"00000000",
          8789 => x"496e7375",
          8790 => x"66666963",
          8791 => x"69656e74",
          8792 => x"206d656d",
          8793 => x"6f72792e",
          8794 => x"0a000000",
          8795 => x"546f6f20",
          8796 => x"6d616e79",
          8797 => x"206f7065",
          8798 => x"6e206669",
          8799 => x"6c65732e",
          8800 => x"0a000000",
          8801 => x"50617261",
          8802 => x"6d657465",
          8803 => x"72732069",
          8804 => x"6e636f72",
          8805 => x"72656374",
          8806 => x"2e0a0000",
          8807 => x"53756363",
          8808 => x"6573732e",
          8809 => x"0a000000",
          8810 => x"556e6b6e",
          8811 => x"6f776e20",
          8812 => x"6572726f",
          8813 => x"722e0a00",
          8814 => x"0a256c75",
          8815 => x"20627974",
          8816 => x"65732025",
          8817 => x"73206174",
          8818 => x"20256c75",
          8819 => x"20627974",
          8820 => x"65732f73",
          8821 => x"65632e0a",
          8822 => x"00000000",
          8823 => x"25303858",
          8824 => x"00000000",
          8825 => x"3a202000",
          8826 => x"25303458",
          8827 => x"00000000",
          8828 => x"20202020",
          8829 => x"20202020",
          8830 => x"00000000",
          8831 => x"25303258",
          8832 => x"00000000",
          8833 => x"20200000",
          8834 => x"207c0000",
          8835 => x"7c0d0a00",
          8836 => x"72656164",
          8837 => x"00000000",
          8838 => x"5a505554",
          8839 => x"41000000",
          8840 => x"0a2a2a20",
          8841 => x"25732028",
          8842 => x"00000000",
          8843 => x"32392f31",
          8844 => x"322f3230",
          8845 => x"31390000",
          8846 => x"76312e34",
          8847 => x"00000000",
          8848 => x"205a5055",
          8849 => x"2c207265",
          8850 => x"76202530",
          8851 => x"32782920",
          8852 => x"25732025",
          8853 => x"73202a2a",
          8854 => x"0a0a0000",
          8855 => x"5a505554",
          8856 => x"4120496e",
          8857 => x"74657272",
          8858 => x"75707420",
          8859 => x"48616e64",
          8860 => x"6c65720a",
          8861 => x"00000000",
          8862 => x"54696d65",
          8863 => x"7220696e",
          8864 => x"74657272",
          8865 => x"7570740a",
          8866 => x"00000000",
          8867 => x"50533220",
          8868 => x"696e7465",
          8869 => x"72727570",
          8870 => x"740a0000",
          8871 => x"494f4354",
          8872 => x"4c205244",
          8873 => x"20696e74",
          8874 => x"65727275",
          8875 => x"70740a00",
          8876 => x"494f4354",
          8877 => x"4c205752",
          8878 => x"20696e74",
          8879 => x"65727275",
          8880 => x"70740a00",
          8881 => x"55415254",
          8882 => x"30205258",
          8883 => x"20696e74",
          8884 => x"65727275",
          8885 => x"70740a00",
          8886 => x"55415254",
          8887 => x"30205458",
          8888 => x"20696e74",
          8889 => x"65727275",
          8890 => x"70740a00",
          8891 => x"55415254",
          8892 => x"31205258",
          8893 => x"20696e74",
          8894 => x"65727275",
          8895 => x"70740a00",
          8896 => x"55415254",
          8897 => x"31205458",
          8898 => x"20696e74",
          8899 => x"65727275",
          8900 => x"70740a00",
          8901 => x"53657474",
          8902 => x"696e6720",
          8903 => x"75702074",
          8904 => x"696d6572",
          8905 => x"2e2e2e0a",
          8906 => x"00000000",
          8907 => x"456e6162",
          8908 => x"6c696e67",
          8909 => x"2074696d",
          8910 => x"65722e2e",
          8911 => x"2e0a0000",
          8912 => x"6175746f",
          8913 => x"65786563",
          8914 => x"2e626174",
          8915 => x"00000000",
          8916 => x"303a0000",
          8917 => x"4661696c",
          8918 => x"65642074",
          8919 => x"6f20696e",
          8920 => x"69746961",
          8921 => x"6c697365",
          8922 => x"20736420",
          8923 => x"63617264",
          8924 => x"20302c20",
          8925 => x"706c6561",
          8926 => x"73652069",
          8927 => x"6e697420",
          8928 => x"6d616e75",
          8929 => x"616c6c79",
          8930 => x"2e0a0000",
          8931 => x"2a200000",
          8932 => x"42616420",
          8933 => x"6469736b",
          8934 => x"20696421",
          8935 => x"0a000000",
          8936 => x"496e6974",
          8937 => x"69616c69",
          8938 => x"7365642e",
          8939 => x"0a000000",
          8940 => x"4661696c",
          8941 => x"65642074",
          8942 => x"6f20696e",
          8943 => x"69746961",
          8944 => x"6c697365",
          8945 => x"2e0a0000",
          8946 => x"72633d25",
          8947 => x"640a0000",
          8948 => x"25753a00",
          8949 => x"436c6561",
          8950 => x"72696e67",
          8951 => x"2e2e2e2e",
          8952 => x"00000000",
          8953 => x"44756d70",
          8954 => x"204d656d",
          8955 => x"6f72790a",
          8956 => x"00000000",
          8957 => x"0a436f6d",
          8958 => x"706c6574",
          8959 => x"652e0a00",
          8960 => x"25303858",
          8961 => x"20253032",
          8962 => x"582d0000",
          8963 => x"3f3f3f0a",
          8964 => x"00000000",
          8965 => x"25303858",
          8966 => x"20253034",
          8967 => x"582d0000",
          8968 => x"25303858",
          8969 => x"20253038",
          8970 => x"582d0000",
          8971 => x"53656172",
          8972 => x"6368696e",
          8973 => x"672e2e0a",
          8974 => x"00000000",
          8975 => x"2530386c",
          8976 => x"782d3e25",
          8977 => x"30386c78",
          8978 => x"0a000000",
          8979 => x"44697361",
          8980 => x"626c696e",
          8981 => x"6720696e",
          8982 => x"74657272",
          8983 => x"75707473",
          8984 => x"0a000000",
          8985 => x"456e6162",
          8986 => x"6c696e67",
          8987 => x"20696e74",
          8988 => x"65727275",
          8989 => x"7074730a",
          8990 => x"00000000",
          8991 => x"44697361",
          8992 => x"626c6564",
          8993 => x"20756172",
          8994 => x"74206669",
          8995 => x"666f0a00",
          8996 => x"456e6162",
          8997 => x"6c696e67",
          8998 => x"20756172",
          8999 => x"74206669",
          9000 => x"666f0a00",
          9001 => x"45786563",
          9002 => x"7574696e",
          9003 => x"6720636f",
          9004 => x"64652040",
          9005 => x"20253038",
          9006 => x"78202e2e",
          9007 => x"2e0a0000",
          9008 => x"43616c6c",
          9009 => x"696e6720",
          9010 => x"636f6465",
          9011 => x"20402025",
          9012 => x"30387820",
          9013 => x"2e2e2e0a",
          9014 => x"00000000",
          9015 => x"43616c6c",
          9016 => x"20726574",
          9017 => x"75726e65",
          9018 => x"6420636f",
          9019 => x"64652028",
          9020 => x"2564292e",
          9021 => x"0a000000",
          9022 => x"52657374",
          9023 => x"61727469",
          9024 => x"6e672061",
          9025 => x"70706c69",
          9026 => x"63617469",
          9027 => x"6f6e2e2e",
          9028 => x"2e0a0000",
          9029 => x"436f6c64",
          9030 => x"20726562",
          9031 => x"6f6f7469",
          9032 => x"6e672e2e",
          9033 => x"2e0a0000",
          9034 => x"5a505500",
          9035 => x"62696e00",
          9036 => x"25643a5c",
          9037 => x"25735c25",
          9038 => x"732e2573",
          9039 => x"00000000",
          9040 => x"25643a5c",
          9041 => x"25735c25",
          9042 => x"73000000",
          9043 => x"25643a5c",
          9044 => x"25730000",
          9045 => x"42616420",
          9046 => x"636f6d6d",
          9047 => x"616e642e",
          9048 => x"0a000000",
          9049 => x"52756e6e",
          9050 => x"696e672e",
          9051 => x"2e2e0a00",
          9052 => x"456e6162",
          9053 => x"6c696e67",
          9054 => x"20696e74",
          9055 => x"65727275",
          9056 => x"7074732e",
          9057 => x"2e2e0a00",
          9058 => x"00000000",
          9059 => x"00000000",
          9060 => x"00007fff",
          9061 => x"00000000",
          9062 => x"00007fff",
          9063 => x"00010000",
          9064 => x"00007fff",
          9065 => x"00010000",
          9066 => x"00810000",
          9067 => x"01000000",
          9068 => x"017fffff",
          9069 => x"00000000",
          9070 => x"00000000",
          9071 => x"00007800",
          9072 => x"00000000",
          9073 => x"05f5e100",
          9074 => x"05f5e100",
          9075 => x"05f5e100",
          9076 => x"00000000",
          9077 => x"01010101",
          9078 => x"01010101",
          9079 => x"01011001",
          9080 => x"01000000",
          9081 => x"00000000",
          9082 => x"01000000",
          9083 => x"00000000",
          9084 => x"00006768",
          9085 => x"01020100",
          9086 => x"00000000",
          9087 => x"00000000",
          9088 => x"00006770",
          9089 => x"01040100",
          9090 => x"00000000",
          9091 => x"00000000",
          9092 => x"00006778",
          9093 => x"01140300",
          9094 => x"00000000",
          9095 => x"00000000",
          9096 => x"00006780",
          9097 => x"012b0300",
          9098 => x"00000000",
          9099 => x"00000000",
          9100 => x"00006788",
          9101 => x"01300300",
          9102 => x"00000000",
          9103 => x"00000000",
          9104 => x"00006790",
          9105 => x"013c0400",
          9106 => x"00000000",
          9107 => x"00000000",
          9108 => x"00006798",
          9109 => x"01400400",
          9110 => x"00000000",
          9111 => x"00000000",
          9112 => x"000067a0",
          9113 => x"01450400",
          9114 => x"00000000",
          9115 => x"00000000",
          9116 => x"000067a8",
          9117 => x"01410400",
          9118 => x"00000000",
          9119 => x"00000000",
          9120 => x"000067ac",
          9121 => x"01420400",
          9122 => x"00000000",
          9123 => x"00000000",
          9124 => x"000067b0",
          9125 => x"01430400",
          9126 => x"00000000",
          9127 => x"00000000",
          9128 => x"000067b4",
          9129 => x"01500500",
          9130 => x"00000000",
          9131 => x"00000000",
          9132 => x"000067b8",
          9133 => x"01510500",
          9134 => x"00000000",
          9135 => x"00000000",
          9136 => x"000067bc",
          9137 => x"01540500",
          9138 => x"00000000",
          9139 => x"00000000",
          9140 => x"000067c0",
          9141 => x"01550500",
          9142 => x"00000000",
          9143 => x"00000000",
          9144 => x"000067c4",
          9145 => x"01790700",
          9146 => x"00000000",
          9147 => x"00000000",
          9148 => x"000067cc",
          9149 => x"01780700",
          9150 => x"00000000",
          9151 => x"00000000",
          9152 => x"000067d0",
          9153 => x"01820800",
          9154 => x"00000000",
          9155 => x"00000000",
          9156 => x"000067d8",
          9157 => x"01830800",
          9158 => x"00000000",
          9159 => x"00000000",
          9160 => x"000067e0",
          9161 => x"01850800",
          9162 => x"00000000",
          9163 => x"00000000",
          9164 => x"000067e8",
          9165 => x"01870800",
          9166 => x"00000000",
          9167 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

