-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e9040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"88738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cb2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8a",
           179 => x"fd2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"80040088",
           281 => x"e2040000",
           282 => x"009fac70",
           283 => x"9fdc278b",
           284 => x"38807170",
           285 => x"8405530c",
           286 => x"88eb0488",
           287 => x"e2519e99",
           288 => x"04940802",
           289 => x"940cfd3d",
           290 => x"0d805394",
           291 => x"088c0508",
           292 => x"52940888",
           293 => x"05085182",
           294 => x"de3f8808",
           295 => x"70880c54",
           296 => x"853d0d94",
           297 => x"0c049408",
           298 => x"02940cfd",
           299 => x"3d0d8153",
           300 => x"94088c05",
           301 => x"08529408",
           302 => x"88050851",
           303 => x"82b93f88",
           304 => x"0870880c",
           305 => x"54853d0d",
           306 => x"940c0494",
           307 => x"0802940c",
           308 => x"f93d0d80",
           309 => x"0b9408fc",
           310 => x"050c9408",
           311 => x"88050880",
           312 => x"25ab3894",
           313 => x"08880508",
           314 => x"30940888",
           315 => x"050c800b",
           316 => x"9408f405",
           317 => x"0c9408fc",
           318 => x"05088838",
           319 => x"810b9408",
           320 => x"f4050c94",
           321 => x"08f40508",
           322 => x"9408fc05",
           323 => x"0c94088c",
           324 => x"05088025",
           325 => x"ab389408",
           326 => x"8c050830",
           327 => x"94088c05",
           328 => x"0c800b94",
           329 => x"08f0050c",
           330 => x"9408fc05",
           331 => x"08883881",
           332 => x"0b9408f0",
           333 => x"050c9408",
           334 => x"f0050894",
           335 => x"08fc050c",
           336 => x"80539408",
           337 => x"8c050852",
           338 => x"94088805",
           339 => x"085181a7",
           340 => x"3f880870",
           341 => x"9408f805",
           342 => x"0c549408",
           343 => x"fc050880",
           344 => x"2e8c3894",
           345 => x"08f80508",
           346 => x"309408f8",
           347 => x"050c9408",
           348 => x"f8050870",
           349 => x"880c5489",
           350 => x"3d0d940c",
           351 => x"04940802",
           352 => x"940cfb3d",
           353 => x"0d800b94",
           354 => x"08fc050c",
           355 => x"94088805",
           356 => x"08802593",
           357 => x"38940888",
           358 => x"05083094",
           359 => x"0888050c",
           360 => x"810b9408",
           361 => x"fc050c94",
           362 => x"088c0508",
           363 => x"80258c38",
           364 => x"94088c05",
           365 => x"08309408",
           366 => x"8c050c81",
           367 => x"5394088c",
           368 => x"05085294",
           369 => x"08880508",
           370 => x"51ad3f88",
           371 => x"08709408",
           372 => x"f8050c54",
           373 => x"9408fc05",
           374 => x"08802e8c",
           375 => x"389408f8",
           376 => x"05083094",
           377 => x"08f8050c",
           378 => x"9408f805",
           379 => x"0870880c",
           380 => x"54873d0d",
           381 => x"940c0494",
           382 => x"0802940c",
           383 => x"fd3d0d81",
           384 => x"0b9408fc",
           385 => x"050c800b",
           386 => x"9408f805",
           387 => x"0c94088c",
           388 => x"05089408",
           389 => x"88050827",
           390 => x"ac389408",
           391 => x"fc050880",
           392 => x"2ea33880",
           393 => x"0b94088c",
           394 => x"05082499",
           395 => x"3894088c",
           396 => x"05081094",
           397 => x"088c050c",
           398 => x"9408fc05",
           399 => x"08109408",
           400 => x"fc050cc9",
           401 => x"399408fc",
           402 => x"0508802e",
           403 => x"80c93894",
           404 => x"088c0508",
           405 => x"94088805",
           406 => x"0826a138",
           407 => x"94088805",
           408 => x"0894088c",
           409 => x"05083194",
           410 => x"0888050c",
           411 => x"9408f805",
           412 => x"089408fc",
           413 => x"05080794",
           414 => x"08f8050c",
           415 => x"9408fc05",
           416 => x"08812a94",
           417 => x"08fc050c",
           418 => x"94088c05",
           419 => x"08812a94",
           420 => x"088c050c",
           421 => x"ffaf3994",
           422 => x"08900508",
           423 => x"802e8f38",
           424 => x"94088805",
           425 => x"08709408",
           426 => x"f4050c51",
           427 => x"8d399408",
           428 => x"f8050870",
           429 => x"9408f405",
           430 => x"0c519408",
           431 => x"f4050888",
           432 => x"0c853d0d",
           433 => x"940c04ff",
           434 => x"3d0d8188",
           435 => x"0b87c092",
           436 => x"8c0c810b",
           437 => x"87c0928c",
           438 => x"0c850b87",
           439 => x"c0988c0c",
           440 => x"87c0928c",
           441 => x"08708206",
           442 => x"51517080",
           443 => x"2e8a3887",
           444 => x"c0988c08",
           445 => x"5170e938",
           446 => x"87c0928c",
           447 => x"08fc8080",
           448 => x"06527193",
           449 => x"3887c098",
           450 => x"8c085170",
           451 => x"802e8838",
           452 => x"710b0b0b",
           453 => x"9fa8340b",
           454 => x"0b0b9fa8",
           455 => x"33880c83",
           456 => x"3d0d04fa",
           457 => x"3d0d787b",
           458 => x"7d565856",
           459 => x"800b0b0b",
           460 => x"0b9fa833",
           461 => x"81065255",
           462 => x"82527075",
           463 => x"2e098106",
           464 => x"819e3885",
           465 => x"0b87c098",
           466 => x"8c0c7987",
           467 => x"c092800c",
           468 => x"840b87c0",
           469 => x"928c0c87",
           470 => x"c0928c08",
           471 => x"70852a70",
           472 => x"81065152",
           473 => x"5370802e",
           474 => x"a73887c0",
           475 => x"92840870",
           476 => x"81ff0676",
           477 => x"79275253",
           478 => x"5173802e",
           479 => x"90387080",
           480 => x"2e8b3871",
           481 => x"76708105",
           482 => x"5834ff14",
           483 => x"54811555",
           484 => x"72a20651",
           485 => x"70802e8b",
           486 => x"3887c098",
           487 => x"8c085170",
           488 => x"ffb53887",
           489 => x"c0988c08",
           490 => x"51709538",
           491 => x"810b87c0",
           492 => x"928c0c87",
           493 => x"c0928c08",
           494 => x"70820651",
           495 => x"5170f438",
           496 => x"8073fc80",
           497 => x"80065252",
           498 => x"70722e09",
           499 => x"81068f38",
           500 => x"87c0988c",
           501 => x"08517072",
           502 => x"2e098106",
           503 => x"83388152",
           504 => x"71880c88",
           505 => x"3d0d04fe",
           506 => x"3d0d7481",
           507 => x"11337133",
           508 => x"71882b07",
           509 => x"880c5351",
           510 => x"843d0d04",
           511 => x"fd3d0d75",
           512 => x"83113382",
           513 => x"12337190",
           514 => x"2b71882b",
           515 => x"07811433",
           516 => x"70720788",
           517 => x"2b753371",
           518 => x"07880c52",
           519 => x"53545654",
           520 => x"52853d0d",
           521 => x"04f93d0d",
           522 => x"790b0b0b",
           523 => x"9fac0857",
           524 => x"57817727",
           525 => x"80ed3876",
           526 => x"88170827",
           527 => x"80e53875",
           528 => x"33557482",
           529 => x"2e893874",
           530 => x"832eae38",
           531 => x"80d53974",
           532 => x"54761083",
           533 => x"fe065376",
           534 => x"882a8c17",
           535 => x"08055288",
           536 => x"3d705255",
           537 => x"fdbd3f88",
           538 => x"08b93874",
           539 => x"51fef83f",
           540 => x"880883ff",
           541 => x"ff0655ad",
           542 => x"39845476",
           543 => x"822b83fc",
           544 => x"06537687",
           545 => x"2a8c1708",
           546 => x"0552883d",
           547 => x"705255fd",
           548 => x"923f8808",
           549 => x"8e387451",
           550 => x"fee23f88",
           551 => x"08f00a06",
           552 => x"55833981",
           553 => x"5574880c",
           554 => x"893d0d04",
           555 => x"fb3d0d0b",
           556 => x"0b0b9fac",
           557 => x"08fe1988",
           558 => x"1208fe05",
           559 => x"55565480",
           560 => x"56747327",
           561 => x"8d388214",
           562 => x"33757129",
           563 => x"94160805",
           564 => x"57537588",
           565 => x"0c873d0d",
           566 => x"04fd3d0d",
           567 => x"7554800b",
           568 => x"0b0b0b9f",
           569 => x"ac087033",
           570 => x"51535371",
           571 => x"832e0981",
           572 => x"068c3894",
           573 => x"1451fdef",
           574 => x"3f880890",
           575 => x"2b539a14",
           576 => x"51fde43f",
           577 => x"880883ff",
           578 => x"ff067307",
           579 => x"880c853d",
           580 => x"0d04fc3d",
           581 => x"0d760b0b",
           582 => x"0b9fac08",
           583 => x"55558075",
           584 => x"23881508",
           585 => x"5372812e",
           586 => x"88388814",
           587 => x"08732685",
           588 => x"388152b0",
           589 => x"39729038",
           590 => x"73335271",
           591 => x"832e0981",
           592 => x"06853890",
           593 => x"14085372",
           594 => x"8c160c72",
           595 => x"802e8b38",
           596 => x"7251fed8",
           597 => x"3f880852",
           598 => x"85399014",
           599 => x"08527190",
           600 => x"160c8052",
           601 => x"71880c86",
           602 => x"3d0d04fa",
           603 => x"3d0d780b",
           604 => x"0b0b9fac",
           605 => x"08712281",
           606 => x"057083ff",
           607 => x"ff065754",
           608 => x"57557380",
           609 => x"2e883890",
           610 => x"15085372",
           611 => x"86388352",
           612 => x"80dc3973",
           613 => x"8f065271",
           614 => x"80cf3881",
           615 => x"1390160c",
           616 => x"8c150853",
           617 => x"728f3883",
           618 => x"0b841722",
           619 => x"57527376",
           620 => x"27bc38b5",
           621 => x"39821633",
           622 => x"ff057484",
           623 => x"2a065271",
           624 => x"a8387251",
           625 => x"fcdf3f81",
           626 => x"52718808",
           627 => x"27a03883",
           628 => x"52880888",
           629 => x"17082796",
           630 => x"3888088c",
           631 => x"160c8808",
           632 => x"51fdc93f",
           633 => x"88089016",
           634 => x"0c737523",
           635 => x"80527188",
           636 => x"0c883d0d",
           637 => x"04f23d0d",
           638 => x"60626458",
           639 => x"5e5c7533",
           640 => x"5574a02e",
           641 => x"09810688",
           642 => x"38811670",
           643 => x"4456ef39",
           644 => x"62703356",
           645 => x"5674af2e",
           646 => x"09810684",
           647 => x"38811643",
           648 => x"800b881d",
           649 => x"0c627033",
           650 => x"5155749f",
           651 => x"268f387b",
           652 => x"51fddf3f",
           653 => x"88085680",
           654 => x"7d3482d3",
           655 => x"39933d84",
           656 => x"1d087058",
           657 => x"5a5f8a55",
           658 => x"a0767081",
           659 => x"055834ff",
           660 => x"155574ff",
           661 => x"2e098106",
           662 => x"ef388070",
           663 => x"595b887f",
           664 => x"085f5a7a",
           665 => x"811c7081",
           666 => x"ff066013",
           667 => x"703370af",
           668 => x"327030a0",
           669 => x"73277180",
           670 => x"25075151",
           671 => x"525b535d",
           672 => x"57557480",
           673 => x"c73876ae",
           674 => x"2e098106",
           675 => x"83388155",
           676 => x"777a2775",
           677 => x"07557480",
           678 => x"2e9f3879",
           679 => x"88327030",
           680 => x"78ae3270",
           681 => x"30707307",
           682 => x"9f2a5351",
           683 => x"57515675",
           684 => x"9b388858",
           685 => x"8b5affab",
           686 => x"39778119",
           687 => x"7081ff06",
           688 => x"721c535a",
           689 => x"57557675",
           690 => x"34ff9839",
           691 => x"7a1e7f0c",
           692 => x"805576a0",
           693 => x"26833881",
           694 => x"55748b1a",
           695 => x"347b51fc",
           696 => x"b13f8808",
           697 => x"80ef38a0",
           698 => x"547b2270",
           699 => x"852b83e0",
           700 => x"06545590",
           701 => x"1c08527c",
           702 => x"51f8a83f",
           703 => x"88085788",
           704 => x"0880fb38",
           705 => x"7c335574",
           706 => x"802e80ee",
           707 => x"388b1d33",
           708 => x"70832a70",
           709 => x"81065156",
           710 => x"5674b238",
           711 => x"8b7d841e",
           712 => x"08880859",
           713 => x"5b5b58ff",
           714 => x"185877ff",
           715 => x"2e9a3879",
           716 => x"7081055b",
           717 => x"33797081",
           718 => x"055b3371",
           719 => x"71315256",
           720 => x"5675802e",
           721 => x"e2388639",
           722 => x"75802e92",
           723 => x"387b51fc",
           724 => x"9a3fff8e",
           725 => x"39880856",
           726 => x"8808b438",
           727 => x"83397656",
           728 => x"841c088b",
           729 => x"11335155",
           730 => x"74a5388b",
           731 => x"1d337084",
           732 => x"2a708106",
           733 => x"51565674",
           734 => x"89388356",
           735 => x"92398156",
           736 => x"8e397c51",
           737 => x"fad33f88",
           738 => x"08881d0c",
           739 => x"fdaf3975",
           740 => x"880c903d",
           741 => x"0d04f93d",
           742 => x"0d797b59",
           743 => x"57825483",
           744 => x"fe537752",
           745 => x"7651f6fb",
           746 => x"3f835688",
           747 => x"0880e738",
           748 => x"7651f8b3",
           749 => x"3f880883",
           750 => x"ffff0655",
           751 => x"82567482",
           752 => x"d4d52e09",
           753 => x"810680ce",
           754 => x"387554b6",
           755 => x"53775276",
           756 => x"51f6d03f",
           757 => x"88085688",
           758 => x"08943876",
           759 => x"51f8883f",
           760 => x"880883ff",
           761 => x"ff065574",
           762 => x"8182c62e",
           763 => x"a9388254",
           764 => x"80d25377",
           765 => x"527651f6",
           766 => x"aa3f8808",
           767 => x"56880894",
           768 => x"387651f7",
           769 => x"e23f8808",
           770 => x"83ffff06",
           771 => x"55748182",
           772 => x"c62e8338",
           773 => x"81567588",
           774 => x"0c893d0d",
           775 => x"04ed3d0d",
           776 => x"6559800b",
           777 => x"0b0b0b9f",
           778 => x"ac0cf59b",
           779 => x"3f880881",
           780 => x"06558256",
           781 => x"7482f238",
           782 => x"7475538d",
           783 => x"3d705357",
           784 => x"5afed33f",
           785 => x"880881ff",
           786 => x"06577681",
           787 => x"2e098106",
           788 => x"b3389054",
           789 => x"83be5374",
           790 => x"527551f5",
           791 => x"c63f8808",
           792 => x"ab388d3d",
           793 => x"33557480",
           794 => x"2eac3895",
           795 => x"3de40551",
           796 => x"f78a3f88",
           797 => x"08880853",
           798 => x"76525afe",
           799 => x"993f8808",
           800 => x"81ff0657",
           801 => x"76832e09",
           802 => x"81068638",
           803 => x"81568299",
           804 => x"3976802e",
           805 => x"86388656",
           806 => x"828f39a4",
           807 => x"548d5379",
           808 => x"527551f4",
           809 => x"fe3f8156",
           810 => x"880881fd",
           811 => x"38953de5",
           812 => x"0551f6b3",
           813 => x"3f880883",
           814 => x"ffff0658",
           815 => x"778c3895",
           816 => x"3df30551",
           817 => x"f6b63f88",
           818 => x"085802af",
           819 => x"05337871",
           820 => x"29028805",
           821 => x"ad057054",
           822 => x"52595bf6",
           823 => x"8a3f8808",
           824 => x"83ffff06",
           825 => x"7a058c1a",
           826 => x"0c8c3d33",
           827 => x"821a3495",
           828 => x"3de00551",
           829 => x"f5f13f88",
           830 => x"08841a23",
           831 => x"953de205",
           832 => x"51f5e43f",
           833 => x"880883ff",
           834 => x"ff065675",
           835 => x"8c38953d",
           836 => x"ef0551f5",
           837 => x"e73f8808",
           838 => x"567a51f5",
           839 => x"ca3f8808",
           840 => x"83ffff06",
           841 => x"76713179",
           842 => x"31841b22",
           843 => x"70842a82",
           844 => x"1d335672",
           845 => x"71315559",
           846 => x"5c5155ee",
           847 => x"c43f8808",
           848 => x"82057088",
           849 => x"1b0c8808",
           850 => x"e08a0556",
           851 => x"567483df",
           852 => x"fe268338",
           853 => x"825783ff",
           854 => x"f6762785",
           855 => x"38835789",
           856 => x"39865676",
           857 => x"802e80c1",
           858 => x"38767934",
           859 => x"76832e09",
           860 => x"81069038",
           861 => x"953dfb05",
           862 => x"51f5813f",
           863 => x"8808901a",
           864 => x"0c88398c",
           865 => x"19081890",
           866 => x"1a0c7983",
           867 => x"ffff068c",
           868 => x"1a081971",
           869 => x"842a0594",
           870 => x"1b0c5580",
           871 => x"0b811a34",
           872 => x"780b0b0b",
           873 => x"9fac0c80",
           874 => x"5675880c",
           875 => x"953d0d04",
           876 => x"ea3d0d0b",
           877 => x"0b0b9fac",
           878 => x"08558554",
           879 => x"74802e80",
           880 => x"df38800b",
           881 => x"81163498",
           882 => x"3de01145",
           883 => x"6954893d",
           884 => x"705457ec",
           885 => x"0551f89d",
           886 => x"3f880854",
           887 => x"880880c0",
           888 => x"38883d33",
           889 => x"5473802e",
           890 => x"933802a7",
           891 => x"05337084",
           892 => x"2a708106",
           893 => x"51555773",
           894 => x"802e8538",
           895 => x"8354a139",
           896 => x"7551f5d5",
           897 => x"3f8808a0",
           898 => x"160c983d",
           899 => x"dc0551f3",
           900 => x"eb3f8808",
           901 => x"9c160c73",
           902 => x"98160c81",
           903 => x"0b811634",
           904 => x"73880c98",
           905 => x"3d0d04f6",
           906 => x"3d0d7d7f",
           907 => x"7e0b0b0b",
           908 => x"9fac0859",
           909 => x"5b5c5880",
           910 => x"7b0c8557",
           911 => x"75802e81",
           912 => x"d1388116",
           913 => x"33810655",
           914 => x"84577480",
           915 => x"2e81c338",
           916 => x"91397481",
           917 => x"17348639",
           918 => x"800b8117",
           919 => x"34815781",
           920 => x"b1399c16",
           921 => x"08981708",
           922 => x"31557478",
           923 => x"27833874",
           924 => x"5877802e",
           925 => x"819a3898",
           926 => x"16087083",
           927 => x"ff065657",
           928 => x"7480c738",
           929 => x"821633ff",
           930 => x"0577892a",
           931 => x"067081ff",
           932 => x"065b5579",
           933 => x"9e387687",
           934 => x"38a01608",
           935 => x"558b39a4",
           936 => x"160851f3",
           937 => x"803f8808",
           938 => x"55817527",
           939 => x"ffaa3874",
           940 => x"a4170ca4",
           941 => x"160851f3",
           942 => x"f33f8808",
           943 => x"55880880",
           944 => x"2eff8f38",
           945 => x"88081aa8",
           946 => x"170c9816",
           947 => x"0883ff06",
           948 => x"84807131",
           949 => x"51557775",
           950 => x"27833877",
           951 => x"55745498",
           952 => x"160883ff",
           953 => x"0653a816",
           954 => x"08527851",
           955 => x"f0b53f88",
           956 => x"08fee538",
           957 => x"98160815",
           958 => x"98170c77",
           959 => x"75317b08",
           960 => x"167c0c58",
           961 => x"78802efe",
           962 => x"e8387419",
           963 => x"59fee239",
           964 => x"80577688",
           965 => x"0c8c3d0d",
           966 => x"04fb3d0d",
           967 => x"9b9086e4",
           968 => x"0b87c094",
           969 => x"8c0c9b90",
           970 => x"86e40b87",
           971 => x"c0949c0c",
           972 => x"8c80830b",
           973 => x"87c09484",
           974 => x"0c8c8083",
           975 => x"0b87c094",
           976 => x"940c9fb0",
           977 => x"51f9d63f",
           978 => x"8808b838",
           979 => x"9f9851fc",
           980 => x"df3f8808",
           981 => x"ae38a080",
           982 => x"0b880887",
           983 => x"c098880c",
           984 => x"55873dfc",
           985 => x"05538480",
           986 => x"527451fd",
           987 => x"ba3f8808",
           988 => x"8d387554",
           989 => x"73802e86",
           990 => x"38731555",
           991 => x"e439a080",
           992 => x"54730480",
           993 => x"54fb3900",
           994 => x"00ffffff",
           995 => x"ff00ffff",
           996 => x"ffff00ff",
           997 => x"ffffff00",
           998 => x"424f4f54",
           999 => x"54494e59",
          1000 => x"2e524f4d",
          1001 => x"00000000",
          1002 => x"01000000",
          2048 => x"0b0b0b88",
          2049 => x"800b0b0b",
          2050 => x"0b8eae04",
          2051 => x"ffffffff",
          2052 => x"ffffffff",
          2053 => x"ffffffff",
          2054 => x"ffffffff",
          2055 => x"ffffffff",
          2056 => x"0b0b0b88",
          2057 => x"80040b0b",
          2058 => x"0b888404",
          2059 => x"0b0b0b88",
          2060 => x"94040b0b",
          2061 => x"0b88a404",
          2062 => x"0b0b0b88",
          2063 => x"b4040b0b",
          2064 => x"0b88c404",
          2065 => x"0b0b0b88",
          2066 => x"d4040b0b",
          2067 => x"0b88e404",
          2068 => x"0b0b0b88",
          2069 => x"f4040b0b",
          2070 => x"0b898404",
          2071 => x"0b0b0b89",
          2072 => x"94040b0b",
          2073 => x"0b89a404",
          2074 => x"0b0b0b89",
          2075 => x"b4040b0b",
          2076 => x"0b89c404",
          2077 => x"0b0b0b89",
          2078 => x"d4040b0b",
          2079 => x"0b89e404",
          2080 => x"0b0b0b89",
          2081 => x"f4040b0b",
          2082 => x"0b8a8404",
          2083 => x"0b0b0b8a",
          2084 => x"94040b0b",
          2085 => x"0b8aa504",
          2086 => x"0b0b0b8a",
          2087 => x"b6040b0b",
          2088 => x"0b8ac704",
          2089 => x"0b0b0b8a",
          2090 => x"d8040b0b",
          2091 => x"0b8ae904",
          2092 => x"0b0b0b8a",
          2093 => x"fa040b0b",
          2094 => x"0b8b8b04",
          2095 => x"0b0b0b8b",
          2096 => x"9c040b0b",
          2097 => x"0b8bad04",
          2098 => x"0b0b0b8b",
          2099 => x"be040b0b",
          2100 => x"0b8bcf04",
          2101 => x"0b0b0b8b",
          2102 => x"e0040b0b",
          2103 => x"0b8bf104",
          2104 => x"0b0b0b8c",
          2105 => x"82040b0b",
          2106 => x"0b8c9304",
          2107 => x"0b0b0b8c",
          2108 => x"a4040b0b",
          2109 => x"0b8cb504",
          2110 => x"0b0b0b8c",
          2111 => x"c6040b0b",
          2112 => x"0b8cd704",
          2113 => x"0b0b0b8c",
          2114 => x"e8040b0b",
          2115 => x"0b8cf904",
          2116 => x"0b0b0b8d",
          2117 => x"8a040b0b",
          2118 => x"0b8d9b04",
          2119 => x"0b0b0b8d",
          2120 => x"ac040b0b",
          2121 => x"0b8dbd04",
          2122 => x"0b0b0b8d",
          2123 => x"cd040b0b",
          2124 => x"0b8ddd04",
          2125 => x"0b0b0b8d",
          2126 => x"ed040b0b",
          2127 => x"0b8dfd04",
          2128 => x"0b0b0b8e",
          2129 => x"8d040b0b",
          2130 => x"0b8e9d04",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"00000000",
          2137 => x"00000000",
          2138 => x"00000000",
          2139 => x"00000000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"00000000",
          2145 => x"00000000",
          2146 => x"00000000",
          2147 => x"00000000",
          2148 => x"00000000",
          2149 => x"00000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"00000000",
          2153 => x"00000000",
          2154 => x"00000000",
          2155 => x"00000000",
          2156 => x"00000000",
          2157 => x"00000000",
          2158 => x"00000000",
          2159 => x"00000000",
          2160 => x"00000000",
          2161 => x"00000000",
          2162 => x"00000000",
          2163 => x"00000000",
          2164 => x"00000000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"00000000",
          2169 => x"00000000",
          2170 => x"00000000",
          2171 => x"00000000",
          2172 => x"00000000",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"00000000",
          2177 => x"00000000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"00000000",
          2185 => x"00000000",
          2186 => x"00000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"00000000",
          2193 => x"00000000",
          2194 => x"00000000",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"00000000",
          2201 => x"00000000",
          2202 => x"00000000",
          2203 => x"00000000",
          2204 => x"00000000",
          2205 => x"00000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"00000000",
          2209 => x"00000000",
          2210 => x"00000000",
          2211 => x"00000000",
          2212 => x"00000000",
          2213 => x"00000000",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"00000000",
          2217 => x"00000000",
          2218 => x"00000000",
          2219 => x"00000000",
          2220 => x"00000000",
          2221 => x"00000000",
          2222 => x"00000000",
          2223 => x"00000000",
          2224 => x"00000000",
          2225 => x"00000000",
          2226 => x"00000000",
          2227 => x"00000000",
          2228 => x"00000000",
          2229 => x"00000000",
          2230 => x"00000000",
          2231 => x"00000000",
          2232 => x"00000000",
          2233 => x"00000000",
          2234 => x"00000000",
          2235 => x"00000000",
          2236 => x"00000000",
          2237 => x"00000000",
          2238 => x"00000000",
          2239 => x"00000000",
          2240 => x"00000000",
          2241 => x"00000000",
          2242 => x"00000000",
          2243 => x"00000000",
          2244 => x"00000000",
          2245 => x"00000000",
          2246 => x"00000000",
          2247 => x"00000000",
          2248 => x"00000000",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"00000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"00000000",
          2265 => x"00000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"00000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"00000000",
          2281 => x"00000000",
          2282 => x"00000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"00000000",
          2297 => x"00000000",
          2298 => x"00000000",
          2299 => x"00000000",
          2300 => x"00000000",
          2301 => x"00000000",
          2302 => x"00000000",
          2303 => x"00000000",
          2304 => x"00888004",
          2305 => x"81cbe00c",
          2306 => x"98f62d81",
          2307 => x"cbe00888",
          2308 => x"80809004",
          2309 => x"81cbe00c",
          2310 => x"a3a62d81",
          2311 => x"cbe00888",
          2312 => x"80809004",
          2313 => x"81cbe00c",
          2314 => x"a3e52d81",
          2315 => x"cbe00888",
          2316 => x"80809004",
          2317 => x"81cbe00c",
          2318 => x"a4832d81",
          2319 => x"cbe00888",
          2320 => x"80809004",
          2321 => x"81cbe00c",
          2322 => x"aac12d81",
          2323 => x"cbe00888",
          2324 => x"80809004",
          2325 => x"81cbe00c",
          2326 => x"abbf2d81",
          2327 => x"cbe00888",
          2328 => x"80809004",
          2329 => x"81cbe00c",
          2330 => x"a4a62d81",
          2331 => x"cbe00888",
          2332 => x"80809004",
          2333 => x"81cbe00c",
          2334 => x"abdc2d81",
          2335 => x"cbe00888",
          2336 => x"80809004",
          2337 => x"81cbe00c",
          2338 => x"adce2d81",
          2339 => x"cbe00888",
          2340 => x"80809004",
          2341 => x"81cbe00c",
          2342 => x"a9e72d81",
          2343 => x"cbe00888",
          2344 => x"80809004",
          2345 => x"81cbe00c",
          2346 => x"a9fd2d81",
          2347 => x"cbe00888",
          2348 => x"80809004",
          2349 => x"81cbe00c",
          2350 => x"aaa12d81",
          2351 => x"cbe00888",
          2352 => x"80809004",
          2353 => x"81cbe00c",
          2354 => x"9b832d81",
          2355 => x"cbe00888",
          2356 => x"80809004",
          2357 => x"81cbe00c",
          2358 => x"9bd42d81",
          2359 => x"cbe00888",
          2360 => x"80809004",
          2361 => x"81cbe00c",
          2362 => x"93f02d81",
          2363 => x"cbe00888",
          2364 => x"80809004",
          2365 => x"81cbe00c",
          2366 => x"95a52d81",
          2367 => x"cbe00888",
          2368 => x"80809004",
          2369 => x"81cbe00c",
          2370 => x"96d82d81",
          2371 => x"cbe00888",
          2372 => x"80809004",
          2373 => x"81cbe00c",
          2374 => x"80e0832d",
          2375 => x"81cbe008",
          2376 => x"88808090",
          2377 => x"0481cbe0",
          2378 => x"0c80ecf4",
          2379 => x"2d81cbe0",
          2380 => x"08888080",
          2381 => x"900481cb",
          2382 => x"e00c80e4",
          2383 => x"e82d81cb",
          2384 => x"e0088880",
          2385 => x"80900481",
          2386 => x"cbe00c80",
          2387 => x"e7e52d81",
          2388 => x"cbe00888",
          2389 => x"80809004",
          2390 => x"81cbe00c",
          2391 => x"80f2832d",
          2392 => x"81cbe008",
          2393 => x"88808090",
          2394 => x"0481cbe0",
          2395 => x"0c80fae3",
          2396 => x"2d81cbe0",
          2397 => x"08888080",
          2398 => x"900481cb",
          2399 => x"e00c80eb",
          2400 => x"d62d81cb",
          2401 => x"e0088880",
          2402 => x"80900481",
          2403 => x"cbe00c80",
          2404 => x"f5a22d81",
          2405 => x"cbe00888",
          2406 => x"80809004",
          2407 => x"81cbe00c",
          2408 => x"80f6c12d",
          2409 => x"81cbe008",
          2410 => x"88808090",
          2411 => x"0481cbe0",
          2412 => x"0c80f6e0",
          2413 => x"2d81cbe0",
          2414 => x"08888080",
          2415 => x"900481cb",
          2416 => x"e00c80fe",
          2417 => x"ca2d81cb",
          2418 => x"e0088880",
          2419 => x"80900481",
          2420 => x"cbe00c80",
          2421 => x"fcb02d81",
          2422 => x"cbe00888",
          2423 => x"80809004",
          2424 => x"81cbe00c",
          2425 => x"81819e2d",
          2426 => x"81cbe008",
          2427 => x"88808090",
          2428 => x"0481cbe0",
          2429 => x"0c80f7e4",
          2430 => x"2d81cbe0",
          2431 => x"08888080",
          2432 => x"900481cb",
          2433 => x"e00c8184",
          2434 => x"9e2d81cb",
          2435 => x"e0088880",
          2436 => x"80900481",
          2437 => x"cbe00c81",
          2438 => x"859f2d81",
          2439 => x"cbe00888",
          2440 => x"80809004",
          2441 => x"81cbe00c",
          2442 => x"80edd42d",
          2443 => x"81cbe008",
          2444 => x"88808090",
          2445 => x"0481cbe0",
          2446 => x"0c80edad",
          2447 => x"2d81cbe0",
          2448 => x"08888080",
          2449 => x"900481cb",
          2450 => x"e00c80ee",
          2451 => x"d82d81cb",
          2452 => x"e0088880",
          2453 => x"80900481",
          2454 => x"cbe00c80",
          2455 => x"f8bb2d81",
          2456 => x"cbe00888",
          2457 => x"80809004",
          2458 => x"81cbe00c",
          2459 => x"8186902d",
          2460 => x"81cbe008",
          2461 => x"88808090",
          2462 => x"0481cbe0",
          2463 => x"0c81889a",
          2464 => x"2d81cbe0",
          2465 => x"08888080",
          2466 => x"900481cb",
          2467 => x"e00c818b",
          2468 => x"dc2d81cb",
          2469 => x"e0088880",
          2470 => x"80900481",
          2471 => x"cbe00c80",
          2472 => x"dfa22d81",
          2473 => x"cbe00888",
          2474 => x"80809004",
          2475 => x"81cbe00c",
          2476 => x"818ec82d",
          2477 => x"81cbe008",
          2478 => x"88808090",
          2479 => x"0481cbe0",
          2480 => x"0cb0dd2d",
          2481 => x"81cbe008",
          2482 => x"88808090",
          2483 => x"0481cbe0",
          2484 => x"0cb2c72d",
          2485 => x"81cbe008",
          2486 => x"88808090",
          2487 => x"0481cbe0",
          2488 => x"0cb4ab2d",
          2489 => x"81cbe008",
          2490 => x"88808090",
          2491 => x"0481cbe0",
          2492 => x"0c94992d",
          2493 => x"81cbe008",
          2494 => x"88808090",
          2495 => x"0481cbe0",
          2496 => x"0c94fb2d",
          2497 => x"81cbe008",
          2498 => x"88808090",
          2499 => x"0481cbe0",
          2500 => x"0c97e82d",
          2501 => x"81cbe008",
          2502 => x"88808090",
          2503 => x"0481cbe0",
          2504 => x"0c819ae9",
          2505 => x"2d81cbe0",
          2506 => x"08888080",
          2507 => x"900481cb",
          2508 => x"d47081e2",
          2509 => x"d8278e38",
          2510 => x"80717084",
          2511 => x"05530c0b",
          2512 => x"0b0b8eb1",
          2513 => x"04888051",
          2514 => x"81b4bd04",
          2515 => x"3c0481cb",
          2516 => x"e0080281",
          2517 => x"cbe00cfd",
          2518 => x"3d0d8053",
          2519 => x"81cbe008",
          2520 => x"8c050852",
          2521 => x"81cbe008",
          2522 => x"88050851",
          2523 => x"80c53f81",
          2524 => x"cbd40870",
          2525 => x"81cbd40c",
          2526 => x"54853d0d",
          2527 => x"81cbe00c",
          2528 => x"0481cbe0",
          2529 => x"080281cb",
          2530 => x"e00cfd3d",
          2531 => x"0d815381",
          2532 => x"cbe0088c",
          2533 => x"05085281",
          2534 => x"cbe00888",
          2535 => x"05085193",
          2536 => x"3f81cbd4",
          2537 => x"087081cb",
          2538 => x"d40c5485",
          2539 => x"3d0d81cb",
          2540 => x"e00c0481",
          2541 => x"cbe00802",
          2542 => x"81cbe00c",
          2543 => x"fd3d0d81",
          2544 => x"0b81cbe0",
          2545 => x"08fc050c",
          2546 => x"800b81cb",
          2547 => x"e008f805",
          2548 => x"0c81cbe0",
          2549 => x"088c0508",
          2550 => x"81cbe008",
          2551 => x"88050827",
          2552 => x"b93881cb",
          2553 => x"e008fc05",
          2554 => x"08802eae",
          2555 => x"38800b81",
          2556 => x"cbe0088c",
          2557 => x"050824a2",
          2558 => x"3881cbe0",
          2559 => x"088c0508",
          2560 => x"1081cbe0",
          2561 => x"088c050c",
          2562 => x"81cbe008",
          2563 => x"fc050810",
          2564 => x"81cbe008",
          2565 => x"fc050cff",
          2566 => x"b83981cb",
          2567 => x"e008fc05",
          2568 => x"08802e80",
          2569 => x"e13881cb",
          2570 => x"e0088c05",
          2571 => x"0881cbe0",
          2572 => x"08880508",
          2573 => x"26ad3881",
          2574 => x"cbe00888",
          2575 => x"050881cb",
          2576 => x"e0088c05",
          2577 => x"083181cb",
          2578 => x"e0088805",
          2579 => x"0c81cbe0",
          2580 => x"08f80508",
          2581 => x"81cbe008",
          2582 => x"fc050807",
          2583 => x"81cbe008",
          2584 => x"f8050c81",
          2585 => x"cbe008fc",
          2586 => x"0508812a",
          2587 => x"81cbe008",
          2588 => x"fc050c81",
          2589 => x"cbe0088c",
          2590 => x"0508812a",
          2591 => x"81cbe008",
          2592 => x"8c050cff",
          2593 => x"953981cb",
          2594 => x"e0089005",
          2595 => x"08802e93",
          2596 => x"3881cbe0",
          2597 => x"08880508",
          2598 => x"7081cbe0",
          2599 => x"08f4050c",
          2600 => x"51913981",
          2601 => x"cbe008f8",
          2602 => x"05087081",
          2603 => x"cbe008f4",
          2604 => x"050c5181",
          2605 => x"cbe008f4",
          2606 => x"050881cb",
          2607 => x"d40c853d",
          2608 => x"0d81cbe0",
          2609 => x"0c04fc3d",
          2610 => x"0d767971",
          2611 => x"028c059f",
          2612 => x"05335755",
          2613 => x"53558372",
          2614 => x"278a3874",
          2615 => x"83065170",
          2616 => x"802ea438",
          2617 => x"ff125271",
          2618 => x"ff2e9338",
          2619 => x"73737081",
          2620 => x"055534ff",
          2621 => x"125271ff",
          2622 => x"2e098106",
          2623 => x"ef387481",
          2624 => x"cbd40c86",
          2625 => x"3d0d0474",
          2626 => x"74882b75",
          2627 => x"07707190",
          2628 => x"2b075154",
          2629 => x"518f7227",
          2630 => x"a5387271",
          2631 => x"70840553",
          2632 => x"0c727170",
          2633 => x"8405530c",
          2634 => x"72717084",
          2635 => x"05530c72",
          2636 => x"71708405",
          2637 => x"530cf012",
          2638 => x"52718f26",
          2639 => x"dd388372",
          2640 => x"27903872",
          2641 => x"71708405",
          2642 => x"530cfc12",
          2643 => x"52718326",
          2644 => x"f2387053",
          2645 => x"ff8e39fb",
          2646 => x"3d0d7779",
          2647 => x"70720783",
          2648 => x"06535452",
          2649 => x"70933871",
          2650 => x"73730854",
          2651 => x"56547173",
          2652 => x"082e80c6",
          2653 => x"38737554",
          2654 => x"52713370",
          2655 => x"81ff0652",
          2656 => x"5470802e",
          2657 => x"9d387233",
          2658 => x"5570752e",
          2659 => x"09810695",
          2660 => x"38811281",
          2661 => x"14713370",
          2662 => x"81ff0654",
          2663 => x"56545270",
          2664 => x"e5387233",
          2665 => x"557381ff",
          2666 => x"067581ff",
          2667 => x"06717131",
          2668 => x"81cbd40c",
          2669 => x"5252873d",
          2670 => x"0d047109",
          2671 => x"70f7fbfd",
          2672 => x"ff140670",
          2673 => x"f8848281",
          2674 => x"80065151",
          2675 => x"51709738",
          2676 => x"84148416",
          2677 => x"71085456",
          2678 => x"54717508",
          2679 => x"2edc3873",
          2680 => x"755452ff",
          2681 => x"9439800b",
          2682 => x"81cbd40c",
          2683 => x"873d0d04",
          2684 => x"fe3d0d80",
          2685 => x"52835371",
          2686 => x"882b5287",
          2687 => x"863f81cb",
          2688 => x"d40881ff",
          2689 => x"067207ff",
          2690 => x"14545272",
          2691 => x"8025e838",
          2692 => x"7181cbd4",
          2693 => x"0c843d0d",
          2694 => x"04fb3d0d",
          2695 => x"77700870",
          2696 => x"53535671",
          2697 => x"802e80ca",
          2698 => x"38713351",
          2699 => x"70a02e09",
          2700 => x"81068638",
          2701 => x"811252f1",
          2702 => x"39715384",
          2703 => x"39811353",
          2704 => x"80733370",
          2705 => x"81ff0653",
          2706 => x"555570a0",
          2707 => x"2e833881",
          2708 => x"5570802e",
          2709 => x"843874e5",
          2710 => x"387381ff",
          2711 => x"065170a0",
          2712 => x"2e098106",
          2713 => x"88388073",
          2714 => x"70810555",
          2715 => x"3472760c",
          2716 => x"71517081",
          2717 => x"cbd40c87",
          2718 => x"3d0d04fc",
          2719 => x"3d0d7653",
          2720 => x"7208802e",
          2721 => x"9138863d",
          2722 => x"fc055272",
          2723 => x"5198bf3f",
          2724 => x"81cbd408",
          2725 => x"85388053",
          2726 => x"83397453",
          2727 => x"7281cbd4",
          2728 => x"0c863d0d",
          2729 => x"04fc3d0d",
          2730 => x"76821133",
          2731 => x"ff055253",
          2732 => x"8152708b",
          2733 => x"26819838",
          2734 => x"831333ff",
          2735 => x"05518252",
          2736 => x"709e2681",
          2737 => x"8a388413",
          2738 => x"33518352",
          2739 => x"70972680",
          2740 => x"fe388513",
          2741 => x"33518452",
          2742 => x"70bb2680",
          2743 => x"f2388613",
          2744 => x"33518552",
          2745 => x"70bb2680",
          2746 => x"e6388813",
          2747 => x"22558652",
          2748 => x"7487e726",
          2749 => x"80d9388a",
          2750 => x"13225487",
          2751 => x"527387e7",
          2752 => x"2680cc38",
          2753 => x"810b87c0",
          2754 => x"989c0c72",
          2755 => x"2287c098",
          2756 => x"bc0c8213",
          2757 => x"3387c098",
          2758 => x"b80c8313",
          2759 => x"3387c098",
          2760 => x"b40c8413",
          2761 => x"3387c098",
          2762 => x"b00c8513",
          2763 => x"3387c098",
          2764 => x"ac0c8613",
          2765 => x"3387c098",
          2766 => x"a80c7487",
          2767 => x"c098a40c",
          2768 => x"7387c098",
          2769 => x"a00c800b",
          2770 => x"87c0989c",
          2771 => x"0c805271",
          2772 => x"81cbd40c",
          2773 => x"863d0d04",
          2774 => x"f33d0d7f",
          2775 => x"5b87c098",
          2776 => x"9c5d817d",
          2777 => x"0c87c098",
          2778 => x"bc085e7d",
          2779 => x"7b2387c0",
          2780 => x"98b8085a",
          2781 => x"79821c34",
          2782 => x"87c098b4",
          2783 => x"085a7983",
          2784 => x"1c3487c0",
          2785 => x"98b0085a",
          2786 => x"79841c34",
          2787 => x"87c098ac",
          2788 => x"085a7985",
          2789 => x"1c3487c0",
          2790 => x"98a8085a",
          2791 => x"79861c34",
          2792 => x"87c098a4",
          2793 => x"085c7b88",
          2794 => x"1c2387c0",
          2795 => x"98a0085a",
          2796 => x"798a1c23",
          2797 => x"807d0c79",
          2798 => x"83ffff06",
          2799 => x"597b83ff",
          2800 => x"ff065886",
          2801 => x"1b335785",
          2802 => x"1b335684",
          2803 => x"1b335583",
          2804 => x"1b335482",
          2805 => x"1b33537d",
          2806 => x"83ffff06",
          2807 => x"5281b688",
          2808 => x"5192843f",
          2809 => x"8f3d0d04",
          2810 => x"ff3d0d02",
          2811 => x"8f053370",
          2812 => x"30709f2a",
          2813 => x"51525270",
          2814 => x"0b0b81c8",
          2815 => x"bc34833d",
          2816 => x"0d04fb3d",
          2817 => x"0d770b0b",
          2818 => x"81c8bc33",
          2819 => x"7081ff06",
          2820 => x"57555687",
          2821 => x"c0948451",
          2822 => x"74802e86",
          2823 => x"3887c094",
          2824 => x"94517008",
          2825 => x"70962a70",
          2826 => x"81065354",
          2827 => x"5270802e",
          2828 => x"8c387191",
          2829 => x"2a708106",
          2830 => x"515170d7",
          2831 => x"38728132",
          2832 => x"70810651",
          2833 => x"5170802e",
          2834 => x"8d387193",
          2835 => x"2a708106",
          2836 => x"515170ff",
          2837 => x"be387381",
          2838 => x"ff065187",
          2839 => x"c0948052",
          2840 => x"70802e86",
          2841 => x"3887c094",
          2842 => x"90527572",
          2843 => x"0c7581cb",
          2844 => x"d40c873d",
          2845 => x"0d04fb3d",
          2846 => x"0d029f05",
          2847 => x"330b0b81",
          2848 => x"c8bc3370",
          2849 => x"81ff0657",
          2850 => x"555687c0",
          2851 => x"94845174",
          2852 => x"802e8638",
          2853 => x"87c09494",
          2854 => x"51700870",
          2855 => x"962a7081",
          2856 => x"06535452",
          2857 => x"70802e8c",
          2858 => x"3871912a",
          2859 => x"70810651",
          2860 => x"5170d738",
          2861 => x"72813270",
          2862 => x"81065151",
          2863 => x"70802e8d",
          2864 => x"3871932a",
          2865 => x"70810651",
          2866 => x"5170ffbe",
          2867 => x"387381ff",
          2868 => x"065187c0",
          2869 => x"94805270",
          2870 => x"802e8638",
          2871 => x"87c09490",
          2872 => x"5275720c",
          2873 => x"873d0d04",
          2874 => x"f93d0d79",
          2875 => x"54807433",
          2876 => x"7081ff06",
          2877 => x"53535770",
          2878 => x"772e80fe",
          2879 => x"387181ff",
          2880 => x"0681150b",
          2881 => x"0b81c8bc",
          2882 => x"337081ff",
          2883 => x"06595755",
          2884 => x"5887c094",
          2885 => x"84517580",
          2886 => x"2e863887",
          2887 => x"c0949451",
          2888 => x"70087096",
          2889 => x"2a708106",
          2890 => x"53545270",
          2891 => x"802e8c38",
          2892 => x"71912a70",
          2893 => x"81065151",
          2894 => x"70d73872",
          2895 => x"81327081",
          2896 => x"06515170",
          2897 => x"802e8d38",
          2898 => x"71932a70",
          2899 => x"81065151",
          2900 => x"70ffbe38",
          2901 => x"7481ff06",
          2902 => x"5187c094",
          2903 => x"80527080",
          2904 => x"2e863887",
          2905 => x"c0949052",
          2906 => x"77720c81",
          2907 => x"17743370",
          2908 => x"81ff0653",
          2909 => x"535770ff",
          2910 => x"84387681",
          2911 => x"cbd40c89",
          2912 => x"3d0d04fe",
          2913 => x"3d0d0b0b",
          2914 => x"81c8bc33",
          2915 => x"7081ff06",
          2916 => x"545287c0",
          2917 => x"94845172",
          2918 => x"802e8638",
          2919 => x"87c09494",
          2920 => x"51700870",
          2921 => x"822a7081",
          2922 => x"06515151",
          2923 => x"70802ee2",
          2924 => x"387181ff",
          2925 => x"065187c0",
          2926 => x"94805270",
          2927 => x"802e8638",
          2928 => x"87c09490",
          2929 => x"52710870",
          2930 => x"81ff0681",
          2931 => x"cbd40c51",
          2932 => x"843d0d04",
          2933 => x"fe3d0d0b",
          2934 => x"0b81c8bc",
          2935 => x"337081ff",
          2936 => x"06525387",
          2937 => x"c0948452",
          2938 => x"70802e86",
          2939 => x"3887c094",
          2940 => x"94527108",
          2941 => x"70822a70",
          2942 => x"81065151",
          2943 => x"51ff5270",
          2944 => x"802ea038",
          2945 => x"7281ff06",
          2946 => x"5187c094",
          2947 => x"80527080",
          2948 => x"2e863887",
          2949 => x"c0949052",
          2950 => x"71087098",
          2951 => x"2b70982c",
          2952 => x"51535171",
          2953 => x"81cbd40c",
          2954 => x"843d0d04",
          2955 => x"ff3d0d87",
          2956 => x"c09e8008",
          2957 => x"709c2a8a",
          2958 => x"06515170",
          2959 => x"802e8393",
          2960 => x"3887c09e",
          2961 => x"9c0881c8",
          2962 => x"c00c87c0",
          2963 => x"9ea00881",
          2964 => x"c8c40c87",
          2965 => x"c09e8c08",
          2966 => x"81c8c80c",
          2967 => x"87c09e90",
          2968 => x"0881c8cc",
          2969 => x"0c87c09e",
          2970 => x"940881c8",
          2971 => x"d00c87c0",
          2972 => x"9e980881",
          2973 => x"c8d40c87",
          2974 => x"c09ea408",
          2975 => x"81c8d80c",
          2976 => x"87c09ea8",
          2977 => x"0881c8dc",
          2978 => x"0c87c09e",
          2979 => x"ac0881c8",
          2980 => x"e00c87c0",
          2981 => x"9e800851",
          2982 => x"7081c8e4",
          2983 => x"2387c09e",
          2984 => x"840881c8",
          2985 => x"e80c810b",
          2986 => x"81c8ec34",
          2987 => x"800b87c0",
          2988 => x"9e880870",
          2989 => x"a0800651",
          2990 => x"52527080",
          2991 => x"2e833881",
          2992 => x"527181c8",
          2993 => x"ed34800b",
          2994 => x"87c09e88",
          2995 => x"08708180",
          2996 => x"80065152",
          2997 => x"5270802e",
          2998 => x"83388152",
          2999 => x"7181c8ee",
          3000 => x"34800b87",
          3001 => x"c09e8808",
          3002 => x"7080c080",
          3003 => x"06515252",
          3004 => x"70802e83",
          3005 => x"38815271",
          3006 => x"81c8ef34",
          3007 => x"800b87c0",
          3008 => x"9e880870",
          3009 => x"90800651",
          3010 => x"52527080",
          3011 => x"2e833881",
          3012 => x"527181c8",
          3013 => x"f034800b",
          3014 => x"87c09e88",
          3015 => x"08708880",
          3016 => x"06515252",
          3017 => x"70802e83",
          3018 => x"38815271",
          3019 => x"81c8f134",
          3020 => x"800b87c0",
          3021 => x"9e880870",
          3022 => x"84800651",
          3023 => x"52527080",
          3024 => x"2e833881",
          3025 => x"527181c8",
          3026 => x"f234800b",
          3027 => x"87c09e88",
          3028 => x"08708280",
          3029 => x"06515252",
          3030 => x"70802e83",
          3031 => x"38815271",
          3032 => x"81c8f334",
          3033 => x"800b87c0",
          3034 => x"9e880870",
          3035 => x"81800651",
          3036 => x"52527080",
          3037 => x"2e833881",
          3038 => x"527181c8",
          3039 => x"f43487c0",
          3040 => x"9e880870",
          3041 => x"80e00670",
          3042 => x"862c5151",
          3043 => x"517081c8",
          3044 => x"f534800b",
          3045 => x"87c09e88",
          3046 => x"08709006",
          3047 => x"51525270",
          3048 => x"802e8338",
          3049 => x"81527181",
          3050 => x"c8f63480",
          3051 => x"0b87c09e",
          3052 => x"88087088",
          3053 => x"06515252",
          3054 => x"70802e83",
          3055 => x"38815271",
          3056 => x"81c8f734",
          3057 => x"87c09e88",
          3058 => x"08708706",
          3059 => x"51517081",
          3060 => x"c8f83483",
          3061 => x"3d0d04fd",
          3062 => x"3d0d81b6",
          3063 => x"a05184a3",
          3064 => x"3f81c8ec",
          3065 => x"33547380",
          3066 => x"2e883881",
          3067 => x"b6b45184",
          3068 => x"923f81b6",
          3069 => x"c851848b",
          3070 => x"3f81c8ed",
          3071 => x"33547380",
          3072 => x"2e923881",
          3073 => x"c8c40853",
          3074 => x"81c8c008",
          3075 => x"5281b6e0",
          3076 => x"5189d43f",
          3077 => x"81c8ee33",
          3078 => x"5473802e",
          3079 => x"923881c8",
          3080 => x"cc085381",
          3081 => x"c8c80852",
          3082 => x"81b78851",
          3083 => x"89b93f81",
          3084 => x"c8ef3354",
          3085 => x"738b3881",
          3086 => x"c8f03354",
          3087 => x"73802e92",
          3088 => x"3881c8d4",
          3089 => x"085381c8",
          3090 => x"d0085281",
          3091 => x"b7ac5189",
          3092 => x"963f81c8",
          3093 => x"f1335473",
          3094 => x"802e8838",
          3095 => x"81b7d051",
          3096 => x"83a13f81",
          3097 => x"c8f23354",
          3098 => x"73802e88",
          3099 => x"3881b7dc",
          3100 => x"5183903f",
          3101 => x"81c8f333",
          3102 => x"5473802e",
          3103 => x"883881b7",
          3104 => x"e85182ff",
          3105 => x"3f81c8f4",
          3106 => x"33547380",
          3107 => x"2e8d3881",
          3108 => x"c8f53352",
          3109 => x"81b7f451",
          3110 => x"88cd3f81",
          3111 => x"c8f63354",
          3112 => x"73802e88",
          3113 => x"3881b894",
          3114 => x"5182d83f",
          3115 => x"81c8f733",
          3116 => x"5473802e",
          3117 => x"8d3881c8",
          3118 => x"f8335281",
          3119 => x"b8b05188",
          3120 => x"a63f81b8",
          3121 => x"cc5182bb",
          3122 => x"3f81c8d8",
          3123 => x"085281b8",
          3124 => x"d8518893",
          3125 => x"3f81c8dc",
          3126 => x"085281b9",
          3127 => x"80518887",
          3128 => x"3f81c8e0",
          3129 => x"085281b9",
          3130 => x"a85187fb",
          3131 => x"3f81c8e4",
          3132 => x"225281b9",
          3133 => x"d05187ef",
          3134 => x"3f81c8e8",
          3135 => x"085281b9",
          3136 => x"f85187e3",
          3137 => x"3f853d0d",
          3138 => x"04fe3d0d",
          3139 => x"02920533",
          3140 => x"ff055271",
          3141 => x"8426ac38",
          3142 => x"7184290b",
          3143 => x"0b81b5a4",
          3144 => x"05527108",
          3145 => x"0481baa0",
          3146 => x"519d3981",
          3147 => x"baa85197",
          3148 => x"3981bab0",
          3149 => x"51913981",
          3150 => x"bab8518b",
          3151 => x"3981babc",
          3152 => x"51853981",
          3153 => x"bac451f7",
          3154 => x"9f3f843d",
          3155 => x"0d047188",
          3156 => x"800c0480",
          3157 => x"0b87c096",
          3158 => x"840c04ff",
          3159 => x"3d0d87c0",
          3160 => x"96847008",
          3161 => x"52528072",
          3162 => x"0c707407",
          3163 => x"7081c8fc",
          3164 => x"0c720c83",
          3165 => x"3d0d04ff",
          3166 => x"3d0d87c0",
          3167 => x"96847008",
          3168 => x"81c8fc0c",
          3169 => x"5280720c",
          3170 => x"73097081",
          3171 => x"c8fc0806",
          3172 => x"7081c8fc",
          3173 => x"0c730c51",
          3174 => x"833d0d04",
          3175 => x"81c8fc08",
          3176 => x"87c09684",
          3177 => x"0c04fe3d",
          3178 => x"0d029305",
          3179 => x"3353728a",
          3180 => x"2e098106",
          3181 => x"85388d51",
          3182 => x"ed3f81cb",
          3183 => x"ec085271",
          3184 => x"802e9038",
          3185 => x"72723481",
          3186 => x"cbec0881",
          3187 => x"0581cbec",
          3188 => x"0c8f3981",
          3189 => x"cbe40852",
          3190 => x"71802e85",
          3191 => x"38725171",
          3192 => x"2d843d0d",
          3193 => x"04fe3d0d",
          3194 => x"02970533",
          3195 => x"81cbe408",
          3196 => x"7681cbe4",
          3197 => x"0c5451ff",
          3198 => x"ad3f7281",
          3199 => x"cbe40c84",
          3200 => x"3d0d04fd",
          3201 => x"3d0d7554",
          3202 => x"73337081",
          3203 => x"ff065353",
          3204 => x"71802e8e",
          3205 => x"387281ff",
          3206 => x"06518114",
          3207 => x"54ff873f",
          3208 => x"e739853d",
          3209 => x"0d04fc3d",
          3210 => x"0d7781cb",
          3211 => x"e4087881",
          3212 => x"cbe40c56",
          3213 => x"54733370",
          3214 => x"81ff0653",
          3215 => x"5371802e",
          3216 => x"8e387281",
          3217 => x"ff065181",
          3218 => x"1454feda",
          3219 => x"3fe73974",
          3220 => x"81cbe40c",
          3221 => x"863d0d04",
          3222 => x"ec3d0d66",
          3223 => x"68595978",
          3224 => x"7081055a",
          3225 => x"33567580",
          3226 => x"2e84f838",
          3227 => x"75a52e09",
          3228 => x"810682de",
          3229 => x"3880707a",
          3230 => x"7081055c",
          3231 => x"33585b5b",
          3232 => x"75b02e09",
          3233 => x"81068538",
          3234 => x"815a8b39",
          3235 => x"75ad2e09",
          3236 => x"81068a38",
          3237 => x"825a7870",
          3238 => x"81055a33",
          3239 => x"5675aa2e",
          3240 => x"09810692",
          3241 => x"38778419",
          3242 => x"71087b70",
          3243 => x"81055d33",
          3244 => x"595d5953",
          3245 => x"9d39d016",
          3246 => x"53728926",
          3247 => x"95387a88",
          3248 => x"297b1005",
          3249 => x"7605d005",
          3250 => x"79708105",
          3251 => x"5b33575b",
          3252 => x"e5397580",
          3253 => x"ec327030",
          3254 => x"70720780",
          3255 => x"257880cc",
          3256 => x"32703070",
          3257 => x"72078025",
          3258 => x"73075354",
          3259 => x"58515553",
          3260 => x"73802e8c",
          3261 => x"38798407",
          3262 => x"79708105",
          3263 => x"5b33575a",
          3264 => x"75802e83",
          3265 => x"de387554",
          3266 => x"80e07627",
          3267 => x"8938e016",
          3268 => x"7081ff06",
          3269 => x"55537380",
          3270 => x"cf2e81aa",
          3271 => x"387380cf",
          3272 => x"24a23873",
          3273 => x"80c32e81",
          3274 => x"8e387380",
          3275 => x"c3248b38",
          3276 => x"7380c22e",
          3277 => x"818c3881",
          3278 => x"99397380",
          3279 => x"c42e818a",
          3280 => x"38818f39",
          3281 => x"7380d52e",
          3282 => x"81803873",
          3283 => x"80d5248a",
          3284 => x"387380d3",
          3285 => x"2e8e3880",
          3286 => x"f9397380",
          3287 => x"d82e80ee",
          3288 => x"3880ef39",
          3289 => x"77841971",
          3290 => x"08565953",
          3291 => x"80743354",
          3292 => x"5572752e",
          3293 => x"8d388115",
          3294 => x"70157033",
          3295 => x"51545572",
          3296 => x"f5387981",
          3297 => x"2a569039",
          3298 => x"74811656",
          3299 => x"53727b27",
          3300 => x"8f38a051",
          3301 => x"fc903f75",
          3302 => x"81065372",
          3303 => x"802ee938",
          3304 => x"7351fcdf",
          3305 => x"3f748116",
          3306 => x"5653727b",
          3307 => x"27fdb038",
          3308 => x"a051fbf2",
          3309 => x"3fef3977",
          3310 => x"84198312",
          3311 => x"33535953",
          3312 => x"9339825c",
          3313 => x"9539885c",
          3314 => x"91398a5c",
          3315 => x"8d39905c",
          3316 => x"89397551",
          3317 => x"fbd03ffd",
          3318 => x"86397982",
          3319 => x"2a708106",
          3320 => x"51537280",
          3321 => x"2e883877",
          3322 => x"84195953",
          3323 => x"86398418",
          3324 => x"78545872",
          3325 => x"087480c4",
          3326 => x"32703070",
          3327 => x"72078025",
          3328 => x"51555555",
          3329 => x"7480258d",
          3330 => x"3872802e",
          3331 => x"88387430",
          3332 => x"7a90075b",
          3333 => x"55800b8f",
          3334 => x"3d5e577b",
          3335 => x"527451e6",
          3336 => x"e03f81cb",
          3337 => x"d40881ff",
          3338 => x"067c5375",
          3339 => x"5254e69e",
          3340 => x"3f81cbd4",
          3341 => x"08558974",
          3342 => x"279238a7",
          3343 => x"14537580",
          3344 => x"f82e8438",
          3345 => x"87145372",
          3346 => x"81ff0654",
          3347 => x"b0145372",
          3348 => x"7d708105",
          3349 => x"5f348117",
          3350 => x"75307077",
          3351 => x"079f2a51",
          3352 => x"5457769f",
          3353 => x"26853872",
          3354 => x"ffb13879",
          3355 => x"842a7081",
          3356 => x"06515372",
          3357 => x"802e8e38",
          3358 => x"963d7705",
          3359 => x"e00553ad",
          3360 => x"73348117",
          3361 => x"57767a81",
          3362 => x"065455b0",
          3363 => x"54728338",
          3364 => x"a0547981",
          3365 => x"2a708106",
          3366 => x"5456729f",
          3367 => x"38811755",
          3368 => x"767b2797",
          3369 => x"387351f9",
          3370 => x"fd3f7581",
          3371 => x"0653728b",
          3372 => x"38748116",
          3373 => x"56537a73",
          3374 => x"26eb3896",
          3375 => x"3d7705e0",
          3376 => x"0553ff17",
          3377 => x"ff147033",
          3378 => x"535457f9",
          3379 => x"d93f76f2",
          3380 => x"38748116",
          3381 => x"5653727b",
          3382 => x"27fb8438",
          3383 => x"a051f9c6",
          3384 => x"3fef3996",
          3385 => x"3d0d04fd",
          3386 => x"3d0d863d",
          3387 => x"70708405",
          3388 => x"52085552",
          3389 => x"7351fae0",
          3390 => x"3f853d0d",
          3391 => x"04fe3d0d",
          3392 => x"7481cbec",
          3393 => x"0c853d88",
          3394 => x"05527551",
          3395 => x"faca3f81",
          3396 => x"cbec0853",
          3397 => x"80733480",
          3398 => x"0b81cbec",
          3399 => x"0c843d0d",
          3400 => x"04fd3d0d",
          3401 => x"81cbe408",
          3402 => x"7681cbe4",
          3403 => x"0c873d88",
          3404 => x"05537752",
          3405 => x"53faa13f",
          3406 => x"7281cbe4",
          3407 => x"0c853d0d",
          3408 => x"04fb3d0d",
          3409 => x"777981cb",
          3410 => x"e8087056",
          3411 => x"54575580",
          3412 => x"5471802e",
          3413 => x"80e03881",
          3414 => x"cbe80852",
          3415 => x"712d81cb",
          3416 => x"d40881ff",
          3417 => x"06537280",
          3418 => x"2e80cb38",
          3419 => x"728d2eb9",
          3420 => x"38728832",
          3421 => x"70307080",
          3422 => x"25515152",
          3423 => x"73802e8b",
          3424 => x"3871802e",
          3425 => x"8638ff14",
          3426 => x"5497399f",
          3427 => x"7325c838",
          3428 => x"ff165273",
          3429 => x"7225c038",
          3430 => x"74145272",
          3431 => x"72348114",
          3432 => x"547251f8",
          3433 => x"813fffaf",
          3434 => x"39731552",
          3435 => x"8072348a",
          3436 => x"51f7f33f",
          3437 => x"81537281",
          3438 => x"cbd40c87",
          3439 => x"3d0d04fe",
          3440 => x"3d0d81cb",
          3441 => x"e8087581",
          3442 => x"cbe80c77",
          3443 => x"53765253",
          3444 => x"feef3f72",
          3445 => x"81cbe80c",
          3446 => x"843d0d04",
          3447 => x"f83d0d7a",
          3448 => x"7c5a5680",
          3449 => x"707a0c58",
          3450 => x"75087033",
          3451 => x"555373a0",
          3452 => x"2e098106",
          3453 => x"87388113",
          3454 => x"760ced39",
          3455 => x"73ad2e09",
          3456 => x"81068e38",
          3457 => x"81760811",
          3458 => x"770c7608",
          3459 => x"70335654",
          3460 => x"5873b02e",
          3461 => x"09810680",
          3462 => x"c2387508",
          3463 => x"8105760c",
          3464 => x"75087033",
          3465 => x"55537380",
          3466 => x"e22e8b38",
          3467 => x"90577380",
          3468 => x"f82e8538",
          3469 => x"8f398257",
          3470 => x"8113760c",
          3471 => x"75087033",
          3472 => x"5553ac39",
          3473 => x"8155a074",
          3474 => x"2780fa38",
          3475 => x"d0145380",
          3476 => x"55885789",
          3477 => x"73279838",
          3478 => x"80eb39d0",
          3479 => x"14538055",
          3480 => x"72892680",
          3481 => x"e0388639",
          3482 => x"805580d9",
          3483 => x"398a5780",
          3484 => x"55a07427",
          3485 => x"80c23880",
          3486 => x"e0742789",
          3487 => x"38e01470",
          3488 => x"81ff0655",
          3489 => x"53d01470",
          3490 => x"81ff0655",
          3491 => x"53907427",
          3492 => x"8e38f914",
          3493 => x"7081ff06",
          3494 => x"55538974",
          3495 => x"27ca3873",
          3496 => x"7727c538",
          3497 => x"74772914",
          3498 => x"76088105",
          3499 => x"770c7608",
          3500 => x"70335654",
          3501 => x"55ffba39",
          3502 => x"77802e84",
          3503 => x"38743055",
          3504 => x"74790c81",
          3505 => x"557481cb",
          3506 => x"d40c8a3d",
          3507 => x"0d04f83d",
          3508 => x"0d7a7c5a",
          3509 => x"5680707a",
          3510 => x"0c587508",
          3511 => x"70335553",
          3512 => x"73a02e09",
          3513 => x"81068738",
          3514 => x"8113760c",
          3515 => x"ed3973ad",
          3516 => x"2e098106",
          3517 => x"8e388176",
          3518 => x"0811770c",
          3519 => x"76087033",
          3520 => x"56545873",
          3521 => x"b02e0981",
          3522 => x"0680c238",
          3523 => x"75088105",
          3524 => x"760c7508",
          3525 => x"70335553",
          3526 => x"7380e22e",
          3527 => x"8b389057",
          3528 => x"7380f82e",
          3529 => x"85388f39",
          3530 => x"82578113",
          3531 => x"760c7508",
          3532 => x"70335553",
          3533 => x"ac398155",
          3534 => x"a0742780",
          3535 => x"fa38d014",
          3536 => x"53805588",
          3537 => x"57897327",
          3538 => x"983880eb",
          3539 => x"39d01453",
          3540 => x"80557289",
          3541 => x"2680e038",
          3542 => x"86398055",
          3543 => x"80d9398a",
          3544 => x"578055a0",
          3545 => x"742780c2",
          3546 => x"3880e074",
          3547 => x"278938e0",
          3548 => x"147081ff",
          3549 => x"065553d0",
          3550 => x"147081ff",
          3551 => x"06555390",
          3552 => x"74278e38",
          3553 => x"f9147081",
          3554 => x"ff065553",
          3555 => x"897427ca",
          3556 => x"38737727",
          3557 => x"c5387477",
          3558 => x"29147608",
          3559 => x"8105770c",
          3560 => x"76087033",
          3561 => x"565455ff",
          3562 => x"ba397780",
          3563 => x"2e843874",
          3564 => x"30557479",
          3565 => x"0c815574",
          3566 => x"81cbd40c",
          3567 => x"8a3d0d04",
          3568 => x"ff3d0d02",
          3569 => x"8f053351",
          3570 => x"81527072",
          3571 => x"26873881",
          3572 => x"c9801133",
          3573 => x"527181cb",
          3574 => x"d40c833d",
          3575 => x"0d04fc3d",
          3576 => x"0d029b05",
          3577 => x"33028405",
          3578 => x"9f053356",
          3579 => x"53835172",
          3580 => x"812680e0",
          3581 => x"3872842b",
          3582 => x"87c0928c",
          3583 => x"11535188",
          3584 => x"5474802e",
          3585 => x"84388188",
          3586 => x"5473720c",
          3587 => x"87c0928c",
          3588 => x"11518171",
          3589 => x"0c850b87",
          3590 => x"c0988c0c",
          3591 => x"70527108",
          3592 => x"70820651",
          3593 => x"5170802e",
          3594 => x"8a3887c0",
          3595 => x"988c0851",
          3596 => x"70ec3871",
          3597 => x"08fc8080",
          3598 => x"06527192",
          3599 => x"3887c098",
          3600 => x"8c085170",
          3601 => x"802e8738",
          3602 => x"7181c980",
          3603 => x"143481c9",
          3604 => x"80133351",
          3605 => x"7081cbd4",
          3606 => x"0c863d0d",
          3607 => x"04f33d0d",
          3608 => x"60626402",
          3609 => x"8c05bf05",
          3610 => x"33574058",
          3611 => x"5b837452",
          3612 => x"5afecd3f",
          3613 => x"81cbd408",
          3614 => x"81067a54",
          3615 => x"527181be",
          3616 => x"38717275",
          3617 => x"842b87c0",
          3618 => x"92801187",
          3619 => x"c0928c12",
          3620 => x"87c09284",
          3621 => x"13415a40",
          3622 => x"575a5885",
          3623 => x"0b87c098",
          3624 => x"8c0c767d",
          3625 => x"0c84760c",
          3626 => x"75087085",
          3627 => x"2a708106",
          3628 => x"51535471",
          3629 => x"802e8e38",
          3630 => x"7b085271",
          3631 => x"7b708105",
          3632 => x"5d348119",
          3633 => x"598074a2",
          3634 => x"06535371",
          3635 => x"732e8338",
          3636 => x"81537883",
          3637 => x"ff268f38",
          3638 => x"72802e8a",
          3639 => x"3887c098",
          3640 => x"8c085271",
          3641 => x"c33887c0",
          3642 => x"988c0852",
          3643 => x"71802e87",
          3644 => x"38788480",
          3645 => x"2e993881",
          3646 => x"760c87c0",
          3647 => x"928c1553",
          3648 => x"72087082",
          3649 => x"06515271",
          3650 => x"f738ff1a",
          3651 => x"5a8d3984",
          3652 => x"80178119",
          3653 => x"7081ff06",
          3654 => x"5a535779",
          3655 => x"802e9038",
          3656 => x"73fc8080",
          3657 => x"06527187",
          3658 => x"387d7826",
          3659 => x"feed3873",
          3660 => x"fc808006",
          3661 => x"5271802e",
          3662 => x"83388152",
          3663 => x"71537281",
          3664 => x"cbd40c8f",
          3665 => x"3d0d04f3",
          3666 => x"3d0d6062",
          3667 => x"64028c05",
          3668 => x"bf053357",
          3669 => x"40585b83",
          3670 => x"59807452",
          3671 => x"58fce13f",
          3672 => x"81cbd408",
          3673 => x"81067954",
          3674 => x"5271782e",
          3675 => x"09810681",
          3676 => x"b1387774",
          3677 => x"842b87c0",
          3678 => x"92801187",
          3679 => x"c0928c12",
          3680 => x"87c09284",
          3681 => x"1340595f",
          3682 => x"565a850b",
          3683 => x"87c0988c",
          3684 => x"0c767d0c",
          3685 => x"82760c80",
          3686 => x"58750870",
          3687 => x"842a7081",
          3688 => x"06515354",
          3689 => x"71802e8c",
          3690 => x"387a7081",
          3691 => x"055c337c",
          3692 => x"0c811858",
          3693 => x"73812a70",
          3694 => x"81065152",
          3695 => x"71802e8a",
          3696 => x"3887c098",
          3697 => x"8c085271",
          3698 => x"d03887c0",
          3699 => x"988c0852",
          3700 => x"71802e87",
          3701 => x"38778480",
          3702 => x"2e993881",
          3703 => x"760c87c0",
          3704 => x"928c1553",
          3705 => x"72087082",
          3706 => x"06515271",
          3707 => x"f738ff19",
          3708 => x"598d3981",
          3709 => x"1a7081ff",
          3710 => x"06848019",
          3711 => x"595b5278",
          3712 => x"802e9038",
          3713 => x"73fc8080",
          3714 => x"06527187",
          3715 => x"387d7a26",
          3716 => x"fef83873",
          3717 => x"fc808006",
          3718 => x"5271802e",
          3719 => x"83388152",
          3720 => x"71537281",
          3721 => x"cbd40c8f",
          3722 => x"3d0d04f6",
          3723 => x"3d0d7e02",
          3724 => x"8405b305",
          3725 => x"33028805",
          3726 => x"b7053371",
          3727 => x"54545657",
          3728 => x"fafe3f81",
          3729 => x"cbd40881",
          3730 => x"06538354",
          3731 => x"7280fe38",
          3732 => x"850b87c0",
          3733 => x"988c0c81",
          3734 => x"5671762e",
          3735 => x"80dc3871",
          3736 => x"76249338",
          3737 => x"74842b87",
          3738 => x"c0928c11",
          3739 => x"54547180",
          3740 => x"2e8d3880",
          3741 => x"d4397183",
          3742 => x"2e80c638",
          3743 => x"80cb3972",
          3744 => x"0870812a",
          3745 => x"70810651",
          3746 => x"51527180",
          3747 => x"2e8a3887",
          3748 => x"c0988c08",
          3749 => x"5271e838",
          3750 => x"87c0988c",
          3751 => x"08527196",
          3752 => x"3881730c",
          3753 => x"87c0928c",
          3754 => x"14537208",
          3755 => x"70820651",
          3756 => x"5271f738",
          3757 => x"96398056",
          3758 => x"92398880",
          3759 => x"0a770c85",
          3760 => x"39818077",
          3761 => x"0c725683",
          3762 => x"39845675",
          3763 => x"547381cb",
          3764 => x"d40c8c3d",
          3765 => x"0d04fe3d",
          3766 => x"0d748111",
          3767 => x"33713371",
          3768 => x"882b0781",
          3769 => x"cbd40c53",
          3770 => x"51843d0d",
          3771 => x"04fd3d0d",
          3772 => x"75831133",
          3773 => x"82123371",
          3774 => x"902b7188",
          3775 => x"2b078114",
          3776 => x"33707207",
          3777 => x"882b7533",
          3778 => x"710781cb",
          3779 => x"d40c5253",
          3780 => x"54565452",
          3781 => x"853d0d04",
          3782 => x"ff3d0d73",
          3783 => x"02840592",
          3784 => x"05225252",
          3785 => x"70727081",
          3786 => x"05543470",
          3787 => x"882a5170",
          3788 => x"7234833d",
          3789 => x"0d04ff3d",
          3790 => x"0d737552",
          3791 => x"52707270",
          3792 => x"81055434",
          3793 => x"70882a51",
          3794 => x"70727081",
          3795 => x"05543470",
          3796 => x"882a5170",
          3797 => x"72708105",
          3798 => x"54347088",
          3799 => x"2a517072",
          3800 => x"34833d0d",
          3801 => x"04fe3d0d",
          3802 => x"76757754",
          3803 => x"54517080",
          3804 => x"2e923871",
          3805 => x"70810553",
          3806 => x"33737081",
          3807 => x"055534ff",
          3808 => x"1151eb39",
          3809 => x"843d0d04",
          3810 => x"fe3d0d75",
          3811 => x"77765452",
          3812 => x"53727270",
          3813 => x"81055434",
          3814 => x"ff115170",
          3815 => x"f438843d",
          3816 => x"0d04fc3d",
          3817 => x"0d787779",
          3818 => x"56565374",
          3819 => x"70810556",
          3820 => x"33747081",
          3821 => x"05563371",
          3822 => x"7131ff16",
          3823 => x"56525252",
          3824 => x"72802e86",
          3825 => x"3871802e",
          3826 => x"e2387181",
          3827 => x"cbd40c86",
          3828 => x"3d0d04fe",
          3829 => x"3d0d7476",
          3830 => x"54518939",
          3831 => x"71732e8a",
          3832 => x"38811151",
          3833 => x"70335271",
          3834 => x"f3387033",
          3835 => x"81cbd40c",
          3836 => x"843d0d04",
          3837 => x"800b81cb",
          3838 => x"d40c0480",
          3839 => x"0b81cbd4",
          3840 => x"0c04f73d",
          3841 => x"0d7b5680",
          3842 => x"0b831733",
          3843 => x"565a747a",
          3844 => x"2e80d638",
          3845 => x"8154b016",
          3846 => x"0853b416",
          3847 => x"70538117",
          3848 => x"335259fa",
          3849 => x"a23f81cb",
          3850 => x"d4087a2e",
          3851 => x"098106b7",
          3852 => x"3881cbd4",
          3853 => x"08831734",
          3854 => x"b0160870",
          3855 => x"a4180831",
          3856 => x"9c180859",
          3857 => x"56587477",
          3858 => x"279f3882",
          3859 => x"16335574",
          3860 => x"822e0981",
          3861 => x"06933881",
          3862 => x"54761853",
          3863 => x"78528116",
          3864 => x"3351f9e3",
          3865 => x"3f833981",
          3866 => x"5a7981cb",
          3867 => x"d40c8b3d",
          3868 => x"0d04fa3d",
          3869 => x"0d787a56",
          3870 => x"56805774",
          3871 => x"b017082e",
          3872 => x"af387551",
          3873 => x"fefc3f81",
          3874 => x"cbd40857",
          3875 => x"81cbd408",
          3876 => x"9f388154",
          3877 => x"7453b416",
          3878 => x"52811633",
          3879 => x"51f7be3f",
          3880 => x"81cbd408",
          3881 => x"802e8538",
          3882 => x"ff558157",
          3883 => x"74b0170c",
          3884 => x"7681cbd4",
          3885 => x"0c883d0d",
          3886 => x"04f83d0d",
          3887 => x"7a705257",
          3888 => x"fec03f81",
          3889 => x"cbd40858",
          3890 => x"81cbd408",
          3891 => x"81913876",
          3892 => x"33557483",
          3893 => x"2e098106",
          3894 => x"80f03884",
          3895 => x"17335978",
          3896 => x"812e0981",
          3897 => x"0680e338",
          3898 => x"84805381",
          3899 => x"cbd40852",
          3900 => x"b4177052",
          3901 => x"56fd913f",
          3902 => x"82d4d552",
          3903 => x"84b21751",
          3904 => x"fc963f84",
          3905 => x"8b85a4d2",
          3906 => x"527551fc",
          3907 => x"a93f868a",
          3908 => x"85e4f252",
          3909 => x"84981751",
          3910 => x"fc9c3f90",
          3911 => x"17085284",
          3912 => x"9c1751fc",
          3913 => x"913f8c17",
          3914 => x"085284a0",
          3915 => x"1751fc86",
          3916 => x"3fa01708",
          3917 => x"810570b0",
          3918 => x"190c7955",
          3919 => x"53755281",
          3920 => x"173351f8",
          3921 => x"823f7784",
          3922 => x"18348053",
          3923 => x"80528117",
          3924 => x"3351f9d7",
          3925 => x"3f81cbd4",
          3926 => x"08802e83",
          3927 => x"38815877",
          3928 => x"81cbd40c",
          3929 => x"8a3d0d04",
          3930 => x"fb3d0d77",
          3931 => x"fe1a9812",
          3932 => x"08fe0555",
          3933 => x"56548056",
          3934 => x"7473278d",
          3935 => x"388a1422",
          3936 => x"757129ac",
          3937 => x"16080557",
          3938 => x"537581cb",
          3939 => x"d40c873d",
          3940 => x"0d04f93d",
          3941 => x"0d7a7a70",
          3942 => x"08565457",
          3943 => x"81772781",
          3944 => x"df387698",
          3945 => x"15082781",
          3946 => x"d738ff74",
          3947 => x"33545872",
          3948 => x"822e80f5",
          3949 => x"38728224",
          3950 => x"89387281",
          3951 => x"2e8d3881",
          3952 => x"bf397283",
          3953 => x"2e818e38",
          3954 => x"81b63976",
          3955 => x"812a1770",
          3956 => x"892aa416",
          3957 => x"08055374",
          3958 => x"5255fd96",
          3959 => x"3f81cbd4",
          3960 => x"08819f38",
          3961 => x"7483ff06",
          3962 => x"14b41133",
          3963 => x"81177089",
          3964 => x"2aa41808",
          3965 => x"05557654",
          3966 => x"575753fc",
          3967 => x"f53f81cb",
          3968 => x"d40880fe",
          3969 => x"387483ff",
          3970 => x"0614b411",
          3971 => x"3370882b",
          3972 => x"78077981",
          3973 => x"0671842a",
          3974 => x"5c525851",
          3975 => x"537280e2",
          3976 => x"38759fff",
          3977 => x"065880da",
          3978 => x"3976882a",
          3979 => x"a4150805",
          3980 => x"527351fc",
          3981 => x"bd3f81cb",
          3982 => x"d40880c6",
          3983 => x"38761083",
          3984 => x"fe067405",
          3985 => x"b40551f9",
          3986 => x"8d3f81cb",
          3987 => x"d40883ff",
          3988 => x"ff0658ae",
          3989 => x"3976872a",
          3990 => x"a4150805",
          3991 => x"527351fc",
          3992 => x"913f81cb",
          3993 => x"d4089b38",
          3994 => x"76822b83",
          3995 => x"fc067405",
          3996 => x"b40551f8",
          3997 => x"f83f81cb",
          3998 => x"d408f00a",
          3999 => x"06588339",
          4000 => x"81587781",
          4001 => x"cbd40c89",
          4002 => x"3d0d04f8",
          4003 => x"3d0d7a7c",
          4004 => x"7e5a5856",
          4005 => x"82598177",
          4006 => x"27829e38",
          4007 => x"76981708",
          4008 => x"27829638",
          4009 => x"75335372",
          4010 => x"792e819d",
          4011 => x"38727924",
          4012 => x"89387281",
          4013 => x"2e8d3882",
          4014 => x"80397283",
          4015 => x"2e81b838",
          4016 => x"81f73976",
          4017 => x"812a1770",
          4018 => x"892aa418",
          4019 => x"08055376",
          4020 => x"5255fb9e",
          4021 => x"3f81cbd4",
          4022 => x"085981cb",
          4023 => x"d40881d9",
          4024 => x"387483ff",
          4025 => x"0616b405",
          4026 => x"81167881",
          4027 => x"06595654",
          4028 => x"77537680",
          4029 => x"2e8f3877",
          4030 => x"842b9ff0",
          4031 => x"0674338f",
          4032 => x"06710751",
          4033 => x"53727434",
          4034 => x"810b8317",
          4035 => x"3474892a",
          4036 => x"a4170805",
          4037 => x"527551fa",
          4038 => x"d93f81cb",
          4039 => x"d4085981",
          4040 => x"cbd40881",
          4041 => x"94387483",
          4042 => x"ff0616b4",
          4043 => x"0578842a",
          4044 => x"5454768f",
          4045 => x"3877882a",
          4046 => x"743381f0",
          4047 => x"06718f06",
          4048 => x"07515372",
          4049 => x"743480ec",
          4050 => x"3976882a",
          4051 => x"a4170805",
          4052 => x"527551fa",
          4053 => x"9d3f81cb",
          4054 => x"d4085981",
          4055 => x"cbd40880",
          4056 => x"d8387783",
          4057 => x"ffff0652",
          4058 => x"761083fe",
          4059 => x"067605b4",
          4060 => x"0551f7a4",
          4061 => x"3fbe3976",
          4062 => x"872aa417",
          4063 => x"08055275",
          4064 => x"51f9ef3f",
          4065 => x"81cbd408",
          4066 => x"5981cbd4",
          4067 => x"08ab3877",
          4068 => x"f00a0677",
          4069 => x"822b83fc",
          4070 => x"067018b4",
          4071 => x"05705451",
          4072 => x"5454f6c9",
          4073 => x"3f81cbd4",
          4074 => x"088f0a06",
          4075 => x"74075272",
          4076 => x"51f7833f",
          4077 => x"810b8317",
          4078 => x"347881cb",
          4079 => x"d40c8a3d",
          4080 => x"0d04f83d",
          4081 => x"0d7a7c7e",
          4082 => x"72085956",
          4083 => x"56598175",
          4084 => x"27a43874",
          4085 => x"98170827",
          4086 => x"9d387380",
          4087 => x"2eaa38ff",
          4088 => x"53735275",
          4089 => x"51fda43f",
          4090 => x"81cbd408",
          4091 => x"5481cbd4",
          4092 => x"0880f238",
          4093 => x"93398254",
          4094 => x"80eb3981",
          4095 => x"5480e639",
          4096 => x"81cbd408",
          4097 => x"5480de39",
          4098 => x"74527851",
          4099 => x"fb843f81",
          4100 => x"cbd40858",
          4101 => x"81cbd408",
          4102 => x"802e80c7",
          4103 => x"3881cbd4",
          4104 => x"08812ed2",
          4105 => x"3881cbd4",
          4106 => x"08ff2ecf",
          4107 => x"38805374",
          4108 => x"527551fc",
          4109 => x"d63f81cb",
          4110 => x"d408c538",
          4111 => x"981608fe",
          4112 => x"11901808",
          4113 => x"57555774",
          4114 => x"74279038",
          4115 => x"81159017",
          4116 => x"0c841633",
          4117 => x"81075473",
          4118 => x"84173477",
          4119 => x"55767826",
          4120 => x"ffa63880",
          4121 => x"547381cb",
          4122 => x"d40c8a3d",
          4123 => x"0d04f63d",
          4124 => x"0d7c7e71",
          4125 => x"08595b5b",
          4126 => x"7995388c",
          4127 => x"17085877",
          4128 => x"802e8838",
          4129 => x"98170878",
          4130 => x"26b23881",
          4131 => x"58ae3979",
          4132 => x"527a51f9",
          4133 => x"fd3f8155",
          4134 => x"7481cbd4",
          4135 => x"082782e0",
          4136 => x"3881cbd4",
          4137 => x"085581cb",
          4138 => x"d408ff2e",
          4139 => x"82d23898",
          4140 => x"170881cb",
          4141 => x"d4082682",
          4142 => x"c7387958",
          4143 => x"90170870",
          4144 => x"56547380",
          4145 => x"2e82b938",
          4146 => x"777a2e09",
          4147 => x"810680e2",
          4148 => x"38811a56",
          4149 => x"98170876",
          4150 => x"26833882",
          4151 => x"5675527a",
          4152 => x"51f9af3f",
          4153 => x"805981cb",
          4154 => x"d408812e",
          4155 => x"09810686",
          4156 => x"3881cbd4",
          4157 => x"085981cb",
          4158 => x"d4080970",
          4159 => x"30707207",
          4160 => x"8025707c",
          4161 => x"0781cbd4",
          4162 => x"08545151",
          4163 => x"55557381",
          4164 => x"ef3881cb",
          4165 => x"d408802e",
          4166 => x"95388c17",
          4167 => x"08548174",
          4168 => x"27903873",
          4169 => x"98180827",
          4170 => x"89387358",
          4171 => x"85397580",
          4172 => x"db387756",
          4173 => x"81165698",
          4174 => x"17087626",
          4175 => x"89388256",
          4176 => x"75782681",
          4177 => x"ac387552",
          4178 => x"7a51f8c6",
          4179 => x"3f81cbd4",
          4180 => x"08802eb8",
          4181 => x"38805981",
          4182 => x"cbd40881",
          4183 => x"2e098106",
          4184 => x"863881cb",
          4185 => x"d4085981",
          4186 => x"cbd40809",
          4187 => x"70307072",
          4188 => x"07802570",
          4189 => x"7c075151",
          4190 => x"55557380",
          4191 => x"f8387578",
          4192 => x"2e098106",
          4193 => x"ffae3873",
          4194 => x"5580f539",
          4195 => x"ff537552",
          4196 => x"7651f9f7",
          4197 => x"3f81cbd4",
          4198 => x"0881cbd4",
          4199 => x"08307081",
          4200 => x"cbd40807",
          4201 => x"80255155",
          4202 => x"5579802e",
          4203 => x"94387380",
          4204 => x"2e8f3875",
          4205 => x"53795276",
          4206 => x"51f9d03f",
          4207 => x"81cbd408",
          4208 => x"5574a538",
          4209 => x"758c180c",
          4210 => x"981708fe",
          4211 => x"05901808",
          4212 => x"56547474",
          4213 => x"268638ff",
          4214 => x"1590180c",
          4215 => x"84173381",
          4216 => x"07547384",
          4217 => x"18349739",
          4218 => x"ff567481",
          4219 => x"2e90388c",
          4220 => x"3980558c",
          4221 => x"3981cbd4",
          4222 => x"08558539",
          4223 => x"81567555",
          4224 => x"7481cbd4",
          4225 => x"0c8c3d0d",
          4226 => x"04f83d0d",
          4227 => x"7a705255",
          4228 => x"f3f03f81",
          4229 => x"cbd40858",
          4230 => x"815681cb",
          4231 => x"d40880d8",
          4232 => x"387b5274",
          4233 => x"51f6c13f",
          4234 => x"81cbd408",
          4235 => x"81cbd408",
          4236 => x"b0170c59",
          4237 => x"84805377",
          4238 => x"52b41570",
          4239 => x"5257f2c8",
          4240 => x"3f775684",
          4241 => x"39811656",
          4242 => x"8a152258",
          4243 => x"75782797",
          4244 => x"38815475",
          4245 => x"19537652",
          4246 => x"81153351",
          4247 => x"ede93f81",
          4248 => x"cbd40880",
          4249 => x"2edf388a",
          4250 => x"15227632",
          4251 => x"70307072",
          4252 => x"07709f2a",
          4253 => x"53515656",
          4254 => x"7581cbd4",
          4255 => x"0c8a3d0d",
          4256 => x"04f83d0d",
          4257 => x"7a7c7108",
          4258 => x"58565774",
          4259 => x"f0800a26",
          4260 => x"80f13874",
          4261 => x"9f065372",
          4262 => x"80e93874",
          4263 => x"90180c88",
          4264 => x"17085473",
          4265 => x"aa387533",
          4266 => x"53827327",
          4267 => x"8838a816",
          4268 => x"0854739b",
          4269 => x"3874852a",
          4270 => x"53820b88",
          4271 => x"17225a58",
          4272 => x"72792780",
          4273 => x"fe38a816",
          4274 => x"0898180c",
          4275 => x"80cd398a",
          4276 => x"16227089",
          4277 => x"2b545872",
          4278 => x"7526b238",
          4279 => x"73527651",
          4280 => x"f5b03f81",
          4281 => x"cbd40854",
          4282 => x"81cbd408",
          4283 => x"ff2ebd38",
          4284 => x"810b81cb",
          4285 => x"d408278b",
          4286 => x"38981608",
          4287 => x"81cbd408",
          4288 => x"26853882",
          4289 => x"58bd3974",
          4290 => x"733155cb",
          4291 => x"39735275",
          4292 => x"51f4d53f",
          4293 => x"81cbd408",
          4294 => x"98180c73",
          4295 => x"94180c98",
          4296 => x"17085382",
          4297 => x"5872802e",
          4298 => x"9a388539",
          4299 => x"81589439",
          4300 => x"74892a13",
          4301 => x"98180c74",
          4302 => x"83ff0616",
          4303 => x"b4059c18",
          4304 => x"0c805877",
          4305 => x"81cbd40c",
          4306 => x"8a3d0d04",
          4307 => x"f83d0d7a",
          4308 => x"70089012",
          4309 => x"08a00559",
          4310 => x"5754f080",
          4311 => x"0a772786",
          4312 => x"38800b98",
          4313 => x"150c9814",
          4314 => x"08538455",
          4315 => x"72802e81",
          4316 => x"cb387683",
          4317 => x"ff065877",
          4318 => x"81b53881",
          4319 => x"1398150c",
          4320 => x"94140855",
          4321 => x"74923876",
          4322 => x"852a8817",
          4323 => x"22565374",
          4324 => x"7326819b",
          4325 => x"3880c039",
          4326 => x"8a1622ff",
          4327 => x"0577892a",
          4328 => x"06537281",
          4329 => x"8a387452",
          4330 => x"7351f3e6",
          4331 => x"3f81cbd4",
          4332 => x"08538255",
          4333 => x"810b81cb",
          4334 => x"d4082780",
          4335 => x"ff388155",
          4336 => x"81cbd408",
          4337 => x"ff2e80f4",
          4338 => x"38981608",
          4339 => x"81cbd408",
          4340 => x"2680ca38",
          4341 => x"7b8a3877",
          4342 => x"98150c84",
          4343 => x"5580dd39",
          4344 => x"94140852",
          4345 => x"7351f986",
          4346 => x"3f81cbd4",
          4347 => x"08538755",
          4348 => x"81cbd408",
          4349 => x"802e80c4",
          4350 => x"38825581",
          4351 => x"cbd40881",
          4352 => x"2eba3881",
          4353 => x"5581cbd4",
          4354 => x"08ff2eb0",
          4355 => x"3881cbd4",
          4356 => x"08527551",
          4357 => x"fbf33f81",
          4358 => x"cbd408a0",
          4359 => x"38729415",
          4360 => x"0c725275",
          4361 => x"51f2c13f",
          4362 => x"81cbd408",
          4363 => x"98150c76",
          4364 => x"90150c77",
          4365 => x"16b4059c",
          4366 => x"150c8055",
          4367 => x"7481cbd4",
          4368 => x"0c8a3d0d",
          4369 => x"04f73d0d",
          4370 => x"7b7d7108",
          4371 => x"5b5b5780",
          4372 => x"527651fc",
          4373 => x"ac3f81cb",
          4374 => x"d4085481",
          4375 => x"cbd40880",
          4376 => x"ec3881cb",
          4377 => x"d4085698",
          4378 => x"17085278",
          4379 => x"51f0833f",
          4380 => x"81cbd408",
          4381 => x"5481cbd4",
          4382 => x"0880d238",
          4383 => x"81cbd408",
          4384 => x"9c180870",
          4385 => x"33515458",
          4386 => x"7281e52e",
          4387 => x"09810683",
          4388 => x"38815881",
          4389 => x"cbd40855",
          4390 => x"72833881",
          4391 => x"55777507",
          4392 => x"5372802e",
          4393 => x"8e388116",
          4394 => x"56757a2e",
          4395 => x"09810688",
          4396 => x"38a53981",
          4397 => x"cbd40856",
          4398 => x"81527651",
          4399 => x"fd8e3f81",
          4400 => x"cbd40854",
          4401 => x"81cbd408",
          4402 => x"802eff9b",
          4403 => x"3873842e",
          4404 => x"09810683",
          4405 => x"38875473",
          4406 => x"81cbd40c",
          4407 => x"8b3d0d04",
          4408 => x"fd3d0d76",
          4409 => x"9a115254",
          4410 => x"ebec3f81",
          4411 => x"cbd40883",
          4412 => x"ffff0676",
          4413 => x"70335153",
          4414 => x"5371832e",
          4415 => x"09810690",
          4416 => x"38941451",
          4417 => x"ebd03f81",
          4418 => x"cbd40890",
          4419 => x"2b730753",
          4420 => x"7281cbd4",
          4421 => x"0c853d0d",
          4422 => x"04fc3d0d",
          4423 => x"77797083",
          4424 => x"ffff0654",
          4425 => x"9a125355",
          4426 => x"55ebed3f",
          4427 => x"76703351",
          4428 => x"5372832e",
          4429 => x"0981068b",
          4430 => x"3873902a",
          4431 => x"52941551",
          4432 => x"ebd63f86",
          4433 => x"3d0d04f7",
          4434 => x"3d0d7b7d",
          4435 => x"5b558475",
          4436 => x"085a5898",
          4437 => x"1508802e",
          4438 => x"818a3898",
          4439 => x"15085278",
          4440 => x"51ee8f3f",
          4441 => x"81cbd408",
          4442 => x"5881cbd4",
          4443 => x"0880f538",
          4444 => x"9c150870",
          4445 => x"33555373",
          4446 => x"86388458",
          4447 => x"80e6398b",
          4448 => x"133370bf",
          4449 => x"067081ff",
          4450 => x"06585153",
          4451 => x"72861634",
          4452 => x"81cbd408",
          4453 => x"537381e5",
          4454 => x"2e833881",
          4455 => x"5373ae2e",
          4456 => x"a9388170",
          4457 => x"74065457",
          4458 => x"72802e9e",
          4459 => x"38758f2e",
          4460 => x"993881cb",
          4461 => x"d40876df",
          4462 => x"06545472",
          4463 => x"882e0981",
          4464 => x"06833876",
          4465 => x"54737a2e",
          4466 => x"a0388052",
          4467 => x"7451fafc",
          4468 => x"3f81cbd4",
          4469 => x"085881cb",
          4470 => x"d4088938",
          4471 => x"981508fe",
          4472 => x"fa388639",
          4473 => x"800b9816",
          4474 => x"0c7781cb",
          4475 => x"d40c8b3d",
          4476 => x"0d04fb3d",
          4477 => x"0d777008",
          4478 => x"57548152",
          4479 => x"7351fcc5",
          4480 => x"3f81cbd4",
          4481 => x"085581cb",
          4482 => x"d408b438",
          4483 => x"98140852",
          4484 => x"7551ecde",
          4485 => x"3f81cbd4",
          4486 => x"085581cb",
          4487 => x"d408a038",
          4488 => x"a05381cb",
          4489 => x"d408529c",
          4490 => x"140851ea",
          4491 => x"db3f8b53",
          4492 => x"a014529c",
          4493 => x"140851ea",
          4494 => x"ac3f810b",
          4495 => x"83173474",
          4496 => x"81cbd40c",
          4497 => x"873d0d04",
          4498 => x"fd3d0d75",
          4499 => x"70089812",
          4500 => x"08547053",
          4501 => x"5553ec9a",
          4502 => x"3f81cbd4",
          4503 => x"088d389c",
          4504 => x"130853e5",
          4505 => x"7334810b",
          4506 => x"83153485",
          4507 => x"3d0d04fa",
          4508 => x"3d0d787a",
          4509 => x"5757800b",
          4510 => x"89173498",
          4511 => x"1708802e",
          4512 => x"81823880",
          4513 => x"70891855",
          4514 => x"55559c17",
          4515 => x"08147033",
          4516 => x"81165651",
          4517 => x"5271a02e",
          4518 => x"a8387185",
          4519 => x"2e098106",
          4520 => x"843881e5",
          4521 => x"5273892e",
          4522 => x"0981068b",
          4523 => x"38ae7370",
          4524 => x"81055534",
          4525 => x"81155571",
          4526 => x"73708105",
          4527 => x"55348115",
          4528 => x"558a7427",
          4529 => x"c5387515",
          4530 => x"88055280",
          4531 => x"0b811334",
          4532 => x"9c170852",
          4533 => x"8b123388",
          4534 => x"17349c17",
          4535 => x"089c1152",
          4536 => x"52e88a3f",
          4537 => x"81cbd408",
          4538 => x"760c9612",
          4539 => x"51e7e73f",
          4540 => x"81cbd408",
          4541 => x"86172398",
          4542 => x"1251e7da",
          4543 => x"3f81cbd4",
          4544 => x"08841723",
          4545 => x"883d0d04",
          4546 => x"f33d0d7f",
          4547 => x"70085e5b",
          4548 => x"80617033",
          4549 => x"51555573",
          4550 => x"af2e8338",
          4551 => x"81557380",
          4552 => x"dc2e9138",
          4553 => x"74802e8c",
          4554 => x"38941d08",
          4555 => x"881c0caa",
          4556 => x"39811541",
          4557 => x"80617033",
          4558 => x"56565673",
          4559 => x"af2e0981",
          4560 => x"06833881",
          4561 => x"567380dc",
          4562 => x"32703070",
          4563 => x"80257807",
          4564 => x"51515473",
          4565 => x"dc387388",
          4566 => x"1c0c6070",
          4567 => x"33515473",
          4568 => x"9f269638",
          4569 => x"ff800bab",
          4570 => x"1c348052",
          4571 => x"7a51f691",
          4572 => x"3f81cbd4",
          4573 => x"08558598",
          4574 => x"39913d61",
          4575 => x"a01d5c5a",
          4576 => x"5e8b53a0",
          4577 => x"527951e7",
          4578 => x"ff3f8070",
          4579 => x"59578879",
          4580 => x"33555c73",
          4581 => x"ae2e0981",
          4582 => x"0680d438",
          4583 => x"78187033",
          4584 => x"811a71ae",
          4585 => x"32703070",
          4586 => x"9f2a7382",
          4587 => x"26075151",
          4588 => x"535a5754",
          4589 => x"738c3879",
          4590 => x"17547574",
          4591 => x"34811757",
          4592 => x"db3975af",
          4593 => x"32703070",
          4594 => x"9f2a5151",
          4595 => x"547580dc",
          4596 => x"2e8c3873",
          4597 => x"802e8738",
          4598 => x"75a02682",
          4599 => x"bd387719",
          4600 => x"7e0ca454",
          4601 => x"a0762782",
          4602 => x"bd38a054",
          4603 => x"82b83978",
          4604 => x"18703381",
          4605 => x"1a5a5754",
          4606 => x"a0762781",
          4607 => x"fc3875af",
          4608 => x"32703077",
          4609 => x"80dc3270",
          4610 => x"30728025",
          4611 => x"71802507",
          4612 => x"51515651",
          4613 => x"5573802e",
          4614 => x"ac388439",
          4615 => x"81185880",
          4616 => x"781a7033",
          4617 => x"51555573",
          4618 => x"af2e0981",
          4619 => x"06833881",
          4620 => x"557380dc",
          4621 => x"32703070",
          4622 => x"80257707",
          4623 => x"51515473",
          4624 => x"db3881b5",
          4625 => x"3975ae2e",
          4626 => x"09810683",
          4627 => x"38815476",
          4628 => x"7c277407",
          4629 => x"5473802e",
          4630 => x"a2387b8b",
          4631 => x"32703077",
          4632 => x"ae327030",
          4633 => x"72802571",
          4634 => x"9f2a0753",
          4635 => x"51565155",
          4636 => x"7481a738",
          4637 => x"88578b5c",
          4638 => x"fef53975",
          4639 => x"982b5473",
          4640 => x"80258c38",
          4641 => x"7580ff06",
          4642 => x"81bbb011",
          4643 => x"33575475",
          4644 => x"51e6e13f",
          4645 => x"81cbd408",
          4646 => x"802eb238",
          4647 => x"78187033",
          4648 => x"811a7154",
          4649 => x"5a5654e6",
          4650 => x"d23f81cb",
          4651 => x"d408802e",
          4652 => x"80e838ff",
          4653 => x"1c547674",
          4654 => x"2780df38",
          4655 => x"79175475",
          4656 => x"74348117",
          4657 => x"7a115557",
          4658 => x"747434a7",
          4659 => x"39755281",
          4660 => x"bad051e5",
          4661 => x"fe3f81cb",
          4662 => x"d408bf38",
          4663 => x"ff9f1654",
          4664 => x"73992689",
          4665 => x"38e01670",
          4666 => x"81ff0657",
          4667 => x"54791754",
          4668 => x"75743481",
          4669 => x"1757fdf7",
          4670 => x"3977197e",
          4671 => x"0c76802e",
          4672 => x"99387933",
          4673 => x"547381e5",
          4674 => x"2e098106",
          4675 => x"8438857a",
          4676 => x"348454a0",
          4677 => x"76278f38",
          4678 => x"8b398655",
          4679 => x"81f23984",
          4680 => x"5680f339",
          4681 => x"8054738b",
          4682 => x"1b34807b",
          4683 => x"0858527a",
          4684 => x"51f2ce3f",
          4685 => x"81cbd408",
          4686 => x"5681cbd4",
          4687 => x"0880d738",
          4688 => x"981b0852",
          4689 => x"7651e6aa",
          4690 => x"3f81cbd4",
          4691 => x"085681cb",
          4692 => x"d40880c2",
          4693 => x"389c1b08",
          4694 => x"70335555",
          4695 => x"73802eff",
          4696 => x"be388b15",
          4697 => x"33bf0654",
          4698 => x"73861c34",
          4699 => x"8b153370",
          4700 => x"832a7081",
          4701 => x"06515558",
          4702 => x"7392388b",
          4703 => x"53795274",
          4704 => x"51e49f3f",
          4705 => x"81cbd408",
          4706 => x"802e8b38",
          4707 => x"75527a51",
          4708 => x"f3ba3fff",
          4709 => x"9f3975ab",
          4710 => x"1c335755",
          4711 => x"74802ebb",
          4712 => x"3874842e",
          4713 => x"09810680",
          4714 => x"e7387585",
          4715 => x"2a708106",
          4716 => x"77822a58",
          4717 => x"51547380",
          4718 => x"2e963875",
          4719 => x"81065473",
          4720 => x"802efbb5",
          4721 => x"38ff800b",
          4722 => x"ab1c3480",
          4723 => x"5580c139",
          4724 => x"75810654",
          4725 => x"73ba3885",
          4726 => x"55b63975",
          4727 => x"822a7081",
          4728 => x"06515473",
          4729 => x"ab38861b",
          4730 => x"3370842a",
          4731 => x"70810651",
          4732 => x"55557380",
          4733 => x"2ee13890",
          4734 => x"1b0883ff",
          4735 => x"061db405",
          4736 => x"527c51f5",
          4737 => x"db3f81cb",
          4738 => x"d408881c",
          4739 => x"0cfaea39",
          4740 => x"7481cbd4",
          4741 => x"0c8f3d0d",
          4742 => x"04f63d0d",
          4743 => x"7c5bff7b",
          4744 => x"08707173",
          4745 => x"55595c55",
          4746 => x"5973802e",
          4747 => x"81c63875",
          4748 => x"70810557",
          4749 => x"3370a026",
          4750 => x"525271ba",
          4751 => x"2e8d3870",
          4752 => x"ee3871ba",
          4753 => x"2e098106",
          4754 => x"81a53873",
          4755 => x"33d01170",
          4756 => x"81ff0651",
          4757 => x"52537089",
          4758 => x"26913882",
          4759 => x"147381ff",
          4760 => x"06d00556",
          4761 => x"5271762e",
          4762 => x"80f73880",
          4763 => x"0b81bba0",
          4764 => x"59557708",
          4765 => x"7a555776",
          4766 => x"70810558",
          4767 => x"33747081",
          4768 => x"055633ff",
          4769 => x"9f125353",
          4770 => x"53709926",
          4771 => x"8938e013",
          4772 => x"7081ff06",
          4773 => x"5451ff9f",
          4774 => x"12517099",
          4775 => x"268938e0",
          4776 => x"127081ff",
          4777 => x"06535172",
          4778 => x"30709f2a",
          4779 => x"51517272",
          4780 => x"2e098106",
          4781 => x"853870ff",
          4782 => x"be387230",
          4783 => x"74773270",
          4784 => x"30707207",
          4785 => x"9f2a739f",
          4786 => x"2a075354",
          4787 => x"54517080",
          4788 => x"2e8f3881",
          4789 => x"15841959",
          4790 => x"55837525",
          4791 => x"ff94388b",
          4792 => x"39748324",
          4793 => x"86387476",
          4794 => x"7c0c5978",
          4795 => x"51863981",
          4796 => x"cc843351",
          4797 => x"7081cbd4",
          4798 => x"0c8c3d0d",
          4799 => x"04fa3d0d",
          4800 => x"7856800b",
          4801 => x"831734ff",
          4802 => x"0bb0170c",
          4803 => x"79527551",
          4804 => x"e2e03f84",
          4805 => x"5581cbd4",
          4806 => x"08818038",
          4807 => x"84b21651",
          4808 => x"dfb43f81",
          4809 => x"cbd40883",
          4810 => x"ffff0654",
          4811 => x"83557382",
          4812 => x"d4d52e09",
          4813 => x"810680e3",
          4814 => x"38800bb4",
          4815 => x"17335657",
          4816 => x"7481e92e",
          4817 => x"09810683",
          4818 => x"38815774",
          4819 => x"81eb3270",
          4820 => x"30708025",
          4821 => x"79075151",
          4822 => x"54738a38",
          4823 => x"7481e82e",
          4824 => x"098106b5",
          4825 => x"38835381",
          4826 => x"bae05280",
          4827 => x"ea1651e0",
          4828 => x"b13f81cb",
          4829 => x"d4085581",
          4830 => x"cbd40880",
          4831 => x"2e9d3885",
          4832 => x"5381bae4",
          4833 => x"52818616",
          4834 => x"51e0973f",
          4835 => x"81cbd408",
          4836 => x"5581cbd4",
          4837 => x"08802e83",
          4838 => x"38825574",
          4839 => x"81cbd40c",
          4840 => x"883d0d04",
          4841 => x"f23d0d61",
          4842 => x"02840580",
          4843 => x"cb053358",
          4844 => x"5580750c",
          4845 => x"6051fce1",
          4846 => x"3f81cbd4",
          4847 => x"08588b56",
          4848 => x"800b81cb",
          4849 => x"d4082486",
          4850 => x"fc3881cb",
          4851 => x"d4088429",
          4852 => x"81cbf005",
          4853 => x"70085553",
          4854 => x"8c567380",
          4855 => x"2e86e638",
          4856 => x"73750c76",
          4857 => x"81fe0674",
          4858 => x"33545772",
          4859 => x"802eae38",
          4860 => x"81143351",
          4861 => x"d7ca3f81",
          4862 => x"cbd40881",
          4863 => x"ff067081",
          4864 => x"06545572",
          4865 => x"98387680",
          4866 => x"2e86b838",
          4867 => x"74822a70",
          4868 => x"81065153",
          4869 => x"8a567286",
          4870 => x"ac3886a7",
          4871 => x"39807434",
          4872 => x"77811534",
          4873 => x"81528114",
          4874 => x"3351d7b2",
          4875 => x"3f81cbd4",
          4876 => x"0881ff06",
          4877 => x"70810654",
          4878 => x"55835672",
          4879 => x"86873876",
          4880 => x"802e8f38",
          4881 => x"74822a70",
          4882 => x"81065153",
          4883 => x"8a567285",
          4884 => x"f4388070",
          4885 => x"5374525b",
          4886 => x"fda33f81",
          4887 => x"cbd40881",
          4888 => x"ff065776",
          4889 => x"822e0981",
          4890 => x"0680e238",
          4891 => x"8c3d7456",
          4892 => x"58835683",
          4893 => x"f6153370",
          4894 => x"58537280",
          4895 => x"2e8d3883",
          4896 => x"fa1551dc",
          4897 => x"e83f81cb",
          4898 => x"d4085776",
          4899 => x"78708405",
          4900 => x"5a0cff16",
          4901 => x"90165656",
          4902 => x"758025d7",
          4903 => x"38800b8d",
          4904 => x"3d545672",
          4905 => x"70840554",
          4906 => x"085b8357",
          4907 => x"7a802e95",
          4908 => x"387a5273",
          4909 => x"51fcc63f",
          4910 => x"81cbd408",
          4911 => x"81ff0657",
          4912 => x"81772789",
          4913 => x"38811656",
          4914 => x"837627d7",
          4915 => x"38815676",
          4916 => x"842e84f1",
          4917 => x"388d5676",
          4918 => x"812684e9",
          4919 => x"38bf1451",
          4920 => x"dbf43f81",
          4921 => x"cbd40883",
          4922 => x"ffff0653",
          4923 => x"7284802e",
          4924 => x"09810684",
          4925 => x"d03880ca",
          4926 => x"1451dbda",
          4927 => x"3f81cbd4",
          4928 => x"0883ffff",
          4929 => x"0658778d",
          4930 => x"3880d814",
          4931 => x"51dbde3f",
          4932 => x"81cbd408",
          4933 => x"58779c15",
          4934 => x"0c80c414",
          4935 => x"33821534",
          4936 => x"80c41433",
          4937 => x"ff117081",
          4938 => x"ff065154",
          4939 => x"558d5672",
          4940 => x"81268491",
          4941 => x"387481ff",
          4942 => x"06787129",
          4943 => x"80c11633",
          4944 => x"52595372",
          4945 => x"8a152372",
          4946 => x"802e8b38",
          4947 => x"ff137306",
          4948 => x"5372802e",
          4949 => x"86388d56",
          4950 => x"83eb3980",
          4951 => x"c51451da",
          4952 => x"f53f81cb",
          4953 => x"d4085381",
          4954 => x"cbd40888",
          4955 => x"1523728f",
          4956 => x"06578d56",
          4957 => x"7683ce38",
          4958 => x"80c71451",
          4959 => x"dad83f81",
          4960 => x"cbd40883",
          4961 => x"ffff0655",
          4962 => x"748d3880",
          4963 => x"d41451da",
          4964 => x"dc3f81cb",
          4965 => x"d4085580",
          4966 => x"c21451da",
          4967 => x"b93f81cb",
          4968 => x"d40883ff",
          4969 => x"ff06538d",
          4970 => x"5672802e",
          4971 => x"83973888",
          4972 => x"14227814",
          4973 => x"71842a05",
          4974 => x"5a5a7875",
          4975 => x"26838638",
          4976 => x"8a142252",
          4977 => x"74793151",
          4978 => x"ffb3833f",
          4979 => x"81cbd408",
          4980 => x"5581cbd4",
          4981 => x"08802e82",
          4982 => x"ec3881cb",
          4983 => x"d40880ff",
          4984 => x"fffff526",
          4985 => x"83388357",
          4986 => x"7483fff5",
          4987 => x"26833882",
          4988 => x"57749ff5",
          4989 => x"26853881",
          4990 => x"5789398d",
          4991 => x"5676802e",
          4992 => x"82c33882",
          4993 => x"15709816",
          4994 => x"0c7ba016",
          4995 => x"0c731c70",
          4996 => x"a4170c7a",
          4997 => x"1dac170c",
          4998 => x"54557683",
          4999 => x"2e098106",
          5000 => x"af3880de",
          5001 => x"1451d9ae",
          5002 => x"3f81cbd4",
          5003 => x"0883ffff",
          5004 => x"06538d56",
          5005 => x"72828e38",
          5006 => x"79828a38",
          5007 => x"80e01451",
          5008 => x"d9ab3f81",
          5009 => x"cbd408a8",
          5010 => x"150c7482",
          5011 => x"2b53a239",
          5012 => x"8d567980",
          5013 => x"2e81ee38",
          5014 => x"7713a815",
          5015 => x"0c741553",
          5016 => x"76822e8d",
          5017 => x"38741015",
          5018 => x"70812a76",
          5019 => x"81060551",
          5020 => x"5383ff13",
          5021 => x"892a538d",
          5022 => x"56729c15",
          5023 => x"082681c5",
          5024 => x"38ff0b90",
          5025 => x"150cff0b",
          5026 => x"8c150cff",
          5027 => x"800b8415",
          5028 => x"3476832e",
          5029 => x"09810681",
          5030 => x"923880e4",
          5031 => x"1451d8b6",
          5032 => x"3f81cbd4",
          5033 => x"0883ffff",
          5034 => x"06537281",
          5035 => x"2e098106",
          5036 => x"80f93881",
          5037 => x"1b527351",
          5038 => x"dbb83f81",
          5039 => x"cbd40880",
          5040 => x"ea3881cb",
          5041 => x"d4088415",
          5042 => x"3484b214",
          5043 => x"51d8873f",
          5044 => x"81cbd408",
          5045 => x"83ffff06",
          5046 => x"537282d4",
          5047 => x"d52e0981",
          5048 => x"0680c838",
          5049 => x"b41451d8",
          5050 => x"843f81cb",
          5051 => x"d408848b",
          5052 => x"85a4d22e",
          5053 => x"098106b3",
          5054 => x"38849814",
          5055 => x"51d7ee3f",
          5056 => x"81cbd408",
          5057 => x"868a85e4",
          5058 => x"f22e0981",
          5059 => x"069d3884",
          5060 => x"9c1451d7",
          5061 => x"d83f81cb",
          5062 => x"d4089015",
          5063 => x"0c84a014",
          5064 => x"51d7ca3f",
          5065 => x"81cbd408",
          5066 => x"8c150c76",
          5067 => x"743481cc",
          5068 => x"80228105",
          5069 => x"537281cc",
          5070 => x"80237286",
          5071 => x"1523800b",
          5072 => x"94150c80",
          5073 => x"567581cb",
          5074 => x"d40c903d",
          5075 => x"0d04fb3d",
          5076 => x"0d775489",
          5077 => x"5573802e",
          5078 => x"b9387308",
          5079 => x"5372802e",
          5080 => x"b1387233",
          5081 => x"5271802e",
          5082 => x"a9388613",
          5083 => x"22841522",
          5084 => x"57527176",
          5085 => x"2e098106",
          5086 => x"99388113",
          5087 => x"3351d0c0",
          5088 => x"3f81cbd4",
          5089 => x"08810652",
          5090 => x"71883871",
          5091 => x"74085455",
          5092 => x"83398053",
          5093 => x"7873710c",
          5094 => x"527481cb",
          5095 => x"d40c873d",
          5096 => x"0d04fa3d",
          5097 => x"0d02ab05",
          5098 => x"337a5889",
          5099 => x"3dfc0552",
          5100 => x"56f4e63f",
          5101 => x"8b54800b",
          5102 => x"81cbd408",
          5103 => x"24bc3881",
          5104 => x"cbd40884",
          5105 => x"2981cbf0",
          5106 => x"05700855",
          5107 => x"5573802e",
          5108 => x"84388074",
          5109 => x"34785473",
          5110 => x"802e8438",
          5111 => x"80743478",
          5112 => x"750c7554",
          5113 => x"75802e92",
          5114 => x"38805389",
          5115 => x"3d705384",
          5116 => x"0551f7b0",
          5117 => x"3f81cbd4",
          5118 => x"08547381",
          5119 => x"cbd40c88",
          5120 => x"3d0d04eb",
          5121 => x"3d0d6702",
          5122 => x"840580e7",
          5123 => x"05335959",
          5124 => x"89547880",
          5125 => x"2e84c838",
          5126 => x"77bf0670",
          5127 => x"54983dd0",
          5128 => x"0553993d",
          5129 => x"84055258",
          5130 => x"f6fa3f81",
          5131 => x"cbd40855",
          5132 => x"81cbd408",
          5133 => x"84a4387a",
          5134 => x"5c68528c",
          5135 => x"3d705256",
          5136 => x"edc63f81",
          5137 => x"cbd40855",
          5138 => x"81cbd408",
          5139 => x"92380280",
          5140 => x"d7053370",
          5141 => x"982b5557",
          5142 => x"73802583",
          5143 => x"38865577",
          5144 => x"9c065473",
          5145 => x"802e81ab",
          5146 => x"3874802e",
          5147 => x"95387484",
          5148 => x"2e098106",
          5149 => x"aa387551",
          5150 => x"eaf83f81",
          5151 => x"cbd40855",
          5152 => x"9e3902b2",
          5153 => x"05339106",
          5154 => x"547381b8",
          5155 => x"3877822a",
          5156 => x"70810651",
          5157 => x"5473802e",
          5158 => x"8e388855",
          5159 => x"83bc3977",
          5160 => x"88075874",
          5161 => x"83b43877",
          5162 => x"832a7081",
          5163 => x"06515473",
          5164 => x"802e81af",
          5165 => x"3862527a",
          5166 => x"51e8a53f",
          5167 => x"81cbd408",
          5168 => x"568288b2",
          5169 => x"0a52628e",
          5170 => x"0551d4ea",
          5171 => x"3f6254a0",
          5172 => x"0b8b1534",
          5173 => x"80536252",
          5174 => x"7a51e8bd",
          5175 => x"3f805262",
          5176 => x"9c0551d4",
          5177 => x"d13f7a54",
          5178 => x"810b8315",
          5179 => x"3475802e",
          5180 => x"80f1387a",
          5181 => x"b0110851",
          5182 => x"54805375",
          5183 => x"52973dd4",
          5184 => x"0551ddbe",
          5185 => x"3f81cbd4",
          5186 => x"085581cb",
          5187 => x"d40882ca",
          5188 => x"38b73974",
          5189 => x"82c43802",
          5190 => x"b2053370",
          5191 => x"842a7081",
          5192 => x"06515556",
          5193 => x"73802e86",
          5194 => x"38845582",
          5195 => x"ad397781",
          5196 => x"2a708106",
          5197 => x"51547380",
          5198 => x"2ea93875",
          5199 => x"81065473",
          5200 => x"802ea038",
          5201 => x"87558292",
          5202 => x"3973527a",
          5203 => x"51d6a33f",
          5204 => x"81cbd408",
          5205 => x"7bff188c",
          5206 => x"120c5555",
          5207 => x"81cbd408",
          5208 => x"81f83877",
          5209 => x"832a7081",
          5210 => x"06515473",
          5211 => x"802e8638",
          5212 => x"7780c007",
          5213 => x"587ab011",
          5214 => x"08a01b0c",
          5215 => x"63a41b0c",
          5216 => x"63537052",
          5217 => x"57e6d93f",
          5218 => x"81cbd408",
          5219 => x"81cbd408",
          5220 => x"881b0c63",
          5221 => x"9c05525a",
          5222 => x"d2d33f81",
          5223 => x"cbd40881",
          5224 => x"cbd4088c",
          5225 => x"1b0c777a",
          5226 => x"0c568617",
          5227 => x"22841a23",
          5228 => x"77901a34",
          5229 => x"800b911a",
          5230 => x"34800b9c",
          5231 => x"1a0c800b",
          5232 => x"941a0c77",
          5233 => x"852a7081",
          5234 => x"06515473",
          5235 => x"802e818d",
          5236 => x"3881cbd4",
          5237 => x"08802e81",
          5238 => x"843881cb",
          5239 => x"d408941a",
          5240 => x"0c8a1722",
          5241 => x"70892b7b",
          5242 => x"525957a8",
          5243 => x"39765278",
          5244 => x"51d79f3f",
          5245 => x"81cbd408",
          5246 => x"5781cbd4",
          5247 => x"08812683",
          5248 => x"38825581",
          5249 => x"cbd408ff",
          5250 => x"2e098106",
          5251 => x"83387955",
          5252 => x"75783156",
          5253 => x"74307076",
          5254 => x"07802551",
          5255 => x"54777627",
          5256 => x"8a388170",
          5257 => x"7506555a",
          5258 => x"73c33876",
          5259 => x"981a0c74",
          5260 => x"a9387583",
          5261 => x"ff065473",
          5262 => x"802ea238",
          5263 => x"76527a51",
          5264 => x"d6a63f81",
          5265 => x"cbd40885",
          5266 => x"3882558e",
          5267 => x"3975892a",
          5268 => x"81cbd408",
          5269 => x"059c1a0c",
          5270 => x"84398079",
          5271 => x"0c745473",
          5272 => x"81cbd40c",
          5273 => x"973d0d04",
          5274 => x"f23d0d60",
          5275 => x"63656440",
          5276 => x"405d5980",
          5277 => x"7e0c903d",
          5278 => x"fc055278",
          5279 => x"51f9cf3f",
          5280 => x"81cbd408",
          5281 => x"5581cbd4",
          5282 => x"088a3891",
          5283 => x"19335574",
          5284 => x"802e8638",
          5285 => x"745682c4",
          5286 => x"39901933",
          5287 => x"81065587",
          5288 => x"5674802e",
          5289 => x"82b63895",
          5290 => x"39820b91",
          5291 => x"1a348256",
          5292 => x"82aa3981",
          5293 => x"0b911a34",
          5294 => x"815682a0",
          5295 => x"398c1908",
          5296 => x"941a0831",
          5297 => x"55747c27",
          5298 => x"8338745c",
          5299 => x"7b802e82",
          5300 => x"89389419",
          5301 => x"087083ff",
          5302 => x"06565674",
          5303 => x"81b2387e",
          5304 => x"8a1122ff",
          5305 => x"0577892a",
          5306 => x"065b5579",
          5307 => x"a8387587",
          5308 => x"38881908",
          5309 => x"558f3998",
          5310 => x"19085278",
          5311 => x"51d5933f",
          5312 => x"81cbd408",
          5313 => x"55817527",
          5314 => x"ff9f3874",
          5315 => x"ff2effa3",
          5316 => x"3874981a",
          5317 => x"0c981908",
          5318 => x"527e51d4",
          5319 => x"cb3f81cb",
          5320 => x"d408802e",
          5321 => x"ff833881",
          5322 => x"cbd4081a",
          5323 => x"7c892a59",
          5324 => x"5777802e",
          5325 => x"80d63877",
          5326 => x"1a7f8a11",
          5327 => x"22585c55",
          5328 => x"75752785",
          5329 => x"38757a31",
          5330 => x"58775476",
          5331 => x"537c5281",
          5332 => x"1b3351ca",
          5333 => x"883f81cb",
          5334 => x"d408fed7",
          5335 => x"387e8311",
          5336 => x"33565674",
          5337 => x"802e9f38",
          5338 => x"b0160877",
          5339 => x"31557478",
          5340 => x"27943884",
          5341 => x"8053b416",
          5342 => x"52b01608",
          5343 => x"7731892b",
          5344 => x"7d0551cf",
          5345 => x"e03f7789",
          5346 => x"2b56b939",
          5347 => x"769c1a0c",
          5348 => x"94190883",
          5349 => x"ff068480",
          5350 => x"71315755",
          5351 => x"7b762783",
          5352 => x"387b569c",
          5353 => x"1908527e",
          5354 => x"51d1c73f",
          5355 => x"81cbd408",
          5356 => x"fe813875",
          5357 => x"53941908",
          5358 => x"83ff061f",
          5359 => x"b405527c",
          5360 => x"51cfa23f",
          5361 => x"7b76317e",
          5362 => x"08177f0c",
          5363 => x"761e941b",
          5364 => x"0818941c",
          5365 => x"0c5e5cfd",
          5366 => x"f3398056",
          5367 => x"7581cbd4",
          5368 => x"0c903d0d",
          5369 => x"04f23d0d",
          5370 => x"60636564",
          5371 => x"40405d58",
          5372 => x"807e0c90",
          5373 => x"3dfc0552",
          5374 => x"7751f6d2",
          5375 => x"3f81cbd4",
          5376 => x"085581cb",
          5377 => x"d4088a38",
          5378 => x"91183355",
          5379 => x"74802e86",
          5380 => x"38745683",
          5381 => x"b8399018",
          5382 => x"3370812a",
          5383 => x"70810651",
          5384 => x"56568756",
          5385 => x"74802e83",
          5386 => x"a4389539",
          5387 => x"820b9119",
          5388 => x"34825683",
          5389 => x"9839810b",
          5390 => x"91193481",
          5391 => x"56838e39",
          5392 => x"9418087c",
          5393 => x"11565674",
          5394 => x"76278438",
          5395 => x"75095c7b",
          5396 => x"802e82ec",
          5397 => x"38941808",
          5398 => x"7083ff06",
          5399 => x"56567481",
          5400 => x"fd387e8a",
          5401 => x"1122ff05",
          5402 => x"77892a06",
          5403 => x"5c557abf",
          5404 => x"38758c38",
          5405 => x"88180855",
          5406 => x"749c387a",
          5407 => x"52853998",
          5408 => x"18085277",
          5409 => x"51d7e73f",
          5410 => x"81cbd408",
          5411 => x"5581cbd4",
          5412 => x"08802e82",
          5413 => x"ab387481",
          5414 => x"2eff9138",
          5415 => x"74ff2eff",
          5416 => x"95387498",
          5417 => x"190c8818",
          5418 => x"08853874",
          5419 => x"88190c7e",
          5420 => x"55b01508",
          5421 => x"9c19082e",
          5422 => x"0981068d",
          5423 => x"387451ce",
          5424 => x"c13f81cb",
          5425 => x"d408feee",
          5426 => x"38981808",
          5427 => x"527e51d1",
          5428 => x"973f81cb",
          5429 => x"d408802e",
          5430 => x"fed23881",
          5431 => x"cbd4081b",
          5432 => x"7c892a5a",
          5433 => x"5778802e",
          5434 => x"80d53878",
          5435 => x"1b7f8a11",
          5436 => x"22585b55",
          5437 => x"75752785",
          5438 => x"38757b31",
          5439 => x"59785476",
          5440 => x"537c5281",
          5441 => x"1a3351c8",
          5442 => x"be3f81cb",
          5443 => x"d408fea6",
          5444 => x"387eb011",
          5445 => x"08783156",
          5446 => x"56747927",
          5447 => x"9b388480",
          5448 => x"53b01608",
          5449 => x"7731892b",
          5450 => x"7d0552b4",
          5451 => x"1651ccb5",
          5452 => x"3f7e5580",
          5453 => x"0b831634",
          5454 => x"78892b56",
          5455 => x"80db398c",
          5456 => x"18089419",
          5457 => x"08269338",
          5458 => x"7e51cdb6",
          5459 => x"3f81cbd4",
          5460 => x"08fde338",
          5461 => x"7e77b012",
          5462 => x"0c55769c",
          5463 => x"190c9418",
          5464 => x"0883ff06",
          5465 => x"84807131",
          5466 => x"57557b76",
          5467 => x"2783387b",
          5468 => x"569c1808",
          5469 => x"527e51cd",
          5470 => x"f93f81cb",
          5471 => x"d408fdb6",
          5472 => x"3875537c",
          5473 => x"52941808",
          5474 => x"83ff061f",
          5475 => x"b40551cb",
          5476 => x"d43f7e55",
          5477 => x"810b8316",
          5478 => x"347b7631",
          5479 => x"7e08177f",
          5480 => x"0c761e94",
          5481 => x"1a081870",
          5482 => x"941c0c8c",
          5483 => x"1b085858",
          5484 => x"5e5c7476",
          5485 => x"27833875",
          5486 => x"55748c19",
          5487 => x"0cfd9039",
          5488 => x"90183380",
          5489 => x"c0075574",
          5490 => x"90193480",
          5491 => x"567581cb",
          5492 => x"d40c903d",
          5493 => x"0d04f83d",
          5494 => x"0d7a8b3d",
          5495 => x"fc055370",
          5496 => x"5256f2ea",
          5497 => x"3f81cbd4",
          5498 => x"085781cb",
          5499 => x"d40880fb",
          5500 => x"38901633",
          5501 => x"70862a70",
          5502 => x"81065155",
          5503 => x"5573802e",
          5504 => x"80e938a0",
          5505 => x"16085278",
          5506 => x"51cce73f",
          5507 => x"81cbd408",
          5508 => x"5781cbd4",
          5509 => x"0880d438",
          5510 => x"a416088b",
          5511 => x"1133a007",
          5512 => x"5555738b",
          5513 => x"16348816",
          5514 => x"08537452",
          5515 => x"750851dd",
          5516 => x"e83f8c16",
          5517 => x"08529c15",
          5518 => x"51c9fb3f",
          5519 => x"8288b20a",
          5520 => x"52961551",
          5521 => x"c9f03f76",
          5522 => x"52921551",
          5523 => x"c9ca3f78",
          5524 => x"54810b83",
          5525 => x"15347851",
          5526 => x"ccdf3f81",
          5527 => x"cbd40890",
          5528 => x"173381bf",
          5529 => x"06555773",
          5530 => x"90173476",
          5531 => x"81cbd40c",
          5532 => x"8a3d0d04",
          5533 => x"fc3d0d76",
          5534 => x"705254fe",
          5535 => x"d93f81cb",
          5536 => x"d4085381",
          5537 => x"cbd4089c",
          5538 => x"38863dfc",
          5539 => x"05527351",
          5540 => x"f1bc3f81",
          5541 => x"cbd40853",
          5542 => x"81cbd408",
          5543 => x"873881cb",
          5544 => x"d408740c",
          5545 => x"7281cbd4",
          5546 => x"0c863d0d",
          5547 => x"04ff3d0d",
          5548 => x"843d51e6",
          5549 => x"e43f8b52",
          5550 => x"800b81cb",
          5551 => x"d408248b",
          5552 => x"3881cbd4",
          5553 => x"0881cc84",
          5554 => x"34805271",
          5555 => x"81cbd40c",
          5556 => x"833d0d04",
          5557 => x"ef3d0d80",
          5558 => x"53933dd0",
          5559 => x"0552943d",
          5560 => x"51e9c13f",
          5561 => x"81cbd408",
          5562 => x"5581cbd4",
          5563 => x"0880e038",
          5564 => x"76586352",
          5565 => x"933dd405",
          5566 => x"51e08d3f",
          5567 => x"81cbd408",
          5568 => x"5581cbd4",
          5569 => x"08bc3802",
          5570 => x"80c70533",
          5571 => x"70982b55",
          5572 => x"56738025",
          5573 => x"8938767a",
          5574 => x"94120c54",
          5575 => x"b23902a2",
          5576 => x"05337084",
          5577 => x"2a708106",
          5578 => x"51555673",
          5579 => x"802e9e38",
          5580 => x"767f5370",
          5581 => x"5254dba8",
          5582 => x"3f81cbd4",
          5583 => x"0894150c",
          5584 => x"8e3981cb",
          5585 => x"d408842e",
          5586 => x"09810683",
          5587 => x"38855574",
          5588 => x"81cbd40c",
          5589 => x"933d0d04",
          5590 => x"e43d0d6f",
          5591 => x"6f5b5b80",
          5592 => x"7a348053",
          5593 => x"9e3dffb8",
          5594 => x"05529f3d",
          5595 => x"51e8b53f",
          5596 => x"81cbd408",
          5597 => x"5781cbd4",
          5598 => x"0882fc38",
          5599 => x"7b437a7c",
          5600 => x"94110847",
          5601 => x"55586454",
          5602 => x"73802e81",
          5603 => x"ed38a052",
          5604 => x"933d7052",
          5605 => x"55d5ea3f",
          5606 => x"81cbd408",
          5607 => x"5781cbd4",
          5608 => x"0882d438",
          5609 => x"68527b51",
          5610 => x"c9c83f81",
          5611 => x"cbd40857",
          5612 => x"81cbd408",
          5613 => x"82c13869",
          5614 => x"527b51da",
          5615 => x"a33f81cb",
          5616 => x"d4084576",
          5617 => x"527451d5",
          5618 => x"b83f81cb",
          5619 => x"d4085781",
          5620 => x"cbd40882",
          5621 => x"a2388052",
          5622 => x"7451daeb",
          5623 => x"3f81cbd4",
          5624 => x"085781cb",
          5625 => x"d408a438",
          5626 => x"69527b51",
          5627 => x"d9f23f73",
          5628 => x"81cbd408",
          5629 => x"2ea63876",
          5630 => x"527451d6",
          5631 => x"cf3f81cb",
          5632 => x"d4085781",
          5633 => x"cbd40880",
          5634 => x"2ecc3876",
          5635 => x"842e0981",
          5636 => x"06863882",
          5637 => x"5781e039",
          5638 => x"7681dc38",
          5639 => x"9e3dffbc",
          5640 => x"05527451",
          5641 => x"dcc93f76",
          5642 => x"903d7811",
          5643 => x"81113351",
          5644 => x"565a5673",
          5645 => x"802e9138",
          5646 => x"02b90555",
          5647 => x"81168116",
          5648 => x"70335656",
          5649 => x"5673f538",
          5650 => x"81165473",
          5651 => x"78268190",
          5652 => x"3875802e",
          5653 => x"99387816",
          5654 => x"810555ff",
          5655 => x"186f11ff",
          5656 => x"18ff1858",
          5657 => x"58555874",
          5658 => x"33743475",
          5659 => x"ee38ff18",
          5660 => x"6f115558",
          5661 => x"af7434fe",
          5662 => x"8d39777b",
          5663 => x"2e098106",
          5664 => x"8a38ff18",
          5665 => x"6f115558",
          5666 => x"af743480",
          5667 => x"0b81cc84",
          5668 => x"33708429",
          5669 => x"81bba005",
          5670 => x"70087033",
          5671 => x"525c5656",
          5672 => x"5673762e",
          5673 => x"8d388116",
          5674 => x"701a7033",
          5675 => x"51555673",
          5676 => x"f5388216",
          5677 => x"54737826",
          5678 => x"a7388055",
          5679 => x"74762791",
          5680 => x"38741954",
          5681 => x"73337a70",
          5682 => x"81055c34",
          5683 => x"811555ec",
          5684 => x"39ba7a70",
          5685 => x"81055c34",
          5686 => x"74ff2e09",
          5687 => x"81068538",
          5688 => x"91579439",
          5689 => x"6e188119",
          5690 => x"59547333",
          5691 => x"7a708105",
          5692 => x"5c347a78",
          5693 => x"26ee3880",
          5694 => x"7a347681",
          5695 => x"cbd40c9e",
          5696 => x"3d0d04f7",
          5697 => x"3d0d7b7d",
          5698 => x"8d3dfc05",
          5699 => x"54715357",
          5700 => x"55ecbb3f",
          5701 => x"81cbd408",
          5702 => x"5381cbd4",
          5703 => x"0882fa38",
          5704 => x"91153353",
          5705 => x"7282f238",
          5706 => x"8c150854",
          5707 => x"73762792",
          5708 => x"38901533",
          5709 => x"70812a70",
          5710 => x"81065154",
          5711 => x"57728338",
          5712 => x"73569415",
          5713 => x"08548070",
          5714 => x"94170c58",
          5715 => x"75782e82",
          5716 => x"9738798a",
          5717 => x"11227089",
          5718 => x"2b595153",
          5719 => x"73782eb7",
          5720 => x"387652ff",
          5721 => x"1651ff9b",
          5722 => x"e53f81cb",
          5723 => x"d408ff15",
          5724 => x"78547053",
          5725 => x"5553ff9b",
          5726 => x"d53f81cb",
          5727 => x"d4087326",
          5728 => x"96387630",
          5729 => x"70750670",
          5730 => x"94180c77",
          5731 => x"71319818",
          5732 => x"08575851",
          5733 => x"53b13988",
          5734 => x"15085473",
          5735 => x"a6387352",
          5736 => x"7451cdca",
          5737 => x"3f81cbd4",
          5738 => x"085481cb",
          5739 => x"d408812e",
          5740 => x"819a3881",
          5741 => x"cbd408ff",
          5742 => x"2e819b38",
          5743 => x"81cbd408",
          5744 => x"88160c73",
          5745 => x"98160c73",
          5746 => x"802e819c",
          5747 => x"38767627",
          5748 => x"80dc3875",
          5749 => x"77319416",
          5750 => x"08189417",
          5751 => x"0c901633",
          5752 => x"70812a70",
          5753 => x"81065155",
          5754 => x"5a567280",
          5755 => x"2e9a3873",
          5756 => x"527451cc",
          5757 => x"f93f81cb",
          5758 => x"d4085481",
          5759 => x"cbd40894",
          5760 => x"3881cbd4",
          5761 => x"0856a739",
          5762 => x"73527451",
          5763 => x"c7843f81",
          5764 => x"cbd40854",
          5765 => x"73ff2ebe",
          5766 => x"38817427",
          5767 => x"af387953",
          5768 => x"73981408",
          5769 => x"27a63873",
          5770 => x"98160cff",
          5771 => x"a0399415",
          5772 => x"08169416",
          5773 => x"0c7583ff",
          5774 => x"06537280",
          5775 => x"2eaa3873",
          5776 => x"527951c6",
          5777 => x"a33f81cb",
          5778 => x"d4089438",
          5779 => x"820b9116",
          5780 => x"34825380",
          5781 => x"c439810b",
          5782 => x"91163481",
          5783 => x"53bb3975",
          5784 => x"892a81cb",
          5785 => x"d4080558",
          5786 => x"94150854",
          5787 => x"8c150874",
          5788 => x"27903873",
          5789 => x"8c160c90",
          5790 => x"153380c0",
          5791 => x"07537290",
          5792 => x"16347383",
          5793 => x"ff065372",
          5794 => x"802e8c38",
          5795 => x"779c1608",
          5796 => x"2e853877",
          5797 => x"9c160c80",
          5798 => x"537281cb",
          5799 => x"d40c8b3d",
          5800 => x"0d04f93d",
          5801 => x"0d795689",
          5802 => x"5475802e",
          5803 => x"818a3880",
          5804 => x"53893dfc",
          5805 => x"05528a3d",
          5806 => x"840551e1",
          5807 => x"e73f81cb",
          5808 => x"d4085581",
          5809 => x"cbd40880",
          5810 => x"ea387776",
          5811 => x"0c7a5275",
          5812 => x"51d8b53f",
          5813 => x"81cbd408",
          5814 => x"5581cbd4",
          5815 => x"0880c338",
          5816 => x"ab163370",
          5817 => x"982b5557",
          5818 => x"807424a2",
          5819 => x"38861633",
          5820 => x"70842a70",
          5821 => x"81065155",
          5822 => x"5773802e",
          5823 => x"ad389c16",
          5824 => x"08527751",
          5825 => x"d3da3f81",
          5826 => x"cbd40888",
          5827 => x"170c7754",
          5828 => x"86142284",
          5829 => x"17237452",
          5830 => x"7551cee5",
          5831 => x"3f81cbd4",
          5832 => x"08557484",
          5833 => x"2e098106",
          5834 => x"85388555",
          5835 => x"86397480",
          5836 => x"2e843880",
          5837 => x"760c7454",
          5838 => x"7381cbd4",
          5839 => x"0c893d0d",
          5840 => x"04fc3d0d",
          5841 => x"76873dfc",
          5842 => x"05537052",
          5843 => x"53e7ff3f",
          5844 => x"81cbd408",
          5845 => x"873881cb",
          5846 => x"d408730c",
          5847 => x"863d0d04",
          5848 => x"fb3d0d77",
          5849 => x"79893dfc",
          5850 => x"05547153",
          5851 => x"5654e7de",
          5852 => x"3f81cbd4",
          5853 => x"085381cb",
          5854 => x"d40880df",
          5855 => x"38749338",
          5856 => x"81cbd408",
          5857 => x"527351cd",
          5858 => x"f83f81cb",
          5859 => x"d4085380",
          5860 => x"ca3981cb",
          5861 => x"d4085273",
          5862 => x"51d3ac3f",
          5863 => x"81cbd408",
          5864 => x"5381cbd4",
          5865 => x"08842e09",
          5866 => x"81068538",
          5867 => x"80538739",
          5868 => x"81cbd408",
          5869 => x"a6387452",
          5870 => x"7351d5b3",
          5871 => x"3f725273",
          5872 => x"51cf893f",
          5873 => x"81cbd408",
          5874 => x"84327030",
          5875 => x"7072079f",
          5876 => x"2c7081cb",
          5877 => x"d4080651",
          5878 => x"51545472",
          5879 => x"81cbd40c",
          5880 => x"873d0d04",
          5881 => x"ee3d0d65",
          5882 => x"57805389",
          5883 => x"3d705396",
          5884 => x"3d5256df",
          5885 => x"af3f81cb",
          5886 => x"d4085581",
          5887 => x"cbd408b2",
          5888 => x"38645275",
          5889 => x"51d6813f",
          5890 => x"81cbd408",
          5891 => x"5581cbd4",
          5892 => x"08a03802",
          5893 => x"80cb0533",
          5894 => x"70982b55",
          5895 => x"58738025",
          5896 => x"85388655",
          5897 => x"8d397680",
          5898 => x"2e883876",
          5899 => x"527551d4",
          5900 => x"be3f7481",
          5901 => x"cbd40c94",
          5902 => x"3d0d04f0",
          5903 => x"3d0d6365",
          5904 => x"555c8053",
          5905 => x"923dec05",
          5906 => x"52933d51",
          5907 => x"ded63f81",
          5908 => x"cbd4085b",
          5909 => x"81cbd408",
          5910 => x"8280387c",
          5911 => x"740c7308",
          5912 => x"981108fe",
          5913 => x"11901308",
          5914 => x"59565855",
          5915 => x"75742691",
          5916 => x"38757c0c",
          5917 => x"81e43981",
          5918 => x"5b81cc39",
          5919 => x"825b81c7",
          5920 => x"3981cbd4",
          5921 => x"08753355",
          5922 => x"5973812e",
          5923 => x"098106bf",
          5924 => x"3882755f",
          5925 => x"57765292",
          5926 => x"3df00551",
          5927 => x"c1f43f81",
          5928 => x"cbd408ff",
          5929 => x"2ed13881",
          5930 => x"cbd40881",
          5931 => x"2ece3881",
          5932 => x"cbd40830",
          5933 => x"7081cbd4",
          5934 => x"08078025",
          5935 => x"7a058119",
          5936 => x"7f53595a",
          5937 => x"54981408",
          5938 => x"7726ca38",
          5939 => x"80f939a4",
          5940 => x"150881cb",
          5941 => x"d4085758",
          5942 => x"75983877",
          5943 => x"5281187d",
          5944 => x"5258ffbf",
          5945 => x"8d3f81cb",
          5946 => x"d4085b81",
          5947 => x"cbd40880",
          5948 => x"d6387c70",
          5949 => x"337712ff",
          5950 => x"1a5d5256",
          5951 => x"5474822e",
          5952 => x"0981069e",
          5953 => x"38b41451",
          5954 => x"ffbbcb3f",
          5955 => x"81cbd408",
          5956 => x"83ffff06",
          5957 => x"70307080",
          5958 => x"251b8219",
          5959 => x"595b5154",
          5960 => x"9b39b414",
          5961 => x"51ffbbc5",
          5962 => x"3f81cbd4",
          5963 => x"08f00a06",
          5964 => x"70307080",
          5965 => x"251b8419",
          5966 => x"595b5154",
          5967 => x"7583ff06",
          5968 => x"7a585679",
          5969 => x"ff923878",
          5970 => x"7c0c7c79",
          5971 => x"90120c84",
          5972 => x"11338107",
          5973 => x"56547484",
          5974 => x"15347a81",
          5975 => x"cbd40c92",
          5976 => x"3d0d04f9",
          5977 => x"3d0d798a",
          5978 => x"3dfc0553",
          5979 => x"705257e3",
          5980 => x"dd3f81cb",
          5981 => x"d4085681",
          5982 => x"cbd40881",
          5983 => x"a8389117",
          5984 => x"33567581",
          5985 => x"a0389017",
          5986 => x"3370812a",
          5987 => x"70810651",
          5988 => x"55558755",
          5989 => x"73802e81",
          5990 => x"8e389417",
          5991 => x"0854738c",
          5992 => x"18082781",
          5993 => x"8038739b",
          5994 => x"3881cbd4",
          5995 => x"08538817",
          5996 => x"08527651",
          5997 => x"c48c3f81",
          5998 => x"cbd40874",
          5999 => x"88190c56",
          6000 => x"80c93998",
          6001 => x"17085276",
          6002 => x"51ffbfc6",
          6003 => x"3f81cbd4",
          6004 => x"08ff2e09",
          6005 => x"81068338",
          6006 => x"815681cb",
          6007 => x"d408812e",
          6008 => x"09810685",
          6009 => x"388256a3",
          6010 => x"3975a038",
          6011 => x"775481cb",
          6012 => x"d4089815",
          6013 => x"08279438",
          6014 => x"98170853",
          6015 => x"81cbd408",
          6016 => x"527651c3",
          6017 => x"bd3f81cb",
          6018 => x"d4085694",
          6019 => x"17088c18",
          6020 => x"0c901733",
          6021 => x"80c00754",
          6022 => x"73901834",
          6023 => x"75802e85",
          6024 => x"38759118",
          6025 => x"34755574",
          6026 => x"81cbd40c",
          6027 => x"893d0d04",
          6028 => x"e23d0d82",
          6029 => x"53a03dff",
          6030 => x"a40552a1",
          6031 => x"3d51dae4",
          6032 => x"3f81cbd4",
          6033 => x"085581cb",
          6034 => x"d40881f5",
          6035 => x"387845a1",
          6036 => x"3d085295",
          6037 => x"3d705258",
          6038 => x"d1ae3f81",
          6039 => x"cbd40855",
          6040 => x"81cbd408",
          6041 => x"81db3802",
          6042 => x"80fb0533",
          6043 => x"70852a70",
          6044 => x"81065155",
          6045 => x"56865573",
          6046 => x"81c73875",
          6047 => x"982b5480",
          6048 => x"742481bd",
          6049 => x"380280d6",
          6050 => x"05337081",
          6051 => x"06585487",
          6052 => x"557681ad",
          6053 => x"386b5278",
          6054 => x"51ccc53f",
          6055 => x"81cbd408",
          6056 => x"74842a70",
          6057 => x"81065155",
          6058 => x"5673802e",
          6059 => x"80d43878",
          6060 => x"5481cbd4",
          6061 => x"08941508",
          6062 => x"2e818638",
          6063 => x"735a81cb",
          6064 => x"d4085c76",
          6065 => x"528a3d70",
          6066 => x"5254c7b5",
          6067 => x"3f81cbd4",
          6068 => x"085581cb",
          6069 => x"d40880e9",
          6070 => x"3881cbd4",
          6071 => x"08527351",
          6072 => x"cce53f81",
          6073 => x"cbd40855",
          6074 => x"81cbd408",
          6075 => x"86388755",
          6076 => x"80cf3981",
          6077 => x"cbd40884",
          6078 => x"2e883881",
          6079 => x"cbd40880",
          6080 => x"c0387751",
          6081 => x"cec23f81",
          6082 => x"cbd40881",
          6083 => x"cbd40830",
          6084 => x"7081cbd4",
          6085 => x"08078025",
          6086 => x"51555575",
          6087 => x"802e9438",
          6088 => x"73802e8f",
          6089 => x"38805375",
          6090 => x"527751c1",
          6091 => x"953f81cb",
          6092 => x"d4085574",
          6093 => x"8c387851",
          6094 => x"ffbafe3f",
          6095 => x"81cbd408",
          6096 => x"557481cb",
          6097 => x"d40ca03d",
          6098 => x"0d04e93d",
          6099 => x"0d825399",
          6100 => x"3dc00552",
          6101 => x"9a3d51d8",
          6102 => x"cb3f81cb",
          6103 => x"d4085481",
          6104 => x"cbd40882",
          6105 => x"b038785e",
          6106 => x"69528e3d",
          6107 => x"705258cf",
          6108 => x"973f81cb",
          6109 => x"d4085481",
          6110 => x"cbd40886",
          6111 => x"38885482",
          6112 => x"943981cb",
          6113 => x"d408842e",
          6114 => x"09810682",
          6115 => x"88380280",
          6116 => x"df053370",
          6117 => x"852a8106",
          6118 => x"51558654",
          6119 => x"7481f638",
          6120 => x"785a7452",
          6121 => x"8a3d7052",
          6122 => x"57c1c33f",
          6123 => x"81cbd408",
          6124 => x"75555681",
          6125 => x"cbd40883",
          6126 => x"38875481",
          6127 => x"cbd40881",
          6128 => x"2e098106",
          6129 => x"83388254",
          6130 => x"81cbd408",
          6131 => x"ff2e0981",
          6132 => x"06863881",
          6133 => x"5481b439",
          6134 => x"7381b038",
          6135 => x"81cbd408",
          6136 => x"527851c4",
          6137 => x"a43f81cb",
          6138 => x"d4085481",
          6139 => x"cbd40881",
          6140 => x"9a388b53",
          6141 => x"a052b419",
          6142 => x"51ffb78c",
          6143 => x"3f7854ae",
          6144 => x"0bb41534",
          6145 => x"7854900b",
          6146 => x"bf153482",
          6147 => x"88b20a52",
          6148 => x"80ca1951",
          6149 => x"ffb69f3f",
          6150 => x"755378b4",
          6151 => x"115351c9",
          6152 => x"f83fa053",
          6153 => x"78b41153",
          6154 => x"80d40551",
          6155 => x"ffb6b63f",
          6156 => x"7854ae0b",
          6157 => x"80d51534",
          6158 => x"7f537880",
          6159 => x"d4115351",
          6160 => x"c9d73f78",
          6161 => x"54810b83",
          6162 => x"15347751",
          6163 => x"cba43f81",
          6164 => x"cbd40854",
          6165 => x"81cbd408",
          6166 => x"b2388288",
          6167 => x"b20a5264",
          6168 => x"960551ff",
          6169 => x"b5d03f75",
          6170 => x"53645278",
          6171 => x"51c9aa3f",
          6172 => x"6454900b",
          6173 => x"8b153478",
          6174 => x"54810b83",
          6175 => x"15347851",
          6176 => x"ffb8b63f",
          6177 => x"81cbd408",
          6178 => x"548b3980",
          6179 => x"53755276",
          6180 => x"51ffbeae",
          6181 => x"3f7381cb",
          6182 => x"d40c993d",
          6183 => x"0d04da3d",
          6184 => x"0da93d84",
          6185 => x"0551d2f1",
          6186 => x"3f8253a8",
          6187 => x"3dff8405",
          6188 => x"52a93d51",
          6189 => x"d5ee3f81",
          6190 => x"cbd40855",
          6191 => x"81cbd408",
          6192 => x"82d33878",
          6193 => x"4da93d08",
          6194 => x"529d3d70",
          6195 => x"5258ccb8",
          6196 => x"3f81cbd4",
          6197 => x"085581cb",
          6198 => x"d40882b9",
          6199 => x"3802819b",
          6200 => x"053381a0",
          6201 => x"06548655",
          6202 => x"7382aa38",
          6203 => x"a053a43d",
          6204 => x"0852a83d",
          6205 => x"ff880551",
          6206 => x"ffb4ea3f",
          6207 => x"ac537752",
          6208 => x"923d7052",
          6209 => x"54ffb4dd",
          6210 => x"3faa3d08",
          6211 => x"527351cb",
          6212 => x"f73f81cb",
          6213 => x"d4085581",
          6214 => x"cbd40895",
          6215 => x"38636f2e",
          6216 => x"09810688",
          6217 => x"3865a23d",
          6218 => x"082e9238",
          6219 => x"885581e5",
          6220 => x"3981cbd4",
          6221 => x"08842e09",
          6222 => x"810681b8",
          6223 => x"387351c9",
          6224 => x"b13f81cb",
          6225 => x"d4085581",
          6226 => x"cbd40881",
          6227 => x"c8386856",
          6228 => x"9353a83d",
          6229 => x"ff950552",
          6230 => x"8d1651ff",
          6231 => x"b4873f02",
          6232 => x"af05338b",
          6233 => x"17348b16",
          6234 => x"3370842a",
          6235 => x"70810651",
          6236 => x"55557389",
          6237 => x"3874a007",
          6238 => x"54738b17",
          6239 => x"34785481",
          6240 => x"0b831534",
          6241 => x"8b163370",
          6242 => x"842a7081",
          6243 => x"06515555",
          6244 => x"73802e80",
          6245 => x"e5386e64",
          6246 => x"2e80df38",
          6247 => x"75527851",
          6248 => x"c6be3f81",
          6249 => x"cbd40852",
          6250 => x"7851ffb7",
          6251 => x"bb3f8255",
          6252 => x"81cbd408",
          6253 => x"802e80dd",
          6254 => x"3881cbd4",
          6255 => x"08527851",
          6256 => x"ffb5af3f",
          6257 => x"81cbd408",
          6258 => x"7980d411",
          6259 => x"58585581",
          6260 => x"cbd40880",
          6261 => x"c0388116",
          6262 => x"335473ae",
          6263 => x"2e098106",
          6264 => x"99386353",
          6265 => x"75527651",
          6266 => x"c6af3f78",
          6267 => x"54810b83",
          6268 => x"15348739",
          6269 => x"81cbd408",
          6270 => x"9c387751",
          6271 => x"c8ca3f81",
          6272 => x"cbd40855",
          6273 => x"81cbd408",
          6274 => x"8c387851",
          6275 => x"ffb5aa3f",
          6276 => x"81cbd408",
          6277 => x"557481cb",
          6278 => x"d40ca83d",
          6279 => x"0d04ed3d",
          6280 => x"0d0280db",
          6281 => x"05330284",
          6282 => x"0580df05",
          6283 => x"33575782",
          6284 => x"53953dd0",
          6285 => x"0552963d",
          6286 => x"51d2e93f",
          6287 => x"81cbd408",
          6288 => x"5581cbd4",
          6289 => x"0880cf38",
          6290 => x"785a6552",
          6291 => x"953dd405",
          6292 => x"51c9b53f",
          6293 => x"81cbd408",
          6294 => x"5581cbd4",
          6295 => x"08b83802",
          6296 => x"80cf0533",
          6297 => x"81a00654",
          6298 => x"865573aa",
          6299 => x"3875a706",
          6300 => x"6171098b",
          6301 => x"12337106",
          6302 => x"7a740607",
          6303 => x"51575556",
          6304 => x"748b1534",
          6305 => x"7854810b",
          6306 => x"83153478",
          6307 => x"51ffb4a9",
          6308 => x"3f81cbd4",
          6309 => x"08557481",
          6310 => x"cbd40c95",
          6311 => x"3d0d04ef",
          6312 => x"3d0d6456",
          6313 => x"8253933d",
          6314 => x"d0055294",
          6315 => x"3d51d1f4",
          6316 => x"3f81cbd4",
          6317 => x"085581cb",
          6318 => x"d40880cb",
          6319 => x"38765863",
          6320 => x"52933dd4",
          6321 => x"0551c8c0",
          6322 => x"3f81cbd4",
          6323 => x"085581cb",
          6324 => x"d408b438",
          6325 => x"0280c705",
          6326 => x"3381a006",
          6327 => x"54865573",
          6328 => x"a6388416",
          6329 => x"22861722",
          6330 => x"71902b07",
          6331 => x"5354961f",
          6332 => x"51ffb0c2",
          6333 => x"3f765481",
          6334 => x"0b831534",
          6335 => x"7651ffb3",
          6336 => x"b83f81cb",
          6337 => x"d4085574",
          6338 => x"81cbd40c",
          6339 => x"933d0d04",
          6340 => x"ea3d0d69",
          6341 => x"6b5c5a80",
          6342 => x"53983dd0",
          6343 => x"0552993d",
          6344 => x"51d1813f",
          6345 => x"81cbd408",
          6346 => x"81cbd408",
          6347 => x"307081cb",
          6348 => x"d4080780",
          6349 => x"25515557",
          6350 => x"79802e81",
          6351 => x"85388170",
          6352 => x"75065555",
          6353 => x"73802e80",
          6354 => x"f9387b5d",
          6355 => x"805f8052",
          6356 => x"8d3d7052",
          6357 => x"54ffbea9",
          6358 => x"3f81cbd4",
          6359 => x"085781cb",
          6360 => x"d40880d1",
          6361 => x"38745273",
          6362 => x"51c3dc3f",
          6363 => x"81cbd408",
          6364 => x"5781cbd4",
          6365 => x"08bf3881",
          6366 => x"cbd40881",
          6367 => x"cbd40865",
          6368 => x"5b595678",
          6369 => x"1881197b",
          6370 => x"18565955",
          6371 => x"74337434",
          6372 => x"8116568a",
          6373 => x"7827ec38",
          6374 => x"8b56751a",
          6375 => x"54807434",
          6376 => x"75802e9e",
          6377 => x"38ff1670",
          6378 => x"1b703351",
          6379 => x"555673a0",
          6380 => x"2ee8388e",
          6381 => x"3976842e",
          6382 => x"09810686",
          6383 => x"38807a34",
          6384 => x"80577630",
          6385 => x"70780780",
          6386 => x"2551547a",
          6387 => x"802e80c1",
          6388 => x"3873802e",
          6389 => x"bc387ba0",
          6390 => x"11085351",
          6391 => x"ffb1933f",
          6392 => x"81cbd408",
          6393 => x"5781cbd4",
          6394 => x"08a7387b",
          6395 => x"70335555",
          6396 => x"80c35673",
          6397 => x"832e8b38",
          6398 => x"80e45673",
          6399 => x"842e8338",
          6400 => x"a7567515",
          6401 => x"b40551ff",
          6402 => x"ade33f81",
          6403 => x"cbd4087b",
          6404 => x"0c7681cb",
          6405 => x"d40c983d",
          6406 => x"0d04e63d",
          6407 => x"0d82539c",
          6408 => x"3dffb805",
          6409 => x"529d3d51",
          6410 => x"cefa3f81",
          6411 => x"cbd40881",
          6412 => x"cbd40856",
          6413 => x"5481cbd4",
          6414 => x"08839838",
          6415 => x"8b53a052",
          6416 => x"8b3d7052",
          6417 => x"59ffaec0",
          6418 => x"3f736d70",
          6419 => x"337081ff",
          6420 => x"06525755",
          6421 => x"579f7427",
          6422 => x"81bc3878",
          6423 => x"587481ff",
          6424 => x"066d8105",
          6425 => x"4e705255",
          6426 => x"ffaf893f",
          6427 => x"81cbd408",
          6428 => x"802ea538",
          6429 => x"6c703370",
          6430 => x"535754ff",
          6431 => x"aefd3f81",
          6432 => x"cbd40880",
          6433 => x"2e8d3874",
          6434 => x"882b7607",
          6435 => x"6d81054e",
          6436 => x"55863981",
          6437 => x"cbd40855",
          6438 => x"ff9f1570",
          6439 => x"83ffff06",
          6440 => x"51547399",
          6441 => x"268a38e0",
          6442 => x"157083ff",
          6443 => x"ff065654",
          6444 => x"80ff7527",
          6445 => x"873881ba",
          6446 => x"b0153355",
          6447 => x"74802ea3",
          6448 => x"38745281",
          6449 => x"bcb051ff",
          6450 => x"ae893f81",
          6451 => x"cbd40893",
          6452 => x"3881ff75",
          6453 => x"27883876",
          6454 => x"89268838",
          6455 => x"8b398a77",
          6456 => x"27863886",
          6457 => x"5581ec39",
          6458 => x"81ff7527",
          6459 => x"8f387488",
          6460 => x"2a547378",
          6461 => x"7081055a",
          6462 => x"34811757",
          6463 => x"74787081",
          6464 => x"055a3481",
          6465 => x"176d7033",
          6466 => x"7081ff06",
          6467 => x"52575557",
          6468 => x"739f26fe",
          6469 => x"c8388b3d",
          6470 => x"33548655",
          6471 => x"7381e52e",
          6472 => x"81b13876",
          6473 => x"802e9938",
          6474 => x"02a70555",
          6475 => x"76157033",
          6476 => x"515473a0",
          6477 => x"2e098106",
          6478 => x"8738ff17",
          6479 => x"5776ed38",
          6480 => x"79418043",
          6481 => x"8052913d",
          6482 => x"705255ff",
          6483 => x"bab33f81",
          6484 => x"cbd40854",
          6485 => x"81cbd408",
          6486 => x"80f73881",
          6487 => x"527451ff",
          6488 => x"bfe53f81",
          6489 => x"cbd40854",
          6490 => x"81cbd408",
          6491 => x"8d387680",
          6492 => x"c4386754",
          6493 => x"e5743480",
          6494 => x"c63981cb",
          6495 => x"d408842e",
          6496 => x"09810680",
          6497 => x"cc388054",
          6498 => x"76742e80",
          6499 => x"c4388152",
          6500 => x"7451ffbd",
          6501 => x"b03f81cb",
          6502 => x"d4085481",
          6503 => x"cbd408b1",
          6504 => x"38a05381",
          6505 => x"cbd40852",
          6506 => x"6751ffab",
          6507 => x"db3f6754",
          6508 => x"880b8b15",
          6509 => x"348b5378",
          6510 => x"526751ff",
          6511 => x"aba73f79",
          6512 => x"54810b83",
          6513 => x"15347951",
          6514 => x"ffadee3f",
          6515 => x"81cbd408",
          6516 => x"54735574",
          6517 => x"81cbd40c",
          6518 => x"9c3d0d04",
          6519 => x"f23d0d60",
          6520 => x"62028805",
          6521 => x"80cb0533",
          6522 => x"933dfc05",
          6523 => x"55725440",
          6524 => x"5e5ad2da",
          6525 => x"3f81cbd4",
          6526 => x"085881cb",
          6527 => x"d40882bd",
          6528 => x"38911a33",
          6529 => x"587782b5",
          6530 => x"387c802e",
          6531 => x"97388c1a",
          6532 => x"08597890",
          6533 => x"38901a33",
          6534 => x"70812a70",
          6535 => x"81065155",
          6536 => x"55739038",
          6537 => x"87548297",
          6538 => x"39825882",
          6539 => x"90398158",
          6540 => x"828b397e",
          6541 => x"8a112270",
          6542 => x"892b7055",
          6543 => x"7f545656",
          6544 => x"56ff828a",
          6545 => x"3fff147d",
          6546 => x"06703070",
          6547 => x"72079f2a",
          6548 => x"81cbd408",
          6549 => x"058c1908",
          6550 => x"7c405a5d",
          6551 => x"55558177",
          6552 => x"27883898",
          6553 => x"16087726",
          6554 => x"83388257",
          6555 => x"76775659",
          6556 => x"80567452",
          6557 => x"7951ffae",
          6558 => x"993f8115",
          6559 => x"7f555598",
          6560 => x"14087526",
          6561 => x"83388255",
          6562 => x"81cbd408",
          6563 => x"812eff99",
          6564 => x"3881cbd4",
          6565 => x"08ff2eff",
          6566 => x"953881cb",
          6567 => x"d4088e38",
          6568 => x"81165675",
          6569 => x"7b2e0981",
          6570 => x"06873893",
          6571 => x"39745980",
          6572 => x"5674772e",
          6573 => x"098106ff",
          6574 => x"b9388758",
          6575 => x"80ff397d",
          6576 => x"802eba38",
          6577 => x"787b5555",
          6578 => x"7a802eb4",
          6579 => x"38811556",
          6580 => x"73812e09",
          6581 => x"81068338",
          6582 => x"ff567553",
          6583 => x"74527e51",
          6584 => x"ffafa83f",
          6585 => x"81cbd408",
          6586 => x"5881cbd4",
          6587 => x"0880ce38",
          6588 => x"748116ff",
          6589 => x"1656565c",
          6590 => x"73d33884",
          6591 => x"39ff195c",
          6592 => x"7e7c8c12",
          6593 => x"0c557d80",
          6594 => x"2eb33878",
          6595 => x"881b0c7c",
          6596 => x"8c1b0c90",
          6597 => x"1a3380c0",
          6598 => x"07547390",
          6599 => x"1b349815",
          6600 => x"08fe0590",
          6601 => x"16085754",
          6602 => x"75742691",
          6603 => x"38757b31",
          6604 => x"90160c84",
          6605 => x"15338107",
          6606 => x"54738416",
          6607 => x"34775473",
          6608 => x"81cbd40c",
          6609 => x"903d0d04",
          6610 => x"e93d0d6b",
          6611 => x"6d028805",
          6612 => x"80eb0533",
          6613 => x"9d3d545a",
          6614 => x"5c59c5bd",
          6615 => x"3f8b5680",
          6616 => x"0b81cbd4",
          6617 => x"08248bf8",
          6618 => x"3881cbd4",
          6619 => x"08842981",
          6620 => x"cbf00570",
          6621 => x"08515574",
          6622 => x"802e8438",
          6623 => x"80753481",
          6624 => x"cbd40881",
          6625 => x"ff065f81",
          6626 => x"527e51ff",
          6627 => x"a0d03f81",
          6628 => x"cbd40881",
          6629 => x"ff067081",
          6630 => x"06565783",
          6631 => x"56748bc0",
          6632 => x"3876822a",
          6633 => x"70810651",
          6634 => x"558a5674",
          6635 => x"8bb23899",
          6636 => x"3dfc0553",
          6637 => x"83527e51",
          6638 => x"ffa4f03f",
          6639 => x"81cbd408",
          6640 => x"99386755",
          6641 => x"74802e92",
          6642 => x"38748280",
          6643 => x"80268b38",
          6644 => x"ff157506",
          6645 => x"5574802e",
          6646 => x"83388148",
          6647 => x"78802e87",
          6648 => x"38848079",
          6649 => x"26923878",
          6650 => x"81800a26",
          6651 => x"8b38ff19",
          6652 => x"79065574",
          6653 => x"802e8638",
          6654 => x"93568ae4",
          6655 => x"3978892a",
          6656 => x"6e892a70",
          6657 => x"892b7759",
          6658 => x"4843597a",
          6659 => x"83388156",
          6660 => x"61307080",
          6661 => x"25770751",
          6662 => x"55915674",
          6663 => x"8ac23899",
          6664 => x"3df80553",
          6665 => x"81527e51",
          6666 => x"ffa4803f",
          6667 => x"815681cb",
          6668 => x"d4088aac",
          6669 => x"3877832a",
          6670 => x"70770681",
          6671 => x"cbd40843",
          6672 => x"56457483",
          6673 => x"38bf4166",
          6674 => x"558e5660",
          6675 => x"75268a90",
          6676 => x"38746131",
          6677 => x"70485580",
          6678 => x"ff75278a",
          6679 => x"83389356",
          6680 => x"78818026",
          6681 => x"89fa3877",
          6682 => x"812a7081",
          6683 => x"06564374",
          6684 => x"802e9538",
          6685 => x"77870655",
          6686 => x"74822e83",
          6687 => x"8d387781",
          6688 => x"06557480",
          6689 => x"2e838338",
          6690 => x"77810655",
          6691 => x"9356825e",
          6692 => x"74802e89",
          6693 => x"cb38785a",
          6694 => x"7d832e09",
          6695 => x"810680e1",
          6696 => x"3878ae38",
          6697 => x"66912a57",
          6698 => x"810b81bc",
          6699 => x"d422565a",
          6700 => x"74802e9d",
          6701 => x"38747726",
          6702 => x"983881bc",
          6703 => x"d4567910",
          6704 => x"82177022",
          6705 => x"57575a74",
          6706 => x"802e8638",
          6707 => x"767527ee",
          6708 => x"38795266",
          6709 => x"51fefcf6",
          6710 => x"3f81cbd4",
          6711 => x"08842984",
          6712 => x"87057089",
          6713 => x"2a5e55a0",
          6714 => x"5c800b81",
          6715 => x"cbd408fc",
          6716 => x"808a0556",
          6717 => x"44fdfff0",
          6718 => x"0a752780",
          6719 => x"ec3888d3",
          6720 => x"3978ae38",
          6721 => x"668c2a57",
          6722 => x"810b81bc",
          6723 => x"c422565a",
          6724 => x"74802e9d",
          6725 => x"38747726",
          6726 => x"983881bc",
          6727 => x"c4567910",
          6728 => x"82177022",
          6729 => x"57575a74",
          6730 => x"802e8638",
          6731 => x"767527ee",
          6732 => x"38795266",
          6733 => x"51fefc96",
          6734 => x"3f81cbd4",
          6735 => x"08108405",
          6736 => x"5781cbd4",
          6737 => x"089ff526",
          6738 => x"9638810b",
          6739 => x"81cbd408",
          6740 => x"1081cbd4",
          6741 => x"08057111",
          6742 => x"722a8305",
          6743 => x"59565e83",
          6744 => x"ff17892a",
          6745 => x"5d815ca0",
          6746 => x"44601c7d",
          6747 => x"11650569",
          6748 => x"7012ff05",
          6749 => x"71307072",
          6750 => x"0674315c",
          6751 => x"52595759",
          6752 => x"407d832e",
          6753 => x"09810689",
          6754 => x"38761c60",
          6755 => x"18415c84",
          6756 => x"39761d5d",
          6757 => x"79902918",
          6758 => x"70623168",
          6759 => x"58515574",
          6760 => x"762687af",
          6761 => x"38757c31",
          6762 => x"7d317a53",
          6763 => x"70653152",
          6764 => x"55fefb9a",
          6765 => x"3f81cbd4",
          6766 => x"08587d83",
          6767 => x"2e098106",
          6768 => x"9b3881cb",
          6769 => x"d40883ff",
          6770 => x"f52680dd",
          6771 => x"38788783",
          6772 => x"3879812a",
          6773 => x"5978fdbe",
          6774 => x"3886f839",
          6775 => x"7d822e09",
          6776 => x"810680c5",
          6777 => x"3883fff5",
          6778 => x"0b81cbd4",
          6779 => x"0827a038",
          6780 => x"788f3879",
          6781 => x"1a557480",
          6782 => x"c0268638",
          6783 => x"7459fd96",
          6784 => x"39628106",
          6785 => x"5574802e",
          6786 => x"8f38835e",
          6787 => x"fd883981",
          6788 => x"cbd4089f",
          6789 => x"f5269238",
          6790 => x"7886b838",
          6791 => x"791a5981",
          6792 => x"807927fc",
          6793 => x"f13886ab",
          6794 => x"3980557d",
          6795 => x"812e0981",
          6796 => x"0683387d",
          6797 => x"559ff578",
          6798 => x"278b3874",
          6799 => x"8106558e",
          6800 => x"5674869c",
          6801 => x"38848053",
          6802 => x"80527a51",
          6803 => x"ffa2b93f",
          6804 => x"8b5381ba",
          6805 => x"ec527a51",
          6806 => x"ffa28a3f",
          6807 => x"8480528b",
          6808 => x"1b51ffa1",
          6809 => x"b33f798d",
          6810 => x"1c347b83",
          6811 => x"ffff0652",
          6812 => x"8e1b51ff",
          6813 => x"a1a23f81",
          6814 => x"0b901c34",
          6815 => x"7d833270",
          6816 => x"3070962a",
          6817 => x"84800654",
          6818 => x"5155911b",
          6819 => x"51ffa188",
          6820 => x"3f665574",
          6821 => x"83ffff26",
          6822 => x"90387483",
          6823 => x"ffff0652",
          6824 => x"931b51ff",
          6825 => x"a0f23f8a",
          6826 => x"397452a0",
          6827 => x"1b51ffa1",
          6828 => x"853ff80b",
          6829 => x"951c34bf",
          6830 => x"52981b51",
          6831 => x"ffa0d93f",
          6832 => x"81ff529a",
          6833 => x"1b51ffa0",
          6834 => x"cf3f6052",
          6835 => x"9c1b51ff",
          6836 => x"a0e43f7d",
          6837 => x"832e0981",
          6838 => x"0680cb38",
          6839 => x"8288b20a",
          6840 => x"5280c31b",
          6841 => x"51ffa0ce",
          6842 => x"3f7c52a4",
          6843 => x"1b51ffa0",
          6844 => x"c53f8252",
          6845 => x"ac1b51ff",
          6846 => x"a0bc3f81",
          6847 => x"52b01b51",
          6848 => x"ffa0953f",
          6849 => x"8652b21b",
          6850 => x"51ffa08c",
          6851 => x"3fff800b",
          6852 => x"80c01c34",
          6853 => x"a90b80c2",
          6854 => x"1c349353",
          6855 => x"81baf852",
          6856 => x"80c71b51",
          6857 => x"ae398288",
          6858 => x"b20a52a7",
          6859 => x"1b51ffa0",
          6860 => x"853f7c83",
          6861 => x"ffff0652",
          6862 => x"961b51ff",
          6863 => x"9fda3fff",
          6864 => x"800ba41c",
          6865 => x"34a90ba6",
          6866 => x"1c349353",
          6867 => x"81bb8c52",
          6868 => x"ab1b51ff",
          6869 => x"a08f3f82",
          6870 => x"d4d55283",
          6871 => x"fe1b7052",
          6872 => x"59ff9fb4",
          6873 => x"3f815460",
          6874 => x"537a527e",
          6875 => x"51ff9bd7",
          6876 => x"3f815681",
          6877 => x"cbd40883",
          6878 => x"e7387d83",
          6879 => x"2e098106",
          6880 => x"80ee3875",
          6881 => x"54608605",
          6882 => x"537a527e",
          6883 => x"51ff9bb7",
          6884 => x"3f848053",
          6885 => x"80527a51",
          6886 => x"ff9fed3f",
          6887 => x"848b85a4",
          6888 => x"d2527a51",
          6889 => x"ff9f8f3f",
          6890 => x"868a85e4",
          6891 => x"f25283e4",
          6892 => x"1b51ff9f",
          6893 => x"813fff18",
          6894 => x"5283e81b",
          6895 => x"51ff9ef6",
          6896 => x"3f825283",
          6897 => x"ec1b51ff",
          6898 => x"9eec3f82",
          6899 => x"d4d55278",
          6900 => x"51ff9ec4",
          6901 => x"3f755460",
          6902 => x"8705537a",
          6903 => x"527e51ff",
          6904 => x"9ae53f75",
          6905 => x"54601653",
          6906 => x"7a527e51",
          6907 => x"ff9ad83f",
          6908 => x"65538052",
          6909 => x"7a51ff9f",
          6910 => x"8f3f7f56",
          6911 => x"80587d83",
          6912 => x"2e098106",
          6913 => x"9a38f852",
          6914 => x"7a51ff9e",
          6915 => x"a93fff52",
          6916 => x"841b51ff",
          6917 => x"9ea03ff0",
          6918 => x"0a52881b",
          6919 => x"51913987",
          6920 => x"fffff855",
          6921 => x"7d812e83",
          6922 => x"38f85574",
          6923 => x"527a51ff",
          6924 => x"9e843f7c",
          6925 => x"55615774",
          6926 => x"62268338",
          6927 => x"74577654",
          6928 => x"75537a52",
          6929 => x"7e51ff99",
          6930 => x"fe3f81cb",
          6931 => x"d4088287",
          6932 => x"38848053",
          6933 => x"81cbd408",
          6934 => x"527a51ff",
          6935 => x"9eaa3f76",
          6936 => x"16757831",
          6937 => x"565674cd",
          6938 => x"38811858",
          6939 => x"77802eff",
          6940 => x"8d387955",
          6941 => x"7d832e83",
          6942 => x"38635561",
          6943 => x"57746226",
          6944 => x"83387457",
          6945 => x"76547553",
          6946 => x"7a527e51",
          6947 => x"ff99b83f",
          6948 => x"81cbd408",
          6949 => x"81c13876",
          6950 => x"16757831",
          6951 => x"565674db",
          6952 => x"388c567d",
          6953 => x"832e9338",
          6954 => x"86566683",
          6955 => x"ffff268a",
          6956 => x"3884567d",
          6957 => x"822e8338",
          6958 => x"81566481",
          6959 => x"06587780",
          6960 => x"fe388480",
          6961 => x"5377527a",
          6962 => x"51ff9dbc",
          6963 => x"3f82d4d5",
          6964 => x"527851ff",
          6965 => x"9cc23f83",
          6966 => x"be1b5577",
          6967 => x"7534810b",
          6968 => x"81163481",
          6969 => x"0b821634",
          6970 => x"77831634",
          6971 => x"75841634",
          6972 => x"60670556",
          6973 => x"80fdc152",
          6974 => x"7551fef4",
          6975 => x"d13ffe0b",
          6976 => x"85163481",
          6977 => x"cbd40882",
          6978 => x"2abf0756",
          6979 => x"75861634",
          6980 => x"81cbd408",
          6981 => x"87163460",
          6982 => x"5283c61b",
          6983 => x"51ff9c96",
          6984 => x"3f665283",
          6985 => x"ca1b51ff",
          6986 => x"9c8c3f81",
          6987 => x"5477537a",
          6988 => x"527e51ff",
          6989 => x"98913f81",
          6990 => x"5681cbd4",
          6991 => x"08a23880",
          6992 => x"5380527e",
          6993 => x"51ff99e3",
          6994 => x"3f815681",
          6995 => x"cbd40890",
          6996 => x"3889398e",
          6997 => x"568a3981",
          6998 => x"56863981",
          6999 => x"cbd40856",
          7000 => x"7581cbd4",
          7001 => x"0c993d0d",
          7002 => x"04ff3d0d",
          7003 => x"73527193",
          7004 => x"26818e38",
          7005 => x"71842981",
          7006 => x"b5b80552",
          7007 => x"71080481",
          7008 => x"bdec5181",
          7009 => x"803981bd",
          7010 => x"f85180f9",
          7011 => x"3981be8c",
          7012 => x"5180f239",
          7013 => x"81bea051",
          7014 => x"80eb3981",
          7015 => x"beb05180",
          7016 => x"e43981be",
          7017 => x"c05180dd",
          7018 => x"3981bed4",
          7019 => x"5180d639",
          7020 => x"81bee451",
          7021 => x"80cf3981",
          7022 => x"befc5180",
          7023 => x"c83981bf",
          7024 => x"945180c1",
          7025 => x"3981bfac",
          7026 => x"51bb3981",
          7027 => x"bfc851b5",
          7028 => x"3981bfdc",
          7029 => x"51af3981",
          7030 => x"c08851a9",
          7031 => x"3981c09c",
          7032 => x"51a33981",
          7033 => x"c0bc519d",
          7034 => x"3981c0d0",
          7035 => x"51973981",
          7036 => x"c0e85191",
          7037 => x"3981c180",
          7038 => x"518b3981",
          7039 => x"c1985185",
          7040 => x"3981c1a4",
          7041 => x"51ff87fb",
          7042 => x"3f833d0d",
          7043 => x"04fb3d0d",
          7044 => x"77795656",
          7045 => x"7487e726",
          7046 => x"8a387452",
          7047 => x"7587e829",
          7048 => x"51913987",
          7049 => x"e8527451",
          7050 => x"fef2a33f",
          7051 => x"81cbd408",
          7052 => x"527551fe",
          7053 => x"f2983f81",
          7054 => x"cbd40854",
          7055 => x"79537552",
          7056 => x"81c1b451",
          7057 => x"ff8da03f",
          7058 => x"873d0d04",
          7059 => x"f53d0d7d",
          7060 => x"7f61028c",
          7061 => x"0580c705",
          7062 => x"33737315",
          7063 => x"665f5d5a",
          7064 => x"5a5c5c5c",
          7065 => x"785281c1",
          7066 => x"d851ff8c",
          7067 => x"fa3f81c1",
          7068 => x"e051ff87",
          7069 => x"8e3f8055",
          7070 => x"74772780",
          7071 => x"fc387990",
          7072 => x"2e893879",
          7073 => x"a02ea738",
          7074 => x"80c63974",
          7075 => x"16537278",
          7076 => x"278e3872",
          7077 => x"225281c1",
          7078 => x"e451ff8c",
          7079 => x"ca3f8939",
          7080 => x"81c1f051",
          7081 => x"ff86dc3f",
          7082 => x"82155580",
          7083 => x"c3397416",
          7084 => x"53727827",
          7085 => x"8e387208",
          7086 => x"5281c1d8",
          7087 => x"51ff8ca7",
          7088 => x"3f893981",
          7089 => x"c1ec51ff",
          7090 => x"86b93f84",
          7091 => x"1555a139",
          7092 => x"74165372",
          7093 => x"78278e38",
          7094 => x"72335281",
          7095 => x"c1f851ff",
          7096 => x"8c853f89",
          7097 => x"3981c280",
          7098 => x"51ff8697",
          7099 => x"3f811555",
          7100 => x"a051fefa",
          7101 => x"8d3fff80",
          7102 => x"3981c284",
          7103 => x"51ff8683",
          7104 => x"3f805574",
          7105 => x"7727aa38",
          7106 => x"74167033",
          7107 => x"79722652",
          7108 => x"55539f74",
          7109 => x"27903872",
          7110 => x"802e8b38",
          7111 => x"7380fe26",
          7112 => x"85387351",
          7113 => x"8339a051",
          7114 => x"fef9d73f",
          7115 => x"811555d3",
          7116 => x"3981c288",
          7117 => x"51ff85cb",
          7118 => x"3f761677",
          7119 => x"1a5a56fe",
          7120 => x"fd923f81",
          7121 => x"cbd40898",
          7122 => x"2b70982c",
          7123 => x"515574a0",
          7124 => x"2e098106",
          7125 => x"a538fefc",
          7126 => x"fb3f81cb",
          7127 => x"d408982b",
          7128 => x"70982c70",
          7129 => x"a0327030",
          7130 => x"7072079f",
          7131 => x"2a515656",
          7132 => x"5155749b",
          7133 => x"2e8c3872",
          7134 => x"dd38749b",
          7135 => x"2e098106",
          7136 => x"85388053",
          7137 => x"8c397a1c",
          7138 => x"53727626",
          7139 => x"fdd638ff",
          7140 => x"537281cb",
          7141 => x"d40c8d3d",
          7142 => x"0d04ec3d",
          7143 => x"0d660284",
          7144 => x"0580e305",
          7145 => x"33697230",
          7146 => x"70740780",
          7147 => x"257087ff",
          7148 => x"74270751",
          7149 => x"51585a5b",
          7150 => x"56935774",
          7151 => x"80fb3881",
          7152 => x"5375528c",
          7153 => x"3d705257",
          7154 => x"c0b93f81",
          7155 => x"cbd40856",
          7156 => x"81cbd408",
          7157 => x"b83881cb",
          7158 => x"d40887c0",
          7159 => x"98880c81",
          7160 => x"cbd40859",
          7161 => x"963dd405",
          7162 => x"54848053",
          7163 => x"77527651",
          7164 => x"c4f63f81",
          7165 => x"cbd40856",
          7166 => x"81cbd408",
          7167 => x"90387a55",
          7168 => x"74802e89",
          7169 => x"38741975",
          7170 => x"195959d8",
          7171 => x"39963dd8",
          7172 => x"0551cce0",
          7173 => x"3f753070",
          7174 => x"77078025",
          7175 => x"51557980",
          7176 => x"2e953874",
          7177 => x"802e9038",
          7178 => x"81c28c53",
          7179 => x"87c09888",
          7180 => x"08527851",
          7181 => x"fbd73f75",
          7182 => x"577681cb",
          7183 => x"d40c963d",
          7184 => x"0d04f93d",
          7185 => x"0d7b0284",
          7186 => x"05b30533",
          7187 => x"5758ff57",
          7188 => x"80537a52",
          7189 => x"7951fec2",
          7190 => x"3f81cbd4",
          7191 => x"08a43875",
          7192 => x"802e8838",
          7193 => x"75812e98",
          7194 => x"38983960",
          7195 => x"557f5481",
          7196 => x"cbd4537e",
          7197 => x"527d5177",
          7198 => x"2d81cbd4",
          7199 => x"08578339",
          7200 => x"77047681",
          7201 => x"cbd40c89",
          7202 => x"3d0d04fc",
          7203 => x"3d0d029b",
          7204 => x"053381c2",
          7205 => x"945381c2",
          7206 => x"9c5255ff",
          7207 => x"88c93f81",
          7208 => x"c8e42251",
          7209 => x"ff80e23f",
          7210 => x"81c2a854",
          7211 => x"81c2b453",
          7212 => x"81c8e533",
          7213 => x"5281c2bc",
          7214 => x"51ff88ab",
          7215 => x"3f74802e",
          7216 => x"8538fefe",
          7217 => x"923f863d",
          7218 => x"0d04fe3d",
          7219 => x"0d87c096",
          7220 => x"800853ff",
          7221 => x"80fd3f81",
          7222 => x"51fef68c",
          7223 => x"3f81c2d8",
          7224 => x"51fef884",
          7225 => x"3f8051fe",
          7226 => x"f5fe3f72",
          7227 => x"812a7081",
          7228 => x"06515271",
          7229 => x"802e9538",
          7230 => x"8151fef5",
          7231 => x"eb3f81c2",
          7232 => x"f451fef7",
          7233 => x"e33f8051",
          7234 => x"fef5dd3f",
          7235 => x"72822a70",
          7236 => x"81065152",
          7237 => x"71802e95",
          7238 => x"388151fe",
          7239 => x"f5ca3f81",
          7240 => x"c38851fe",
          7241 => x"f7c23f80",
          7242 => x"51fef5bc",
          7243 => x"3f72832a",
          7244 => x"70810651",
          7245 => x"5271802e",
          7246 => x"95388151",
          7247 => x"fef5a93f",
          7248 => x"81c39851",
          7249 => x"fef7a13f",
          7250 => x"8051fef5",
          7251 => x"9b3f7284",
          7252 => x"2a708106",
          7253 => x"51527180",
          7254 => x"2e953881",
          7255 => x"51fef588",
          7256 => x"3f81c3ac",
          7257 => x"51fef780",
          7258 => x"3f8051fe",
          7259 => x"f4fa3f72",
          7260 => x"852a7081",
          7261 => x"06515271",
          7262 => x"802e9538",
          7263 => x"8151fef4",
          7264 => x"e73f81c3",
          7265 => x"c051fef6",
          7266 => x"df3f8051",
          7267 => x"fef4d93f",
          7268 => x"72862a70",
          7269 => x"81065152",
          7270 => x"71802e95",
          7271 => x"388151fe",
          7272 => x"f4c63f81",
          7273 => x"c3d451fe",
          7274 => x"f6be3f80",
          7275 => x"51fef4b8",
          7276 => x"3f72872a",
          7277 => x"70810651",
          7278 => x"5271802e",
          7279 => x"95388151",
          7280 => x"fef4a53f",
          7281 => x"81c3e851",
          7282 => x"fef69d3f",
          7283 => x"8051fef4",
          7284 => x"973f7288",
          7285 => x"2a708106",
          7286 => x"51527180",
          7287 => x"2e953881",
          7288 => x"51fef484",
          7289 => x"3f81c3fc",
          7290 => x"51fef5fc",
          7291 => x"3f8051fe",
          7292 => x"f3f63ffe",
          7293 => x"ffa63f84",
          7294 => x"3d0d04fa",
          7295 => x"3d0d7870",
          7296 => x"08705555",
          7297 => x"5773802e",
          7298 => x"80f0388e",
          7299 => x"3973770c",
          7300 => x"85153353",
          7301 => x"80e43981",
          7302 => x"14548074",
          7303 => x"337081ff",
          7304 => x"06575753",
          7305 => x"74a02e83",
          7306 => x"38815374",
          7307 => x"802e8438",
          7308 => x"72e53875",
          7309 => x"81ff0653",
          7310 => x"72a02e09",
          7311 => x"81068838",
          7312 => x"80747081",
          7313 => x"05563480",
          7314 => x"56759029",
          7315 => x"81c98405",
          7316 => x"77085370",
          7317 => x"085255fe",
          7318 => x"edfd3f81",
          7319 => x"cbd4088b",
          7320 => x"38841533",
          7321 => x"5372812e",
          7322 => x"ffa33881",
          7323 => x"167081ff",
          7324 => x"06575394",
          7325 => x"7627d238",
          7326 => x"ff537281",
          7327 => x"cbd40c88",
          7328 => x"3d0d04cb",
          7329 => x"3d0d8070",
          7330 => x"7181e2d4",
          7331 => x"0c5e5c81",
          7332 => x"527b51ff",
          7333 => x"8ac83f81",
          7334 => x"cbd40881",
          7335 => x"ff065978",
          7336 => x"7c2e0981",
          7337 => x"06a23881",
          7338 => x"c4bc5299",
          7339 => x"3d705259",
          7340 => x"ff84ca3f",
          7341 => x"7b537852",
          7342 => x"81cd8451",
          7343 => x"ffb9e33f",
          7344 => x"81cbd408",
          7345 => x"7c2e8838",
          7346 => x"81c4c051",
          7347 => x"8ee83981",
          7348 => x"705e5c81",
          7349 => x"c4f851fe",
          7350 => x"fea93f99",
          7351 => x"3d70465a",
          7352 => x"80f85380",
          7353 => x"527951fe",
          7354 => x"ebdc3f80",
          7355 => x"f8526451",
          7356 => x"ff84ce3f",
          7357 => x"b73dfef8",
          7358 => x"0551fdff",
          7359 => x"3f81cbd4",
          7360 => x"08902b70",
          7361 => x"902c5159",
          7362 => x"7880c32e",
          7363 => x"8a9b3878",
          7364 => x"80c32480",
          7365 => x"dc3878ab",
          7366 => x"2e83bc38",
          7367 => x"78ab24a4",
          7368 => x"3878822e",
          7369 => x"81af3878",
          7370 => x"82248a38",
          7371 => x"78802eff",
          7372 => x"a2388d88",
          7373 => x"3978842e",
          7374 => x"82823878",
          7375 => x"942e82ad",
          7376 => x"388cf939",
          7377 => x"7880c02e",
          7378 => x"858a3878",
          7379 => x"80c02490",
          7380 => x"3878b02e",
          7381 => x"83a93878",
          7382 => x"bc2e848b",
          7383 => x"388cdd39",
          7384 => x"7880c12e",
          7385 => x"86eb3878",
          7386 => x"80c22e88",
          7387 => x"8c388ccc",
          7388 => x"397880f8",
          7389 => x"2e8bba38",
          7390 => x"7880f824",
          7391 => x"a9387880",
          7392 => x"d12e8ae2",
          7393 => x"387880d1",
          7394 => x"248b3878",
          7395 => x"80d02e8a",
          7396 => x"c4388ca8",
          7397 => x"397880d4",
          7398 => x"2e8adc38",
          7399 => x"7880d52e",
          7400 => x"8af2388c",
          7401 => x"97397881",
          7402 => x"832e8bfc",
          7403 => x"38788183",
          7404 => x"24923878",
          7405 => x"80f92e8b",
          7406 => x"9d387881",
          7407 => x"822e8bd9",
          7408 => x"388bf939",
          7409 => x"7881852e",
          7410 => x"8beb3878",
          7411 => x"81872efe",
          7412 => x"82388be8",
          7413 => x"39b73dfe",
          7414 => x"f41153fe",
          7415 => x"f80551ff",
          7416 => x"83fa3f81",
          7417 => x"cbd40888",
          7418 => x"3881c4fc",
          7419 => x"518cc739",
          7420 => x"b73dfef0",
          7421 => x"1153fef8",
          7422 => x"0551ff83",
          7423 => x"df3f81cb",
          7424 => x"d408802e",
          7425 => x"88388163",
          7426 => x"25833880",
          7427 => x"430280cb",
          7428 => x"05335202",
          7429 => x"80cf0533",
          7430 => x"51ff87c2",
          7431 => x"3f81cbd4",
          7432 => x"0881ff06",
          7433 => x"59788e38",
          7434 => x"81c58c51",
          7435 => x"fefbd43f",
          7436 => x"815dfd9f",
          7437 => x"3981c59c",
          7438 => x"5189d239",
          7439 => x"b73dfef4",
          7440 => x"1153fef8",
          7441 => x"0551ff83",
          7442 => x"933f81cb",
          7443 => x"d408802e",
          7444 => x"fd813880",
          7445 => x"53805202",
          7446 => x"80cf0533",
          7447 => x"51ff8bcb",
          7448 => x"3f81cbd4",
          7449 => x"085281c5",
          7450 => x"b4518aa6",
          7451 => x"39b73dfe",
          7452 => x"f41153fe",
          7453 => x"f80551ff",
          7454 => x"82e23f81",
          7455 => x"cbd40880",
          7456 => x"2e873863",
          7457 => x"8926fccb",
          7458 => x"38b73dfe",
          7459 => x"f01153fe",
          7460 => x"f80551ff",
          7461 => x"82c63f81",
          7462 => x"cbd40886",
          7463 => x"3881cbd4",
          7464 => x"08436353",
          7465 => x"81c5bc52",
          7466 => x"7951ff80",
          7467 => x"d03f0280",
          7468 => x"cb053353",
          7469 => x"79526384",
          7470 => x"b42981cd",
          7471 => x"840551ff",
          7472 => x"b5e03f81",
          7473 => x"cbd40881",
          7474 => x"933881c5",
          7475 => x"8c51fefa",
          7476 => x"b23f815c",
          7477 => x"fbfd39b7",
          7478 => x"3dfef805",
          7479 => x"51feeab9",
          7480 => x"3f81cbd4",
          7481 => x"08b83dfe",
          7482 => x"f805525b",
          7483 => x"feeb8c3f",
          7484 => x"815381cb",
          7485 => x"d408527a",
          7486 => x"51f59f3f",
          7487 => x"80d539b7",
          7488 => x"3dfef805",
          7489 => x"51feea91",
          7490 => x"3f81cbd4",
          7491 => x"08b83dfe",
          7492 => x"f805525b",
          7493 => x"feeae43f",
          7494 => x"81cbd408",
          7495 => x"b83dfef8",
          7496 => x"05525afe",
          7497 => x"ead53f81",
          7498 => x"cbd408b8",
          7499 => x"3dfef805",
          7500 => x"5259feea",
          7501 => x"c63f81c8",
          7502 => x"c05881cc",
          7503 => x"88578056",
          7504 => x"805581cb",
          7505 => x"d40881ff",
          7506 => x"06547853",
          7507 => x"79527a51",
          7508 => x"f5f03f81",
          7509 => x"cbd40880",
          7510 => x"2efaf838",
          7511 => x"81cbd408",
          7512 => x"51f0863f",
          7513 => x"faed39b7",
          7514 => x"3dfef411",
          7515 => x"53fef805",
          7516 => x"51ff80e8",
          7517 => x"3f81cbd4",
          7518 => x"08802efa",
          7519 => x"d638b73d",
          7520 => x"fef01153",
          7521 => x"fef80551",
          7522 => x"ff80d13f",
          7523 => x"81cbd408",
          7524 => x"802efabf",
          7525 => x"38b73dfe",
          7526 => x"ec1153fe",
          7527 => x"f80551ff",
          7528 => x"80ba3f81",
          7529 => x"cbd40886",
          7530 => x"3881cbd4",
          7531 => x"084281c5",
          7532 => x"c051fef8",
          7533 => x"ce3f6363",
          7534 => x"5c5a797b",
          7535 => x"278f3861",
          7536 => x"59787a70",
          7537 => x"84055c0c",
          7538 => x"7a7a26f5",
          7539 => x"3881c588",
          7540 => x"5186ba39",
          7541 => x"b73dfef4",
          7542 => x"1153fef8",
          7543 => x"0551feff",
          7544 => x"fb3f81cb",
          7545 => x"d40880c4",
          7546 => x"3881c8ed",
          7547 => x"33597880",
          7548 => x"2e883881",
          7549 => x"c8c00844",
          7550 => x"b33981c8",
          7551 => x"ee335978",
          7552 => x"802e8838",
          7553 => x"81c8c808",
          7554 => x"44a23981",
          7555 => x"c8ef3359",
          7556 => x"788b3881",
          7557 => x"c8f03359",
          7558 => x"78802e88",
          7559 => x"3881c8d0",
          7560 => x"08448939",
          7561 => x"81c8e008",
          7562 => x"fc800544",
          7563 => x"b73dfef0",
          7564 => x"1153fef8",
          7565 => x"0551feff",
          7566 => x"a33f81cb",
          7567 => x"d40880c3",
          7568 => x"3881c8ed",
          7569 => x"33597880",
          7570 => x"2e883881",
          7571 => x"c8c40843",
          7572 => x"b23981c8",
          7573 => x"ee335978",
          7574 => x"802e8838",
          7575 => x"81c8cc08",
          7576 => x"43a13981",
          7577 => x"c8ef3359",
          7578 => x"788b3881",
          7579 => x"c8f03359",
          7580 => x"78802e88",
          7581 => x"3881c8d4",
          7582 => x"08438839",
          7583 => x"81c8e008",
          7584 => x"880543b7",
          7585 => x"3dfeec11",
          7586 => x"53fef805",
          7587 => x"51fefecc",
          7588 => x"3f81cbd4",
          7589 => x"08802e9b",
          7590 => x"3880625b",
          7591 => x"5979882e",
          7592 => x"83388159",
          7593 => x"79902e8d",
          7594 => x"3878802e",
          7595 => x"883879a0",
          7596 => x"2e833888",
          7597 => x"4281c5cc",
          7598 => x"51fef6c7",
          7599 => x"3fa05563",
          7600 => x"54615362",
          7601 => x"526351ef",
          7602 => x"833f81c5",
          7603 => x"dc5184bd",
          7604 => x"39b73dfe",
          7605 => x"f41153fe",
          7606 => x"f80551fe",
          7607 => x"fdfe3f81",
          7608 => x"cbd40880",
          7609 => x"2ef7ec38",
          7610 => x"b73dfef0",
          7611 => x"1153fef8",
          7612 => x"0551fefd",
          7613 => x"e73f81cb",
          7614 => x"d408802e",
          7615 => x"a5386359",
          7616 => x"0280cb05",
          7617 => x"33793463",
          7618 => x"810544b7",
          7619 => x"3dfef011",
          7620 => x"53fef805",
          7621 => x"51fefdc4",
          7622 => x"3f81cbd4",
          7623 => x"08e038f7",
          7624 => x"b2396370",
          7625 => x"33545281",
          7626 => x"c5e851fe",
          7627 => x"fbb93f80",
          7628 => x"f8527951",
          7629 => x"fefc8a3f",
          7630 => x"79457933",
          7631 => x"5978ae2e",
          7632 => x"f791389f",
          7633 => x"7927a038",
          7634 => x"b73dfef0",
          7635 => x"1153fef8",
          7636 => x"0551fefd",
          7637 => x"873f81cb",
          7638 => x"d408802e",
          7639 => x"91386359",
          7640 => x"0280cb05",
          7641 => x"33793463",
          7642 => x"810544ff",
          7643 => x"b53981c5",
          7644 => x"f451fef5",
          7645 => x"8e3fffaa",
          7646 => x"39b73dfe",
          7647 => x"e81153fe",
          7648 => x"f80551fe",
          7649 => x"fec83f81",
          7650 => x"cbd40880",
          7651 => x"2ef6c438",
          7652 => x"b73dfee4",
          7653 => x"1153fef8",
          7654 => x"0551fefe",
          7655 => x"b13f81cb",
          7656 => x"d408802e",
          7657 => x"a6386059",
          7658 => x"02be0522",
          7659 => x"79708205",
          7660 => x"5b237841",
          7661 => x"b73dfee4",
          7662 => x"1153fef8",
          7663 => x"0551fefe",
          7664 => x"8d3f81cb",
          7665 => x"d408df38",
          7666 => x"f6893960",
          7667 => x"70225452",
          7668 => x"81c5fc51",
          7669 => x"fefa903f",
          7670 => x"80f85279",
          7671 => x"51fefae1",
          7672 => x"3f794579",
          7673 => x"335978ae",
          7674 => x"2ef5e838",
          7675 => x"789f2687",
          7676 => x"38608405",
          7677 => x"41d539b7",
          7678 => x"3dfee411",
          7679 => x"53fef805",
          7680 => x"51fefdca",
          7681 => x"3f81cbd4",
          7682 => x"08802e92",
          7683 => x"38605902",
          7684 => x"be052279",
          7685 => x"7082055b",
          7686 => x"237841ff",
          7687 => x"ae3981c5",
          7688 => x"f451fef3",
          7689 => x"de3fffa3",
          7690 => x"39b73dfe",
          7691 => x"e81153fe",
          7692 => x"f80551fe",
          7693 => x"fd983f81",
          7694 => x"cbd40880",
          7695 => x"2ef59438",
          7696 => x"b73dfee4",
          7697 => x"1153fef8",
          7698 => x"0551fefd",
          7699 => x"813f81cb",
          7700 => x"d408802e",
          7701 => x"a1386060",
          7702 => x"710c5960",
          7703 => x"840541b7",
          7704 => x"3dfee411",
          7705 => x"53fef805",
          7706 => x"51fefce2",
          7707 => x"3f81cbd4",
          7708 => x"08e438f4",
          7709 => x"de396070",
          7710 => x"08545281",
          7711 => x"c68851fe",
          7712 => x"f8e53f80",
          7713 => x"f8527951",
          7714 => x"fef9b63f",
          7715 => x"79457933",
          7716 => x"5978ae2e",
          7717 => x"f4bd389f",
          7718 => x"7927a838",
          7719 => x"b73dfee4",
          7720 => x"1153fef8",
          7721 => x"0551fefc",
          7722 => x"a53f81cb",
          7723 => x"d408802e",
          7724 => x"99387f53",
          7725 => x"605281c6",
          7726 => x"8851fef8",
          7727 => x"aa3f6060",
          7728 => x"710c5960",
          7729 => x"840541ff",
          7730 => x"ad3981c5",
          7731 => x"f451fef2",
          7732 => x"b23fffa2",
          7733 => x"3981c694",
          7734 => x"51fef2a7",
          7735 => x"3f8251fe",
          7736 => x"f1953ff3",
          7737 => x"ee3981c6",
          7738 => x"ac51fef2",
          7739 => x"963fa251",
          7740 => x"fef0e83f",
          7741 => x"f3dd3984",
          7742 => x"80810b87",
          7743 => x"c094840c",
          7744 => x"8480810b",
          7745 => x"87c09494",
          7746 => x"0c81c6c4",
          7747 => x"51fef1f3",
          7748 => x"3ff3c039",
          7749 => x"81c6d851",
          7750 => x"fef1e83f",
          7751 => x"8c80830b",
          7752 => x"87c09484",
          7753 => x"0c8c8083",
          7754 => x"0b87c094",
          7755 => x"940cf3a3",
          7756 => x"39b73dfe",
          7757 => x"f41153fe",
          7758 => x"f80551fe",
          7759 => x"f99e3f81",
          7760 => x"cbd40880",
          7761 => x"2ef38c38",
          7762 => x"635281c6",
          7763 => x"ec51fef7",
          7764 => x"963f6359",
          7765 => x"7804b73d",
          7766 => x"fef41153",
          7767 => x"fef80551",
          7768 => x"fef8f93f",
          7769 => x"81cbd408",
          7770 => x"802ef2e7",
          7771 => x"38635281",
          7772 => x"c78851fe",
          7773 => x"f6f13f63",
          7774 => x"59782d81",
          7775 => x"cbd4085e",
          7776 => x"81cbd408",
          7777 => x"802ef2cb",
          7778 => x"3881cbd4",
          7779 => x"085281c7",
          7780 => x"a451fef6",
          7781 => x"d23ff2bb",
          7782 => x"3981c7c0",
          7783 => x"51fef0e3",
          7784 => x"3ffeccdc",
          7785 => x"3ff2ac39",
          7786 => x"81c7dc51",
          7787 => x"fef0d43f",
          7788 => x"8059ffa0",
          7789 => x"39feec9f",
          7790 => x"3ff29839",
          7791 => x"64703351",
          7792 => x"5978802e",
          7793 => x"f28d387b",
          7794 => x"802e80d2",
          7795 => x"387c802e",
          7796 => x"80cc38b7",
          7797 => x"3dfef805",
          7798 => x"51fee0bd",
          7799 => x"3f81c7f0",
          7800 => x"5681cbd4",
          7801 => x"085581c7",
          7802 => x"f4548053",
          7803 => x"81c7f852",
          7804 => x"a33d7052",
          7805 => x"5afef685",
          7806 => x"3f81c8c0",
          7807 => x"5881cc88",
          7808 => x"57805664",
          7809 => x"81114681",
          7810 => x"05558054",
          7811 => x"81800a53",
          7812 => x"81800a52",
          7813 => x"7951ecaa",
          7814 => x"3f81cbd4",
          7815 => x"085e7c81",
          7816 => x"327c8132",
          7817 => x"0759788a",
          7818 => x"387dff2e",
          7819 => x"098106f1",
          7820 => x"a23881c8",
          7821 => x"8851fef5",
          7822 => x"ae3ff197",
          7823 => x"39803d0d",
          7824 => x"800b81cc",
          7825 => x"88349b90",
          7826 => x"86e40b87",
          7827 => x"c0948c0c",
          7828 => x"9b9086e4",
          7829 => x"0b87c094",
          7830 => x"9c0c8c80",
          7831 => x"830b87c0",
          7832 => x"94840c8c",
          7833 => x"80830b87",
          7834 => x"c094940c",
          7835 => x"98820b81",
          7836 => x"cbe40c9b",
          7837 => x"830b81cb",
          7838 => x"e80cfee7",
          7839 => x"af3ffeed",
          7840 => x"d23f81c8",
          7841 => x"9851fee4",
          7842 => x"df3f81c8",
          7843 => x"a451feee",
          7844 => x"f23f81a1",
          7845 => x"ca51feed",
          7846 => x"b53f8151",
          7847 => x"ebed3fef",
          7848 => x"e23f8004",
          7849 => x"00001125",
          7850 => x"0000112b",
          7851 => x"00001131",
          7852 => x"00001137",
          7853 => x"0000113d",
          7854 => x"00004dfb",
          7855 => x"00004d7f",
          7856 => x"00004d86",
          7857 => x"00004d8d",
          7858 => x"00004d94",
          7859 => x"00004d9b",
          7860 => x"00004da2",
          7861 => x"00004da9",
          7862 => x"00004db0",
          7863 => x"00004db7",
          7864 => x"00004dbe",
          7865 => x"00004dc5",
          7866 => x"00004dcb",
          7867 => x"00004dd1",
          7868 => x"00004dd7",
          7869 => x"00004ddd",
          7870 => x"00004de3",
          7871 => x"00004de9",
          7872 => x"00004def",
          7873 => x"00004df5",
          7874 => x"25642f25",
          7875 => x"642f2564",
          7876 => x"2025643a",
          7877 => x"25643a25",
          7878 => x"642e2564",
          7879 => x"25640a00",
          7880 => x"536f4320",
          7881 => x"436f6e66",
          7882 => x"69677572",
          7883 => x"6174696f",
          7884 => x"6e000000",
          7885 => x"20286672",
          7886 => x"6f6d2053",
          7887 => x"6f432063",
          7888 => x"6f6e6669",
          7889 => x"67290000",
          7890 => x"3a0a4465",
          7891 => x"76696365",
          7892 => x"7320696d",
          7893 => x"706c656d",
          7894 => x"656e7465",
          7895 => x"643a0a00",
          7896 => x"20202020",
          7897 => x"494e534e",
          7898 => x"20425241",
          7899 => x"4d202853",
          7900 => x"74617274",
          7901 => x"3d253038",
          7902 => x"582c2053",
          7903 => x"697a653d",
          7904 => x"25303858",
          7905 => x"292e0a00",
          7906 => x"20202020",
          7907 => x"4252414d",
          7908 => x"20285374",
          7909 => x"6172743d",
          7910 => x"25303858",
          7911 => x"2c205369",
          7912 => x"7a653d25",
          7913 => x"30385829",
          7914 => x"2e0a0000",
          7915 => x"20202020",
          7916 => x"52414d20",
          7917 => x"28537461",
          7918 => x"72743d25",
          7919 => x"3038582c",
          7920 => x"2053697a",
          7921 => x"653d2530",
          7922 => x"3858292e",
          7923 => x"0a000000",
          7924 => x"20202020",
          7925 => x"494f4354",
          7926 => x"4c0a0000",
          7927 => x"20202020",
          7928 => x"5053320a",
          7929 => x"00000000",
          7930 => x"20202020",
          7931 => x"5350490a",
          7932 => x"00000000",
          7933 => x"20202020",
          7934 => x"53442043",
          7935 => x"61726420",
          7936 => x"28446576",
          7937 => x"69636573",
          7938 => x"3d253032",
          7939 => x"58292e0a",
          7940 => x"00000000",
          7941 => x"20202020",
          7942 => x"494e5445",
          7943 => x"52525550",
          7944 => x"5420434f",
          7945 => x"4e54524f",
          7946 => x"4c4c4552",
          7947 => x"0a000000",
          7948 => x"20202020",
          7949 => x"54494d45",
          7950 => x"52312028",
          7951 => x"54696d65",
          7952 => x"72733d25",
          7953 => x"30315829",
          7954 => x"2e0a0000",
          7955 => x"41646472",
          7956 => x"65737365",
          7957 => x"733a0a00",
          7958 => x"20202020",
          7959 => x"43505520",
          7960 => x"52657365",
          7961 => x"74205665",
          7962 => x"63746f72",
          7963 => x"20416464",
          7964 => x"72657373",
          7965 => x"203d2025",
          7966 => x"3038580a",
          7967 => x"00000000",
          7968 => x"20202020",
          7969 => x"43505520",
          7970 => x"4d656d6f",
          7971 => x"72792053",
          7972 => x"74617274",
          7973 => x"20416464",
          7974 => x"72657373",
          7975 => x"203d2025",
          7976 => x"3038580a",
          7977 => x"00000000",
          7978 => x"20202020",
          7979 => x"53746163",
          7980 => x"6b205374",
          7981 => x"61727420",
          7982 => x"41646472",
          7983 => x"65737320",
          7984 => x"20202020",
          7985 => x"203d2025",
          7986 => x"3038580a",
          7987 => x"00000000",
          7988 => x"20202020",
          7989 => x"5a505520",
          7990 => x"49642020",
          7991 => x"20202020",
          7992 => x"20202020",
          7993 => x"20202020",
          7994 => x"20202020",
          7995 => x"203d2025",
          7996 => x"3038580a",
          7997 => x"00000000",
          7998 => x"20202020",
          7999 => x"53797374",
          8000 => x"656d2043",
          8001 => x"6c6f636b",
          8002 => x"20467265",
          8003 => x"71202020",
          8004 => x"20202020",
          8005 => x"203d2025",
          8006 => x"3038580a",
          8007 => x"00000000",
          8008 => x"536d616c",
          8009 => x"6c000000",
          8010 => x"4d656469",
          8011 => x"756d0000",
          8012 => x"466c6578",
          8013 => x"00000000",
          8014 => x"45564f00",
          8015 => x"45564f6d",
          8016 => x"696e0000",
          8017 => x"556e6b6e",
          8018 => x"6f776e00",
          8019 => x"53440000",
          8020 => x"222a2b2c",
          8021 => x"3a3b3c3d",
          8022 => x"3e3f5b5d",
          8023 => x"7c7f0000",
          8024 => x"46415400",
          8025 => x"46415433",
          8026 => x"32000000",
          8027 => x"ebfe904d",
          8028 => x"53444f53",
          8029 => x"352e3000",
          8030 => x"4e4f204e",
          8031 => x"414d4520",
          8032 => x"20202046",
          8033 => x"41543332",
          8034 => x"20202000",
          8035 => x"4e4f204e",
          8036 => x"414d4520",
          8037 => x"20202046",
          8038 => x"41542020",
          8039 => x"20202000",
          8040 => x"00005d4c",
          8041 => x"00000000",
          8042 => x"00000000",
          8043 => x"00000000",
          8044 => x"809a4541",
          8045 => x"8e418f80",
          8046 => x"45454549",
          8047 => x"49498e8f",
          8048 => x"9092924f",
          8049 => x"994f5555",
          8050 => x"59999a9b",
          8051 => x"9c9d9e9f",
          8052 => x"41494f55",
          8053 => x"a5a5a6a7",
          8054 => x"a8a9aaab",
          8055 => x"acadaeaf",
          8056 => x"b0b1b2b3",
          8057 => x"b4b5b6b7",
          8058 => x"b8b9babb",
          8059 => x"bcbdbebf",
          8060 => x"c0c1c2c3",
          8061 => x"c4c5c6c7",
          8062 => x"c8c9cacb",
          8063 => x"cccdcecf",
          8064 => x"d0d1d2d3",
          8065 => x"d4d5d6d7",
          8066 => x"d8d9dadb",
          8067 => x"dcdddedf",
          8068 => x"e0e1e2e3",
          8069 => x"e4e5e6e7",
          8070 => x"e8e9eaeb",
          8071 => x"ecedeeef",
          8072 => x"f0f1f2f3",
          8073 => x"f4f5f6f7",
          8074 => x"f8f9fafb",
          8075 => x"fcfdfeff",
          8076 => x"2b2e2c3b",
          8077 => x"3d5b5d2f",
          8078 => x"5c222a3a",
          8079 => x"3c3e3f7c",
          8080 => x"7f000000",
          8081 => x"00010004",
          8082 => x"00100040",
          8083 => x"01000200",
          8084 => x"00000000",
          8085 => x"00010002",
          8086 => x"00040008",
          8087 => x"00100020",
          8088 => x"00000000",
          8089 => x"64696e69",
          8090 => x"74000000",
          8091 => x"64696f63",
          8092 => x"746c0000",
          8093 => x"66696e69",
          8094 => x"74000000",
          8095 => x"666c6f61",
          8096 => x"64000000",
          8097 => x"66657865",
          8098 => x"63000000",
          8099 => x"6d636c65",
          8100 => x"61720000",
          8101 => x"6d64756d",
          8102 => x"70000000",
          8103 => x"6d746573",
          8104 => x"74000000",
          8105 => x"6d656200",
          8106 => x"6d656800",
          8107 => x"6d657700",
          8108 => x"68696400",
          8109 => x"68696500",
          8110 => x"68666400",
          8111 => x"68666500",
          8112 => x"63616c6c",
          8113 => x"00000000",
          8114 => x"6a6d7000",
          8115 => x"72657374",
          8116 => x"61727400",
          8117 => x"72657365",
          8118 => x"74000000",
          8119 => x"696e666f",
          8120 => x"00000000",
          8121 => x"74657374",
          8122 => x"00000000",
          8123 => x"4469736b",
          8124 => x"20457272",
          8125 => x"6f720a00",
          8126 => x"496e7465",
          8127 => x"726e616c",
          8128 => x"20657272",
          8129 => x"6f722e0a",
          8130 => x"00000000",
          8131 => x"4469736b",
          8132 => x"206e6f74",
          8133 => x"20726561",
          8134 => x"64792e0a",
          8135 => x"00000000",
          8136 => x"4e6f2066",
          8137 => x"696c6520",
          8138 => x"666f756e",
          8139 => x"642e0a00",
          8140 => x"4e6f2070",
          8141 => x"61746820",
          8142 => x"666f756e",
          8143 => x"642e0a00",
          8144 => x"496e7661",
          8145 => x"6c696420",
          8146 => x"66696c65",
          8147 => x"6e616d65",
          8148 => x"2e0a0000",
          8149 => x"41636365",
          8150 => x"73732064",
          8151 => x"656e6965",
          8152 => x"642e0a00",
          8153 => x"46696c65",
          8154 => x"20616c72",
          8155 => x"65616479",
          8156 => x"20657869",
          8157 => x"7374732e",
          8158 => x"0a000000",
          8159 => x"46696c65",
          8160 => x"2068616e",
          8161 => x"646c6520",
          8162 => x"696e7661",
          8163 => x"6c69642e",
          8164 => x"0a000000",
          8165 => x"53442069",
          8166 => x"73207772",
          8167 => x"69746520",
          8168 => x"70726f74",
          8169 => x"65637465",
          8170 => x"642e0a00",
          8171 => x"44726976",
          8172 => x"65206e75",
          8173 => x"6d626572",
          8174 => x"20697320",
          8175 => x"696e7661",
          8176 => x"6c69642e",
          8177 => x"0a000000",
          8178 => x"4469736b",
          8179 => x"206e6f74",
          8180 => x"20656e61",
          8181 => x"626c6564",
          8182 => x"2e0a0000",
          8183 => x"4e6f2063",
          8184 => x"6f6d7061",
          8185 => x"7469626c",
          8186 => x"65206669",
          8187 => x"6c657379",
          8188 => x"7374656d",
          8189 => x"20666f75",
          8190 => x"6e64206f",
          8191 => x"6e206469",
          8192 => x"736b2e0a",
          8193 => x"00000000",
          8194 => x"466f726d",
          8195 => x"61742061",
          8196 => x"626f7274",
          8197 => x"65642e0a",
          8198 => x"00000000",
          8199 => x"54696d65",
          8200 => x"6f75742c",
          8201 => x"206f7065",
          8202 => x"72617469",
          8203 => x"6f6e2063",
          8204 => x"616e6365",
          8205 => x"6c6c6564",
          8206 => x"2e0a0000",
          8207 => x"46696c65",
          8208 => x"20697320",
          8209 => x"6c6f636b",
          8210 => x"65642e0a",
          8211 => x"00000000",
          8212 => x"496e7375",
          8213 => x"66666963",
          8214 => x"69656e74",
          8215 => x"206d656d",
          8216 => x"6f72792e",
          8217 => x"0a000000",
          8218 => x"546f6f20",
          8219 => x"6d616e79",
          8220 => x"206f7065",
          8221 => x"6e206669",
          8222 => x"6c65732e",
          8223 => x"0a000000",
          8224 => x"50617261",
          8225 => x"6d657465",
          8226 => x"72732069",
          8227 => x"6e636f72",
          8228 => x"72656374",
          8229 => x"2e0a0000",
          8230 => x"53756363",
          8231 => x"6573732e",
          8232 => x"0a000000",
          8233 => x"556e6b6e",
          8234 => x"6f776e20",
          8235 => x"6572726f",
          8236 => x"722e0a00",
          8237 => x"0a256c75",
          8238 => x"20627974",
          8239 => x"65732025",
          8240 => x"73206174",
          8241 => x"20256c75",
          8242 => x"20627974",
          8243 => x"65732f73",
          8244 => x"65632e0a",
          8245 => x"00000000",
          8246 => x"25303858",
          8247 => x"00000000",
          8248 => x"3a202000",
          8249 => x"25303458",
          8250 => x"00000000",
          8251 => x"20202020",
          8252 => x"20202020",
          8253 => x"00000000",
          8254 => x"25303258",
          8255 => x"00000000",
          8256 => x"20200000",
          8257 => x"207c0000",
          8258 => x"7c0d0a00",
          8259 => x"72656164",
          8260 => x"00000000",
          8261 => x"5a505554",
          8262 => x"41000000",
          8263 => x"0a2a2a20",
          8264 => x"25732028",
          8265 => x"00000000",
          8266 => x"31382f30",
          8267 => x"372f3230",
          8268 => x"31390000",
          8269 => x"76312e33",
          8270 => x"00000000",
          8271 => x"205a5055",
          8272 => x"2c207265",
          8273 => x"76202530",
          8274 => x"32782920",
          8275 => x"25732025",
          8276 => x"73202a2a",
          8277 => x"0a0a0000",
          8278 => x"5a505554",
          8279 => x"4120496e",
          8280 => x"74657272",
          8281 => x"75707420",
          8282 => x"48616e64",
          8283 => x"6c65720a",
          8284 => x"00000000",
          8285 => x"54696d65",
          8286 => x"7220696e",
          8287 => x"74657272",
          8288 => x"7570740a",
          8289 => x"00000000",
          8290 => x"50533220",
          8291 => x"696e7465",
          8292 => x"72727570",
          8293 => x"740a0000",
          8294 => x"494f4354",
          8295 => x"4c205244",
          8296 => x"20696e74",
          8297 => x"65727275",
          8298 => x"70740a00",
          8299 => x"494f4354",
          8300 => x"4c205752",
          8301 => x"20696e74",
          8302 => x"65727275",
          8303 => x"70740a00",
          8304 => x"55415254",
          8305 => x"30205258",
          8306 => x"20696e74",
          8307 => x"65727275",
          8308 => x"70740a00",
          8309 => x"55415254",
          8310 => x"30205458",
          8311 => x"20696e74",
          8312 => x"65727275",
          8313 => x"70740a00",
          8314 => x"55415254",
          8315 => x"31205258",
          8316 => x"20696e74",
          8317 => x"65727275",
          8318 => x"70740a00",
          8319 => x"55415254",
          8320 => x"31205458",
          8321 => x"20696e74",
          8322 => x"65727275",
          8323 => x"70740a00",
          8324 => x"53657474",
          8325 => x"696e6720",
          8326 => x"75702074",
          8327 => x"696d6572",
          8328 => x"2e2e2e0a",
          8329 => x"00000000",
          8330 => x"456e6162",
          8331 => x"6c696e67",
          8332 => x"2074696d",
          8333 => x"65722e2e",
          8334 => x"2e0a0000",
          8335 => x"303a0000",
          8336 => x"4661696c",
          8337 => x"65642074",
          8338 => x"6f20696e",
          8339 => x"69746961",
          8340 => x"6c697365",
          8341 => x"20736420",
          8342 => x"63617264",
          8343 => x"20302c20",
          8344 => x"706c6561",
          8345 => x"73652069",
          8346 => x"6e697420",
          8347 => x"6d616e75",
          8348 => x"616c6c79",
          8349 => x"2e0a0000",
          8350 => x"2a200000",
          8351 => x"42616420",
          8352 => x"6469736b",
          8353 => x"20696421",
          8354 => x"0a000000",
          8355 => x"496e6974",
          8356 => x"69616c69",
          8357 => x"7365642e",
          8358 => x"0a000000",
          8359 => x"4661696c",
          8360 => x"65642074",
          8361 => x"6f20696e",
          8362 => x"69746961",
          8363 => x"6c697365",
          8364 => x"2e0a0000",
          8365 => x"72633d25",
          8366 => x"640a0000",
          8367 => x"25753a00",
          8368 => x"436c6561",
          8369 => x"72696e67",
          8370 => x"2e2e2e00",
          8371 => x"44756d70",
          8372 => x"204d656d",
          8373 => x"6f72790a",
          8374 => x"00000000",
          8375 => x"0a436f6d",
          8376 => x"706c6574",
          8377 => x"652e0a00",
          8378 => x"25303858",
          8379 => x"20253032",
          8380 => x"582d0000",
          8381 => x"3f3f3f0a",
          8382 => x"00000000",
          8383 => x"25303858",
          8384 => x"20253034",
          8385 => x"582d0000",
          8386 => x"25303858",
          8387 => x"20253038",
          8388 => x"582d0000",
          8389 => x"44697361",
          8390 => x"626c696e",
          8391 => x"6720696e",
          8392 => x"74657272",
          8393 => x"75707473",
          8394 => x"0a000000",
          8395 => x"456e6162",
          8396 => x"6c696e67",
          8397 => x"20696e74",
          8398 => x"65727275",
          8399 => x"7074730a",
          8400 => x"00000000",
          8401 => x"44697361",
          8402 => x"626c6564",
          8403 => x"20756172",
          8404 => x"74206669",
          8405 => x"666f0a00",
          8406 => x"456e6162",
          8407 => x"6c696e67",
          8408 => x"20756172",
          8409 => x"74206669",
          8410 => x"666f0a00",
          8411 => x"45786563",
          8412 => x"7574696e",
          8413 => x"6720636f",
          8414 => x"64652040",
          8415 => x"20253038",
          8416 => x"78202e2e",
          8417 => x"2e0a0000",
          8418 => x"43616c6c",
          8419 => x"696e6720",
          8420 => x"636f6465",
          8421 => x"20402025",
          8422 => x"30387820",
          8423 => x"2e2e2e0a",
          8424 => x"00000000",
          8425 => x"43616c6c",
          8426 => x"20726574",
          8427 => x"75726e65",
          8428 => x"6420636f",
          8429 => x"64652028",
          8430 => x"2564292e",
          8431 => x"0a000000",
          8432 => x"52657374",
          8433 => x"61727469",
          8434 => x"6e672061",
          8435 => x"70706c69",
          8436 => x"63617469",
          8437 => x"6f6e2e2e",
          8438 => x"2e0a0000",
          8439 => x"436f6c64",
          8440 => x"20726562",
          8441 => x"6f6f7469",
          8442 => x"6e672e2e",
          8443 => x"2e0a0000",
          8444 => x"5a505500",
          8445 => x"62696e00",
          8446 => x"25643a5c",
          8447 => x"25735c25",
          8448 => x"732e2573",
          8449 => x"00000000",
          8450 => x"42616420",
          8451 => x"636f6d6d",
          8452 => x"616e642e",
          8453 => x"0a000000",
          8454 => x"52756e6e",
          8455 => x"696e672e",
          8456 => x"2e2e0a00",
          8457 => x"456e6162",
          8458 => x"6c696e67",
          8459 => x"20696e74",
          8460 => x"65727275",
          8461 => x"7074732e",
          8462 => x"2e2e0a00",
          8463 => x"00000000",
          8464 => x"00000000",
          8465 => x"00007fff",
          8466 => x"00000000",
          8467 => x"00007fff",
          8468 => x"00010000",
          8469 => x"00007fff",
          8470 => x"00000000",
          8471 => x"00000000",
          8472 => x"00007800",
          8473 => x"00000000",
          8474 => x"05f5e100",
          8475 => x"00010101",
          8476 => x"01010101",
          8477 => x"80010101",
          8478 => x"01000000",
          8479 => x"00000000",
          8480 => x"01000000",
          8481 => x"00005e64",
          8482 => x"01020100",
          8483 => x"00000000",
          8484 => x"00000000",
          8485 => x"00005e6c",
          8486 => x"01040100",
          8487 => x"00000000",
          8488 => x"00000000",
          8489 => x"00005e74",
          8490 => x"01140300",
          8491 => x"00000000",
          8492 => x"00000000",
          8493 => x"00005e7c",
          8494 => x"012b0300",
          8495 => x"00000000",
          8496 => x"00000000",
          8497 => x"00005e84",
          8498 => x"01300300",
          8499 => x"00000000",
          8500 => x"00000000",
          8501 => x"00005e8c",
          8502 => x"013c0400",
          8503 => x"00000000",
          8504 => x"00000000",
          8505 => x"00005e94",
          8506 => x"01400400",
          8507 => x"00000000",
          8508 => x"00000000",
          8509 => x"00005e9c",
          8510 => x"01440400",
          8511 => x"00000000",
          8512 => x"00000000",
          8513 => x"00005ea4",
          8514 => x"01410400",
          8515 => x"00000000",
          8516 => x"00000000",
          8517 => x"00005ea8",
          8518 => x"01420400",
          8519 => x"00000000",
          8520 => x"00000000",
          8521 => x"00005eac",
          8522 => x"01430400",
          8523 => x"00000000",
          8524 => x"00000000",
          8525 => x"00005eb0",
          8526 => x"01500500",
          8527 => x"00000000",
          8528 => x"00000000",
          8529 => x"00005eb4",
          8530 => x"01510500",
          8531 => x"00000000",
          8532 => x"00000000",
          8533 => x"00005eb8",
          8534 => x"01540500",
          8535 => x"00000000",
          8536 => x"00000000",
          8537 => x"00005ebc",
          8538 => x"01550500",
          8539 => x"00000000",
          8540 => x"00000000",
          8541 => x"00005ec0",
          8542 => x"01790700",
          8543 => x"00000000",
          8544 => x"00000000",
          8545 => x"00005ec8",
          8546 => x"01780700",
          8547 => x"00000000",
          8548 => x"00000000",
          8549 => x"00005ecc",
          8550 => x"01820800",
          8551 => x"00000000",
          8552 => x"00000000",
          8553 => x"00005ed4",
          8554 => x"01830800",
          8555 => x"00000000",
          8556 => x"00000000",
          8557 => x"00005edc",
          8558 => x"01850800",
          8559 => x"00000000",
          8560 => x"00000000",
          8561 => x"00005ee4",
          8562 => x"01870800",
          8563 => x"00000000",
          8564 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;


end arch;

