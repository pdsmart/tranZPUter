-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e9040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"88738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cb2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8a",
           179 => x"fd2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"80040088",
           281 => x"e2040000",
           282 => x"009fac70",
           283 => x"9fdc278b",
           284 => x"38807170",
           285 => x"8405530c",
           286 => x"88eb0488",
           287 => x"e2519e99",
           288 => x"04940802",
           289 => x"940cfd3d",
           290 => x"0d805394",
           291 => x"088c0508",
           292 => x"52940888",
           293 => x"05085182",
           294 => x"de3f8808",
           295 => x"70880c54",
           296 => x"853d0d94",
           297 => x"0c049408",
           298 => x"02940cfd",
           299 => x"3d0d8153",
           300 => x"94088c05",
           301 => x"08529408",
           302 => x"88050851",
           303 => x"82b93f88",
           304 => x"0870880c",
           305 => x"54853d0d",
           306 => x"940c0494",
           307 => x"0802940c",
           308 => x"f93d0d80",
           309 => x"0b9408fc",
           310 => x"050c9408",
           311 => x"88050880",
           312 => x"25ab3894",
           313 => x"08880508",
           314 => x"30940888",
           315 => x"050c800b",
           316 => x"9408f405",
           317 => x"0c9408fc",
           318 => x"05088838",
           319 => x"810b9408",
           320 => x"f4050c94",
           321 => x"08f40508",
           322 => x"9408fc05",
           323 => x"0c94088c",
           324 => x"05088025",
           325 => x"ab389408",
           326 => x"8c050830",
           327 => x"94088c05",
           328 => x"0c800b94",
           329 => x"08f0050c",
           330 => x"9408fc05",
           331 => x"08883881",
           332 => x"0b9408f0",
           333 => x"050c9408",
           334 => x"f0050894",
           335 => x"08fc050c",
           336 => x"80539408",
           337 => x"8c050852",
           338 => x"94088805",
           339 => x"085181a7",
           340 => x"3f880870",
           341 => x"9408f805",
           342 => x"0c549408",
           343 => x"fc050880",
           344 => x"2e8c3894",
           345 => x"08f80508",
           346 => x"309408f8",
           347 => x"050c9408",
           348 => x"f8050870",
           349 => x"880c5489",
           350 => x"3d0d940c",
           351 => x"04940802",
           352 => x"940cfb3d",
           353 => x"0d800b94",
           354 => x"08fc050c",
           355 => x"94088805",
           356 => x"08802593",
           357 => x"38940888",
           358 => x"05083094",
           359 => x"0888050c",
           360 => x"810b9408",
           361 => x"fc050c94",
           362 => x"088c0508",
           363 => x"80258c38",
           364 => x"94088c05",
           365 => x"08309408",
           366 => x"8c050c81",
           367 => x"5394088c",
           368 => x"05085294",
           369 => x"08880508",
           370 => x"51ad3f88",
           371 => x"08709408",
           372 => x"f8050c54",
           373 => x"9408fc05",
           374 => x"08802e8c",
           375 => x"389408f8",
           376 => x"05083094",
           377 => x"08f8050c",
           378 => x"9408f805",
           379 => x"0870880c",
           380 => x"54873d0d",
           381 => x"940c0494",
           382 => x"0802940c",
           383 => x"fd3d0d81",
           384 => x"0b9408fc",
           385 => x"050c800b",
           386 => x"9408f805",
           387 => x"0c94088c",
           388 => x"05089408",
           389 => x"88050827",
           390 => x"ac389408",
           391 => x"fc050880",
           392 => x"2ea33880",
           393 => x"0b94088c",
           394 => x"05082499",
           395 => x"3894088c",
           396 => x"05081094",
           397 => x"088c050c",
           398 => x"9408fc05",
           399 => x"08109408",
           400 => x"fc050cc9",
           401 => x"399408fc",
           402 => x"0508802e",
           403 => x"80c93894",
           404 => x"088c0508",
           405 => x"94088805",
           406 => x"0826a138",
           407 => x"94088805",
           408 => x"0894088c",
           409 => x"05083194",
           410 => x"0888050c",
           411 => x"9408f805",
           412 => x"089408fc",
           413 => x"05080794",
           414 => x"08f8050c",
           415 => x"9408fc05",
           416 => x"08812a94",
           417 => x"08fc050c",
           418 => x"94088c05",
           419 => x"08812a94",
           420 => x"088c050c",
           421 => x"ffaf3994",
           422 => x"08900508",
           423 => x"802e8f38",
           424 => x"94088805",
           425 => x"08709408",
           426 => x"f4050c51",
           427 => x"8d399408",
           428 => x"f8050870",
           429 => x"9408f405",
           430 => x"0c519408",
           431 => x"f4050888",
           432 => x"0c853d0d",
           433 => x"940c04ff",
           434 => x"3d0d8188",
           435 => x"0b87c092",
           436 => x"8c0c810b",
           437 => x"87c0928c",
           438 => x"0c850b87",
           439 => x"c0988c0c",
           440 => x"87c0928c",
           441 => x"08708206",
           442 => x"51517080",
           443 => x"2e8a3887",
           444 => x"c0988c08",
           445 => x"5170e938",
           446 => x"87c0928c",
           447 => x"08fc8080",
           448 => x"06527193",
           449 => x"3887c098",
           450 => x"8c085170",
           451 => x"802e8838",
           452 => x"710b0b0b",
           453 => x"9fa8340b",
           454 => x"0b0b9fa8",
           455 => x"33880c83",
           456 => x"3d0d04fa",
           457 => x"3d0d787b",
           458 => x"7d565856",
           459 => x"800b0b0b",
           460 => x"0b9fa833",
           461 => x"81065255",
           462 => x"82527075",
           463 => x"2e098106",
           464 => x"819e3885",
           465 => x"0b87c098",
           466 => x"8c0c7987",
           467 => x"c092800c",
           468 => x"840b87c0",
           469 => x"928c0c87",
           470 => x"c0928c08",
           471 => x"70852a70",
           472 => x"81065152",
           473 => x"5370802e",
           474 => x"a73887c0",
           475 => x"92840870",
           476 => x"81ff0676",
           477 => x"79275253",
           478 => x"5173802e",
           479 => x"90387080",
           480 => x"2e8b3871",
           481 => x"76708105",
           482 => x"5834ff14",
           483 => x"54811555",
           484 => x"72a20651",
           485 => x"70802e8b",
           486 => x"3887c098",
           487 => x"8c085170",
           488 => x"ffb53887",
           489 => x"c0988c08",
           490 => x"51709538",
           491 => x"810b87c0",
           492 => x"928c0c87",
           493 => x"c0928c08",
           494 => x"70820651",
           495 => x"5170f438",
           496 => x"8073fc80",
           497 => x"80065252",
           498 => x"70722e09",
           499 => x"81068f38",
           500 => x"87c0988c",
           501 => x"08517072",
           502 => x"2e098106",
           503 => x"83388152",
           504 => x"71880c88",
           505 => x"3d0d04fe",
           506 => x"3d0d7481",
           507 => x"11337133",
           508 => x"71882b07",
           509 => x"880c5351",
           510 => x"843d0d04",
           511 => x"fd3d0d75",
           512 => x"83113382",
           513 => x"12337190",
           514 => x"2b71882b",
           515 => x"07811433",
           516 => x"70720788",
           517 => x"2b753371",
           518 => x"07880c52",
           519 => x"53545654",
           520 => x"52853d0d",
           521 => x"04f93d0d",
           522 => x"790b0b0b",
           523 => x"9fac0857",
           524 => x"57817727",
           525 => x"80ed3876",
           526 => x"88170827",
           527 => x"80e53875",
           528 => x"33557482",
           529 => x"2e893874",
           530 => x"832eae38",
           531 => x"80d53974",
           532 => x"54761083",
           533 => x"fe065376",
           534 => x"882a8c17",
           535 => x"08055288",
           536 => x"3d705255",
           537 => x"fdbd3f88",
           538 => x"08b93874",
           539 => x"51fef83f",
           540 => x"880883ff",
           541 => x"ff0655ad",
           542 => x"39845476",
           543 => x"822b83fc",
           544 => x"06537687",
           545 => x"2a8c1708",
           546 => x"0552883d",
           547 => x"705255fd",
           548 => x"923f8808",
           549 => x"8e387451",
           550 => x"fee23f88",
           551 => x"08f00a06",
           552 => x"55833981",
           553 => x"5574880c",
           554 => x"893d0d04",
           555 => x"fb3d0d0b",
           556 => x"0b0b9fac",
           557 => x"08fe1988",
           558 => x"1208fe05",
           559 => x"55565480",
           560 => x"56747327",
           561 => x"8d388214",
           562 => x"33757129",
           563 => x"94160805",
           564 => x"57537588",
           565 => x"0c873d0d",
           566 => x"04fd3d0d",
           567 => x"7554800b",
           568 => x"0b0b0b9f",
           569 => x"ac087033",
           570 => x"51535371",
           571 => x"832e0981",
           572 => x"068c3894",
           573 => x"1451fdef",
           574 => x"3f880890",
           575 => x"2b539a14",
           576 => x"51fde43f",
           577 => x"880883ff",
           578 => x"ff067307",
           579 => x"880c853d",
           580 => x"0d04fc3d",
           581 => x"0d760b0b",
           582 => x"0b9fac08",
           583 => x"55558075",
           584 => x"23881508",
           585 => x"5372812e",
           586 => x"88388814",
           587 => x"08732685",
           588 => x"388152b0",
           589 => x"39729038",
           590 => x"73335271",
           591 => x"832e0981",
           592 => x"06853890",
           593 => x"14085372",
           594 => x"8c160c72",
           595 => x"802e8b38",
           596 => x"7251fed8",
           597 => x"3f880852",
           598 => x"85399014",
           599 => x"08527190",
           600 => x"160c8052",
           601 => x"71880c86",
           602 => x"3d0d04fa",
           603 => x"3d0d780b",
           604 => x"0b0b9fac",
           605 => x"08712281",
           606 => x"057083ff",
           607 => x"ff065754",
           608 => x"57557380",
           609 => x"2e883890",
           610 => x"15085372",
           611 => x"86388352",
           612 => x"80dc3973",
           613 => x"8f065271",
           614 => x"80cf3881",
           615 => x"1390160c",
           616 => x"8c150853",
           617 => x"728f3883",
           618 => x"0b841722",
           619 => x"57527376",
           620 => x"27bc38b5",
           621 => x"39821633",
           622 => x"ff057484",
           623 => x"2a065271",
           624 => x"a8387251",
           625 => x"fcdf3f81",
           626 => x"52718808",
           627 => x"27a03883",
           628 => x"52880888",
           629 => x"17082796",
           630 => x"3888088c",
           631 => x"160c8808",
           632 => x"51fdc93f",
           633 => x"88089016",
           634 => x"0c737523",
           635 => x"80527188",
           636 => x"0c883d0d",
           637 => x"04f23d0d",
           638 => x"60626458",
           639 => x"5e5c7533",
           640 => x"5574a02e",
           641 => x"09810688",
           642 => x"38811670",
           643 => x"4456ef39",
           644 => x"62703356",
           645 => x"5674af2e",
           646 => x"09810684",
           647 => x"38811643",
           648 => x"800b881d",
           649 => x"0c627033",
           650 => x"5155749f",
           651 => x"268f387b",
           652 => x"51fddf3f",
           653 => x"88085680",
           654 => x"7d3482d3",
           655 => x"39933d84",
           656 => x"1d087058",
           657 => x"5a5f8a55",
           658 => x"a0767081",
           659 => x"055834ff",
           660 => x"155574ff",
           661 => x"2e098106",
           662 => x"ef388070",
           663 => x"595b887f",
           664 => x"085f5a7a",
           665 => x"811c7081",
           666 => x"ff066013",
           667 => x"703370af",
           668 => x"327030a0",
           669 => x"73277180",
           670 => x"25075151",
           671 => x"525b535d",
           672 => x"57557480",
           673 => x"c73876ae",
           674 => x"2e098106",
           675 => x"83388155",
           676 => x"777a2775",
           677 => x"07557480",
           678 => x"2e9f3879",
           679 => x"88327030",
           680 => x"78ae3270",
           681 => x"30707307",
           682 => x"9f2a5351",
           683 => x"57515675",
           684 => x"9b388858",
           685 => x"8b5affab",
           686 => x"39778119",
           687 => x"7081ff06",
           688 => x"721c535a",
           689 => x"57557675",
           690 => x"34ff9839",
           691 => x"7a1e7f0c",
           692 => x"805576a0",
           693 => x"26833881",
           694 => x"55748b1a",
           695 => x"347b51fc",
           696 => x"b13f8808",
           697 => x"80ef38a0",
           698 => x"547b2270",
           699 => x"852b83e0",
           700 => x"06545590",
           701 => x"1c08527c",
           702 => x"51f8a83f",
           703 => x"88085788",
           704 => x"0880fb38",
           705 => x"7c335574",
           706 => x"802e80ee",
           707 => x"388b1d33",
           708 => x"70832a70",
           709 => x"81065156",
           710 => x"5674b238",
           711 => x"8b7d841e",
           712 => x"08880859",
           713 => x"5b5b58ff",
           714 => x"185877ff",
           715 => x"2e9a3879",
           716 => x"7081055b",
           717 => x"33797081",
           718 => x"055b3371",
           719 => x"71315256",
           720 => x"5675802e",
           721 => x"e2388639",
           722 => x"75802e92",
           723 => x"387b51fc",
           724 => x"9a3fff8e",
           725 => x"39880856",
           726 => x"8808b438",
           727 => x"83397656",
           728 => x"841c088b",
           729 => x"11335155",
           730 => x"74a5388b",
           731 => x"1d337084",
           732 => x"2a708106",
           733 => x"51565674",
           734 => x"89388356",
           735 => x"92398156",
           736 => x"8e397c51",
           737 => x"fad33f88",
           738 => x"08881d0c",
           739 => x"fdaf3975",
           740 => x"880c903d",
           741 => x"0d04f93d",
           742 => x"0d797b59",
           743 => x"57825483",
           744 => x"fe537752",
           745 => x"7651f6fb",
           746 => x"3f835688",
           747 => x"0880e738",
           748 => x"7651f8b3",
           749 => x"3f880883",
           750 => x"ffff0655",
           751 => x"82567482",
           752 => x"d4d52e09",
           753 => x"810680ce",
           754 => x"387554b6",
           755 => x"53775276",
           756 => x"51f6d03f",
           757 => x"88085688",
           758 => x"08943876",
           759 => x"51f8883f",
           760 => x"880883ff",
           761 => x"ff065574",
           762 => x"8182c62e",
           763 => x"a9388254",
           764 => x"80d25377",
           765 => x"527651f6",
           766 => x"aa3f8808",
           767 => x"56880894",
           768 => x"387651f7",
           769 => x"e23f8808",
           770 => x"83ffff06",
           771 => x"55748182",
           772 => x"c62e8338",
           773 => x"81567588",
           774 => x"0c893d0d",
           775 => x"04ed3d0d",
           776 => x"6559800b",
           777 => x"0b0b0b9f",
           778 => x"ac0cf59b",
           779 => x"3f880881",
           780 => x"06558256",
           781 => x"7482f238",
           782 => x"7475538d",
           783 => x"3d705357",
           784 => x"5afed33f",
           785 => x"880881ff",
           786 => x"06577681",
           787 => x"2e098106",
           788 => x"b3389054",
           789 => x"83be5374",
           790 => x"527551f5",
           791 => x"c63f8808",
           792 => x"ab388d3d",
           793 => x"33557480",
           794 => x"2eac3895",
           795 => x"3de40551",
           796 => x"f78a3f88",
           797 => x"08880853",
           798 => x"76525afe",
           799 => x"993f8808",
           800 => x"81ff0657",
           801 => x"76832e09",
           802 => x"81068638",
           803 => x"81568299",
           804 => x"3976802e",
           805 => x"86388656",
           806 => x"828f39a4",
           807 => x"548d5379",
           808 => x"527551f4",
           809 => x"fe3f8156",
           810 => x"880881fd",
           811 => x"38953de5",
           812 => x"0551f6b3",
           813 => x"3f880883",
           814 => x"ffff0658",
           815 => x"778c3895",
           816 => x"3df30551",
           817 => x"f6b63f88",
           818 => x"085802af",
           819 => x"05337871",
           820 => x"29028805",
           821 => x"ad057054",
           822 => x"52595bf6",
           823 => x"8a3f8808",
           824 => x"83ffff06",
           825 => x"7a058c1a",
           826 => x"0c8c3d33",
           827 => x"821a3495",
           828 => x"3de00551",
           829 => x"f5f13f88",
           830 => x"08841a23",
           831 => x"953de205",
           832 => x"51f5e43f",
           833 => x"880883ff",
           834 => x"ff065675",
           835 => x"8c38953d",
           836 => x"ef0551f5",
           837 => x"e73f8808",
           838 => x"567a51f5",
           839 => x"ca3f8808",
           840 => x"83ffff06",
           841 => x"76713179",
           842 => x"31841b22",
           843 => x"70842a82",
           844 => x"1d335672",
           845 => x"71315559",
           846 => x"5c5155ee",
           847 => x"c43f8808",
           848 => x"82057088",
           849 => x"1b0c8808",
           850 => x"e08a0556",
           851 => x"567483df",
           852 => x"fe268338",
           853 => x"825783ff",
           854 => x"f6762785",
           855 => x"38835789",
           856 => x"39865676",
           857 => x"802e80c1",
           858 => x"38767934",
           859 => x"76832e09",
           860 => x"81069038",
           861 => x"953dfb05",
           862 => x"51f5813f",
           863 => x"8808901a",
           864 => x"0c88398c",
           865 => x"19081890",
           866 => x"1a0c7983",
           867 => x"ffff068c",
           868 => x"1a081971",
           869 => x"842a0594",
           870 => x"1b0c5580",
           871 => x"0b811a34",
           872 => x"780b0b0b",
           873 => x"9fac0c80",
           874 => x"5675880c",
           875 => x"953d0d04",
           876 => x"ea3d0d0b",
           877 => x"0b0b9fac",
           878 => x"08558554",
           879 => x"74802e80",
           880 => x"df38800b",
           881 => x"81163498",
           882 => x"3de01145",
           883 => x"6954893d",
           884 => x"705457ec",
           885 => x"0551f89d",
           886 => x"3f880854",
           887 => x"880880c0",
           888 => x"38883d33",
           889 => x"5473802e",
           890 => x"933802a7",
           891 => x"05337084",
           892 => x"2a708106",
           893 => x"51555773",
           894 => x"802e8538",
           895 => x"8354a139",
           896 => x"7551f5d5",
           897 => x"3f8808a0",
           898 => x"160c983d",
           899 => x"dc0551f3",
           900 => x"eb3f8808",
           901 => x"9c160c73",
           902 => x"98160c81",
           903 => x"0b811634",
           904 => x"73880c98",
           905 => x"3d0d04f6",
           906 => x"3d0d7d7f",
           907 => x"7e0b0b0b",
           908 => x"9fac0859",
           909 => x"5b5c5880",
           910 => x"7b0c8557",
           911 => x"75802e81",
           912 => x"d1388116",
           913 => x"33810655",
           914 => x"84577480",
           915 => x"2e81c338",
           916 => x"91397481",
           917 => x"17348639",
           918 => x"800b8117",
           919 => x"34815781",
           920 => x"b1399c16",
           921 => x"08981708",
           922 => x"31557478",
           923 => x"27833874",
           924 => x"5877802e",
           925 => x"819a3898",
           926 => x"16087083",
           927 => x"ff065657",
           928 => x"7480c738",
           929 => x"821633ff",
           930 => x"0577892a",
           931 => x"067081ff",
           932 => x"065b5579",
           933 => x"9e387687",
           934 => x"38a01608",
           935 => x"558b39a4",
           936 => x"160851f3",
           937 => x"803f8808",
           938 => x"55817527",
           939 => x"ffaa3874",
           940 => x"a4170ca4",
           941 => x"160851f3",
           942 => x"f33f8808",
           943 => x"55880880",
           944 => x"2eff8f38",
           945 => x"88081aa8",
           946 => x"170c9816",
           947 => x"0883ff06",
           948 => x"84807131",
           949 => x"51557775",
           950 => x"27833877",
           951 => x"55745498",
           952 => x"160883ff",
           953 => x"0653a816",
           954 => x"08527851",
           955 => x"f0b53f88",
           956 => x"08fee538",
           957 => x"98160815",
           958 => x"98170c77",
           959 => x"75317b08",
           960 => x"167c0c58",
           961 => x"78802efe",
           962 => x"e8387419",
           963 => x"59fee239",
           964 => x"80577688",
           965 => x"0c8c3d0d",
           966 => x"04fb3d0d",
           967 => x"9b9086e4",
           968 => x"0b87c094",
           969 => x"8c0c9b90",
           970 => x"86e40b87",
           971 => x"c0949c0c",
           972 => x"8c80830b",
           973 => x"87c09484",
           974 => x"0c8c8083",
           975 => x"0b87c094",
           976 => x"940c9fb0",
           977 => x"51f9d63f",
           978 => x"8808b838",
           979 => x"9f9851fc",
           980 => x"df3f8808",
           981 => x"ae38a080",
           982 => x"0b880887",
           983 => x"c098880c",
           984 => x"55873dfc",
           985 => x"05538480",
           986 => x"527451fd",
           987 => x"ba3f8808",
           988 => x"8d387554",
           989 => x"73802e86",
           990 => x"38731555",
           991 => x"e439a080",
           992 => x"54730480",
           993 => x"54fb3900",
           994 => x"00ffffff",
           995 => x"ff00ffff",
           996 => x"ffff00ff",
           997 => x"ffffff00",
           998 => x"424f4f54",
           999 => x"54494e59",
          1000 => x"2e524f4d",
          1001 => x"00000000",
          1002 => x"01000000",
          2048 => x"0b0b0b92",
          2049 => x"d8040000",
          2050 => x"00000000",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b92",
          2121 => x"bc040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b929f",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b81bc",
          2210 => x"dc738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"92a40400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b0b93",
          2219 => x"dd2d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b0b95",
          2227 => x"c92d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"94040b0b",
          2317 => x"0b8ca304",
          2318 => x"0b0b0b8c",
          2319 => x"b2040b0b",
          2320 => x"0b8cc104",
          2321 => x"0b0b0b8c",
          2322 => x"d0040b0b",
          2323 => x"0b8cdf04",
          2324 => x"0b0b0b8c",
          2325 => x"ee040b0b",
          2326 => x"0b8cfd04",
          2327 => x"0b0b0b8d",
          2328 => x"8c040b0b",
          2329 => x"0b8d9b04",
          2330 => x"0b0b0b8d",
          2331 => x"aa040b0b",
          2332 => x"0b8db904",
          2333 => x"0b0b0b8d",
          2334 => x"c8040b0b",
          2335 => x"0b8dd704",
          2336 => x"0b0b0b8d",
          2337 => x"e6040b0b",
          2338 => x"0b8df504",
          2339 => x"0b0b0b8e",
          2340 => x"84040b0b",
          2341 => x"0b8e9404",
          2342 => x"0b0b0b8e",
          2343 => x"a4040b0b",
          2344 => x"0b8eb404",
          2345 => x"0b0b0b8e",
          2346 => x"c4040b0b",
          2347 => x"0b8ed404",
          2348 => x"0b0b0b8e",
          2349 => x"e4040b0b",
          2350 => x"0b8ef404",
          2351 => x"0b0b0b8f",
          2352 => x"84040b0b",
          2353 => x"0b8f9404",
          2354 => x"0b0b0b8f",
          2355 => x"a4040b0b",
          2356 => x"0b8fb404",
          2357 => x"0b0b0b8f",
          2358 => x"c4040b0b",
          2359 => x"0b8fd404",
          2360 => x"0b0b0b8f",
          2361 => x"e4040b0b",
          2362 => x"0b8ff404",
          2363 => x"0b0b0b90",
          2364 => x"84040b0b",
          2365 => x"0b909404",
          2366 => x"0b0b0b90",
          2367 => x"a4040b0b",
          2368 => x"0b90b404",
          2369 => x"0b0b0b90",
          2370 => x"c4040b0b",
          2371 => x"0b90d404",
          2372 => x"0b0b0b90",
          2373 => x"e4040b0b",
          2374 => x"0b90f404",
          2375 => x"0b0b0b91",
          2376 => x"84040b0b",
          2377 => x"0b919404",
          2378 => x"0b0b0b91",
          2379 => x"a3040b0b",
          2380 => x"0b91b204",
          2381 => x"0b0b0b91",
          2382 => x"c1040b0b",
          2383 => x"0b91d004",
          2384 => x"0b0b0b91",
          2385 => x"df040b0b",
          2386 => x"0b91ee04",
          2387 => x"ffffffff",
          2388 => x"ffffffff",
          2389 => x"ffffffff",
          2390 => x"ffffffff",
          2391 => x"ffffffff",
          2392 => x"ffffffff",
          2393 => x"ffffffff",
          2394 => x"ffffffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0481d390",
          2434 => x"0ca0ae2d",
          2435 => x"81d39008",
          2436 => x"82809004",
          2437 => x"81d3900c",
          2438 => x"aadc2d81",
          2439 => x"d3900882",
          2440 => x"80900481",
          2441 => x"d3900cab",
          2442 => x"9b2d81d3",
          2443 => x"90088280",
          2444 => x"900481d3",
          2445 => x"900cabb9",
          2446 => x"2d81d390",
          2447 => x"08828090",
          2448 => x"0481d390",
          2449 => x"0cb1f72d",
          2450 => x"81d39008",
          2451 => x"82809004",
          2452 => x"81d3900c",
          2453 => x"b2f52d81",
          2454 => x"d3900882",
          2455 => x"80900481",
          2456 => x"d3900cab",
          2457 => x"dc2d81d3",
          2458 => x"90088280",
          2459 => x"900481d3",
          2460 => x"900cb392",
          2461 => x"2d81d390",
          2462 => x"08828090",
          2463 => x"0481d390",
          2464 => x"0cb5842d",
          2465 => x"81d39008",
          2466 => x"82809004",
          2467 => x"81d3900c",
          2468 => x"b19d2d81",
          2469 => x"d3900882",
          2470 => x"80900481",
          2471 => x"d3900cb1",
          2472 => x"b32d81d3",
          2473 => x"90088280",
          2474 => x"900481d3",
          2475 => x"900cb1d7",
          2476 => x"2d81d390",
          2477 => x"08828090",
          2478 => x"0481d390",
          2479 => x"0ca2bb2d",
          2480 => x"81d39008",
          2481 => x"82809004",
          2482 => x"81d3900c",
          2483 => x"a38c2d81",
          2484 => x"d3900882",
          2485 => x"80900481",
          2486 => x"d3900c9b",
          2487 => x"a82d81d3",
          2488 => x"90088280",
          2489 => x"900481d3",
          2490 => x"900c9cdd",
          2491 => x"2d81d390",
          2492 => x"08828090",
          2493 => x"0481d390",
          2494 => x"0c9e902d",
          2495 => x"81d39008",
          2496 => x"82809004",
          2497 => x"81d3900c",
          2498 => x"80e7b92d",
          2499 => x"81d39008",
          2500 => x"82809004",
          2501 => x"81d3900c",
          2502 => x"80f4aa2d",
          2503 => x"81d39008",
          2504 => x"82809004",
          2505 => x"81d3900c",
          2506 => x"80ec9e2d",
          2507 => x"81d39008",
          2508 => x"82809004",
          2509 => x"81d3900c",
          2510 => x"80ef9b2d",
          2511 => x"81d39008",
          2512 => x"82809004",
          2513 => x"81d3900c",
          2514 => x"80f9b92d",
          2515 => x"81d39008",
          2516 => x"82809004",
          2517 => x"81d3900c",
          2518 => x"8182992d",
          2519 => x"81d39008",
          2520 => x"82809004",
          2521 => x"81d3900c",
          2522 => x"80f38c2d",
          2523 => x"81d39008",
          2524 => x"82809004",
          2525 => x"81d3900c",
          2526 => x"80fcd82d",
          2527 => x"81d39008",
          2528 => x"82809004",
          2529 => x"81d3900c",
          2530 => x"80fdf72d",
          2531 => x"81d39008",
          2532 => x"82809004",
          2533 => x"81d3900c",
          2534 => x"80fe962d",
          2535 => x"81d39008",
          2536 => x"82809004",
          2537 => x"81d3900c",
          2538 => x"8186802d",
          2539 => x"81d39008",
          2540 => x"82809004",
          2541 => x"81d3900c",
          2542 => x"8183e62d",
          2543 => x"81d39008",
          2544 => x"82809004",
          2545 => x"81d3900c",
          2546 => x"8188d42d",
          2547 => x"81d39008",
          2548 => x"82809004",
          2549 => x"81d3900c",
          2550 => x"80ff9a2d",
          2551 => x"81d39008",
          2552 => x"82809004",
          2553 => x"81d3900c",
          2554 => x"818bd42d",
          2555 => x"81d39008",
          2556 => x"82809004",
          2557 => x"81d3900c",
          2558 => x"818cd52d",
          2559 => x"81d39008",
          2560 => x"82809004",
          2561 => x"81d3900c",
          2562 => x"80f58a2d",
          2563 => x"81d39008",
          2564 => x"82809004",
          2565 => x"81d3900c",
          2566 => x"80f4e32d",
          2567 => x"81d39008",
          2568 => x"82809004",
          2569 => x"81d3900c",
          2570 => x"80f68e2d",
          2571 => x"81d39008",
          2572 => x"82809004",
          2573 => x"81d3900c",
          2574 => x"80fff12d",
          2575 => x"81d39008",
          2576 => x"82809004",
          2577 => x"81d3900c",
          2578 => x"818dc62d",
          2579 => x"81d39008",
          2580 => x"82809004",
          2581 => x"81d3900c",
          2582 => x"818fd02d",
          2583 => x"81d39008",
          2584 => x"82809004",
          2585 => x"81d3900c",
          2586 => x"8193922d",
          2587 => x"81d39008",
          2588 => x"82809004",
          2589 => x"81d3900c",
          2590 => x"80e6d82d",
          2591 => x"81d39008",
          2592 => x"82809004",
          2593 => x"81d3900c",
          2594 => x"8195fe2d",
          2595 => x"81d39008",
          2596 => x"82809004",
          2597 => x"81d3900c",
          2598 => x"b8932d81",
          2599 => x"d3900882",
          2600 => x"80900481",
          2601 => x"d3900cb9",
          2602 => x"fd2d81d3",
          2603 => x"90088280",
          2604 => x"900481d3",
          2605 => x"900cbbe1",
          2606 => x"2d81d390",
          2607 => x"08828090",
          2608 => x"0481d390",
          2609 => x"0c9bd12d",
          2610 => x"81d39008",
          2611 => x"82809004",
          2612 => x"81d3900c",
          2613 => x"9cb32d81",
          2614 => x"d3900882",
          2615 => x"80900481",
          2616 => x"d3900c9f",
          2617 => x"a02d81d3",
          2618 => x"90088280",
          2619 => x"900481d3",
          2620 => x"900c81a2",
          2621 => x"9f2d81d3",
          2622 => x"90088280",
          2623 => x"90043c04",
          2624 => x"10101010",
          2625 => x"10101010",
          2626 => x"10101010",
          2627 => x"10101010",
          2628 => x"10101010",
          2629 => x"10101010",
          2630 => x"10101010",
          2631 => x"10101053",
          2632 => x"51040000",
          2633 => x"7381ff06",
          2634 => x"73830609",
          2635 => x"81058305",
          2636 => x"1010102b",
          2637 => x"0772fc06",
          2638 => x"0c515104",
          2639 => x"72728072",
          2640 => x"8106ff05",
          2641 => x"09720605",
          2642 => x"71105272",
          2643 => x"0a100a53",
          2644 => x"72ed3851",
          2645 => x"51535104",
          2646 => x"81d38470",
          2647 => x"81ea8827",
          2648 => x"8e388071",
          2649 => x"70840553",
          2650 => x"0c0b0b0b",
          2651 => x"92db048c",
          2652 => x"815181bb",
          2653 => x"f3040081",
          2654 => x"d3900802",
          2655 => x"81d3900c",
          2656 => x"fd3d0d80",
          2657 => x"5381d390",
          2658 => x"088c0508",
          2659 => x"5281d390",
          2660 => x"08880508",
          2661 => x"5183d43f",
          2662 => x"81d38408",
          2663 => x"7081d384",
          2664 => x"0c54853d",
          2665 => x"0d81d390",
          2666 => x"0c0481d3",
          2667 => x"90080281",
          2668 => x"d3900cfd",
          2669 => x"3d0d8153",
          2670 => x"81d39008",
          2671 => x"8c050852",
          2672 => x"81d39008",
          2673 => x"88050851",
          2674 => x"83a13f81",
          2675 => x"d3840870",
          2676 => x"81d3840c",
          2677 => x"54853d0d",
          2678 => x"81d3900c",
          2679 => x"0481d390",
          2680 => x"080281d3",
          2681 => x"900cf93d",
          2682 => x"0d800b81",
          2683 => x"d39008fc",
          2684 => x"050c81d3",
          2685 => x"90088805",
          2686 => x"088025b9",
          2687 => x"3881d390",
          2688 => x"08880508",
          2689 => x"3081d390",
          2690 => x"0888050c",
          2691 => x"800b81d3",
          2692 => x"9008f405",
          2693 => x"0c81d390",
          2694 => x"08fc0508",
          2695 => x"8a38810b",
          2696 => x"81d39008",
          2697 => x"f4050c81",
          2698 => x"d39008f4",
          2699 => x"050881d3",
          2700 => x"9008fc05",
          2701 => x"0c81d390",
          2702 => x"088c0508",
          2703 => x"8025b938",
          2704 => x"81d39008",
          2705 => x"8c050830",
          2706 => x"81d39008",
          2707 => x"8c050c80",
          2708 => x"0b81d390",
          2709 => x"08f0050c",
          2710 => x"81d39008",
          2711 => x"fc05088a",
          2712 => x"38810b81",
          2713 => x"d39008f0",
          2714 => x"050c81d3",
          2715 => x"9008f005",
          2716 => x"0881d390",
          2717 => x"08fc050c",
          2718 => x"805381d3",
          2719 => x"90088c05",
          2720 => x"085281d3",
          2721 => x"90088805",
          2722 => x"085181df",
          2723 => x"3f81d384",
          2724 => x"087081d3",
          2725 => x"9008f805",
          2726 => x"0c5481d3",
          2727 => x"9008fc05",
          2728 => x"08802e90",
          2729 => x"3881d390",
          2730 => x"08f80508",
          2731 => x"3081d390",
          2732 => x"08f8050c",
          2733 => x"81d39008",
          2734 => x"f8050870",
          2735 => x"81d3840c",
          2736 => x"54893d0d",
          2737 => x"81d3900c",
          2738 => x"0481d390",
          2739 => x"080281d3",
          2740 => x"900cfb3d",
          2741 => x"0d800b81",
          2742 => x"d39008fc",
          2743 => x"050c81d3",
          2744 => x"90088805",
          2745 => x"08802599",
          2746 => x"3881d390",
          2747 => x"08880508",
          2748 => x"3081d390",
          2749 => x"0888050c",
          2750 => x"810b81d3",
          2751 => x"9008fc05",
          2752 => x"0c81d390",
          2753 => x"088c0508",
          2754 => x"80259038",
          2755 => x"81d39008",
          2756 => x"8c050830",
          2757 => x"81d39008",
          2758 => x"8c050c81",
          2759 => x"5381d390",
          2760 => x"088c0508",
          2761 => x"5281d390",
          2762 => x"08880508",
          2763 => x"51bd3f81",
          2764 => x"d3840870",
          2765 => x"81d39008",
          2766 => x"f8050c54",
          2767 => x"81d39008",
          2768 => x"fc050880",
          2769 => x"2e903881",
          2770 => x"d39008f8",
          2771 => x"05083081",
          2772 => x"d39008f8",
          2773 => x"050c81d3",
          2774 => x"9008f805",
          2775 => x"087081d3",
          2776 => x"840c5487",
          2777 => x"3d0d81d3",
          2778 => x"900c0481",
          2779 => x"d3900802",
          2780 => x"81d3900c",
          2781 => x"fd3d0d81",
          2782 => x"0b81d390",
          2783 => x"08fc050c",
          2784 => x"800b81d3",
          2785 => x"9008f805",
          2786 => x"0c81d390",
          2787 => x"088c0508",
          2788 => x"81d39008",
          2789 => x"88050827",
          2790 => x"b93881d3",
          2791 => x"9008fc05",
          2792 => x"08802eae",
          2793 => x"38800b81",
          2794 => x"d390088c",
          2795 => x"050824a2",
          2796 => x"3881d390",
          2797 => x"088c0508",
          2798 => x"1081d390",
          2799 => x"088c050c",
          2800 => x"81d39008",
          2801 => x"fc050810",
          2802 => x"81d39008",
          2803 => x"fc050cff",
          2804 => x"b83981d3",
          2805 => x"9008fc05",
          2806 => x"08802e80",
          2807 => x"e13881d3",
          2808 => x"90088c05",
          2809 => x"0881d390",
          2810 => x"08880508",
          2811 => x"26ad3881",
          2812 => x"d3900888",
          2813 => x"050881d3",
          2814 => x"90088c05",
          2815 => x"083181d3",
          2816 => x"90088805",
          2817 => x"0c81d390",
          2818 => x"08f80508",
          2819 => x"81d39008",
          2820 => x"fc050807",
          2821 => x"81d39008",
          2822 => x"f8050c81",
          2823 => x"d39008fc",
          2824 => x"0508812a",
          2825 => x"81d39008",
          2826 => x"fc050c81",
          2827 => x"d390088c",
          2828 => x"0508812a",
          2829 => x"81d39008",
          2830 => x"8c050cff",
          2831 => x"953981d3",
          2832 => x"90089005",
          2833 => x"08802e93",
          2834 => x"3881d390",
          2835 => x"08880508",
          2836 => x"7081d390",
          2837 => x"08f4050c",
          2838 => x"51913981",
          2839 => x"d39008f8",
          2840 => x"05087081",
          2841 => x"d39008f4",
          2842 => x"050c5181",
          2843 => x"d39008f4",
          2844 => x"050881d3",
          2845 => x"840c853d",
          2846 => x"0d81d390",
          2847 => x"0c04fc3d",
          2848 => x"0d767971",
          2849 => x"028c059f",
          2850 => x"05335755",
          2851 => x"53558372",
          2852 => x"278a3874",
          2853 => x"83065170",
          2854 => x"802ea438",
          2855 => x"ff125271",
          2856 => x"ff2e9338",
          2857 => x"73737081",
          2858 => x"055534ff",
          2859 => x"125271ff",
          2860 => x"2e098106",
          2861 => x"ef387481",
          2862 => x"d3840c86",
          2863 => x"3d0d0474",
          2864 => x"74882b75",
          2865 => x"07707190",
          2866 => x"2b075154",
          2867 => x"518f7227",
          2868 => x"a5387271",
          2869 => x"70840553",
          2870 => x"0c727170",
          2871 => x"8405530c",
          2872 => x"72717084",
          2873 => x"05530c72",
          2874 => x"71708405",
          2875 => x"530cf012",
          2876 => x"52718f26",
          2877 => x"dd388372",
          2878 => x"27903872",
          2879 => x"71708405",
          2880 => x"530cfc12",
          2881 => x"52718326",
          2882 => x"f2387053",
          2883 => x"ff8e39fb",
          2884 => x"3d0d7779",
          2885 => x"70720783",
          2886 => x"06535452",
          2887 => x"70933871",
          2888 => x"73730854",
          2889 => x"56547173",
          2890 => x"082e80c6",
          2891 => x"38737554",
          2892 => x"52713370",
          2893 => x"81ff0652",
          2894 => x"5470802e",
          2895 => x"9d387233",
          2896 => x"5570752e",
          2897 => x"09810695",
          2898 => x"38811281",
          2899 => x"14713370",
          2900 => x"81ff0654",
          2901 => x"56545270",
          2902 => x"e5387233",
          2903 => x"557381ff",
          2904 => x"067581ff",
          2905 => x"06717131",
          2906 => x"81d3840c",
          2907 => x"5252873d",
          2908 => x"0d047109",
          2909 => x"70f7fbfd",
          2910 => x"ff140670",
          2911 => x"f8848281",
          2912 => x"80065151",
          2913 => x"51709738",
          2914 => x"84148416",
          2915 => x"71085456",
          2916 => x"54717508",
          2917 => x"2edc3873",
          2918 => x"755452ff",
          2919 => x"9439800b",
          2920 => x"81d3840c",
          2921 => x"873d0d04",
          2922 => x"fe3d0d80",
          2923 => x"52835371",
          2924 => x"882b5287",
          2925 => x"863f81d3",
          2926 => x"840881ff",
          2927 => x"067207ff",
          2928 => x"14545272",
          2929 => x"8025e838",
          2930 => x"7181d384",
          2931 => x"0c843d0d",
          2932 => x"04fb3d0d",
          2933 => x"77700870",
          2934 => x"53535671",
          2935 => x"802e80ca",
          2936 => x"38713351",
          2937 => x"70a02e09",
          2938 => x"81068638",
          2939 => x"811252f1",
          2940 => x"39715384",
          2941 => x"39811353",
          2942 => x"80733370",
          2943 => x"81ff0653",
          2944 => x"555570a0",
          2945 => x"2e833881",
          2946 => x"5570802e",
          2947 => x"843874e5",
          2948 => x"387381ff",
          2949 => x"065170a0",
          2950 => x"2e098106",
          2951 => x"88388073",
          2952 => x"70810555",
          2953 => x"3472760c",
          2954 => x"71517081",
          2955 => x"d3840c87",
          2956 => x"3d0d04fc",
          2957 => x"3d0d7653",
          2958 => x"7208802e",
          2959 => x"9138863d",
          2960 => x"fc055272",
          2961 => x"5198bd3f",
          2962 => x"81d38408",
          2963 => x"85388053",
          2964 => x"83397453",
          2965 => x"7281d384",
          2966 => x"0c863d0d",
          2967 => x"04fc3d0d",
          2968 => x"76821133",
          2969 => x"ff055253",
          2970 => x"8152708b",
          2971 => x"26819838",
          2972 => x"831333ff",
          2973 => x"05518252",
          2974 => x"709e2681",
          2975 => x"8a388413",
          2976 => x"33518352",
          2977 => x"70972680",
          2978 => x"fe388513",
          2979 => x"33518452",
          2980 => x"70bb2680",
          2981 => x"f2388613",
          2982 => x"33518552",
          2983 => x"70bb2680",
          2984 => x"e6388813",
          2985 => x"22558652",
          2986 => x"7487e726",
          2987 => x"80d9388a",
          2988 => x"13225487",
          2989 => x"527387e7",
          2990 => x"2680cc38",
          2991 => x"810b87c0",
          2992 => x"989c0c72",
          2993 => x"2287c098",
          2994 => x"bc0c8213",
          2995 => x"3387c098",
          2996 => x"b80c8313",
          2997 => x"3387c098",
          2998 => x"b40c8413",
          2999 => x"3387c098",
          3000 => x"b00c8513",
          3001 => x"3387c098",
          3002 => x"ac0c8613",
          3003 => x"3387c098",
          3004 => x"a80c7487",
          3005 => x"c098a40c",
          3006 => x"7387c098",
          3007 => x"a00c800b",
          3008 => x"87c0989c",
          3009 => x"0c805271",
          3010 => x"81d3840c",
          3011 => x"863d0d04",
          3012 => x"f33d0d7f",
          3013 => x"5b87c098",
          3014 => x"9c5d817d",
          3015 => x"0c87c098",
          3016 => x"bc085e7d",
          3017 => x"7b2387c0",
          3018 => x"98b8085a",
          3019 => x"79821c34",
          3020 => x"87c098b4",
          3021 => x"085a7983",
          3022 => x"1c3487c0",
          3023 => x"98b0085a",
          3024 => x"79841c34",
          3025 => x"87c098ac",
          3026 => x"085a7985",
          3027 => x"1c3487c0",
          3028 => x"98a8085a",
          3029 => x"79861c34",
          3030 => x"87c098a4",
          3031 => x"085c7b88",
          3032 => x"1c2387c0",
          3033 => x"98a0085a",
          3034 => x"798a1c23",
          3035 => x"807d0c79",
          3036 => x"83ffff06",
          3037 => x"597b83ff",
          3038 => x"ff065886",
          3039 => x"1b335785",
          3040 => x"1b335684",
          3041 => x"1b335583",
          3042 => x"1b335482",
          3043 => x"1b33537d",
          3044 => x"83ffff06",
          3045 => x"5281bdd0",
          3046 => x"5192823f",
          3047 => x"8f3d0d04",
          3048 => x"ff3d0d02",
          3049 => x"8f053370",
          3050 => x"30709f2a",
          3051 => x"51525270",
          3052 => x"0b0b81cf",
          3053 => x"fc34833d",
          3054 => x"0d04fb3d",
          3055 => x"0d770b0b",
          3056 => x"81cffc33",
          3057 => x"7081ff06",
          3058 => x"57555687",
          3059 => x"c0948451",
          3060 => x"74802e86",
          3061 => x"3887c094",
          3062 => x"94517008",
          3063 => x"70962a70",
          3064 => x"81065354",
          3065 => x"5270802e",
          3066 => x"8c387191",
          3067 => x"2a708106",
          3068 => x"515170d7",
          3069 => x"38728132",
          3070 => x"70810651",
          3071 => x"5170802e",
          3072 => x"8d387193",
          3073 => x"2a708106",
          3074 => x"515170ff",
          3075 => x"be387381",
          3076 => x"ff065187",
          3077 => x"c0948052",
          3078 => x"70802e86",
          3079 => x"3887c094",
          3080 => x"90527572",
          3081 => x"0c7581d3",
          3082 => x"840c873d",
          3083 => x"0d04fb3d",
          3084 => x"0d029f05",
          3085 => x"330b0b81",
          3086 => x"cffc3370",
          3087 => x"81ff0657",
          3088 => x"555687c0",
          3089 => x"94845174",
          3090 => x"802e8638",
          3091 => x"87c09494",
          3092 => x"51700870",
          3093 => x"962a7081",
          3094 => x"06535452",
          3095 => x"70802e8c",
          3096 => x"3871912a",
          3097 => x"70810651",
          3098 => x"5170d738",
          3099 => x"72813270",
          3100 => x"81065151",
          3101 => x"70802e8d",
          3102 => x"3871932a",
          3103 => x"70810651",
          3104 => x"5170ffbe",
          3105 => x"387381ff",
          3106 => x"065187c0",
          3107 => x"94805270",
          3108 => x"802e8638",
          3109 => x"87c09490",
          3110 => x"5275720c",
          3111 => x"873d0d04",
          3112 => x"f93d0d79",
          3113 => x"54807433",
          3114 => x"7081ff06",
          3115 => x"53535770",
          3116 => x"772e80fe",
          3117 => x"387181ff",
          3118 => x"0681150b",
          3119 => x"0b81cffc",
          3120 => x"337081ff",
          3121 => x"06595755",
          3122 => x"5887c094",
          3123 => x"84517580",
          3124 => x"2e863887",
          3125 => x"c0949451",
          3126 => x"70087096",
          3127 => x"2a708106",
          3128 => x"53545270",
          3129 => x"802e8c38",
          3130 => x"71912a70",
          3131 => x"81065151",
          3132 => x"70d73872",
          3133 => x"81327081",
          3134 => x"06515170",
          3135 => x"802e8d38",
          3136 => x"71932a70",
          3137 => x"81065151",
          3138 => x"70ffbe38",
          3139 => x"7481ff06",
          3140 => x"5187c094",
          3141 => x"80527080",
          3142 => x"2e863887",
          3143 => x"c0949052",
          3144 => x"77720c81",
          3145 => x"17743370",
          3146 => x"81ff0653",
          3147 => x"535770ff",
          3148 => x"84387681",
          3149 => x"d3840c89",
          3150 => x"3d0d04fe",
          3151 => x"3d0d0b0b",
          3152 => x"81cffc33",
          3153 => x"7081ff06",
          3154 => x"545287c0",
          3155 => x"94845172",
          3156 => x"802e8638",
          3157 => x"87c09494",
          3158 => x"51700870",
          3159 => x"822a7081",
          3160 => x"06515151",
          3161 => x"70802ee2",
          3162 => x"387181ff",
          3163 => x"065187c0",
          3164 => x"94805270",
          3165 => x"802e8638",
          3166 => x"87c09490",
          3167 => x"52710870",
          3168 => x"81ff0681",
          3169 => x"d3840c51",
          3170 => x"843d0d04",
          3171 => x"fe3d0d0b",
          3172 => x"0b81cffc",
          3173 => x"337081ff",
          3174 => x"06525387",
          3175 => x"c0948452",
          3176 => x"70802e86",
          3177 => x"3887c094",
          3178 => x"94527108",
          3179 => x"70822a70",
          3180 => x"81065151",
          3181 => x"51ff5270",
          3182 => x"802ea038",
          3183 => x"7281ff06",
          3184 => x"5187c094",
          3185 => x"80527080",
          3186 => x"2e863887",
          3187 => x"c0949052",
          3188 => x"71087098",
          3189 => x"2b70982c",
          3190 => x"51535171",
          3191 => x"81d3840c",
          3192 => x"843d0d04",
          3193 => x"ff3d0d87",
          3194 => x"c09e8008",
          3195 => x"709c2a8a",
          3196 => x"06515170",
          3197 => x"802e8393",
          3198 => x"3887c09e",
          3199 => x"9c0881d0",
          3200 => x"800c87c0",
          3201 => x"9ea00881",
          3202 => x"d0840c87",
          3203 => x"c09e8c08",
          3204 => x"81d0880c",
          3205 => x"87c09e90",
          3206 => x"0881d08c",
          3207 => x"0c87c09e",
          3208 => x"940881d0",
          3209 => x"900c87c0",
          3210 => x"9e980881",
          3211 => x"d0940c87",
          3212 => x"c09ea408",
          3213 => x"81d0980c",
          3214 => x"87c09ea8",
          3215 => x"0881d09c",
          3216 => x"0c87c09e",
          3217 => x"ac0881d0",
          3218 => x"a00c87c0",
          3219 => x"9e800851",
          3220 => x"7081d0a4",
          3221 => x"2387c09e",
          3222 => x"840881d0",
          3223 => x"a80c810b",
          3224 => x"81d0ac34",
          3225 => x"800b87c0",
          3226 => x"9e880870",
          3227 => x"a0800651",
          3228 => x"52527080",
          3229 => x"2e833881",
          3230 => x"527181d0",
          3231 => x"ad34800b",
          3232 => x"87c09e88",
          3233 => x"08708180",
          3234 => x"80065152",
          3235 => x"5270802e",
          3236 => x"83388152",
          3237 => x"7181d0ae",
          3238 => x"34800b87",
          3239 => x"c09e8808",
          3240 => x"7080c080",
          3241 => x"06515252",
          3242 => x"70802e83",
          3243 => x"38815271",
          3244 => x"81d0af34",
          3245 => x"800b87c0",
          3246 => x"9e880870",
          3247 => x"90800651",
          3248 => x"52527080",
          3249 => x"2e833881",
          3250 => x"527181d0",
          3251 => x"b034800b",
          3252 => x"87c09e88",
          3253 => x"08708880",
          3254 => x"06515252",
          3255 => x"70802e83",
          3256 => x"38815271",
          3257 => x"81d0b134",
          3258 => x"800b87c0",
          3259 => x"9e880870",
          3260 => x"84800651",
          3261 => x"52527080",
          3262 => x"2e833881",
          3263 => x"527181d0",
          3264 => x"b234800b",
          3265 => x"87c09e88",
          3266 => x"08708280",
          3267 => x"06515252",
          3268 => x"70802e83",
          3269 => x"38815271",
          3270 => x"81d0b334",
          3271 => x"800b87c0",
          3272 => x"9e880870",
          3273 => x"81800651",
          3274 => x"52527080",
          3275 => x"2e833881",
          3276 => x"527181d0",
          3277 => x"b43487c0",
          3278 => x"9e880870",
          3279 => x"80e00670",
          3280 => x"862c5151",
          3281 => x"517081d0",
          3282 => x"b534800b",
          3283 => x"87c09e88",
          3284 => x"08709006",
          3285 => x"51525270",
          3286 => x"802e8338",
          3287 => x"81527181",
          3288 => x"d0b63480",
          3289 => x"0b87c09e",
          3290 => x"88087088",
          3291 => x"06515252",
          3292 => x"70802e83",
          3293 => x"38815271",
          3294 => x"81d0b734",
          3295 => x"87c09e88",
          3296 => x"08708706",
          3297 => x"51517081",
          3298 => x"d0b83483",
          3299 => x"3d0d04fd",
          3300 => x"3d0d81bd",
          3301 => x"e85184a1",
          3302 => x"3f81d0ac",
          3303 => x"33547380",
          3304 => x"2e883881",
          3305 => x"bdfc5184",
          3306 => x"903f81be",
          3307 => x"90518489",
          3308 => x"3f81d0ad",
          3309 => x"33547380",
          3310 => x"2e923881",
          3311 => x"d0840853",
          3312 => x"81d08008",
          3313 => x"5281bea8",
          3314 => x"5189d23f",
          3315 => x"81d0ae33",
          3316 => x"5473802e",
          3317 => x"923881d0",
          3318 => x"8c085381",
          3319 => x"d0880852",
          3320 => x"81bed051",
          3321 => x"89b73f81",
          3322 => x"d0af3354",
          3323 => x"738b3881",
          3324 => x"d0b03354",
          3325 => x"73802e92",
          3326 => x"3881d094",
          3327 => x"085381d0",
          3328 => x"90085281",
          3329 => x"bef45189",
          3330 => x"943f81d0",
          3331 => x"b1335473",
          3332 => x"802e8838",
          3333 => x"81bf9851",
          3334 => x"839f3f81",
          3335 => x"d0b23354",
          3336 => x"73802e88",
          3337 => x"3881bfa4",
          3338 => x"51838e3f",
          3339 => x"81d0b333",
          3340 => x"5473802e",
          3341 => x"883881bf",
          3342 => x"b05182fd",
          3343 => x"3f81d0b4",
          3344 => x"33547380",
          3345 => x"2e8d3881",
          3346 => x"d0b53352",
          3347 => x"81bfbc51",
          3348 => x"88cb3f81",
          3349 => x"d0b63354",
          3350 => x"73802e88",
          3351 => x"3881bfdc",
          3352 => x"5182d63f",
          3353 => x"81d0b733",
          3354 => x"5473802e",
          3355 => x"8d3881d0",
          3356 => x"b8335281",
          3357 => x"bff85188",
          3358 => x"a43f81c0",
          3359 => x"945182b9",
          3360 => x"3f81d098",
          3361 => x"085281c0",
          3362 => x"a0518891",
          3363 => x"3f81d09c",
          3364 => x"085281c0",
          3365 => x"c8518885",
          3366 => x"3f81d0a0",
          3367 => x"085281c0",
          3368 => x"f05187f9",
          3369 => x"3f81d0a4",
          3370 => x"225281c1",
          3371 => x"985187ed",
          3372 => x"3f81d0a8",
          3373 => x"085281c1",
          3374 => x"c05187e1",
          3375 => x"3f853d0d",
          3376 => x"04fe3d0d",
          3377 => x"02920533",
          3378 => x"ff055271",
          3379 => x"8426aa38",
          3380 => x"71842981",
          3381 => x"bcec0552",
          3382 => x"71080481",
          3383 => x"c1e8519d",
          3384 => x"3981c1f0",
          3385 => x"51973981",
          3386 => x"c1f85191",
          3387 => x"3981c280",
          3388 => x"518b3981",
          3389 => x"c2845185",
          3390 => x"3981c28c",
          3391 => x"51f7a13f",
          3392 => x"843d0d04",
          3393 => x"7188800c",
          3394 => x"04800b87",
          3395 => x"c096840c",
          3396 => x"04ff3d0d",
          3397 => x"87c09684",
          3398 => x"70085252",
          3399 => x"80720c70",
          3400 => x"74077081",
          3401 => x"d0bc0c72",
          3402 => x"0c833d0d",
          3403 => x"04ff3d0d",
          3404 => x"87c09684",
          3405 => x"700881d0",
          3406 => x"bc0c5280",
          3407 => x"720c7309",
          3408 => x"7081d0bc",
          3409 => x"08067081",
          3410 => x"d0bc0c73",
          3411 => x"0c51833d",
          3412 => x"0d0481d0",
          3413 => x"bc0887c0",
          3414 => x"96840c04",
          3415 => x"fe3d0d02",
          3416 => x"93053353",
          3417 => x"728a2e09",
          3418 => x"81068538",
          3419 => x"8d51ed3f",
          3420 => x"81d39c08",
          3421 => x"5271802e",
          3422 => x"90387272",
          3423 => x"3481d39c",
          3424 => x"08810581",
          3425 => x"d39c0c8f",
          3426 => x"3981d394",
          3427 => x"08527180",
          3428 => x"2e853872",
          3429 => x"51712d84",
          3430 => x"3d0d04fe",
          3431 => x"3d0d0297",
          3432 => x"053381d3",
          3433 => x"94087681",
          3434 => x"d3940c54",
          3435 => x"51ffad3f",
          3436 => x"7281d394",
          3437 => x"0c843d0d",
          3438 => x"04fd3d0d",
          3439 => x"75547333",
          3440 => x"7081ff06",
          3441 => x"53537180",
          3442 => x"2e8e3872",
          3443 => x"81ff0651",
          3444 => x"811454ff",
          3445 => x"873fe739",
          3446 => x"853d0d04",
          3447 => x"fc3d0d77",
          3448 => x"81d39408",
          3449 => x"7881d394",
          3450 => x"0c565473",
          3451 => x"337081ff",
          3452 => x"06535371",
          3453 => x"802e8e38",
          3454 => x"7281ff06",
          3455 => x"51811454",
          3456 => x"feda3fe7",
          3457 => x"397481d3",
          3458 => x"940c863d",
          3459 => x"0d04ec3d",
          3460 => x"0d666859",
          3461 => x"59787081",
          3462 => x"055a3356",
          3463 => x"75802e84",
          3464 => x"f83875a5",
          3465 => x"2e098106",
          3466 => x"82de3880",
          3467 => x"707a7081",
          3468 => x"055c3358",
          3469 => x"5b5b75b0",
          3470 => x"2e098106",
          3471 => x"8538815a",
          3472 => x"8b3975ad",
          3473 => x"2e098106",
          3474 => x"8a38825a",
          3475 => x"78708105",
          3476 => x"5a335675",
          3477 => x"aa2e0981",
          3478 => x"06923877",
          3479 => x"84197108",
          3480 => x"7b708105",
          3481 => x"5d33595d",
          3482 => x"59539d39",
          3483 => x"d0165372",
          3484 => x"89269538",
          3485 => x"7a88297b",
          3486 => x"10057605",
          3487 => x"d0057970",
          3488 => x"81055b33",
          3489 => x"575be539",
          3490 => x"7580ec32",
          3491 => x"70307072",
          3492 => x"07802578",
          3493 => x"80cc3270",
          3494 => x"30707207",
          3495 => x"80257307",
          3496 => x"53545851",
          3497 => x"55537380",
          3498 => x"2e8c3879",
          3499 => x"84077970",
          3500 => x"81055b33",
          3501 => x"575a7580",
          3502 => x"2e83de38",
          3503 => x"755480e0",
          3504 => x"76278938",
          3505 => x"e0167081",
          3506 => x"ff065553",
          3507 => x"7380cf2e",
          3508 => x"81aa3873",
          3509 => x"80cf24a2",
          3510 => x"387380c3",
          3511 => x"2e818e38",
          3512 => x"7380c324",
          3513 => x"8b387380",
          3514 => x"c22e818c",
          3515 => x"38819939",
          3516 => x"7380c42e",
          3517 => x"818a3881",
          3518 => x"8f397380",
          3519 => x"d52e8180",
          3520 => x"387380d5",
          3521 => x"248a3873",
          3522 => x"80d32e8e",
          3523 => x"3880f939",
          3524 => x"7380d82e",
          3525 => x"80ee3880",
          3526 => x"ef397784",
          3527 => x"19710856",
          3528 => x"59538074",
          3529 => x"33545572",
          3530 => x"752e8d38",
          3531 => x"81157015",
          3532 => x"70335154",
          3533 => x"5572f538",
          3534 => x"79812a56",
          3535 => x"90397481",
          3536 => x"16565372",
          3537 => x"7b278f38",
          3538 => x"a051fc90",
          3539 => x"3f758106",
          3540 => x"5372802e",
          3541 => x"e9387351",
          3542 => x"fcdf3f74",
          3543 => x"81165653",
          3544 => x"727b27fd",
          3545 => x"b038a051",
          3546 => x"fbf23fef",
          3547 => x"39778419",
          3548 => x"83123353",
          3549 => x"59539339",
          3550 => x"825c9539",
          3551 => x"885c9139",
          3552 => x"8a5c8d39",
          3553 => x"905c8939",
          3554 => x"7551fbd0",
          3555 => x"3ffd8639",
          3556 => x"79822a70",
          3557 => x"81065153",
          3558 => x"72802e88",
          3559 => x"38778419",
          3560 => x"59538639",
          3561 => x"84187854",
          3562 => x"58720874",
          3563 => x"80c43270",
          3564 => x"30707207",
          3565 => x"80255155",
          3566 => x"55557480",
          3567 => x"258d3872",
          3568 => x"802e8838",
          3569 => x"74307a90",
          3570 => x"075b5580",
          3571 => x"0b8f3d5e",
          3572 => x"577b5274",
          3573 => x"51e3d33f",
          3574 => x"81d38408",
          3575 => x"81ff067c",
          3576 => x"53755254",
          3577 => x"e3913f81",
          3578 => x"d3840855",
          3579 => x"89742792",
          3580 => x"38a71453",
          3581 => x"7580f82e",
          3582 => x"84388714",
          3583 => x"537281ff",
          3584 => x"0654b014",
          3585 => x"53727d70",
          3586 => x"81055f34",
          3587 => x"81177530",
          3588 => x"7077079f",
          3589 => x"2a515457",
          3590 => x"769f2685",
          3591 => x"3872ffb1",
          3592 => x"3879842a",
          3593 => x"70810651",
          3594 => x"5372802e",
          3595 => x"8e38963d",
          3596 => x"7705e005",
          3597 => x"53ad7334",
          3598 => x"81175776",
          3599 => x"7a810654",
          3600 => x"55b05472",
          3601 => x"8338a054",
          3602 => x"79812a70",
          3603 => x"81065456",
          3604 => x"729f3881",
          3605 => x"1755767b",
          3606 => x"27973873",
          3607 => x"51f9fd3f",
          3608 => x"75810653",
          3609 => x"728b3874",
          3610 => x"81165653",
          3611 => x"7a7326eb",
          3612 => x"38963d77",
          3613 => x"05e00553",
          3614 => x"ff17ff14",
          3615 => x"70335354",
          3616 => x"57f9d93f",
          3617 => x"76f23874",
          3618 => x"81165653",
          3619 => x"727b27fb",
          3620 => x"8438a051",
          3621 => x"f9c63fef",
          3622 => x"39963d0d",
          3623 => x"04fd3d0d",
          3624 => x"863d7070",
          3625 => x"84055208",
          3626 => x"55527351",
          3627 => x"fae03f85",
          3628 => x"3d0d04fe",
          3629 => x"3d0d7481",
          3630 => x"d39c0c85",
          3631 => x"3d880552",
          3632 => x"7551faca",
          3633 => x"3f81d39c",
          3634 => x"08538073",
          3635 => x"34800b81",
          3636 => x"d39c0c84",
          3637 => x"3d0d04fd",
          3638 => x"3d0d81d3",
          3639 => x"94087681",
          3640 => x"d3940c87",
          3641 => x"3d880553",
          3642 => x"775253fa",
          3643 => x"a13f7281",
          3644 => x"d3940c85",
          3645 => x"3d0d04fb",
          3646 => x"3d0d7779",
          3647 => x"81d39808",
          3648 => x"70565457",
          3649 => x"55805471",
          3650 => x"802e80e0",
          3651 => x"3881d398",
          3652 => x"0852712d",
          3653 => x"81d38408",
          3654 => x"81ff0653",
          3655 => x"72802e80",
          3656 => x"cb38728d",
          3657 => x"2eb93872",
          3658 => x"88327030",
          3659 => x"70802551",
          3660 => x"51527380",
          3661 => x"2e8b3871",
          3662 => x"802e8638",
          3663 => x"ff145497",
          3664 => x"399f7325",
          3665 => x"c838ff16",
          3666 => x"52737225",
          3667 => x"c0387414",
          3668 => x"52727234",
          3669 => x"81145472",
          3670 => x"51f8813f",
          3671 => x"ffaf3973",
          3672 => x"15528072",
          3673 => x"348a51f7",
          3674 => x"f33f8153",
          3675 => x"7281d384",
          3676 => x"0c873d0d",
          3677 => x"04fe3d0d",
          3678 => x"81d39808",
          3679 => x"7581d398",
          3680 => x"0c775376",
          3681 => x"5253feef",
          3682 => x"3f7281d3",
          3683 => x"980c843d",
          3684 => x"0d04f83d",
          3685 => x"0d7a7c5a",
          3686 => x"5680707a",
          3687 => x"0c587508",
          3688 => x"70335553",
          3689 => x"73a02e09",
          3690 => x"81068738",
          3691 => x"8113760c",
          3692 => x"ed3973ad",
          3693 => x"2e098106",
          3694 => x"8e388176",
          3695 => x"0811770c",
          3696 => x"76087033",
          3697 => x"56545873",
          3698 => x"b02e0981",
          3699 => x"0680c238",
          3700 => x"75088105",
          3701 => x"760c7508",
          3702 => x"70335553",
          3703 => x"7380e22e",
          3704 => x"8b389057",
          3705 => x"7380f82e",
          3706 => x"85388f39",
          3707 => x"82578113",
          3708 => x"760c7508",
          3709 => x"70335553",
          3710 => x"ac398155",
          3711 => x"a0742780",
          3712 => x"fa38d014",
          3713 => x"53805588",
          3714 => x"57897327",
          3715 => x"983880eb",
          3716 => x"39d01453",
          3717 => x"80557289",
          3718 => x"2680e038",
          3719 => x"86398055",
          3720 => x"80d9398a",
          3721 => x"578055a0",
          3722 => x"742780c2",
          3723 => x"3880e074",
          3724 => x"278938e0",
          3725 => x"147081ff",
          3726 => x"065553d0",
          3727 => x"147081ff",
          3728 => x"06555390",
          3729 => x"74278e38",
          3730 => x"f9147081",
          3731 => x"ff065553",
          3732 => x"897427ca",
          3733 => x"38737727",
          3734 => x"c5387477",
          3735 => x"29147608",
          3736 => x"8105770c",
          3737 => x"76087033",
          3738 => x"565455ff",
          3739 => x"ba397780",
          3740 => x"2e843874",
          3741 => x"30557479",
          3742 => x"0c815574",
          3743 => x"81d3840c",
          3744 => x"8a3d0d04",
          3745 => x"f83d0d7a",
          3746 => x"7c5a5680",
          3747 => x"707a0c58",
          3748 => x"75087033",
          3749 => x"555373a0",
          3750 => x"2e098106",
          3751 => x"87388113",
          3752 => x"760ced39",
          3753 => x"73ad2e09",
          3754 => x"81068e38",
          3755 => x"81760811",
          3756 => x"770c7608",
          3757 => x"70335654",
          3758 => x"5873b02e",
          3759 => x"09810680",
          3760 => x"c2387508",
          3761 => x"8105760c",
          3762 => x"75087033",
          3763 => x"55537380",
          3764 => x"e22e8b38",
          3765 => x"90577380",
          3766 => x"f82e8538",
          3767 => x"8f398257",
          3768 => x"8113760c",
          3769 => x"75087033",
          3770 => x"5553ac39",
          3771 => x"8155a074",
          3772 => x"2780fa38",
          3773 => x"d0145380",
          3774 => x"55885789",
          3775 => x"73279838",
          3776 => x"80eb39d0",
          3777 => x"14538055",
          3778 => x"72892680",
          3779 => x"e0388639",
          3780 => x"805580d9",
          3781 => x"398a5780",
          3782 => x"55a07427",
          3783 => x"80c23880",
          3784 => x"e0742789",
          3785 => x"38e01470",
          3786 => x"81ff0655",
          3787 => x"53d01470",
          3788 => x"81ff0655",
          3789 => x"53907427",
          3790 => x"8e38f914",
          3791 => x"7081ff06",
          3792 => x"55538974",
          3793 => x"27ca3873",
          3794 => x"7727c538",
          3795 => x"74772914",
          3796 => x"76088105",
          3797 => x"770c7608",
          3798 => x"70335654",
          3799 => x"55ffba39",
          3800 => x"77802e84",
          3801 => x"38743055",
          3802 => x"74790c81",
          3803 => x"557481d3",
          3804 => x"840c8a3d",
          3805 => x"0d04ff3d",
          3806 => x"0d028f05",
          3807 => x"33518152",
          3808 => x"70722687",
          3809 => x"3881d0c0",
          3810 => x"11335271",
          3811 => x"81d3840c",
          3812 => x"833d0d04",
          3813 => x"fc3d0d02",
          3814 => x"9b053302",
          3815 => x"84059f05",
          3816 => x"33565383",
          3817 => x"51728126",
          3818 => x"80e03872",
          3819 => x"842b87c0",
          3820 => x"928c1153",
          3821 => x"51885474",
          3822 => x"802e8438",
          3823 => x"81885473",
          3824 => x"720c87c0",
          3825 => x"928c1151",
          3826 => x"81710c85",
          3827 => x"0b87c098",
          3828 => x"8c0c7052",
          3829 => x"71087082",
          3830 => x"06515170",
          3831 => x"802e8a38",
          3832 => x"87c0988c",
          3833 => x"085170ec",
          3834 => x"387108fc",
          3835 => x"80800652",
          3836 => x"71923887",
          3837 => x"c0988c08",
          3838 => x"5170802e",
          3839 => x"87387181",
          3840 => x"d0c01434",
          3841 => x"81d0c013",
          3842 => x"33517081",
          3843 => x"d3840c86",
          3844 => x"3d0d04f3",
          3845 => x"3d0d6062",
          3846 => x"64028c05",
          3847 => x"bf053357",
          3848 => x"40585b83",
          3849 => x"74525afe",
          3850 => x"cd3f81d3",
          3851 => x"84088106",
          3852 => x"7a545271",
          3853 => x"81be3871",
          3854 => x"7275842b",
          3855 => x"87c09280",
          3856 => x"1187c092",
          3857 => x"8c1287c0",
          3858 => x"92841341",
          3859 => x"5a40575a",
          3860 => x"58850b87",
          3861 => x"c0988c0c",
          3862 => x"767d0c84",
          3863 => x"760c7508",
          3864 => x"70852a70",
          3865 => x"81065153",
          3866 => x"5471802e",
          3867 => x"8e387b08",
          3868 => x"52717b70",
          3869 => x"81055d34",
          3870 => x"81195980",
          3871 => x"74a20653",
          3872 => x"5371732e",
          3873 => x"83388153",
          3874 => x"7883ff26",
          3875 => x"8f387280",
          3876 => x"2e8a3887",
          3877 => x"c0988c08",
          3878 => x"5271c338",
          3879 => x"87c0988c",
          3880 => x"08527180",
          3881 => x"2e873878",
          3882 => x"84802e99",
          3883 => x"3881760c",
          3884 => x"87c0928c",
          3885 => x"15537208",
          3886 => x"70820651",
          3887 => x"5271f738",
          3888 => x"ff1a5a8d",
          3889 => x"39848017",
          3890 => x"81197081",
          3891 => x"ff065a53",
          3892 => x"5779802e",
          3893 => x"903873fc",
          3894 => x"80800652",
          3895 => x"7187387d",
          3896 => x"7826feed",
          3897 => x"3873fc80",
          3898 => x"80065271",
          3899 => x"802e8338",
          3900 => x"81527153",
          3901 => x"7281d384",
          3902 => x"0c8f3d0d",
          3903 => x"04f33d0d",
          3904 => x"60626402",
          3905 => x"8c05bf05",
          3906 => x"33574058",
          3907 => x"5b835980",
          3908 => x"745258fc",
          3909 => x"e13f81d3",
          3910 => x"84088106",
          3911 => x"79545271",
          3912 => x"782e0981",
          3913 => x"0681b138",
          3914 => x"7774842b",
          3915 => x"87c09280",
          3916 => x"1187c092",
          3917 => x"8c1287c0",
          3918 => x"92841340",
          3919 => x"595f565a",
          3920 => x"850b87c0",
          3921 => x"988c0c76",
          3922 => x"7d0c8276",
          3923 => x"0c805875",
          3924 => x"0870842a",
          3925 => x"70810651",
          3926 => x"53547180",
          3927 => x"2e8c387a",
          3928 => x"7081055c",
          3929 => x"337c0c81",
          3930 => x"18587381",
          3931 => x"2a708106",
          3932 => x"51527180",
          3933 => x"2e8a3887",
          3934 => x"c0988c08",
          3935 => x"5271d038",
          3936 => x"87c0988c",
          3937 => x"08527180",
          3938 => x"2e873877",
          3939 => x"84802e99",
          3940 => x"3881760c",
          3941 => x"87c0928c",
          3942 => x"15537208",
          3943 => x"70820651",
          3944 => x"5271f738",
          3945 => x"ff19598d",
          3946 => x"39811a70",
          3947 => x"81ff0684",
          3948 => x"8019595b",
          3949 => x"5278802e",
          3950 => x"903873fc",
          3951 => x"80800652",
          3952 => x"7187387d",
          3953 => x"7a26fef8",
          3954 => x"3873fc80",
          3955 => x"80065271",
          3956 => x"802e8338",
          3957 => x"81527153",
          3958 => x"7281d384",
          3959 => x"0c8f3d0d",
          3960 => x"04f63d0d",
          3961 => x"7e028405",
          3962 => x"b3053302",
          3963 => x"8805b705",
          3964 => x"33715454",
          3965 => x"5657fafe",
          3966 => x"3f81d384",
          3967 => x"08810653",
          3968 => x"83547280",
          3969 => x"fe38850b",
          3970 => x"87c0988c",
          3971 => x"0c815671",
          3972 => x"762e80dc",
          3973 => x"38717624",
          3974 => x"93387484",
          3975 => x"2b87c092",
          3976 => x"8c115454",
          3977 => x"71802e8d",
          3978 => x"3880d439",
          3979 => x"71832e80",
          3980 => x"c63880cb",
          3981 => x"39720870",
          3982 => x"812a7081",
          3983 => x"06515152",
          3984 => x"71802e8a",
          3985 => x"3887c098",
          3986 => x"8c085271",
          3987 => x"e83887c0",
          3988 => x"988c0852",
          3989 => x"71963881",
          3990 => x"730c87c0",
          3991 => x"928c1453",
          3992 => x"72087082",
          3993 => x"06515271",
          3994 => x"f7389639",
          3995 => x"80569239",
          3996 => x"88800a77",
          3997 => x"0c853981",
          3998 => x"80770c72",
          3999 => x"56833984",
          4000 => x"56755473",
          4001 => x"81d3840c",
          4002 => x"8c3d0d04",
          4003 => x"fe3d0d74",
          4004 => x"81113371",
          4005 => x"3371882b",
          4006 => x"0781d384",
          4007 => x"0c535184",
          4008 => x"3d0d04fd",
          4009 => x"3d0d7583",
          4010 => x"11338212",
          4011 => x"3371902b",
          4012 => x"71882b07",
          4013 => x"81143370",
          4014 => x"7207882b",
          4015 => x"75337107",
          4016 => x"81d3840c",
          4017 => x"52535456",
          4018 => x"5452853d",
          4019 => x"0d04ff3d",
          4020 => x"0d730284",
          4021 => x"05920522",
          4022 => x"52527072",
          4023 => x"70810554",
          4024 => x"3470882a",
          4025 => x"51707234",
          4026 => x"833d0d04",
          4027 => x"ff3d0d73",
          4028 => x"75525270",
          4029 => x"72708105",
          4030 => x"54347088",
          4031 => x"2a517072",
          4032 => x"70810554",
          4033 => x"3470882a",
          4034 => x"51707270",
          4035 => x"81055434",
          4036 => x"70882a51",
          4037 => x"70723483",
          4038 => x"3d0d04fe",
          4039 => x"3d0d7675",
          4040 => x"77545451",
          4041 => x"70802e92",
          4042 => x"38717081",
          4043 => x"05533373",
          4044 => x"70810555",
          4045 => x"34ff1151",
          4046 => x"eb39843d",
          4047 => x"0d04fe3d",
          4048 => x"0d757776",
          4049 => x"54525372",
          4050 => x"72708105",
          4051 => x"5434ff11",
          4052 => x"5170f438",
          4053 => x"843d0d04",
          4054 => x"fc3d0d78",
          4055 => x"77795656",
          4056 => x"53747081",
          4057 => x"05563374",
          4058 => x"70810556",
          4059 => x"33717131",
          4060 => x"ff165652",
          4061 => x"52527280",
          4062 => x"2e863871",
          4063 => x"802ee238",
          4064 => x"7181d384",
          4065 => x"0c863d0d",
          4066 => x"04fe3d0d",
          4067 => x"74765451",
          4068 => x"89397173",
          4069 => x"2e8a3881",
          4070 => x"11517033",
          4071 => x"5271f338",
          4072 => x"703381d3",
          4073 => x"840c843d",
          4074 => x"0d04800b",
          4075 => x"81d3840c",
          4076 => x"04800b81",
          4077 => x"d3840c04",
          4078 => x"f73d0d7b",
          4079 => x"56800b83",
          4080 => x"1733565a",
          4081 => x"747a2e80",
          4082 => x"d6388154",
          4083 => x"b0160853",
          4084 => x"b4167053",
          4085 => x"81173352",
          4086 => x"59faa23f",
          4087 => x"81d38408",
          4088 => x"7a2e0981",
          4089 => x"06b73881",
          4090 => x"d3840883",
          4091 => x"1734b016",
          4092 => x"0870a418",
          4093 => x"08319c18",
          4094 => x"08595658",
          4095 => x"7477279f",
          4096 => x"38821633",
          4097 => x"5574822e",
          4098 => x"09810693",
          4099 => x"38815476",
          4100 => x"18537852",
          4101 => x"81163351",
          4102 => x"f9e33f83",
          4103 => x"39815a79",
          4104 => x"81d3840c",
          4105 => x"8b3d0d04",
          4106 => x"fa3d0d78",
          4107 => x"7a565680",
          4108 => x"5774b017",
          4109 => x"082eaf38",
          4110 => x"7551fefc",
          4111 => x"3f81d384",
          4112 => x"085781d3",
          4113 => x"84089f38",
          4114 => x"81547453",
          4115 => x"b4165281",
          4116 => x"163351f7",
          4117 => x"be3f81d3",
          4118 => x"8408802e",
          4119 => x"8538ff55",
          4120 => x"815774b0",
          4121 => x"170c7681",
          4122 => x"d3840c88",
          4123 => x"3d0d04f8",
          4124 => x"3d0d7a70",
          4125 => x"5257fec0",
          4126 => x"3f81d384",
          4127 => x"085881d3",
          4128 => x"84088191",
          4129 => x"38763355",
          4130 => x"74832e09",
          4131 => x"810680f0",
          4132 => x"38841733",
          4133 => x"5978812e",
          4134 => x"09810680",
          4135 => x"e3388480",
          4136 => x"5381d384",
          4137 => x"0852b417",
          4138 => x"705256fd",
          4139 => x"913f82d4",
          4140 => x"d55284b2",
          4141 => x"1751fc96",
          4142 => x"3f848b85",
          4143 => x"a4d25275",
          4144 => x"51fca93f",
          4145 => x"868a85e4",
          4146 => x"f2528498",
          4147 => x"1751fc9c",
          4148 => x"3f901708",
          4149 => x"52849c17",
          4150 => x"51fc913f",
          4151 => x"8c170852",
          4152 => x"84a01751",
          4153 => x"fc863fa0",
          4154 => x"17088105",
          4155 => x"70b0190c",
          4156 => x"79555375",
          4157 => x"52811733",
          4158 => x"51f8823f",
          4159 => x"77841834",
          4160 => x"80538052",
          4161 => x"81173351",
          4162 => x"f9d73f81",
          4163 => x"d3840880",
          4164 => x"2e833881",
          4165 => x"587781d3",
          4166 => x"840c8a3d",
          4167 => x"0d04fb3d",
          4168 => x"0d77fe1a",
          4169 => x"981208fe",
          4170 => x"05555654",
          4171 => x"80567473",
          4172 => x"278d388a",
          4173 => x"14227571",
          4174 => x"29ac1608",
          4175 => x"05575375",
          4176 => x"81d3840c",
          4177 => x"873d0d04",
          4178 => x"f93d0d7a",
          4179 => x"7a700856",
          4180 => x"54578177",
          4181 => x"2781df38",
          4182 => x"76981508",
          4183 => x"2781d738",
          4184 => x"ff743354",
          4185 => x"5872822e",
          4186 => x"80f53872",
          4187 => x"82248938",
          4188 => x"72812e8d",
          4189 => x"3881bf39",
          4190 => x"72832e81",
          4191 => x"8e3881b6",
          4192 => x"3976812a",
          4193 => x"1770892a",
          4194 => x"a4160805",
          4195 => x"53745255",
          4196 => x"fd963f81",
          4197 => x"d3840881",
          4198 => x"9f387483",
          4199 => x"ff0614b4",
          4200 => x"11338117",
          4201 => x"70892aa4",
          4202 => x"18080555",
          4203 => x"76545757",
          4204 => x"53fcf53f",
          4205 => x"81d38408",
          4206 => x"80fe3874",
          4207 => x"83ff0614",
          4208 => x"b4113370",
          4209 => x"882b7807",
          4210 => x"79810671",
          4211 => x"842a5c52",
          4212 => x"58515372",
          4213 => x"80e23875",
          4214 => x"9fff0658",
          4215 => x"80da3976",
          4216 => x"882aa415",
          4217 => x"08055273",
          4218 => x"51fcbd3f",
          4219 => x"81d38408",
          4220 => x"80c63876",
          4221 => x"1083fe06",
          4222 => x"7405b405",
          4223 => x"51f98d3f",
          4224 => x"81d38408",
          4225 => x"83ffff06",
          4226 => x"58ae3976",
          4227 => x"872aa415",
          4228 => x"08055273",
          4229 => x"51fc913f",
          4230 => x"81d38408",
          4231 => x"9b387682",
          4232 => x"2b83fc06",
          4233 => x"7405b405",
          4234 => x"51f8f83f",
          4235 => x"81d38408",
          4236 => x"f00a0658",
          4237 => x"83398158",
          4238 => x"7781d384",
          4239 => x"0c893d0d",
          4240 => x"04f83d0d",
          4241 => x"7a7c7e5a",
          4242 => x"58568259",
          4243 => x"81772782",
          4244 => x"9e387698",
          4245 => x"17082782",
          4246 => x"96387533",
          4247 => x"5372792e",
          4248 => x"819d3872",
          4249 => x"79248938",
          4250 => x"72812e8d",
          4251 => x"38828039",
          4252 => x"72832e81",
          4253 => x"b83881f7",
          4254 => x"3976812a",
          4255 => x"1770892a",
          4256 => x"a4180805",
          4257 => x"53765255",
          4258 => x"fb9e3f81",
          4259 => x"d3840859",
          4260 => x"81d38408",
          4261 => x"81d93874",
          4262 => x"83ff0616",
          4263 => x"b4058116",
          4264 => x"78810659",
          4265 => x"56547753",
          4266 => x"76802e8f",
          4267 => x"3877842b",
          4268 => x"9ff00674",
          4269 => x"338f0671",
          4270 => x"07515372",
          4271 => x"7434810b",
          4272 => x"83173474",
          4273 => x"892aa417",
          4274 => x"08055275",
          4275 => x"51fad93f",
          4276 => x"81d38408",
          4277 => x"5981d384",
          4278 => x"08819438",
          4279 => x"7483ff06",
          4280 => x"16b40578",
          4281 => x"842a5454",
          4282 => x"768f3877",
          4283 => x"882a7433",
          4284 => x"81f00671",
          4285 => x"8f060751",
          4286 => x"53727434",
          4287 => x"80ec3976",
          4288 => x"882aa417",
          4289 => x"08055275",
          4290 => x"51fa9d3f",
          4291 => x"81d38408",
          4292 => x"5981d384",
          4293 => x"0880d838",
          4294 => x"7783ffff",
          4295 => x"06527610",
          4296 => x"83fe0676",
          4297 => x"05b40551",
          4298 => x"f7a43fbe",
          4299 => x"3976872a",
          4300 => x"a4170805",
          4301 => x"527551f9",
          4302 => x"ef3f81d3",
          4303 => x"84085981",
          4304 => x"d38408ab",
          4305 => x"3877f00a",
          4306 => x"0677822b",
          4307 => x"83fc0670",
          4308 => x"18b40570",
          4309 => x"54515454",
          4310 => x"f6c93f81",
          4311 => x"d384088f",
          4312 => x"0a067407",
          4313 => x"527251f7",
          4314 => x"833f810b",
          4315 => x"83173478",
          4316 => x"81d3840c",
          4317 => x"8a3d0d04",
          4318 => x"f83d0d7a",
          4319 => x"7c7e7208",
          4320 => x"59565659",
          4321 => x"817527a4",
          4322 => x"38749817",
          4323 => x"08279d38",
          4324 => x"73802eaa",
          4325 => x"38ff5373",
          4326 => x"527551fd",
          4327 => x"a43f81d3",
          4328 => x"84085481",
          4329 => x"d3840880",
          4330 => x"f2389339",
          4331 => x"825480eb",
          4332 => x"39815480",
          4333 => x"e63981d3",
          4334 => x"84085480",
          4335 => x"de397452",
          4336 => x"7851fb84",
          4337 => x"3f81d384",
          4338 => x"085881d3",
          4339 => x"8408802e",
          4340 => x"80c73881",
          4341 => x"d3840881",
          4342 => x"2ed23881",
          4343 => x"d38408ff",
          4344 => x"2ecf3880",
          4345 => x"53745275",
          4346 => x"51fcd63f",
          4347 => x"81d38408",
          4348 => x"c5389816",
          4349 => x"08fe1190",
          4350 => x"18085755",
          4351 => x"57747427",
          4352 => x"90388115",
          4353 => x"90170c84",
          4354 => x"16338107",
          4355 => x"54738417",
          4356 => x"34775576",
          4357 => x"7826ffa6",
          4358 => x"38805473",
          4359 => x"81d3840c",
          4360 => x"8a3d0d04",
          4361 => x"f63d0d7c",
          4362 => x"7e710859",
          4363 => x"5b5b7995",
          4364 => x"388c1708",
          4365 => x"5877802e",
          4366 => x"88389817",
          4367 => x"087826b2",
          4368 => x"388158ae",
          4369 => x"3979527a",
          4370 => x"51f9fd3f",
          4371 => x"81557481",
          4372 => x"d3840827",
          4373 => x"82e03881",
          4374 => x"d3840855",
          4375 => x"81d38408",
          4376 => x"ff2e82d2",
          4377 => x"38981708",
          4378 => x"81d38408",
          4379 => x"2682c738",
          4380 => x"79589017",
          4381 => x"08705654",
          4382 => x"73802e82",
          4383 => x"b938777a",
          4384 => x"2e098106",
          4385 => x"80e23881",
          4386 => x"1a569817",
          4387 => x"08762683",
          4388 => x"38825675",
          4389 => x"527a51f9",
          4390 => x"af3f8059",
          4391 => x"81d38408",
          4392 => x"812e0981",
          4393 => x"06863881",
          4394 => x"d3840859",
          4395 => x"81d38408",
          4396 => x"09703070",
          4397 => x"72078025",
          4398 => x"707c0781",
          4399 => x"d3840854",
          4400 => x"51515555",
          4401 => x"7381ef38",
          4402 => x"81d38408",
          4403 => x"802e9538",
          4404 => x"8c170854",
          4405 => x"81742790",
          4406 => x"38739818",
          4407 => x"08278938",
          4408 => x"73588539",
          4409 => x"7580db38",
          4410 => x"77568116",
          4411 => x"56981708",
          4412 => x"76268938",
          4413 => x"82567578",
          4414 => x"2681ac38",
          4415 => x"75527a51",
          4416 => x"f8c63f81",
          4417 => x"d3840880",
          4418 => x"2eb83880",
          4419 => x"5981d384",
          4420 => x"08812e09",
          4421 => x"81068638",
          4422 => x"81d38408",
          4423 => x"5981d384",
          4424 => x"08097030",
          4425 => x"70720780",
          4426 => x"25707c07",
          4427 => x"51515555",
          4428 => x"7380f838",
          4429 => x"75782e09",
          4430 => x"8106ffae",
          4431 => x"38735580",
          4432 => x"f539ff53",
          4433 => x"75527651",
          4434 => x"f9f73f81",
          4435 => x"d3840881",
          4436 => x"d3840830",
          4437 => x"7081d384",
          4438 => x"08078025",
          4439 => x"51555579",
          4440 => x"802e9438",
          4441 => x"73802e8f",
          4442 => x"38755379",
          4443 => x"527651f9",
          4444 => x"d03f81d3",
          4445 => x"84085574",
          4446 => x"a538758c",
          4447 => x"180c9817",
          4448 => x"08fe0590",
          4449 => x"18085654",
          4450 => x"74742686",
          4451 => x"38ff1590",
          4452 => x"180c8417",
          4453 => x"33810754",
          4454 => x"73841834",
          4455 => x"9739ff56",
          4456 => x"74812e90",
          4457 => x"388c3980",
          4458 => x"558c3981",
          4459 => x"d3840855",
          4460 => x"85398156",
          4461 => x"75557481",
          4462 => x"d3840c8c",
          4463 => x"3d0d04f8",
          4464 => x"3d0d7a70",
          4465 => x"5255f3f0",
          4466 => x"3f81d384",
          4467 => x"08588156",
          4468 => x"81d38408",
          4469 => x"80d8387b",
          4470 => x"527451f6",
          4471 => x"c13f81d3",
          4472 => x"840881d3",
          4473 => x"8408b017",
          4474 => x"0c598480",
          4475 => x"537752b4",
          4476 => x"15705257",
          4477 => x"f2c83f77",
          4478 => x"56843981",
          4479 => x"16568a15",
          4480 => x"22587578",
          4481 => x"27973881",
          4482 => x"54751953",
          4483 => x"76528115",
          4484 => x"3351ede9",
          4485 => x"3f81d384",
          4486 => x"08802edf",
          4487 => x"388a1522",
          4488 => x"76327030",
          4489 => x"70720770",
          4490 => x"9f2a5351",
          4491 => x"56567581",
          4492 => x"d3840c8a",
          4493 => x"3d0d04f8",
          4494 => x"3d0d7a7c",
          4495 => x"71085856",
          4496 => x"5774f080",
          4497 => x"0a2680f1",
          4498 => x"38749f06",
          4499 => x"537280e9",
          4500 => x"38749018",
          4501 => x"0c881708",
          4502 => x"5473aa38",
          4503 => x"75335382",
          4504 => x"73278838",
          4505 => x"a8160854",
          4506 => x"739b3874",
          4507 => x"852a5382",
          4508 => x"0b881722",
          4509 => x"5a587279",
          4510 => x"2780fe38",
          4511 => x"a8160898",
          4512 => x"180c80cd",
          4513 => x"398a1622",
          4514 => x"70892b54",
          4515 => x"58727526",
          4516 => x"b2387352",
          4517 => x"7651f5b0",
          4518 => x"3f81d384",
          4519 => x"085481d3",
          4520 => x"8408ff2e",
          4521 => x"bd38810b",
          4522 => x"81d38408",
          4523 => x"278b3898",
          4524 => x"160881d3",
          4525 => x"84082685",
          4526 => x"388258bd",
          4527 => x"39747331",
          4528 => x"55cb3973",
          4529 => x"527551f4",
          4530 => x"d53f81d3",
          4531 => x"84089818",
          4532 => x"0c739418",
          4533 => x"0c981708",
          4534 => x"53825872",
          4535 => x"802e9a38",
          4536 => x"85398158",
          4537 => x"94397489",
          4538 => x"2a139818",
          4539 => x"0c7483ff",
          4540 => x"0616b405",
          4541 => x"9c180c80",
          4542 => x"587781d3",
          4543 => x"840c8a3d",
          4544 => x"0d04f83d",
          4545 => x"0d7a7008",
          4546 => x"901208a0",
          4547 => x"05595754",
          4548 => x"f0800a77",
          4549 => x"27863880",
          4550 => x"0b98150c",
          4551 => x"98140853",
          4552 => x"84557280",
          4553 => x"2e81cb38",
          4554 => x"7683ff06",
          4555 => x"587781b5",
          4556 => x"38811398",
          4557 => x"150c9414",
          4558 => x"08557492",
          4559 => x"3876852a",
          4560 => x"88172256",
          4561 => x"53747326",
          4562 => x"819b3880",
          4563 => x"c0398a16",
          4564 => x"22ff0577",
          4565 => x"892a0653",
          4566 => x"72818a38",
          4567 => x"74527351",
          4568 => x"f3e63f81",
          4569 => x"d3840853",
          4570 => x"8255810b",
          4571 => x"81d38408",
          4572 => x"2780ff38",
          4573 => x"815581d3",
          4574 => x"8408ff2e",
          4575 => x"80f43898",
          4576 => x"160881d3",
          4577 => x"84082680",
          4578 => x"ca387b8a",
          4579 => x"38779815",
          4580 => x"0c845580",
          4581 => x"dd399414",
          4582 => x"08527351",
          4583 => x"f9863f81",
          4584 => x"d3840853",
          4585 => x"875581d3",
          4586 => x"8408802e",
          4587 => x"80c43882",
          4588 => x"5581d384",
          4589 => x"08812eba",
          4590 => x"38815581",
          4591 => x"d38408ff",
          4592 => x"2eb03881",
          4593 => x"d3840852",
          4594 => x"7551fbf3",
          4595 => x"3f81d384",
          4596 => x"08a03872",
          4597 => x"94150c72",
          4598 => x"527551f2",
          4599 => x"c13f81d3",
          4600 => x"84089815",
          4601 => x"0c769015",
          4602 => x"0c7716b4",
          4603 => x"059c150c",
          4604 => x"80557481",
          4605 => x"d3840c8a",
          4606 => x"3d0d04f7",
          4607 => x"3d0d7b7d",
          4608 => x"71085b5b",
          4609 => x"57805276",
          4610 => x"51fcac3f",
          4611 => x"81d38408",
          4612 => x"5481d384",
          4613 => x"0880ec38",
          4614 => x"81d38408",
          4615 => x"56981708",
          4616 => x"527851f0",
          4617 => x"833f81d3",
          4618 => x"84085481",
          4619 => x"d3840880",
          4620 => x"d23881d3",
          4621 => x"84089c18",
          4622 => x"08703351",
          4623 => x"54587281",
          4624 => x"e52e0981",
          4625 => x"06833881",
          4626 => x"5881d384",
          4627 => x"08557283",
          4628 => x"38815577",
          4629 => x"75075372",
          4630 => x"802e8e38",
          4631 => x"81165675",
          4632 => x"7a2e0981",
          4633 => x"068838a5",
          4634 => x"3981d384",
          4635 => x"08568152",
          4636 => x"7651fd8e",
          4637 => x"3f81d384",
          4638 => x"085481d3",
          4639 => x"8408802e",
          4640 => x"ff9b3873",
          4641 => x"842e0981",
          4642 => x"06833887",
          4643 => x"547381d3",
          4644 => x"840c8b3d",
          4645 => x"0d04fd3d",
          4646 => x"0d769a11",
          4647 => x"5254ebec",
          4648 => x"3f81d384",
          4649 => x"0883ffff",
          4650 => x"06767033",
          4651 => x"51535371",
          4652 => x"832e0981",
          4653 => x"06903894",
          4654 => x"1451ebd0",
          4655 => x"3f81d384",
          4656 => x"08902b73",
          4657 => x"07537281",
          4658 => x"d3840c85",
          4659 => x"3d0d04fc",
          4660 => x"3d0d7779",
          4661 => x"7083ffff",
          4662 => x"06549a12",
          4663 => x"535555eb",
          4664 => x"ed3f7670",
          4665 => x"33515372",
          4666 => x"832e0981",
          4667 => x"068b3873",
          4668 => x"902a5294",
          4669 => x"1551ebd6",
          4670 => x"3f863d0d",
          4671 => x"04f73d0d",
          4672 => x"7b7d5b55",
          4673 => x"8475085a",
          4674 => x"58981508",
          4675 => x"802e818a",
          4676 => x"38981508",
          4677 => x"527851ee",
          4678 => x"8f3f81d3",
          4679 => x"84085881",
          4680 => x"d3840880",
          4681 => x"f5389c15",
          4682 => x"08703355",
          4683 => x"53738638",
          4684 => x"845880e6",
          4685 => x"398b1333",
          4686 => x"70bf0670",
          4687 => x"81ff0658",
          4688 => x"51537286",
          4689 => x"163481d3",
          4690 => x"84085373",
          4691 => x"81e52e83",
          4692 => x"38815373",
          4693 => x"ae2ea938",
          4694 => x"81707406",
          4695 => x"54577280",
          4696 => x"2e9e3875",
          4697 => x"8f2e9938",
          4698 => x"81d38408",
          4699 => x"76df0654",
          4700 => x"5472882e",
          4701 => x"09810683",
          4702 => x"38765473",
          4703 => x"7a2ea038",
          4704 => x"80527451",
          4705 => x"fafc3f81",
          4706 => x"d3840858",
          4707 => x"81d38408",
          4708 => x"89389815",
          4709 => x"08fefa38",
          4710 => x"8639800b",
          4711 => x"98160c77",
          4712 => x"81d3840c",
          4713 => x"8b3d0d04",
          4714 => x"fb3d0d77",
          4715 => x"70085754",
          4716 => x"81527351",
          4717 => x"fcc53f81",
          4718 => x"d3840855",
          4719 => x"81d38408",
          4720 => x"b4389814",
          4721 => x"08527551",
          4722 => x"ecde3f81",
          4723 => x"d3840855",
          4724 => x"81d38408",
          4725 => x"a038a053",
          4726 => x"81d38408",
          4727 => x"529c1408",
          4728 => x"51eadb3f",
          4729 => x"8b53a014",
          4730 => x"529c1408",
          4731 => x"51eaac3f",
          4732 => x"810b8317",
          4733 => x"347481d3",
          4734 => x"840c873d",
          4735 => x"0d04fd3d",
          4736 => x"0d757008",
          4737 => x"98120854",
          4738 => x"70535553",
          4739 => x"ec9a3f81",
          4740 => x"d384088d",
          4741 => x"389c1308",
          4742 => x"53e57334",
          4743 => x"810b8315",
          4744 => x"34853d0d",
          4745 => x"04fa3d0d",
          4746 => x"787a5757",
          4747 => x"800b8917",
          4748 => x"34981708",
          4749 => x"802e8182",
          4750 => x"38807089",
          4751 => x"18555555",
          4752 => x"9c170814",
          4753 => x"70338116",
          4754 => x"56515271",
          4755 => x"a02ea838",
          4756 => x"71852e09",
          4757 => x"81068438",
          4758 => x"81e55273",
          4759 => x"892e0981",
          4760 => x"068b38ae",
          4761 => x"73708105",
          4762 => x"55348115",
          4763 => x"55717370",
          4764 => x"81055534",
          4765 => x"8115558a",
          4766 => x"7427c538",
          4767 => x"75158805",
          4768 => x"52800b81",
          4769 => x"13349c17",
          4770 => x"08528b12",
          4771 => x"33881734",
          4772 => x"9c17089c",
          4773 => x"115252e8",
          4774 => x"8a3f81d3",
          4775 => x"8408760c",
          4776 => x"961251e7",
          4777 => x"e73f81d3",
          4778 => x"84088617",
          4779 => x"23981251",
          4780 => x"e7da3f81",
          4781 => x"d3840884",
          4782 => x"1723883d",
          4783 => x"0d04f33d",
          4784 => x"0d7f7008",
          4785 => x"5e5b8061",
          4786 => x"70335155",
          4787 => x"5573af2e",
          4788 => x"83388155",
          4789 => x"7380dc2e",
          4790 => x"91387480",
          4791 => x"2e8c3894",
          4792 => x"1d08881c",
          4793 => x"0caa3981",
          4794 => x"15418061",
          4795 => x"70335656",
          4796 => x"5673af2e",
          4797 => x"09810683",
          4798 => x"38815673",
          4799 => x"80dc3270",
          4800 => x"30708025",
          4801 => x"78075151",
          4802 => x"5473dc38",
          4803 => x"73881c0c",
          4804 => x"60703351",
          4805 => x"54739f26",
          4806 => x"9638ff80",
          4807 => x"0bab1c34",
          4808 => x"80527a51",
          4809 => x"f6913f81",
          4810 => x"d3840855",
          4811 => x"85983991",
          4812 => x"3d61a01d",
          4813 => x"5c5a5e8b",
          4814 => x"53a05279",
          4815 => x"51e7ff3f",
          4816 => x"80705957",
          4817 => x"88793355",
          4818 => x"5c73ae2e",
          4819 => x"09810680",
          4820 => x"d4387818",
          4821 => x"7033811a",
          4822 => x"71ae3270",
          4823 => x"30709f2a",
          4824 => x"73822607",
          4825 => x"5151535a",
          4826 => x"5754738c",
          4827 => x"38791754",
          4828 => x"75743481",
          4829 => x"1757db39",
          4830 => x"75af3270",
          4831 => x"30709f2a",
          4832 => x"51515475",
          4833 => x"80dc2e8c",
          4834 => x"3873802e",
          4835 => x"873875a0",
          4836 => x"2682bd38",
          4837 => x"77197e0c",
          4838 => x"a454a076",
          4839 => x"2782bd38",
          4840 => x"a05482b8",
          4841 => x"39781870",
          4842 => x"33811a5a",
          4843 => x"5754a076",
          4844 => x"2781fc38",
          4845 => x"75af3270",
          4846 => x"307780dc",
          4847 => x"32703072",
          4848 => x"80257180",
          4849 => x"25075151",
          4850 => x"56515573",
          4851 => x"802eac38",
          4852 => x"84398118",
          4853 => x"5880781a",
          4854 => x"70335155",
          4855 => x"5573af2e",
          4856 => x"09810683",
          4857 => x"38815573",
          4858 => x"80dc3270",
          4859 => x"30708025",
          4860 => x"77075151",
          4861 => x"5473db38",
          4862 => x"81b53975",
          4863 => x"ae2e0981",
          4864 => x"06833881",
          4865 => x"54767c27",
          4866 => x"74075473",
          4867 => x"802ea238",
          4868 => x"7b8b3270",
          4869 => x"3077ae32",
          4870 => x"70307280",
          4871 => x"25719f2a",
          4872 => x"07535156",
          4873 => x"51557481",
          4874 => x"a7388857",
          4875 => x"8b5cfef5",
          4876 => x"3975982b",
          4877 => x"54738025",
          4878 => x"8c387580",
          4879 => x"ff0681c2",
          4880 => x"f8113357",
          4881 => x"547551e6",
          4882 => x"e13f81d3",
          4883 => x"8408802e",
          4884 => x"b2387818",
          4885 => x"7033811a",
          4886 => x"71545a56",
          4887 => x"54e6d23f",
          4888 => x"81d38408",
          4889 => x"802e80e8",
          4890 => x"38ff1c54",
          4891 => x"76742780",
          4892 => x"df387917",
          4893 => x"54757434",
          4894 => x"81177a11",
          4895 => x"55577474",
          4896 => x"34a73975",
          4897 => x"5281c298",
          4898 => x"51e5fe3f",
          4899 => x"81d38408",
          4900 => x"bf38ff9f",
          4901 => x"16547399",
          4902 => x"268938e0",
          4903 => x"167081ff",
          4904 => x"06575479",
          4905 => x"17547574",
          4906 => x"34811757",
          4907 => x"fdf73977",
          4908 => x"197e0c76",
          4909 => x"802e9938",
          4910 => x"79335473",
          4911 => x"81e52e09",
          4912 => x"81068438",
          4913 => x"857a3484",
          4914 => x"54a07627",
          4915 => x"8f388b39",
          4916 => x"865581f2",
          4917 => x"39845680",
          4918 => x"f3398054",
          4919 => x"738b1b34",
          4920 => x"807b0858",
          4921 => x"527a51f2",
          4922 => x"ce3f81d3",
          4923 => x"84085681",
          4924 => x"d3840880",
          4925 => x"d738981b",
          4926 => x"08527651",
          4927 => x"e6aa3f81",
          4928 => x"d3840856",
          4929 => x"81d38408",
          4930 => x"80c2389c",
          4931 => x"1b087033",
          4932 => x"55557380",
          4933 => x"2effbe38",
          4934 => x"8b1533bf",
          4935 => x"06547386",
          4936 => x"1c348b15",
          4937 => x"3370832a",
          4938 => x"70810651",
          4939 => x"55587392",
          4940 => x"388b5379",
          4941 => x"527451e4",
          4942 => x"9f3f81d3",
          4943 => x"8408802e",
          4944 => x"8b387552",
          4945 => x"7a51f3ba",
          4946 => x"3fff9f39",
          4947 => x"75ab1c33",
          4948 => x"57557480",
          4949 => x"2ebb3874",
          4950 => x"842e0981",
          4951 => x"0680e738",
          4952 => x"75852a70",
          4953 => x"81067782",
          4954 => x"2a585154",
          4955 => x"73802e96",
          4956 => x"38758106",
          4957 => x"5473802e",
          4958 => x"fbb538ff",
          4959 => x"800bab1c",
          4960 => x"34805580",
          4961 => x"c1397581",
          4962 => x"065473ba",
          4963 => x"388555b6",
          4964 => x"3975822a",
          4965 => x"70810651",
          4966 => x"5473ab38",
          4967 => x"861b3370",
          4968 => x"842a7081",
          4969 => x"06515555",
          4970 => x"73802ee1",
          4971 => x"38901b08",
          4972 => x"83ff061d",
          4973 => x"b405527c",
          4974 => x"51f5db3f",
          4975 => x"81d38408",
          4976 => x"881c0cfa",
          4977 => x"ea397481",
          4978 => x"d3840c8f",
          4979 => x"3d0d04f6",
          4980 => x"3d0d7c5b",
          4981 => x"ff7b0870",
          4982 => x"71735559",
          4983 => x"5c555973",
          4984 => x"802e81c6",
          4985 => x"38757081",
          4986 => x"05573370",
          4987 => x"a0265252",
          4988 => x"71ba2e8d",
          4989 => x"3870ee38",
          4990 => x"71ba2e09",
          4991 => x"810681a5",
          4992 => x"387333d0",
          4993 => x"117081ff",
          4994 => x"06515253",
          4995 => x"70892691",
          4996 => x"38821473",
          4997 => x"81ff06d0",
          4998 => x"05565271",
          4999 => x"762e80f7",
          5000 => x"38800b81",
          5001 => x"c2e85955",
          5002 => x"77087a55",
          5003 => x"57767081",
          5004 => x"05583374",
          5005 => x"70810556",
          5006 => x"33ff9f12",
          5007 => x"53535370",
          5008 => x"99268938",
          5009 => x"e0137081",
          5010 => x"ff065451",
          5011 => x"ff9f1251",
          5012 => x"70992689",
          5013 => x"38e01270",
          5014 => x"81ff0653",
          5015 => x"51723070",
          5016 => x"9f2a5151",
          5017 => x"72722e09",
          5018 => x"81068538",
          5019 => x"70ffbe38",
          5020 => x"72307477",
          5021 => x"32703070",
          5022 => x"72079f2a",
          5023 => x"739f2a07",
          5024 => x"53545451",
          5025 => x"70802e8f",
          5026 => x"38811584",
          5027 => x"19595583",
          5028 => x"7525ff94",
          5029 => x"388b3974",
          5030 => x"83248638",
          5031 => x"74767c0c",
          5032 => x"59785186",
          5033 => x"3981d3b4",
          5034 => x"33517081",
          5035 => x"d3840c8c",
          5036 => x"3d0d04fa",
          5037 => x"3d0d7856",
          5038 => x"800b8317",
          5039 => x"34ff0bb0",
          5040 => x"170c7952",
          5041 => x"7551e2e0",
          5042 => x"3f845581",
          5043 => x"d3840881",
          5044 => x"803884b2",
          5045 => x"1651dfb4",
          5046 => x"3f81d384",
          5047 => x"0883ffff",
          5048 => x"06548355",
          5049 => x"7382d4d5",
          5050 => x"2e098106",
          5051 => x"80e33880",
          5052 => x"0bb41733",
          5053 => x"56577481",
          5054 => x"e92e0981",
          5055 => x"06833881",
          5056 => x"577481eb",
          5057 => x"32703070",
          5058 => x"80257907",
          5059 => x"51515473",
          5060 => x"8a387481",
          5061 => x"e82e0981",
          5062 => x"06b53883",
          5063 => x"5381c2a8",
          5064 => x"5280ea16",
          5065 => x"51e0b13f",
          5066 => x"81d38408",
          5067 => x"5581d384",
          5068 => x"08802e9d",
          5069 => x"38855381",
          5070 => x"c2ac5281",
          5071 => x"861651e0",
          5072 => x"973f81d3",
          5073 => x"84085581",
          5074 => x"d3840880",
          5075 => x"2e833882",
          5076 => x"557481d3",
          5077 => x"840c883d",
          5078 => x"0d04f23d",
          5079 => x"0d610284",
          5080 => x"0580cb05",
          5081 => x"33585580",
          5082 => x"750c6051",
          5083 => x"fce13f81",
          5084 => x"d3840858",
          5085 => x"8b56800b",
          5086 => x"81d38408",
          5087 => x"2486fc38",
          5088 => x"81d38408",
          5089 => x"842981d3",
          5090 => x"a0057008",
          5091 => x"55538c56",
          5092 => x"73802e86",
          5093 => x"e6387375",
          5094 => x"0c7681fe",
          5095 => x"06743354",
          5096 => x"5772802e",
          5097 => x"ae388114",
          5098 => x"3351d7ca",
          5099 => x"3f81d384",
          5100 => x"0881ff06",
          5101 => x"70810654",
          5102 => x"55729838",
          5103 => x"76802e86",
          5104 => x"b8387482",
          5105 => x"2a708106",
          5106 => x"51538a56",
          5107 => x"7286ac38",
          5108 => x"86a73980",
          5109 => x"74347781",
          5110 => x"15348152",
          5111 => x"81143351",
          5112 => x"d7b23f81",
          5113 => x"d3840881",
          5114 => x"ff067081",
          5115 => x"06545583",
          5116 => x"56728687",
          5117 => x"3876802e",
          5118 => x"8f387482",
          5119 => x"2a708106",
          5120 => x"51538a56",
          5121 => x"7285f438",
          5122 => x"80705374",
          5123 => x"525bfda3",
          5124 => x"3f81d384",
          5125 => x"0881ff06",
          5126 => x"5776822e",
          5127 => x"09810680",
          5128 => x"e2388c3d",
          5129 => x"74565883",
          5130 => x"5683f615",
          5131 => x"33705853",
          5132 => x"72802e8d",
          5133 => x"3883fa15",
          5134 => x"51dce83f",
          5135 => x"81d38408",
          5136 => x"57767870",
          5137 => x"84055a0c",
          5138 => x"ff169016",
          5139 => x"56567580",
          5140 => x"25d73880",
          5141 => x"0b8d3d54",
          5142 => x"56727084",
          5143 => x"0554085b",
          5144 => x"83577a80",
          5145 => x"2e95387a",
          5146 => x"527351fc",
          5147 => x"c63f81d3",
          5148 => x"840881ff",
          5149 => x"06578177",
          5150 => x"27893881",
          5151 => x"16568376",
          5152 => x"27d73881",
          5153 => x"5676842e",
          5154 => x"84f1388d",
          5155 => x"56768126",
          5156 => x"84e938bf",
          5157 => x"1451dbf4",
          5158 => x"3f81d384",
          5159 => x"0883ffff",
          5160 => x"06537284",
          5161 => x"802e0981",
          5162 => x"0684d038",
          5163 => x"80ca1451",
          5164 => x"dbda3f81",
          5165 => x"d3840883",
          5166 => x"ffff0658",
          5167 => x"778d3880",
          5168 => x"d81451db",
          5169 => x"de3f81d3",
          5170 => x"84085877",
          5171 => x"9c150c80",
          5172 => x"c4143382",
          5173 => x"153480c4",
          5174 => x"1433ff11",
          5175 => x"7081ff06",
          5176 => x"5154558d",
          5177 => x"56728126",
          5178 => x"84913874",
          5179 => x"81ff0678",
          5180 => x"712980c1",
          5181 => x"16335259",
          5182 => x"53728a15",
          5183 => x"2372802e",
          5184 => x"8b38ff13",
          5185 => x"73065372",
          5186 => x"802e8638",
          5187 => x"8d5683eb",
          5188 => x"3980c514",
          5189 => x"51daf53f",
          5190 => x"81d38408",
          5191 => x"5381d384",
          5192 => x"08881523",
          5193 => x"728f0657",
          5194 => x"8d567683",
          5195 => x"ce3880c7",
          5196 => x"1451dad8",
          5197 => x"3f81d384",
          5198 => x"0883ffff",
          5199 => x"0655748d",
          5200 => x"3880d414",
          5201 => x"51dadc3f",
          5202 => x"81d38408",
          5203 => x"5580c214",
          5204 => x"51dab93f",
          5205 => x"81d38408",
          5206 => x"83ffff06",
          5207 => x"538d5672",
          5208 => x"802e8397",
          5209 => x"38881422",
          5210 => x"78147184",
          5211 => x"2a055a5a",
          5212 => x"78752683",
          5213 => x"86388a14",
          5214 => x"22527479",
          5215 => x"3151ffaf",
          5216 => x"f63f81d3",
          5217 => x"84085581",
          5218 => x"d3840880",
          5219 => x"2e82ec38",
          5220 => x"81d38408",
          5221 => x"80ffffff",
          5222 => x"f5268338",
          5223 => x"83577483",
          5224 => x"fff52683",
          5225 => x"38825774",
          5226 => x"9ff52685",
          5227 => x"38815789",
          5228 => x"398d5676",
          5229 => x"802e82c3",
          5230 => x"38821570",
          5231 => x"98160c7b",
          5232 => x"a0160c73",
          5233 => x"1c70a417",
          5234 => x"0c7a1dac",
          5235 => x"170c5455",
          5236 => x"76832e09",
          5237 => x"8106af38",
          5238 => x"80de1451",
          5239 => x"d9ae3f81",
          5240 => x"d3840883",
          5241 => x"ffff0653",
          5242 => x"8d567282",
          5243 => x"8e387982",
          5244 => x"8a3880e0",
          5245 => x"1451d9ab",
          5246 => x"3f81d384",
          5247 => x"08a8150c",
          5248 => x"74822b53",
          5249 => x"a2398d56",
          5250 => x"79802e81",
          5251 => x"ee387713",
          5252 => x"a8150c74",
          5253 => x"15537682",
          5254 => x"2e8d3874",
          5255 => x"10157081",
          5256 => x"2a768106",
          5257 => x"05515383",
          5258 => x"ff13892a",
          5259 => x"538d5672",
          5260 => x"9c150826",
          5261 => x"81c538ff",
          5262 => x"0b90150c",
          5263 => x"ff0b8c15",
          5264 => x"0cff800b",
          5265 => x"84153476",
          5266 => x"832e0981",
          5267 => x"06819238",
          5268 => x"80e41451",
          5269 => x"d8b63f81",
          5270 => x"d3840883",
          5271 => x"ffff0653",
          5272 => x"72812e09",
          5273 => x"810680f9",
          5274 => x"38811b52",
          5275 => x"7351dbb8",
          5276 => x"3f81d384",
          5277 => x"0880ea38",
          5278 => x"81d38408",
          5279 => x"84153484",
          5280 => x"b21451d8",
          5281 => x"873f81d3",
          5282 => x"840883ff",
          5283 => x"ff065372",
          5284 => x"82d4d52e",
          5285 => x"09810680",
          5286 => x"c838b414",
          5287 => x"51d8843f",
          5288 => x"81d38408",
          5289 => x"848b85a4",
          5290 => x"d22e0981",
          5291 => x"06b33884",
          5292 => x"981451d7",
          5293 => x"ee3f81d3",
          5294 => x"8408868a",
          5295 => x"85e4f22e",
          5296 => x"0981069d",
          5297 => x"38849c14",
          5298 => x"51d7d83f",
          5299 => x"81d38408",
          5300 => x"90150c84",
          5301 => x"a01451d7",
          5302 => x"ca3f81d3",
          5303 => x"84088c15",
          5304 => x"0c767434",
          5305 => x"81d3b022",
          5306 => x"81055372",
          5307 => x"81d3b023",
          5308 => x"72861523",
          5309 => x"800b9415",
          5310 => x"0c805675",
          5311 => x"81d3840c",
          5312 => x"903d0d04",
          5313 => x"fb3d0d77",
          5314 => x"54895573",
          5315 => x"802eb938",
          5316 => x"73085372",
          5317 => x"802eb138",
          5318 => x"72335271",
          5319 => x"802ea938",
          5320 => x"86132284",
          5321 => x"15225752",
          5322 => x"71762e09",
          5323 => x"81069938",
          5324 => x"81133351",
          5325 => x"d0c03f81",
          5326 => x"d3840881",
          5327 => x"06527188",
          5328 => x"38717408",
          5329 => x"54558339",
          5330 => x"80537873",
          5331 => x"710c5274",
          5332 => x"81d3840c",
          5333 => x"873d0d04",
          5334 => x"fa3d0d02",
          5335 => x"ab05337a",
          5336 => x"58893dfc",
          5337 => x"055256f4",
          5338 => x"e63f8b54",
          5339 => x"800b81d3",
          5340 => x"840824bc",
          5341 => x"3881d384",
          5342 => x"08842981",
          5343 => x"d3a00570",
          5344 => x"08555573",
          5345 => x"802e8438",
          5346 => x"80743478",
          5347 => x"5473802e",
          5348 => x"84388074",
          5349 => x"3478750c",
          5350 => x"75547580",
          5351 => x"2e923880",
          5352 => x"53893d70",
          5353 => x"53840551",
          5354 => x"f7b03f81",
          5355 => x"d3840854",
          5356 => x"7381d384",
          5357 => x"0c883d0d",
          5358 => x"04eb3d0d",
          5359 => x"67028405",
          5360 => x"80e70533",
          5361 => x"59598954",
          5362 => x"78802e84",
          5363 => x"c83877bf",
          5364 => x"06705498",
          5365 => x"3dd00553",
          5366 => x"993d8405",
          5367 => x"5258f6fa",
          5368 => x"3f81d384",
          5369 => x"085581d3",
          5370 => x"840884a4",
          5371 => x"387a5c68",
          5372 => x"528c3d70",
          5373 => x"5256edc6",
          5374 => x"3f81d384",
          5375 => x"085581d3",
          5376 => x"84089238",
          5377 => x"0280d705",
          5378 => x"3370982b",
          5379 => x"55577380",
          5380 => x"25833886",
          5381 => x"55779c06",
          5382 => x"5473802e",
          5383 => x"81ab3874",
          5384 => x"802e9538",
          5385 => x"74842e09",
          5386 => x"8106aa38",
          5387 => x"7551eaf8",
          5388 => x"3f81d384",
          5389 => x"08559e39",
          5390 => x"02b20533",
          5391 => x"91065473",
          5392 => x"81b83877",
          5393 => x"822a7081",
          5394 => x"06515473",
          5395 => x"802e8e38",
          5396 => x"885583bc",
          5397 => x"39778807",
          5398 => x"587483b4",
          5399 => x"3877832a",
          5400 => x"70810651",
          5401 => x"5473802e",
          5402 => x"81af3862",
          5403 => x"527a51e8",
          5404 => x"a53f81d3",
          5405 => x"84085682",
          5406 => x"88b20a52",
          5407 => x"628e0551",
          5408 => x"d4ea3f62",
          5409 => x"54a00b8b",
          5410 => x"15348053",
          5411 => x"62527a51",
          5412 => x"e8bd3f80",
          5413 => x"52629c05",
          5414 => x"51d4d13f",
          5415 => x"7a54810b",
          5416 => x"83153475",
          5417 => x"802e80f1",
          5418 => x"387ab011",
          5419 => x"08515480",
          5420 => x"53755297",
          5421 => x"3dd40551",
          5422 => x"ddbe3f81",
          5423 => x"d3840855",
          5424 => x"81d38408",
          5425 => x"82ca38b7",
          5426 => x"397482c4",
          5427 => x"3802b205",
          5428 => x"3370842a",
          5429 => x"70810651",
          5430 => x"55567380",
          5431 => x"2e863884",
          5432 => x"5582ad39",
          5433 => x"77812a70",
          5434 => x"81065154",
          5435 => x"73802ea9",
          5436 => x"38758106",
          5437 => x"5473802e",
          5438 => x"a0388755",
          5439 => x"82923973",
          5440 => x"527a51d6",
          5441 => x"a33f81d3",
          5442 => x"84087bff",
          5443 => x"188c120c",
          5444 => x"555581d3",
          5445 => x"840881f8",
          5446 => x"3877832a",
          5447 => x"70810651",
          5448 => x"5473802e",
          5449 => x"86387780",
          5450 => x"c007587a",
          5451 => x"b01108a0",
          5452 => x"1b0c63a4",
          5453 => x"1b0c6353",
          5454 => x"705257e6",
          5455 => x"d93f81d3",
          5456 => x"840881d3",
          5457 => x"8408881b",
          5458 => x"0c639c05",
          5459 => x"525ad2d3",
          5460 => x"3f81d384",
          5461 => x"0881d384",
          5462 => x"088c1b0c",
          5463 => x"777a0c56",
          5464 => x"86172284",
          5465 => x"1a237790",
          5466 => x"1a34800b",
          5467 => x"911a3480",
          5468 => x"0b9c1a0c",
          5469 => x"800b941a",
          5470 => x"0c77852a",
          5471 => x"70810651",
          5472 => x"5473802e",
          5473 => x"818d3881",
          5474 => x"d3840880",
          5475 => x"2e818438",
          5476 => x"81d38408",
          5477 => x"941a0c8a",
          5478 => x"17227089",
          5479 => x"2b7b5259",
          5480 => x"57a83976",
          5481 => x"527851d7",
          5482 => x"9f3f81d3",
          5483 => x"84085781",
          5484 => x"d3840881",
          5485 => x"26833882",
          5486 => x"5581d384",
          5487 => x"08ff2e09",
          5488 => x"81068338",
          5489 => x"79557578",
          5490 => x"31567430",
          5491 => x"70760780",
          5492 => x"25515477",
          5493 => x"76278a38",
          5494 => x"81707506",
          5495 => x"555a73c3",
          5496 => x"3876981a",
          5497 => x"0c74a938",
          5498 => x"7583ff06",
          5499 => x"5473802e",
          5500 => x"a2387652",
          5501 => x"7a51d6a6",
          5502 => x"3f81d384",
          5503 => x"08853882",
          5504 => x"558e3975",
          5505 => x"892a81d3",
          5506 => x"8408059c",
          5507 => x"1a0c8439",
          5508 => x"80790c74",
          5509 => x"547381d3",
          5510 => x"840c973d",
          5511 => x"0d04f23d",
          5512 => x"0d606365",
          5513 => x"6440405d",
          5514 => x"59807e0c",
          5515 => x"903dfc05",
          5516 => x"527851f9",
          5517 => x"cf3f81d3",
          5518 => x"84085581",
          5519 => x"d384088a",
          5520 => x"38911933",
          5521 => x"5574802e",
          5522 => x"86387456",
          5523 => x"82c43990",
          5524 => x"19338106",
          5525 => x"55875674",
          5526 => x"802e82b6",
          5527 => x"38953982",
          5528 => x"0b911a34",
          5529 => x"825682aa",
          5530 => x"39810b91",
          5531 => x"1a348156",
          5532 => x"82a0398c",
          5533 => x"1908941a",
          5534 => x"08315574",
          5535 => x"7c278338",
          5536 => x"745c7b80",
          5537 => x"2e828938",
          5538 => x"94190870",
          5539 => x"83ff0656",
          5540 => x"567481b2",
          5541 => x"387e8a11",
          5542 => x"22ff0577",
          5543 => x"892a065b",
          5544 => x"5579a838",
          5545 => x"75873888",
          5546 => x"1908558f",
          5547 => x"39981908",
          5548 => x"527851d5",
          5549 => x"933f81d3",
          5550 => x"84085581",
          5551 => x"7527ff9f",
          5552 => x"3874ff2e",
          5553 => x"ffa33874",
          5554 => x"981a0c98",
          5555 => x"1908527e",
          5556 => x"51d4cb3f",
          5557 => x"81d38408",
          5558 => x"802eff83",
          5559 => x"3881d384",
          5560 => x"081a7c89",
          5561 => x"2a595777",
          5562 => x"802e80d6",
          5563 => x"38771a7f",
          5564 => x"8a112258",
          5565 => x"5c557575",
          5566 => x"27853875",
          5567 => x"7a315877",
          5568 => x"5476537c",
          5569 => x"52811b33",
          5570 => x"51ca883f",
          5571 => x"81d38408",
          5572 => x"fed7387e",
          5573 => x"83113356",
          5574 => x"5674802e",
          5575 => x"9f38b016",
          5576 => x"08773155",
          5577 => x"74782794",
          5578 => x"38848053",
          5579 => x"b41652b0",
          5580 => x"16087731",
          5581 => x"892b7d05",
          5582 => x"51cfe03f",
          5583 => x"77892b56",
          5584 => x"b939769c",
          5585 => x"1a0c9419",
          5586 => x"0883ff06",
          5587 => x"84807131",
          5588 => x"57557b76",
          5589 => x"2783387b",
          5590 => x"569c1908",
          5591 => x"527e51d1",
          5592 => x"c73f81d3",
          5593 => x"8408fe81",
          5594 => x"38755394",
          5595 => x"190883ff",
          5596 => x"061fb405",
          5597 => x"527c51cf",
          5598 => x"a23f7b76",
          5599 => x"317e0817",
          5600 => x"7f0c761e",
          5601 => x"941b0818",
          5602 => x"941c0c5e",
          5603 => x"5cfdf339",
          5604 => x"80567581",
          5605 => x"d3840c90",
          5606 => x"3d0d04f2",
          5607 => x"3d0d6063",
          5608 => x"65644040",
          5609 => x"5d58807e",
          5610 => x"0c903dfc",
          5611 => x"05527751",
          5612 => x"f6d23f81",
          5613 => x"d3840855",
          5614 => x"81d38408",
          5615 => x"8a389118",
          5616 => x"33557480",
          5617 => x"2e863874",
          5618 => x"5683b839",
          5619 => x"90183370",
          5620 => x"812a7081",
          5621 => x"06515656",
          5622 => x"87567480",
          5623 => x"2e83a438",
          5624 => x"9539820b",
          5625 => x"91193482",
          5626 => x"56839839",
          5627 => x"810b9119",
          5628 => x"34815683",
          5629 => x"8e399418",
          5630 => x"087c1156",
          5631 => x"56747627",
          5632 => x"84387509",
          5633 => x"5c7b802e",
          5634 => x"82ec3894",
          5635 => x"18087083",
          5636 => x"ff065656",
          5637 => x"7481fd38",
          5638 => x"7e8a1122",
          5639 => x"ff057789",
          5640 => x"2a065c55",
          5641 => x"7abf3875",
          5642 => x"8c388818",
          5643 => x"0855749c",
          5644 => x"387a5285",
          5645 => x"39981808",
          5646 => x"527751d7",
          5647 => x"e73f81d3",
          5648 => x"84085581",
          5649 => x"d3840880",
          5650 => x"2e82ab38",
          5651 => x"74812eff",
          5652 => x"913874ff",
          5653 => x"2eff9538",
          5654 => x"7498190c",
          5655 => x"88180885",
          5656 => x"38748819",
          5657 => x"0c7e55b0",
          5658 => x"15089c19",
          5659 => x"082e0981",
          5660 => x"068d3874",
          5661 => x"51cec13f",
          5662 => x"81d38408",
          5663 => x"feee3898",
          5664 => x"1808527e",
          5665 => x"51d1973f",
          5666 => x"81d38408",
          5667 => x"802efed2",
          5668 => x"3881d384",
          5669 => x"081b7c89",
          5670 => x"2a5a5778",
          5671 => x"802e80d5",
          5672 => x"38781b7f",
          5673 => x"8a112258",
          5674 => x"5b557575",
          5675 => x"27853875",
          5676 => x"7b315978",
          5677 => x"5476537c",
          5678 => x"52811a33",
          5679 => x"51c8be3f",
          5680 => x"81d38408",
          5681 => x"fea6387e",
          5682 => x"b0110878",
          5683 => x"31565674",
          5684 => x"79279b38",
          5685 => x"848053b0",
          5686 => x"16087731",
          5687 => x"892b7d05",
          5688 => x"52b41651",
          5689 => x"ccb53f7e",
          5690 => x"55800b83",
          5691 => x"16347889",
          5692 => x"2b5680db",
          5693 => x"398c1808",
          5694 => x"94190826",
          5695 => x"93387e51",
          5696 => x"cdb63f81",
          5697 => x"d38408fd",
          5698 => x"e3387e77",
          5699 => x"b0120c55",
          5700 => x"769c190c",
          5701 => x"94180883",
          5702 => x"ff068480",
          5703 => x"71315755",
          5704 => x"7b762783",
          5705 => x"387b569c",
          5706 => x"1808527e",
          5707 => x"51cdf93f",
          5708 => x"81d38408",
          5709 => x"fdb63875",
          5710 => x"537c5294",
          5711 => x"180883ff",
          5712 => x"061fb405",
          5713 => x"51cbd43f",
          5714 => x"7e55810b",
          5715 => x"8316347b",
          5716 => x"76317e08",
          5717 => x"177f0c76",
          5718 => x"1e941a08",
          5719 => x"1870941c",
          5720 => x"0c8c1b08",
          5721 => x"58585e5c",
          5722 => x"74762783",
          5723 => x"38755574",
          5724 => x"8c190cfd",
          5725 => x"90399018",
          5726 => x"3380c007",
          5727 => x"55749019",
          5728 => x"34805675",
          5729 => x"81d3840c",
          5730 => x"903d0d04",
          5731 => x"f83d0d7a",
          5732 => x"8b3dfc05",
          5733 => x"53705256",
          5734 => x"f2ea3f81",
          5735 => x"d3840857",
          5736 => x"81d38408",
          5737 => x"80fb3890",
          5738 => x"16337086",
          5739 => x"2a708106",
          5740 => x"51555573",
          5741 => x"802e80e9",
          5742 => x"38a01608",
          5743 => x"527851cc",
          5744 => x"e73f81d3",
          5745 => x"84085781",
          5746 => x"d3840880",
          5747 => x"d438a416",
          5748 => x"088b1133",
          5749 => x"a0075555",
          5750 => x"738b1634",
          5751 => x"88160853",
          5752 => x"74527508",
          5753 => x"51dde83f",
          5754 => x"8c160852",
          5755 => x"9c1551c9",
          5756 => x"fb3f8288",
          5757 => x"b20a5296",
          5758 => x"1551c9f0",
          5759 => x"3f765292",
          5760 => x"1551c9ca",
          5761 => x"3f785481",
          5762 => x"0b831534",
          5763 => x"7851ccdf",
          5764 => x"3f81d384",
          5765 => x"08901733",
          5766 => x"81bf0655",
          5767 => x"57739017",
          5768 => x"347681d3",
          5769 => x"840c8a3d",
          5770 => x"0d04fc3d",
          5771 => x"0d767052",
          5772 => x"54fed93f",
          5773 => x"81d38408",
          5774 => x"5381d384",
          5775 => x"089c3886",
          5776 => x"3dfc0552",
          5777 => x"7351f1bc",
          5778 => x"3f81d384",
          5779 => x"085381d3",
          5780 => x"84088738",
          5781 => x"81d38408",
          5782 => x"740c7281",
          5783 => x"d3840c86",
          5784 => x"3d0d04ff",
          5785 => x"3d0d843d",
          5786 => x"51e6e43f",
          5787 => x"8b52800b",
          5788 => x"81d38408",
          5789 => x"248b3881",
          5790 => x"d3840881",
          5791 => x"d3b43480",
          5792 => x"527181d3",
          5793 => x"840c833d",
          5794 => x"0d04ef3d",
          5795 => x"0d805393",
          5796 => x"3dd00552",
          5797 => x"943d51e9",
          5798 => x"c13f81d3",
          5799 => x"84085581",
          5800 => x"d3840880",
          5801 => x"e0387658",
          5802 => x"6352933d",
          5803 => x"d40551e0",
          5804 => x"8d3f81d3",
          5805 => x"84085581",
          5806 => x"d38408bc",
          5807 => x"380280c7",
          5808 => x"05337098",
          5809 => x"2b555673",
          5810 => x"80258938",
          5811 => x"767a9412",
          5812 => x"0c54b239",
          5813 => x"02a20533",
          5814 => x"70842a70",
          5815 => x"81065155",
          5816 => x"5673802e",
          5817 => x"9e38767f",
          5818 => x"53705254",
          5819 => x"dba83f81",
          5820 => x"d3840894",
          5821 => x"150c8e39",
          5822 => x"81d38408",
          5823 => x"842e0981",
          5824 => x"06833885",
          5825 => x"557481d3",
          5826 => x"840c933d",
          5827 => x"0d04e43d",
          5828 => x"0d6f6f5b",
          5829 => x"5b807a34",
          5830 => x"80539e3d",
          5831 => x"ffb80552",
          5832 => x"9f3d51e8",
          5833 => x"b53f81d3",
          5834 => x"84085781",
          5835 => x"d3840882",
          5836 => x"fc387b43",
          5837 => x"7a7c9411",
          5838 => x"08475558",
          5839 => x"64547380",
          5840 => x"2e81ed38",
          5841 => x"a052933d",
          5842 => x"705255d5",
          5843 => x"ea3f81d3",
          5844 => x"84085781",
          5845 => x"d3840882",
          5846 => x"d4386852",
          5847 => x"7b51c9c8",
          5848 => x"3f81d384",
          5849 => x"085781d3",
          5850 => x"840882c1",
          5851 => x"3869527b",
          5852 => x"51daa33f",
          5853 => x"81d38408",
          5854 => x"45765274",
          5855 => x"51d5b83f",
          5856 => x"81d38408",
          5857 => x"5781d384",
          5858 => x"0882a238",
          5859 => x"80527451",
          5860 => x"daeb3f81",
          5861 => x"d3840857",
          5862 => x"81d38408",
          5863 => x"a4386952",
          5864 => x"7b51d9f2",
          5865 => x"3f7381d3",
          5866 => x"84082ea6",
          5867 => x"38765274",
          5868 => x"51d6cf3f",
          5869 => x"81d38408",
          5870 => x"5781d384",
          5871 => x"08802ecc",
          5872 => x"3876842e",
          5873 => x"09810686",
          5874 => x"38825781",
          5875 => x"e0397681",
          5876 => x"dc389e3d",
          5877 => x"ffbc0552",
          5878 => x"7451dcc9",
          5879 => x"3f76903d",
          5880 => x"78118111",
          5881 => x"3351565a",
          5882 => x"5673802e",
          5883 => x"913802b9",
          5884 => x"05558116",
          5885 => x"81167033",
          5886 => x"56565673",
          5887 => x"f5388116",
          5888 => x"54737826",
          5889 => x"81903875",
          5890 => x"802e9938",
          5891 => x"78168105",
          5892 => x"55ff186f",
          5893 => x"11ff18ff",
          5894 => x"18585855",
          5895 => x"58743374",
          5896 => x"3475ee38",
          5897 => x"ff186f11",
          5898 => x"5558af74",
          5899 => x"34fe8d39",
          5900 => x"777b2e09",
          5901 => x"81068a38",
          5902 => x"ff186f11",
          5903 => x"5558af74",
          5904 => x"34800b81",
          5905 => x"d3b43370",
          5906 => x"842981c2",
          5907 => x"e8057008",
          5908 => x"7033525c",
          5909 => x"56565673",
          5910 => x"762e8d38",
          5911 => x"8116701a",
          5912 => x"70335155",
          5913 => x"5673f538",
          5914 => x"82165473",
          5915 => x"7826a738",
          5916 => x"80557476",
          5917 => x"27913874",
          5918 => x"19547333",
          5919 => x"7a708105",
          5920 => x"5c348115",
          5921 => x"55ec39ba",
          5922 => x"7a708105",
          5923 => x"5c3474ff",
          5924 => x"2e098106",
          5925 => x"85389157",
          5926 => x"94396e18",
          5927 => x"81195954",
          5928 => x"73337a70",
          5929 => x"81055c34",
          5930 => x"7a7826ee",
          5931 => x"38807a34",
          5932 => x"7681d384",
          5933 => x"0c9e3d0d",
          5934 => x"04f73d0d",
          5935 => x"7b7d8d3d",
          5936 => x"fc055471",
          5937 => x"535755ec",
          5938 => x"bb3f81d3",
          5939 => x"84085381",
          5940 => x"d3840882",
          5941 => x"fa389115",
          5942 => x"33537282",
          5943 => x"f2388c15",
          5944 => x"08547376",
          5945 => x"27923890",
          5946 => x"15337081",
          5947 => x"2a708106",
          5948 => x"51545772",
          5949 => x"83387356",
          5950 => x"94150854",
          5951 => x"80709417",
          5952 => x"0c587578",
          5953 => x"2e829738",
          5954 => x"798a1122",
          5955 => x"70892b59",
          5956 => x"51537378",
          5957 => x"2eb73876",
          5958 => x"52ff1651",
          5959 => x"ff98d83f",
          5960 => x"81d38408",
          5961 => x"ff157854",
          5962 => x"70535553",
          5963 => x"ff98c83f",
          5964 => x"81d38408",
          5965 => x"73269638",
          5966 => x"76307075",
          5967 => x"06709418",
          5968 => x"0c777131",
          5969 => x"98180857",
          5970 => x"585153b1",
          5971 => x"39881508",
          5972 => x"5473a638",
          5973 => x"73527451",
          5974 => x"cdca3f81",
          5975 => x"d3840854",
          5976 => x"81d38408",
          5977 => x"812e819a",
          5978 => x"3881d384",
          5979 => x"08ff2e81",
          5980 => x"9b3881d3",
          5981 => x"84088816",
          5982 => x"0c739816",
          5983 => x"0c73802e",
          5984 => x"819c3876",
          5985 => x"762780dc",
          5986 => x"38757731",
          5987 => x"94160818",
          5988 => x"94170c90",
          5989 => x"16337081",
          5990 => x"2a708106",
          5991 => x"51555a56",
          5992 => x"72802e9a",
          5993 => x"38735274",
          5994 => x"51ccf93f",
          5995 => x"81d38408",
          5996 => x"5481d384",
          5997 => x"08943881",
          5998 => x"d3840856",
          5999 => x"a7397352",
          6000 => x"7451c784",
          6001 => x"3f81d384",
          6002 => x"085473ff",
          6003 => x"2ebe3881",
          6004 => x"7427af38",
          6005 => x"79537398",
          6006 => x"140827a6",
          6007 => x"38739816",
          6008 => x"0cffa039",
          6009 => x"94150816",
          6010 => x"94160c75",
          6011 => x"83ff0653",
          6012 => x"72802eaa",
          6013 => x"38735279",
          6014 => x"51c6a33f",
          6015 => x"81d38408",
          6016 => x"9438820b",
          6017 => x"91163482",
          6018 => x"5380c439",
          6019 => x"810b9116",
          6020 => x"348153bb",
          6021 => x"3975892a",
          6022 => x"81d38408",
          6023 => x"05589415",
          6024 => x"08548c15",
          6025 => x"08742790",
          6026 => x"38738c16",
          6027 => x"0c901533",
          6028 => x"80c00753",
          6029 => x"72901634",
          6030 => x"7383ff06",
          6031 => x"5372802e",
          6032 => x"8c38779c",
          6033 => x"16082e85",
          6034 => x"38779c16",
          6035 => x"0c805372",
          6036 => x"81d3840c",
          6037 => x"8b3d0d04",
          6038 => x"f93d0d79",
          6039 => x"56895475",
          6040 => x"802e818a",
          6041 => x"38805389",
          6042 => x"3dfc0552",
          6043 => x"8a3d8405",
          6044 => x"51e1e73f",
          6045 => x"81d38408",
          6046 => x"5581d384",
          6047 => x"0880ea38",
          6048 => x"77760c7a",
          6049 => x"527551d8",
          6050 => x"b53f81d3",
          6051 => x"84085581",
          6052 => x"d3840880",
          6053 => x"c338ab16",
          6054 => x"3370982b",
          6055 => x"55578074",
          6056 => x"24a23886",
          6057 => x"16337084",
          6058 => x"2a708106",
          6059 => x"51555773",
          6060 => x"802ead38",
          6061 => x"9c160852",
          6062 => x"7751d3da",
          6063 => x"3f81d384",
          6064 => x"0888170c",
          6065 => x"77548614",
          6066 => x"22841723",
          6067 => x"74527551",
          6068 => x"cee53f81",
          6069 => x"d3840855",
          6070 => x"74842e09",
          6071 => x"81068538",
          6072 => x"85558639",
          6073 => x"74802e84",
          6074 => x"3880760c",
          6075 => x"74547381",
          6076 => x"d3840c89",
          6077 => x"3d0d04fc",
          6078 => x"3d0d7687",
          6079 => x"3dfc0553",
          6080 => x"705253e7",
          6081 => x"ff3f81d3",
          6082 => x"84088738",
          6083 => x"81d38408",
          6084 => x"730c863d",
          6085 => x"0d04fb3d",
          6086 => x"0d777989",
          6087 => x"3dfc0554",
          6088 => x"71535654",
          6089 => x"e7de3f81",
          6090 => x"d3840853",
          6091 => x"81d38408",
          6092 => x"80df3874",
          6093 => x"933881d3",
          6094 => x"84085273",
          6095 => x"51cdf83f",
          6096 => x"81d38408",
          6097 => x"5380ca39",
          6098 => x"81d38408",
          6099 => x"527351d3",
          6100 => x"ac3f81d3",
          6101 => x"84085381",
          6102 => x"d3840884",
          6103 => x"2e098106",
          6104 => x"85388053",
          6105 => x"873981d3",
          6106 => x"8408a638",
          6107 => x"74527351",
          6108 => x"d5b33f72",
          6109 => x"527351cf",
          6110 => x"893f81d3",
          6111 => x"84088432",
          6112 => x"70307072",
          6113 => x"079f2c70",
          6114 => x"81d38408",
          6115 => x"06515154",
          6116 => x"547281d3",
          6117 => x"840c873d",
          6118 => x"0d04ee3d",
          6119 => x"0d655780",
          6120 => x"53893d70",
          6121 => x"53963d52",
          6122 => x"56dfaf3f",
          6123 => x"81d38408",
          6124 => x"5581d384",
          6125 => x"08b23864",
          6126 => x"527551d6",
          6127 => x"813f81d3",
          6128 => x"84085581",
          6129 => x"d38408a0",
          6130 => x"380280cb",
          6131 => x"05337098",
          6132 => x"2b555873",
          6133 => x"80258538",
          6134 => x"86558d39",
          6135 => x"76802e88",
          6136 => x"38765275",
          6137 => x"51d4be3f",
          6138 => x"7481d384",
          6139 => x"0c943d0d",
          6140 => x"04f03d0d",
          6141 => x"6365555c",
          6142 => x"8053923d",
          6143 => x"ec055293",
          6144 => x"3d51ded6",
          6145 => x"3f81d384",
          6146 => x"085b81d3",
          6147 => x"84088280",
          6148 => x"387c740c",
          6149 => x"73089811",
          6150 => x"08fe1190",
          6151 => x"13085956",
          6152 => x"58557574",
          6153 => x"26913875",
          6154 => x"7c0c81e4",
          6155 => x"39815b81",
          6156 => x"cc39825b",
          6157 => x"81c73981",
          6158 => x"d3840875",
          6159 => x"33555973",
          6160 => x"812e0981",
          6161 => x"06bf3882",
          6162 => x"755f5776",
          6163 => x"52923df0",
          6164 => x"0551c1f4",
          6165 => x"3f81d384",
          6166 => x"08ff2ed1",
          6167 => x"3881d384",
          6168 => x"08812ece",
          6169 => x"3881d384",
          6170 => x"08307081",
          6171 => x"d3840807",
          6172 => x"80257a05",
          6173 => x"81197f53",
          6174 => x"595a5498",
          6175 => x"14087726",
          6176 => x"ca3880f9",
          6177 => x"39a41508",
          6178 => x"81d38408",
          6179 => x"57587598",
          6180 => x"38775281",
          6181 => x"187d5258",
          6182 => x"ffbf8d3f",
          6183 => x"81d38408",
          6184 => x"5b81d384",
          6185 => x"0880d638",
          6186 => x"7c703377",
          6187 => x"12ff1a5d",
          6188 => x"52565474",
          6189 => x"822e0981",
          6190 => x"069e38b4",
          6191 => x"1451ffbb",
          6192 => x"cb3f81d3",
          6193 => x"840883ff",
          6194 => x"ff067030",
          6195 => x"7080251b",
          6196 => x"8219595b",
          6197 => x"51549b39",
          6198 => x"b41451ff",
          6199 => x"bbc53f81",
          6200 => x"d38408f0",
          6201 => x"0a067030",
          6202 => x"7080251b",
          6203 => x"8419595b",
          6204 => x"51547583",
          6205 => x"ff067a58",
          6206 => x"5679ff92",
          6207 => x"38787c0c",
          6208 => x"7c799012",
          6209 => x"0c841133",
          6210 => x"81075654",
          6211 => x"74841534",
          6212 => x"7a81d384",
          6213 => x"0c923d0d",
          6214 => x"04f93d0d",
          6215 => x"798a3dfc",
          6216 => x"05537052",
          6217 => x"57e3dd3f",
          6218 => x"81d38408",
          6219 => x"5681d384",
          6220 => x"0881a838",
          6221 => x"91173356",
          6222 => x"7581a038",
          6223 => x"90173370",
          6224 => x"812a7081",
          6225 => x"06515555",
          6226 => x"87557380",
          6227 => x"2e818e38",
          6228 => x"94170854",
          6229 => x"738c1808",
          6230 => x"27818038",
          6231 => x"739b3881",
          6232 => x"d3840853",
          6233 => x"88170852",
          6234 => x"7651c48c",
          6235 => x"3f81d384",
          6236 => x"08748819",
          6237 => x"0c5680c9",
          6238 => x"39981708",
          6239 => x"527651ff",
          6240 => x"bfc63f81",
          6241 => x"d38408ff",
          6242 => x"2e098106",
          6243 => x"83388156",
          6244 => x"81d38408",
          6245 => x"812e0981",
          6246 => x"06853882",
          6247 => x"56a33975",
          6248 => x"a0387754",
          6249 => x"81d38408",
          6250 => x"98150827",
          6251 => x"94389817",
          6252 => x"085381d3",
          6253 => x"84085276",
          6254 => x"51c3bd3f",
          6255 => x"81d38408",
          6256 => x"56941708",
          6257 => x"8c180c90",
          6258 => x"173380c0",
          6259 => x"07547390",
          6260 => x"18347580",
          6261 => x"2e853875",
          6262 => x"91183475",
          6263 => x"557481d3",
          6264 => x"840c893d",
          6265 => x"0d04e23d",
          6266 => x"0d8253a0",
          6267 => x"3dffa405",
          6268 => x"52a13d51",
          6269 => x"dae43f81",
          6270 => x"d3840855",
          6271 => x"81d38408",
          6272 => x"81f53878",
          6273 => x"45a13d08",
          6274 => x"52953d70",
          6275 => x"5258d1ae",
          6276 => x"3f81d384",
          6277 => x"085581d3",
          6278 => x"840881db",
          6279 => x"380280fb",
          6280 => x"05337085",
          6281 => x"2a708106",
          6282 => x"51555686",
          6283 => x"557381c7",
          6284 => x"3875982b",
          6285 => x"54807424",
          6286 => x"81bd3802",
          6287 => x"80d60533",
          6288 => x"70810658",
          6289 => x"54875576",
          6290 => x"81ad386b",
          6291 => x"527851cc",
          6292 => x"c53f81d3",
          6293 => x"84087484",
          6294 => x"2a708106",
          6295 => x"51555673",
          6296 => x"802e80d4",
          6297 => x"38785481",
          6298 => x"d3840894",
          6299 => x"15082e81",
          6300 => x"8638735a",
          6301 => x"81d38408",
          6302 => x"5c76528a",
          6303 => x"3d705254",
          6304 => x"c7b53f81",
          6305 => x"d3840855",
          6306 => x"81d38408",
          6307 => x"80e93881",
          6308 => x"d3840852",
          6309 => x"7351cce5",
          6310 => x"3f81d384",
          6311 => x"085581d3",
          6312 => x"84088638",
          6313 => x"875580cf",
          6314 => x"3981d384",
          6315 => x"08842e88",
          6316 => x"3881d384",
          6317 => x"0880c038",
          6318 => x"7751cec2",
          6319 => x"3f81d384",
          6320 => x"0881d384",
          6321 => x"08307081",
          6322 => x"d3840807",
          6323 => x"80255155",
          6324 => x"5575802e",
          6325 => x"94387380",
          6326 => x"2e8f3880",
          6327 => x"53755277",
          6328 => x"51c1953f",
          6329 => x"81d38408",
          6330 => x"55748c38",
          6331 => x"7851ffba",
          6332 => x"fe3f81d3",
          6333 => x"84085574",
          6334 => x"81d3840c",
          6335 => x"a03d0d04",
          6336 => x"e93d0d82",
          6337 => x"53993dc0",
          6338 => x"05529a3d",
          6339 => x"51d8cb3f",
          6340 => x"81d38408",
          6341 => x"5481d384",
          6342 => x"0882b038",
          6343 => x"785e6952",
          6344 => x"8e3d7052",
          6345 => x"58cf973f",
          6346 => x"81d38408",
          6347 => x"5481d384",
          6348 => x"08863888",
          6349 => x"54829439",
          6350 => x"81d38408",
          6351 => x"842e0981",
          6352 => x"06828838",
          6353 => x"0280df05",
          6354 => x"3370852a",
          6355 => x"81065155",
          6356 => x"86547481",
          6357 => x"f638785a",
          6358 => x"74528a3d",
          6359 => x"705257c1",
          6360 => x"c33f81d3",
          6361 => x"84087555",
          6362 => x"5681d384",
          6363 => x"08833887",
          6364 => x"5481d384",
          6365 => x"08812e09",
          6366 => x"81068338",
          6367 => x"825481d3",
          6368 => x"8408ff2e",
          6369 => x"09810686",
          6370 => x"38815481",
          6371 => x"b4397381",
          6372 => x"b03881d3",
          6373 => x"84085278",
          6374 => x"51c4a43f",
          6375 => x"81d38408",
          6376 => x"5481d384",
          6377 => x"08819a38",
          6378 => x"8b53a052",
          6379 => x"b41951ff",
          6380 => x"b78c3f78",
          6381 => x"54ae0bb4",
          6382 => x"15347854",
          6383 => x"900bbf15",
          6384 => x"348288b2",
          6385 => x"0a5280ca",
          6386 => x"1951ffb6",
          6387 => x"9f3f7553",
          6388 => x"78b41153",
          6389 => x"51c9f83f",
          6390 => x"a05378b4",
          6391 => x"115380d4",
          6392 => x"0551ffb6",
          6393 => x"b63f7854",
          6394 => x"ae0b80d5",
          6395 => x"15347f53",
          6396 => x"7880d411",
          6397 => x"5351c9d7",
          6398 => x"3f785481",
          6399 => x"0b831534",
          6400 => x"7751cba4",
          6401 => x"3f81d384",
          6402 => x"085481d3",
          6403 => x"8408b238",
          6404 => x"8288b20a",
          6405 => x"52649605",
          6406 => x"51ffb5d0",
          6407 => x"3f755364",
          6408 => x"527851c9",
          6409 => x"aa3f6454",
          6410 => x"900b8b15",
          6411 => x"34785481",
          6412 => x"0b831534",
          6413 => x"7851ffb8",
          6414 => x"b63f81d3",
          6415 => x"8408548b",
          6416 => x"39805375",
          6417 => x"527651ff",
          6418 => x"beae3f73",
          6419 => x"81d3840c",
          6420 => x"993d0d04",
          6421 => x"da3d0da9",
          6422 => x"3d840551",
          6423 => x"d2f13f82",
          6424 => x"53a83dff",
          6425 => x"840552a9",
          6426 => x"3d51d5ee",
          6427 => x"3f81d384",
          6428 => x"085581d3",
          6429 => x"840882d3",
          6430 => x"38784da9",
          6431 => x"3d08529d",
          6432 => x"3d705258",
          6433 => x"ccb83f81",
          6434 => x"d3840855",
          6435 => x"81d38408",
          6436 => x"82b93802",
          6437 => x"819b0533",
          6438 => x"81a00654",
          6439 => x"86557382",
          6440 => x"aa38a053",
          6441 => x"a43d0852",
          6442 => x"a83dff88",
          6443 => x"0551ffb4",
          6444 => x"ea3fac53",
          6445 => x"7752923d",
          6446 => x"705254ff",
          6447 => x"b4dd3faa",
          6448 => x"3d085273",
          6449 => x"51cbf73f",
          6450 => x"81d38408",
          6451 => x"5581d384",
          6452 => x"08953863",
          6453 => x"6f2e0981",
          6454 => x"06883865",
          6455 => x"a23d082e",
          6456 => x"92388855",
          6457 => x"81e53981",
          6458 => x"d3840884",
          6459 => x"2e098106",
          6460 => x"81b83873",
          6461 => x"51c9b13f",
          6462 => x"81d38408",
          6463 => x"5581d384",
          6464 => x"0881c838",
          6465 => x"68569353",
          6466 => x"a83dff95",
          6467 => x"05528d16",
          6468 => x"51ffb487",
          6469 => x"3f02af05",
          6470 => x"338b1734",
          6471 => x"8b163370",
          6472 => x"842a7081",
          6473 => x"06515555",
          6474 => x"73893874",
          6475 => x"a0075473",
          6476 => x"8b173478",
          6477 => x"54810b83",
          6478 => x"15348b16",
          6479 => x"3370842a",
          6480 => x"70810651",
          6481 => x"55557380",
          6482 => x"2e80e538",
          6483 => x"6e642e80",
          6484 => x"df387552",
          6485 => x"7851c6be",
          6486 => x"3f81d384",
          6487 => x"08527851",
          6488 => x"ffb7bb3f",
          6489 => x"825581d3",
          6490 => x"8408802e",
          6491 => x"80dd3881",
          6492 => x"d3840852",
          6493 => x"7851ffb5",
          6494 => x"af3f81d3",
          6495 => x"84087980",
          6496 => x"d4115858",
          6497 => x"5581d384",
          6498 => x"0880c038",
          6499 => x"81163354",
          6500 => x"73ae2e09",
          6501 => x"81069938",
          6502 => x"63537552",
          6503 => x"7651c6af",
          6504 => x"3f785481",
          6505 => x"0b831534",
          6506 => x"873981d3",
          6507 => x"84089c38",
          6508 => x"7751c8ca",
          6509 => x"3f81d384",
          6510 => x"085581d3",
          6511 => x"84088c38",
          6512 => x"7851ffb5",
          6513 => x"aa3f81d3",
          6514 => x"84085574",
          6515 => x"81d3840c",
          6516 => x"a83d0d04",
          6517 => x"ed3d0d02",
          6518 => x"80db0533",
          6519 => x"02840580",
          6520 => x"df053357",
          6521 => x"57825395",
          6522 => x"3dd00552",
          6523 => x"963d51d2",
          6524 => x"e93f81d3",
          6525 => x"84085581",
          6526 => x"d3840880",
          6527 => x"cf38785a",
          6528 => x"6552953d",
          6529 => x"d40551c9",
          6530 => x"b53f81d3",
          6531 => x"84085581",
          6532 => x"d38408b8",
          6533 => x"380280cf",
          6534 => x"053381a0",
          6535 => x"06548655",
          6536 => x"73aa3875",
          6537 => x"a7066171",
          6538 => x"098b1233",
          6539 => x"71067a74",
          6540 => x"06075157",
          6541 => x"5556748b",
          6542 => x"15347854",
          6543 => x"810b8315",
          6544 => x"347851ff",
          6545 => x"b4a93f81",
          6546 => x"d3840855",
          6547 => x"7481d384",
          6548 => x"0c953d0d",
          6549 => x"04ef3d0d",
          6550 => x"64568253",
          6551 => x"933dd005",
          6552 => x"52943d51",
          6553 => x"d1f43f81",
          6554 => x"d3840855",
          6555 => x"81d38408",
          6556 => x"80cb3876",
          6557 => x"58635293",
          6558 => x"3dd40551",
          6559 => x"c8c03f81",
          6560 => x"d3840855",
          6561 => x"81d38408",
          6562 => x"b4380280",
          6563 => x"c7053381",
          6564 => x"a0065486",
          6565 => x"5573a638",
          6566 => x"84162286",
          6567 => x"17227190",
          6568 => x"2b075354",
          6569 => x"961f51ff",
          6570 => x"b0c23f76",
          6571 => x"54810b83",
          6572 => x"15347651",
          6573 => x"ffb3b83f",
          6574 => x"81d38408",
          6575 => x"557481d3",
          6576 => x"840c933d",
          6577 => x"0d04ea3d",
          6578 => x"0d696b5c",
          6579 => x"5a805398",
          6580 => x"3dd00552",
          6581 => x"993d51d1",
          6582 => x"813f81d3",
          6583 => x"840881d3",
          6584 => x"84083070",
          6585 => x"81d38408",
          6586 => x"07802551",
          6587 => x"55577980",
          6588 => x"2e818538",
          6589 => x"81707506",
          6590 => x"55557380",
          6591 => x"2e80f938",
          6592 => x"7b5d805f",
          6593 => x"80528d3d",
          6594 => x"705254ff",
          6595 => x"bea93f81",
          6596 => x"d3840857",
          6597 => x"81d38408",
          6598 => x"80d13874",
          6599 => x"527351c3",
          6600 => x"dc3f81d3",
          6601 => x"84085781",
          6602 => x"d38408bf",
          6603 => x"3881d384",
          6604 => x"0881d384",
          6605 => x"08655b59",
          6606 => x"56781881",
          6607 => x"197b1856",
          6608 => x"59557433",
          6609 => x"74348116",
          6610 => x"568a7827",
          6611 => x"ec388b56",
          6612 => x"751a5480",
          6613 => x"74347580",
          6614 => x"2e9e38ff",
          6615 => x"16701b70",
          6616 => x"33515556",
          6617 => x"73a02ee8",
          6618 => x"388e3976",
          6619 => x"842e0981",
          6620 => x"06863880",
          6621 => x"7a348057",
          6622 => x"76307078",
          6623 => x"07802551",
          6624 => x"547a802e",
          6625 => x"80c13873",
          6626 => x"802ebc38",
          6627 => x"7ba01108",
          6628 => x"5351ffb1",
          6629 => x"933f81d3",
          6630 => x"84085781",
          6631 => x"d38408a7",
          6632 => x"387b7033",
          6633 => x"555580c3",
          6634 => x"5673832e",
          6635 => x"8b3880e4",
          6636 => x"5673842e",
          6637 => x"8338a756",
          6638 => x"7515b405",
          6639 => x"51ffade3",
          6640 => x"3f81d384",
          6641 => x"087b0c76",
          6642 => x"81d3840c",
          6643 => x"983d0d04",
          6644 => x"e63d0d82",
          6645 => x"539c3dff",
          6646 => x"b805529d",
          6647 => x"3d51cefa",
          6648 => x"3f81d384",
          6649 => x"0881d384",
          6650 => x"08565481",
          6651 => x"d3840883",
          6652 => x"98388b53",
          6653 => x"a0528b3d",
          6654 => x"705259ff",
          6655 => x"aec03f73",
          6656 => x"6d703370",
          6657 => x"81ff0652",
          6658 => x"5755579f",
          6659 => x"742781bc",
          6660 => x"38785874",
          6661 => x"81ff066d",
          6662 => x"81054e70",
          6663 => x"5255ffaf",
          6664 => x"893f81d3",
          6665 => x"8408802e",
          6666 => x"a5386c70",
          6667 => x"33705357",
          6668 => x"54ffaefd",
          6669 => x"3f81d384",
          6670 => x"08802e8d",
          6671 => x"3874882b",
          6672 => x"76076d81",
          6673 => x"054e5586",
          6674 => x"3981d384",
          6675 => x"0855ff9f",
          6676 => x"157083ff",
          6677 => x"ff065154",
          6678 => x"7399268a",
          6679 => x"38e01570",
          6680 => x"83ffff06",
          6681 => x"565480ff",
          6682 => x"75278738",
          6683 => x"81c1f815",
          6684 => x"33557480",
          6685 => x"2ea33874",
          6686 => x"5281c3f8",
          6687 => x"51ffae89",
          6688 => x"3f81d384",
          6689 => x"08933881",
          6690 => x"ff752788",
          6691 => x"38768926",
          6692 => x"88388b39",
          6693 => x"8a772786",
          6694 => x"38865581",
          6695 => x"ec3981ff",
          6696 => x"75278f38",
          6697 => x"74882a54",
          6698 => x"73787081",
          6699 => x"055a3481",
          6700 => x"17577478",
          6701 => x"7081055a",
          6702 => x"3481176d",
          6703 => x"70337081",
          6704 => x"ff065257",
          6705 => x"5557739f",
          6706 => x"26fec838",
          6707 => x"8b3d3354",
          6708 => x"86557381",
          6709 => x"e52e81b1",
          6710 => x"3876802e",
          6711 => x"993802a7",
          6712 => x"05557615",
          6713 => x"70335154",
          6714 => x"73a02e09",
          6715 => x"81068738",
          6716 => x"ff175776",
          6717 => x"ed387941",
          6718 => x"80438052",
          6719 => x"913d7052",
          6720 => x"55ffbab3",
          6721 => x"3f81d384",
          6722 => x"085481d3",
          6723 => x"840880f7",
          6724 => x"38815274",
          6725 => x"51ffbfe5",
          6726 => x"3f81d384",
          6727 => x"085481d3",
          6728 => x"84088d38",
          6729 => x"7680c438",
          6730 => x"6754e574",
          6731 => x"3480c639",
          6732 => x"81d38408",
          6733 => x"842e0981",
          6734 => x"0680cc38",
          6735 => x"80547674",
          6736 => x"2e80c438",
          6737 => x"81527451",
          6738 => x"ffbdb03f",
          6739 => x"81d38408",
          6740 => x"5481d384",
          6741 => x"08b138a0",
          6742 => x"5381d384",
          6743 => x"08526751",
          6744 => x"ffabdb3f",
          6745 => x"6754880b",
          6746 => x"8b15348b",
          6747 => x"53785267",
          6748 => x"51ffaba7",
          6749 => x"3f795481",
          6750 => x"0b831534",
          6751 => x"7951ffad",
          6752 => x"ee3f81d3",
          6753 => x"84085473",
          6754 => x"557481d3",
          6755 => x"840c9c3d",
          6756 => x"0d04f23d",
          6757 => x"0d606202",
          6758 => x"880580cb",
          6759 => x"0533933d",
          6760 => x"fc055572",
          6761 => x"54405e5a",
          6762 => x"d2da3f81",
          6763 => x"d3840858",
          6764 => x"81d38408",
          6765 => x"82bd3891",
          6766 => x"1a335877",
          6767 => x"82b5387c",
          6768 => x"802e9738",
          6769 => x"8c1a0859",
          6770 => x"78903890",
          6771 => x"1a337081",
          6772 => x"2a708106",
          6773 => x"51555573",
          6774 => x"90388754",
          6775 => x"82973982",
          6776 => x"58829039",
          6777 => x"8158828b",
          6778 => x"397e8a11",
          6779 => x"2270892b",
          6780 => x"70557f54",
          6781 => x"565656fe",
          6782 => x"fefd3fff",
          6783 => x"147d0670",
          6784 => x"30707207",
          6785 => x"9f2a81d3",
          6786 => x"8408058c",
          6787 => x"19087c40",
          6788 => x"5a5d5555",
          6789 => x"81772788",
          6790 => x"38981608",
          6791 => x"77268338",
          6792 => x"82577677",
          6793 => x"56598056",
          6794 => x"74527951",
          6795 => x"ffae993f",
          6796 => x"81157f55",
          6797 => x"55981408",
          6798 => x"75268338",
          6799 => x"825581d3",
          6800 => x"8408812e",
          6801 => x"ff993881",
          6802 => x"d38408ff",
          6803 => x"2eff9538",
          6804 => x"81d38408",
          6805 => x"8e388116",
          6806 => x"56757b2e",
          6807 => x"09810687",
          6808 => x"38933974",
          6809 => x"59805674",
          6810 => x"772e0981",
          6811 => x"06ffb938",
          6812 => x"875880ff",
          6813 => x"397d802e",
          6814 => x"ba38787b",
          6815 => x"55557a80",
          6816 => x"2eb43881",
          6817 => x"15567381",
          6818 => x"2e098106",
          6819 => x"8338ff56",
          6820 => x"75537452",
          6821 => x"7e51ffaf",
          6822 => x"a83f81d3",
          6823 => x"84085881",
          6824 => x"d3840880",
          6825 => x"ce387481",
          6826 => x"16ff1656",
          6827 => x"565c73d3",
          6828 => x"388439ff",
          6829 => x"195c7e7c",
          6830 => x"8c120c55",
          6831 => x"7d802eb3",
          6832 => x"3878881b",
          6833 => x"0c7c8c1b",
          6834 => x"0c901a33",
          6835 => x"80c00754",
          6836 => x"73901b34",
          6837 => x"981508fe",
          6838 => x"05901608",
          6839 => x"57547574",
          6840 => x"26913875",
          6841 => x"7b319016",
          6842 => x"0c841533",
          6843 => x"81075473",
          6844 => x"84163477",
          6845 => x"547381d3",
          6846 => x"840c903d",
          6847 => x"0d04e93d",
          6848 => x"0d6b6d02",
          6849 => x"880580eb",
          6850 => x"05339d3d",
          6851 => x"545a5c59",
          6852 => x"c5bd3f8b",
          6853 => x"56800b81",
          6854 => x"d3840824",
          6855 => x"8bf83881",
          6856 => x"d3840884",
          6857 => x"2981d3a0",
          6858 => x"05700851",
          6859 => x"5574802e",
          6860 => x"84388075",
          6861 => x"3481d384",
          6862 => x"0881ff06",
          6863 => x"5f81527e",
          6864 => x"51ffa0d0",
          6865 => x"3f81d384",
          6866 => x"0881ff06",
          6867 => x"70810656",
          6868 => x"57835674",
          6869 => x"8bc03876",
          6870 => x"822a7081",
          6871 => x"0651558a",
          6872 => x"56748bb2",
          6873 => x"38993dfc",
          6874 => x"05538352",
          6875 => x"7e51ffa4",
          6876 => x"f03f81d3",
          6877 => x"84089938",
          6878 => x"67557480",
          6879 => x"2e923874",
          6880 => x"82808026",
          6881 => x"8b38ff15",
          6882 => x"75065574",
          6883 => x"802e8338",
          6884 => x"81487880",
          6885 => x"2e873884",
          6886 => x"80792692",
          6887 => x"38788180",
          6888 => x"0a268b38",
          6889 => x"ff197906",
          6890 => x"5574802e",
          6891 => x"86389356",
          6892 => x"8ae43978",
          6893 => x"892a6e89",
          6894 => x"2a70892b",
          6895 => x"77594843",
          6896 => x"597a8338",
          6897 => x"81566130",
          6898 => x"70802577",
          6899 => x"07515591",
          6900 => x"56748ac2",
          6901 => x"38993df8",
          6902 => x"05538152",
          6903 => x"7e51ffa4",
          6904 => x"803f8156",
          6905 => x"81d38408",
          6906 => x"8aac3877",
          6907 => x"832a7077",
          6908 => x"0681d384",
          6909 => x"08435645",
          6910 => x"748338bf",
          6911 => x"4166558e",
          6912 => x"56607526",
          6913 => x"8a903874",
          6914 => x"61317048",
          6915 => x"5580ff75",
          6916 => x"278a8338",
          6917 => x"93567881",
          6918 => x"802689fa",
          6919 => x"3877812a",
          6920 => x"70810656",
          6921 => x"4374802e",
          6922 => x"95387787",
          6923 => x"06557482",
          6924 => x"2e838d38",
          6925 => x"77810655",
          6926 => x"74802e83",
          6927 => x"83387781",
          6928 => x"06559356",
          6929 => x"825e7480",
          6930 => x"2e89cb38",
          6931 => x"785a7d83",
          6932 => x"2e098106",
          6933 => x"80e13878",
          6934 => x"ae386691",
          6935 => x"2a57810b",
          6936 => x"81c49c22",
          6937 => x"565a7480",
          6938 => x"2e9d3874",
          6939 => x"77269838",
          6940 => x"81c49c56",
          6941 => x"79108217",
          6942 => x"70225757",
          6943 => x"5a74802e",
          6944 => x"86387675",
          6945 => x"27ee3879",
          6946 => x"526651fe",
          6947 => x"f9e93f81",
          6948 => x"d3840884",
          6949 => x"29848705",
          6950 => x"70892a5e",
          6951 => x"55a05c80",
          6952 => x"0b81d384",
          6953 => x"08fc808a",
          6954 => x"055644fd",
          6955 => x"fff00a75",
          6956 => x"2780ec38",
          6957 => x"88d33978",
          6958 => x"ae38668c",
          6959 => x"2a57810b",
          6960 => x"81c48c22",
          6961 => x"565a7480",
          6962 => x"2e9d3874",
          6963 => x"77269838",
          6964 => x"81c48c56",
          6965 => x"79108217",
          6966 => x"70225757",
          6967 => x"5a74802e",
          6968 => x"86387675",
          6969 => x"27ee3879",
          6970 => x"526651fe",
          6971 => x"f9893f81",
          6972 => x"d3840810",
          6973 => x"84055781",
          6974 => x"d384089f",
          6975 => x"f5269638",
          6976 => x"810b81d3",
          6977 => x"84081081",
          6978 => x"d3840805",
          6979 => x"7111722a",
          6980 => x"83055956",
          6981 => x"5e83ff17",
          6982 => x"892a5d81",
          6983 => x"5ca04460",
          6984 => x"1c7d1165",
          6985 => x"05697012",
          6986 => x"ff057130",
          6987 => x"70720674",
          6988 => x"315c5259",
          6989 => x"5759407d",
          6990 => x"832e0981",
          6991 => x"06893876",
          6992 => x"1c601841",
          6993 => x"5c843976",
          6994 => x"1d5d7990",
          6995 => x"29187062",
          6996 => x"31685851",
          6997 => x"55747626",
          6998 => x"87af3875",
          6999 => x"7c317d31",
          7000 => x"7a537065",
          7001 => x"315255fe",
          7002 => x"f88d3f81",
          7003 => x"d3840858",
          7004 => x"7d832e09",
          7005 => x"81069b38",
          7006 => x"81d38408",
          7007 => x"83fff526",
          7008 => x"80dd3878",
          7009 => x"87833879",
          7010 => x"812a5978",
          7011 => x"fdbe3886",
          7012 => x"f8397d82",
          7013 => x"2e098106",
          7014 => x"80c53883",
          7015 => x"fff50b81",
          7016 => x"d3840827",
          7017 => x"a038788f",
          7018 => x"38791a55",
          7019 => x"7480c026",
          7020 => x"86387459",
          7021 => x"fd963962",
          7022 => x"81065574",
          7023 => x"802e8f38",
          7024 => x"835efd88",
          7025 => x"3981d384",
          7026 => x"089ff526",
          7027 => x"92387886",
          7028 => x"b838791a",
          7029 => x"59818079",
          7030 => x"27fcf138",
          7031 => x"86ab3980",
          7032 => x"557d812e",
          7033 => x"09810683",
          7034 => x"387d559f",
          7035 => x"f578278b",
          7036 => x"38748106",
          7037 => x"558e5674",
          7038 => x"869c3884",
          7039 => x"80538052",
          7040 => x"7a51ffa2",
          7041 => x"b93f8b53",
          7042 => x"81c2b452",
          7043 => x"7a51ffa2",
          7044 => x"8a3f8480",
          7045 => x"528b1b51",
          7046 => x"ffa1b33f",
          7047 => x"798d1c34",
          7048 => x"7b83ffff",
          7049 => x"06528e1b",
          7050 => x"51ffa1a2",
          7051 => x"3f810b90",
          7052 => x"1c347d83",
          7053 => x"32703070",
          7054 => x"962a8480",
          7055 => x"06545155",
          7056 => x"911b51ff",
          7057 => x"a1883f66",
          7058 => x"557483ff",
          7059 => x"ff269038",
          7060 => x"7483ffff",
          7061 => x"0652931b",
          7062 => x"51ffa0f2",
          7063 => x"3f8a3974",
          7064 => x"52a01b51",
          7065 => x"ffa1853f",
          7066 => x"f80b951c",
          7067 => x"34bf5298",
          7068 => x"1b51ffa0",
          7069 => x"d93f81ff",
          7070 => x"529a1b51",
          7071 => x"ffa0cf3f",
          7072 => x"60529c1b",
          7073 => x"51ffa0e4",
          7074 => x"3f7d832e",
          7075 => x"09810680",
          7076 => x"cb388288",
          7077 => x"b20a5280",
          7078 => x"c31b51ff",
          7079 => x"a0ce3f7c",
          7080 => x"52a41b51",
          7081 => x"ffa0c53f",
          7082 => x"8252ac1b",
          7083 => x"51ffa0bc",
          7084 => x"3f8152b0",
          7085 => x"1b51ffa0",
          7086 => x"953f8652",
          7087 => x"b21b51ff",
          7088 => x"a08c3fff",
          7089 => x"800b80c0",
          7090 => x"1c34a90b",
          7091 => x"80c21c34",
          7092 => x"935381c2",
          7093 => x"c05280c7",
          7094 => x"1b51ae39",
          7095 => x"8288b20a",
          7096 => x"52a71b51",
          7097 => x"ffa0853f",
          7098 => x"7c83ffff",
          7099 => x"0652961b",
          7100 => x"51ff9fda",
          7101 => x"3fff800b",
          7102 => x"a41c34a9",
          7103 => x"0ba61c34",
          7104 => x"935381c2",
          7105 => x"d452ab1b",
          7106 => x"51ffa08f",
          7107 => x"3f82d4d5",
          7108 => x"5283fe1b",
          7109 => x"705259ff",
          7110 => x"9fb43f81",
          7111 => x"5460537a",
          7112 => x"527e51ff",
          7113 => x"9bd73f81",
          7114 => x"5681d384",
          7115 => x"0883e738",
          7116 => x"7d832e09",
          7117 => x"810680ee",
          7118 => x"38755460",
          7119 => x"8605537a",
          7120 => x"527e51ff",
          7121 => x"9bb73f84",
          7122 => x"80538052",
          7123 => x"7a51ff9f",
          7124 => x"ed3f848b",
          7125 => x"85a4d252",
          7126 => x"7a51ff9f",
          7127 => x"8f3f868a",
          7128 => x"85e4f252",
          7129 => x"83e41b51",
          7130 => x"ff9f813f",
          7131 => x"ff185283",
          7132 => x"e81b51ff",
          7133 => x"9ef63f82",
          7134 => x"5283ec1b",
          7135 => x"51ff9eec",
          7136 => x"3f82d4d5",
          7137 => x"527851ff",
          7138 => x"9ec43f75",
          7139 => x"54608705",
          7140 => x"537a527e",
          7141 => x"51ff9ae5",
          7142 => x"3f755460",
          7143 => x"16537a52",
          7144 => x"7e51ff9a",
          7145 => x"d83f6553",
          7146 => x"80527a51",
          7147 => x"ff9f8f3f",
          7148 => x"7f568058",
          7149 => x"7d832e09",
          7150 => x"81069a38",
          7151 => x"f8527a51",
          7152 => x"ff9ea93f",
          7153 => x"ff52841b",
          7154 => x"51ff9ea0",
          7155 => x"3ff00a52",
          7156 => x"881b5191",
          7157 => x"3987ffff",
          7158 => x"f8557d81",
          7159 => x"2e8338f8",
          7160 => x"5574527a",
          7161 => x"51ff9e84",
          7162 => x"3f7c5561",
          7163 => x"57746226",
          7164 => x"83387457",
          7165 => x"76547553",
          7166 => x"7a527e51",
          7167 => x"ff99fe3f",
          7168 => x"81d38408",
          7169 => x"82873884",
          7170 => x"805381d3",
          7171 => x"8408527a",
          7172 => x"51ff9eaa",
          7173 => x"3f761675",
          7174 => x"78315656",
          7175 => x"74cd3881",
          7176 => x"18587780",
          7177 => x"2eff8d38",
          7178 => x"79557d83",
          7179 => x"2e833863",
          7180 => x"55615774",
          7181 => x"62268338",
          7182 => x"74577654",
          7183 => x"75537a52",
          7184 => x"7e51ff99",
          7185 => x"b83f81d3",
          7186 => x"840881c1",
          7187 => x"38761675",
          7188 => x"78315656",
          7189 => x"74db388c",
          7190 => x"567d832e",
          7191 => x"93388656",
          7192 => x"6683ffff",
          7193 => x"268a3884",
          7194 => x"567d822e",
          7195 => x"83388156",
          7196 => x"64810658",
          7197 => x"7780fe38",
          7198 => x"84805377",
          7199 => x"527a51ff",
          7200 => x"9dbc3f82",
          7201 => x"d4d55278",
          7202 => x"51ff9cc2",
          7203 => x"3f83be1b",
          7204 => x"55777534",
          7205 => x"810b8116",
          7206 => x"34810b82",
          7207 => x"16347783",
          7208 => x"16347584",
          7209 => x"16346067",
          7210 => x"055680fd",
          7211 => x"c1527551",
          7212 => x"fef1c43f",
          7213 => x"fe0b8516",
          7214 => x"3481d384",
          7215 => x"08822abf",
          7216 => x"07567586",
          7217 => x"163481d3",
          7218 => x"84088716",
          7219 => x"34605283",
          7220 => x"c61b51ff",
          7221 => x"9c963f66",
          7222 => x"5283ca1b",
          7223 => x"51ff9c8c",
          7224 => x"3f815477",
          7225 => x"537a527e",
          7226 => x"51ff9891",
          7227 => x"3f815681",
          7228 => x"d38408a2",
          7229 => x"38805380",
          7230 => x"527e51ff",
          7231 => x"99e33f81",
          7232 => x"5681d384",
          7233 => x"08903889",
          7234 => x"398e568a",
          7235 => x"39815686",
          7236 => x"3981d384",
          7237 => x"08567581",
          7238 => x"d3840c99",
          7239 => x"3d0d04ff",
          7240 => x"3d0d7352",
          7241 => x"71932681",
          7242 => x"8e387184",
          7243 => x"2981bd80",
          7244 => x"05527108",
          7245 => x"0481c5ac",
          7246 => x"51818039",
          7247 => x"81c5b851",
          7248 => x"80f93981",
          7249 => x"c5cc5180",
          7250 => x"f23981c5",
          7251 => x"e05180eb",
          7252 => x"3981c5f0",
          7253 => x"5180e439",
          7254 => x"81c68051",
          7255 => x"80dd3981",
          7256 => x"c6945180",
          7257 => x"d63981c6",
          7258 => x"a45180cf",
          7259 => x"3981c6bc",
          7260 => x"5180c839",
          7261 => x"81c6d451",
          7262 => x"80c13981",
          7263 => x"c6ec51bb",
          7264 => x"3981c788",
          7265 => x"51b53981",
          7266 => x"c79c51af",
          7267 => x"3981c7c8",
          7268 => x"51a93981",
          7269 => x"c7dc51a3",
          7270 => x"3981c7fc",
          7271 => x"519d3981",
          7272 => x"c8905197",
          7273 => x"3981c8a8",
          7274 => x"51913981",
          7275 => x"c8c0518b",
          7276 => x"3981c8d8",
          7277 => x"51853981",
          7278 => x"c8e451ff",
          7279 => x"87fb3f83",
          7280 => x"3d0d04fb",
          7281 => x"3d0d7779",
          7282 => x"56567487",
          7283 => x"e7268a38",
          7284 => x"74527587",
          7285 => x"e8295191",
          7286 => x"3987e852",
          7287 => x"7451feef",
          7288 => x"963f81d3",
          7289 => x"84085275",
          7290 => x"51feef8b",
          7291 => x"3f81d384",
          7292 => x"08547953",
          7293 => x"755281c8",
          7294 => x"f451ff8d",
          7295 => x"a03f873d",
          7296 => x"0d04f53d",
          7297 => x"0d7d7f61",
          7298 => x"028c0580",
          7299 => x"c7053373",
          7300 => x"7315665f",
          7301 => x"5d5a5a5c",
          7302 => x"5c5c7852",
          7303 => x"81c99851",
          7304 => x"ff8cfa3f",
          7305 => x"81c9a051",
          7306 => x"ff878e3f",
          7307 => x"80557477",
          7308 => x"2780fc38",
          7309 => x"79902e89",
          7310 => x"3879a02e",
          7311 => x"a73880c6",
          7312 => x"39741653",
          7313 => x"7278278e",
          7314 => x"38722252",
          7315 => x"81c9a451",
          7316 => x"ff8cca3f",
          7317 => x"893981c9",
          7318 => x"b051ff86",
          7319 => x"dc3f8215",
          7320 => x"5580c339",
          7321 => x"74165372",
          7322 => x"78278e38",
          7323 => x"72085281",
          7324 => x"c99851ff",
          7325 => x"8ca73f89",
          7326 => x"3981c9ac",
          7327 => x"51ff86b9",
          7328 => x"3f841555",
          7329 => x"a1397416",
          7330 => x"53727827",
          7331 => x"8e387233",
          7332 => x"5281c9b8",
          7333 => x"51ff8c85",
          7334 => x"3f893981",
          7335 => x"c9c051ff",
          7336 => x"86973f81",
          7337 => x"1555a051",
          7338 => x"fefa8f3f",
          7339 => x"ff803981",
          7340 => x"c9c451ff",
          7341 => x"86833f80",
          7342 => x"55747727",
          7343 => x"aa387416",
          7344 => x"70337972",
          7345 => x"26525553",
          7346 => x"9f742790",
          7347 => x"3872802e",
          7348 => x"8b387380",
          7349 => x"fe268538",
          7350 => x"73518339",
          7351 => x"a051fef9",
          7352 => x"d93f8115",
          7353 => x"55d33981",
          7354 => x"c9c851ff",
          7355 => x"85cb3f76",
          7356 => x"16771a5a",
          7357 => x"56fefd94",
          7358 => x"3f81d384",
          7359 => x"08982b70",
          7360 => x"982c5155",
          7361 => x"74a02e09",
          7362 => x"8106a538",
          7363 => x"fefcfd3f",
          7364 => x"81d38408",
          7365 => x"982b7098",
          7366 => x"2c70a032",
          7367 => x"70307072",
          7368 => x"079f2a51",
          7369 => x"56565155",
          7370 => x"749b2e8c",
          7371 => x"3872dd38",
          7372 => x"749b2e09",
          7373 => x"81068538",
          7374 => x"80538c39",
          7375 => x"7a1c5372",
          7376 => x"7626fdd6",
          7377 => x"38ff5372",
          7378 => x"81d3840c",
          7379 => x"8d3d0d04",
          7380 => x"ec3d0d66",
          7381 => x"02840580",
          7382 => x"e3053369",
          7383 => x"72307074",
          7384 => x"07802570",
          7385 => x"87ff7427",
          7386 => x"07515158",
          7387 => x"5a5b5693",
          7388 => x"577480fb",
          7389 => x"38815375",
          7390 => x"528c3d70",
          7391 => x"5257c0b9",
          7392 => x"3f81d384",
          7393 => x"085681d3",
          7394 => x"8408b838",
          7395 => x"81d38408",
          7396 => x"87c09888",
          7397 => x"0c81d384",
          7398 => x"0859963d",
          7399 => x"d4055484",
          7400 => x"80537752",
          7401 => x"7651c4f6",
          7402 => x"3f81d384",
          7403 => x"085681d3",
          7404 => x"84089038",
          7405 => x"7a557480",
          7406 => x"2e893874",
          7407 => x"19751959",
          7408 => x"59d83996",
          7409 => x"3dd80551",
          7410 => x"cce03f75",
          7411 => x"30707707",
          7412 => x"80255155",
          7413 => x"79802e95",
          7414 => x"3874802e",
          7415 => x"903881c9",
          7416 => x"cc5387c0",
          7417 => x"98880852",
          7418 => x"7851fbd7",
          7419 => x"3f755776",
          7420 => x"81d3840c",
          7421 => x"963d0d04",
          7422 => x"f93d0d7b",
          7423 => x"028405b3",
          7424 => x"05335758",
          7425 => x"ff578053",
          7426 => x"7a527951",
          7427 => x"fec23f81",
          7428 => x"d38408a4",
          7429 => x"3875802e",
          7430 => x"88387581",
          7431 => x"2e983898",
          7432 => x"3960557f",
          7433 => x"5481d384",
          7434 => x"537e527d",
          7435 => x"51772d81",
          7436 => x"d3840857",
          7437 => x"83397704",
          7438 => x"7681d384",
          7439 => x"0c893d0d",
          7440 => x"04fc3d0d",
          7441 => x"029b0533",
          7442 => x"81c9d453",
          7443 => x"81c9dc52",
          7444 => x"55ff88c9",
          7445 => x"3f81d0a4",
          7446 => x"2251ff80",
          7447 => x"e43f81c9",
          7448 => x"e85481c9",
          7449 => x"f45381d0",
          7450 => x"a5335281",
          7451 => x"c9fc51ff",
          7452 => x"88ab3f74",
          7453 => x"802e8538",
          7454 => x"fefe943f",
          7455 => x"863d0d04",
          7456 => x"fe3d0d87",
          7457 => x"c0968008",
          7458 => x"53ff80fd",
          7459 => x"3f8151fe",
          7460 => x"f68e3f81",
          7461 => x"ca9851fe",
          7462 => x"f8863f80",
          7463 => x"51fef680",
          7464 => x"3f72812a",
          7465 => x"70810651",
          7466 => x"5271802e",
          7467 => x"95388151",
          7468 => x"fef5ed3f",
          7469 => x"81cab451",
          7470 => x"fef7e53f",
          7471 => x"8051fef5",
          7472 => x"df3f7282",
          7473 => x"2a708106",
          7474 => x"51527180",
          7475 => x"2e953881",
          7476 => x"51fef5cc",
          7477 => x"3f81cac8",
          7478 => x"51fef7c4",
          7479 => x"3f8051fe",
          7480 => x"f5be3f72",
          7481 => x"832a7081",
          7482 => x"06515271",
          7483 => x"802e9538",
          7484 => x"8151fef5",
          7485 => x"ab3f81ca",
          7486 => x"d851fef7",
          7487 => x"a33f8051",
          7488 => x"fef59d3f",
          7489 => x"72842a70",
          7490 => x"81065152",
          7491 => x"71802e95",
          7492 => x"388151fe",
          7493 => x"f58a3f81",
          7494 => x"caec51fe",
          7495 => x"f7823f80",
          7496 => x"51fef4fc",
          7497 => x"3f72852a",
          7498 => x"70810651",
          7499 => x"5271802e",
          7500 => x"95388151",
          7501 => x"fef4e93f",
          7502 => x"81cb8051",
          7503 => x"fef6e13f",
          7504 => x"8051fef4",
          7505 => x"db3f7286",
          7506 => x"2a708106",
          7507 => x"51527180",
          7508 => x"2e953881",
          7509 => x"51fef4c8",
          7510 => x"3f81cb94",
          7511 => x"51fef6c0",
          7512 => x"3f8051fe",
          7513 => x"f4ba3f72",
          7514 => x"872a7081",
          7515 => x"06515271",
          7516 => x"802e9538",
          7517 => x"8151fef4",
          7518 => x"a73f81cb",
          7519 => x"a851fef6",
          7520 => x"9f3f8051",
          7521 => x"fef4993f",
          7522 => x"72882a70",
          7523 => x"81065152",
          7524 => x"71802e95",
          7525 => x"388151fe",
          7526 => x"f4863f81",
          7527 => x"cbbc51fe",
          7528 => x"f5fe3f80",
          7529 => x"51fef3f8",
          7530 => x"3ffeffa6",
          7531 => x"3f843d0d",
          7532 => x"04fa3d0d",
          7533 => x"78700870",
          7534 => x"55555773",
          7535 => x"802e80f0",
          7536 => x"388e3973",
          7537 => x"770c8515",
          7538 => x"335380e4",
          7539 => x"39811454",
          7540 => x"80743370",
          7541 => x"81ff0657",
          7542 => x"575374a0",
          7543 => x"2e833881",
          7544 => x"5374802e",
          7545 => x"843872e5",
          7546 => x"387581ff",
          7547 => x"065372a0",
          7548 => x"2e098106",
          7549 => x"88388074",
          7550 => x"70810556",
          7551 => x"34805675",
          7552 => x"902981d0",
          7553 => x"c4057708",
          7554 => x"53700852",
          7555 => x"55feedff",
          7556 => x"3f81d384",
          7557 => x"088b3884",
          7558 => x"15335372",
          7559 => x"812effa3",
          7560 => x"38811670",
          7561 => x"81ff0657",
          7562 => x"53937627",
          7563 => x"d238ff53",
          7564 => x"7281d384",
          7565 => x"0c883d0d",
          7566 => x"04cb3d0d",
          7567 => x"80707181",
          7568 => x"ea840c5e",
          7569 => x"5c81527b",
          7570 => x"51ff8ac8",
          7571 => x"3f81d384",
          7572 => x"0881ff06",
          7573 => x"59787c2e",
          7574 => x"098106a2",
          7575 => x"3881cbfc",
          7576 => x"52993d70",
          7577 => x"5259ff84",
          7578 => x"ca3f7b53",
          7579 => x"785281d4",
          7580 => x"b451ffb9",
          7581 => x"e33f81d3",
          7582 => x"84087c2e",
          7583 => x"883881cc",
          7584 => x"80518ee8",
          7585 => x"3981705e",
          7586 => x"5c81ccb8",
          7587 => x"51fefea9",
          7588 => x"3f993d70",
          7589 => x"465a80f8",
          7590 => x"53805279",
          7591 => x"51feebde",
          7592 => x"3f80f852",
          7593 => x"6451ff84",
          7594 => x"ce3fb73d",
          7595 => x"fef80551",
          7596 => x"fdff3f81",
          7597 => x"d3840890",
          7598 => x"2b70902c",
          7599 => x"51597880",
          7600 => x"c32e8a9b",
          7601 => x"387880c3",
          7602 => x"2480dc38",
          7603 => x"78ab2e83",
          7604 => x"bc3878ab",
          7605 => x"24a43878",
          7606 => x"822e81af",
          7607 => x"38788224",
          7608 => x"8a387880",
          7609 => x"2effa238",
          7610 => x"8d883978",
          7611 => x"842e8282",
          7612 => x"3878942e",
          7613 => x"82ad388c",
          7614 => x"f9397880",
          7615 => x"c02e858a",
          7616 => x"387880c0",
          7617 => x"24903878",
          7618 => x"b02e83a9",
          7619 => x"3878bc2e",
          7620 => x"848b388c",
          7621 => x"dd397880",
          7622 => x"c12e86eb",
          7623 => x"387880c2",
          7624 => x"2e888c38",
          7625 => x"8ccc3978",
          7626 => x"80f82e8b",
          7627 => x"ba387880",
          7628 => x"f824a938",
          7629 => x"7880d12e",
          7630 => x"8ae23878",
          7631 => x"80d1248b",
          7632 => x"387880d0",
          7633 => x"2e8ac438",
          7634 => x"8ca83978",
          7635 => x"80d42e8a",
          7636 => x"dc387880",
          7637 => x"d52e8af2",
          7638 => x"388c9739",
          7639 => x"7881832e",
          7640 => x"8bfc3878",
          7641 => x"81832492",
          7642 => x"387880f9",
          7643 => x"2e8b9d38",
          7644 => x"7881822e",
          7645 => x"8bd9388b",
          7646 => x"f9397881",
          7647 => x"852e8beb",
          7648 => x"38788187",
          7649 => x"2efe8238",
          7650 => x"8be839b7",
          7651 => x"3dfef411",
          7652 => x"53fef805",
          7653 => x"51ff83fa",
          7654 => x"3f81d384",
          7655 => x"08883881",
          7656 => x"ccbc518c",
          7657 => x"c739b73d",
          7658 => x"fef01153",
          7659 => x"fef80551",
          7660 => x"ff83df3f",
          7661 => x"81d38408",
          7662 => x"802e8838",
          7663 => x"81632583",
          7664 => x"38804302",
          7665 => x"80cb0533",
          7666 => x"520280cf",
          7667 => x"053351ff",
          7668 => x"87c23f81",
          7669 => x"d3840881",
          7670 => x"ff065978",
          7671 => x"8e3881cc",
          7672 => x"cc51fefb",
          7673 => x"d43f815d",
          7674 => x"fd9f3981",
          7675 => x"ccdc5189",
          7676 => x"d239b73d",
          7677 => x"fef41153",
          7678 => x"fef80551",
          7679 => x"ff83933f",
          7680 => x"81d38408",
          7681 => x"802efd81",
          7682 => x"38805380",
          7683 => x"520280cf",
          7684 => x"053351ff",
          7685 => x"8bcb3f81",
          7686 => x"d3840852",
          7687 => x"81ccf451",
          7688 => x"8aa639b7",
          7689 => x"3dfef411",
          7690 => x"53fef805",
          7691 => x"51ff82e2",
          7692 => x"3f81d384",
          7693 => x"08802e87",
          7694 => x"38638926",
          7695 => x"fccb38b7",
          7696 => x"3dfef011",
          7697 => x"53fef805",
          7698 => x"51ff82c6",
          7699 => x"3f81d384",
          7700 => x"08863881",
          7701 => x"d3840843",
          7702 => x"635381cc",
          7703 => x"fc527951",
          7704 => x"ff80d03f",
          7705 => x"0280cb05",
          7706 => x"33537952",
          7707 => x"6384b429",
          7708 => x"81d4b405",
          7709 => x"51ffb5e0",
          7710 => x"3f81d384",
          7711 => x"08819338",
          7712 => x"81cccc51",
          7713 => x"fefab23f",
          7714 => x"815cfbfd",
          7715 => x"39b73dfe",
          7716 => x"f80551fe",
          7717 => x"eabb3f81",
          7718 => x"d38408b8",
          7719 => x"3dfef805",
          7720 => x"525bfeeb",
          7721 => x"8e3f8153",
          7722 => x"81d38408",
          7723 => x"527a51f5",
          7724 => x"9f3f80d5",
          7725 => x"39b73dfe",
          7726 => x"f80551fe",
          7727 => x"ea933f81",
          7728 => x"d38408b8",
          7729 => x"3dfef805",
          7730 => x"525bfeea",
          7731 => x"e63f81d3",
          7732 => x"8408b83d",
          7733 => x"fef80552",
          7734 => x"5afeead7",
          7735 => x"3f81d384",
          7736 => x"08b83dfe",
          7737 => x"f8055259",
          7738 => x"feeac83f",
          7739 => x"81d08058",
          7740 => x"81d3b857",
          7741 => x"80568055",
          7742 => x"81d38408",
          7743 => x"81ff0654",
          7744 => x"78537952",
          7745 => x"7a51f5f0",
          7746 => x"3f81d384",
          7747 => x"08802efa",
          7748 => x"f83881d3",
          7749 => x"840851f0",
          7750 => x"863ffaed",
          7751 => x"39b73dfe",
          7752 => x"f41153fe",
          7753 => x"f80551ff",
          7754 => x"80e83f81",
          7755 => x"d3840880",
          7756 => x"2efad638",
          7757 => x"b73dfef0",
          7758 => x"1153fef8",
          7759 => x"0551ff80",
          7760 => x"d13f81d3",
          7761 => x"8408802e",
          7762 => x"fabf38b7",
          7763 => x"3dfeec11",
          7764 => x"53fef805",
          7765 => x"51ff80ba",
          7766 => x"3f81d384",
          7767 => x"08863881",
          7768 => x"d3840842",
          7769 => x"81cd8051",
          7770 => x"fef8ce3f",
          7771 => x"63635c5a",
          7772 => x"797b278f",
          7773 => x"38615978",
          7774 => x"7a708405",
          7775 => x"5c0c7a7a",
          7776 => x"26f53881",
          7777 => x"ccc85186",
          7778 => x"ba39b73d",
          7779 => x"fef41153",
          7780 => x"fef80551",
          7781 => x"fefffb3f",
          7782 => x"81d38408",
          7783 => x"80c43881",
          7784 => x"d0ad3359",
          7785 => x"78802e88",
          7786 => x"3881d080",
          7787 => x"0844b339",
          7788 => x"81d0ae33",
          7789 => x"5978802e",
          7790 => x"883881d0",
          7791 => x"880844a2",
          7792 => x"3981d0af",
          7793 => x"3359788b",
          7794 => x"3881d0b0",
          7795 => x"33597880",
          7796 => x"2e883881",
          7797 => x"d0900844",
          7798 => x"893981d0",
          7799 => x"a008fc80",
          7800 => x"0544b73d",
          7801 => x"fef01153",
          7802 => x"fef80551",
          7803 => x"feffa33f",
          7804 => x"81d38408",
          7805 => x"80c33881",
          7806 => x"d0ad3359",
          7807 => x"78802e88",
          7808 => x"3881d084",
          7809 => x"0843b239",
          7810 => x"81d0ae33",
          7811 => x"5978802e",
          7812 => x"883881d0",
          7813 => x"8c0843a1",
          7814 => x"3981d0af",
          7815 => x"3359788b",
          7816 => x"3881d0b0",
          7817 => x"33597880",
          7818 => x"2e883881",
          7819 => x"d0940843",
          7820 => x"883981d0",
          7821 => x"a0088805",
          7822 => x"43b73dfe",
          7823 => x"ec1153fe",
          7824 => x"f80551fe",
          7825 => x"fecc3f81",
          7826 => x"d3840880",
          7827 => x"2e9b3880",
          7828 => x"625b5979",
          7829 => x"882e8338",
          7830 => x"81597990",
          7831 => x"2e8d3878",
          7832 => x"802e8838",
          7833 => x"79a02e83",
          7834 => x"38884281",
          7835 => x"cd8c51fe",
          7836 => x"f6c73fa0",
          7837 => x"55635461",
          7838 => x"53625263",
          7839 => x"51ef833f",
          7840 => x"81cd9c51",
          7841 => x"84bd39b7",
          7842 => x"3dfef411",
          7843 => x"53fef805",
          7844 => x"51fefdfe",
          7845 => x"3f81d384",
          7846 => x"08802ef7",
          7847 => x"ec38b73d",
          7848 => x"fef01153",
          7849 => x"fef80551",
          7850 => x"fefde73f",
          7851 => x"81d38408",
          7852 => x"802ea538",
          7853 => x"63590280",
          7854 => x"cb053379",
          7855 => x"34638105",
          7856 => x"44b73dfe",
          7857 => x"f01153fe",
          7858 => x"f80551fe",
          7859 => x"fdc43f81",
          7860 => x"d38408e0",
          7861 => x"38f7b239",
          7862 => x"63703354",
          7863 => x"5281cda8",
          7864 => x"51fefbb9",
          7865 => x"3f80f852",
          7866 => x"7951fefc",
          7867 => x"8a3f7945",
          7868 => x"79335978",
          7869 => x"ae2ef791",
          7870 => x"389f7927",
          7871 => x"a038b73d",
          7872 => x"fef01153",
          7873 => x"fef80551",
          7874 => x"fefd873f",
          7875 => x"81d38408",
          7876 => x"802e9138",
          7877 => x"63590280",
          7878 => x"cb053379",
          7879 => x"34638105",
          7880 => x"44ffb539",
          7881 => x"81cdb451",
          7882 => x"fef58e3f",
          7883 => x"ffaa39b7",
          7884 => x"3dfee811",
          7885 => x"53fef805",
          7886 => x"51fefec8",
          7887 => x"3f81d384",
          7888 => x"08802ef6",
          7889 => x"c438b73d",
          7890 => x"fee41153",
          7891 => x"fef80551",
          7892 => x"fefeb13f",
          7893 => x"81d38408",
          7894 => x"802ea638",
          7895 => x"605902be",
          7896 => x"05227970",
          7897 => x"82055b23",
          7898 => x"7841b73d",
          7899 => x"fee41153",
          7900 => x"fef80551",
          7901 => x"fefe8d3f",
          7902 => x"81d38408",
          7903 => x"df38f689",
          7904 => x"39607022",
          7905 => x"545281cd",
          7906 => x"bc51fefa",
          7907 => x"903f80f8",
          7908 => x"527951fe",
          7909 => x"fae13f79",
          7910 => x"45793359",
          7911 => x"78ae2ef5",
          7912 => x"e838789f",
          7913 => x"26873860",
          7914 => x"840541d5",
          7915 => x"39b73dfe",
          7916 => x"e41153fe",
          7917 => x"f80551fe",
          7918 => x"fdca3f81",
          7919 => x"d3840880",
          7920 => x"2e923860",
          7921 => x"5902be05",
          7922 => x"22797082",
          7923 => x"055b2378",
          7924 => x"41ffae39",
          7925 => x"81cdb451",
          7926 => x"fef3de3f",
          7927 => x"ffa339b7",
          7928 => x"3dfee811",
          7929 => x"53fef805",
          7930 => x"51fefd98",
          7931 => x"3f81d384",
          7932 => x"08802ef5",
          7933 => x"9438b73d",
          7934 => x"fee41153",
          7935 => x"fef80551",
          7936 => x"fefd813f",
          7937 => x"81d38408",
          7938 => x"802ea138",
          7939 => x"6060710c",
          7940 => x"59608405",
          7941 => x"41b73dfe",
          7942 => x"e41153fe",
          7943 => x"f80551fe",
          7944 => x"fce23f81",
          7945 => x"d38408e4",
          7946 => x"38f4de39",
          7947 => x"60700854",
          7948 => x"5281cdc8",
          7949 => x"51fef8e5",
          7950 => x"3f80f852",
          7951 => x"7951fef9",
          7952 => x"b63f7945",
          7953 => x"79335978",
          7954 => x"ae2ef4bd",
          7955 => x"389f7927",
          7956 => x"a838b73d",
          7957 => x"fee41153",
          7958 => x"fef80551",
          7959 => x"fefca53f",
          7960 => x"81d38408",
          7961 => x"802e9938",
          7962 => x"7f536052",
          7963 => x"81cdc851",
          7964 => x"fef8aa3f",
          7965 => x"6060710c",
          7966 => x"59608405",
          7967 => x"41ffad39",
          7968 => x"81cdb451",
          7969 => x"fef2b23f",
          7970 => x"ffa23981",
          7971 => x"cdd451fe",
          7972 => x"f2a73f82",
          7973 => x"51fef195",
          7974 => x"3ff3ee39",
          7975 => x"81cdec51",
          7976 => x"fef2963f",
          7977 => x"a251fef0",
          7978 => x"e83ff3dd",
          7979 => x"39848081",
          7980 => x"0b87c094",
          7981 => x"840c8480",
          7982 => x"810b87c0",
          7983 => x"94940c81",
          7984 => x"ce8451fe",
          7985 => x"f1f33ff3",
          7986 => x"c03981ce",
          7987 => x"9851fef1",
          7988 => x"e83f8c80",
          7989 => x"830b87c0",
          7990 => x"94840c8c",
          7991 => x"80830b87",
          7992 => x"c094940c",
          7993 => x"f3a339b7",
          7994 => x"3dfef411",
          7995 => x"53fef805",
          7996 => x"51fef99e",
          7997 => x"3f81d384",
          7998 => x"08802ef3",
          7999 => x"8c386352",
          8000 => x"81ceac51",
          8001 => x"fef7963f",
          8002 => x"63597804",
          8003 => x"b73dfef4",
          8004 => x"1153fef8",
          8005 => x"0551fef8",
          8006 => x"f93f81d3",
          8007 => x"8408802e",
          8008 => x"f2e73863",
          8009 => x"5281cec8",
          8010 => x"51fef6f1",
          8011 => x"3f635978",
          8012 => x"2d81d384",
          8013 => x"085e81d3",
          8014 => x"8408802e",
          8015 => x"f2cb3881",
          8016 => x"d3840852",
          8017 => x"81cee451",
          8018 => x"fef6d23f",
          8019 => x"f2bb3981",
          8020 => x"cf8051fe",
          8021 => x"f0e33ffe",
          8022 => x"c5a63ff2",
          8023 => x"ac3981cf",
          8024 => x"9c51fef0",
          8025 => x"d43f8059",
          8026 => x"ffa039fe",
          8027 => x"eca13ff2",
          8028 => x"98396470",
          8029 => x"33515978",
          8030 => x"802ef28d",
          8031 => x"387b802e",
          8032 => x"80d2387c",
          8033 => x"802e80cc",
          8034 => x"38b73dfe",
          8035 => x"f80551fe",
          8036 => x"e0bf3f81",
          8037 => x"cfb05681",
          8038 => x"d3840855",
          8039 => x"81cfb454",
          8040 => x"805381cf",
          8041 => x"b852a33d",
          8042 => x"70525afe",
          8043 => x"f6853f81",
          8044 => x"d0805881",
          8045 => x"d3b85780",
          8046 => x"56648111",
          8047 => x"46810555",
          8048 => x"80548280",
          8049 => x"80538280",
          8050 => x"80527951",
          8051 => x"ecaa3f81",
          8052 => x"d384085e",
          8053 => x"7c81327c",
          8054 => x"81320759",
          8055 => x"788a387d",
          8056 => x"ff2e0981",
          8057 => x"06f1a238",
          8058 => x"81cfc851",
          8059 => x"fef5ae3f",
          8060 => x"f1973980",
          8061 => x"3d0d800b",
          8062 => x"81d3b834",
          8063 => x"9b9086e4",
          8064 => x"0b87c094",
          8065 => x"8c0c9b90",
          8066 => x"86e40b87",
          8067 => x"c0949c0c",
          8068 => x"8c80830b",
          8069 => x"87c09484",
          8070 => x"0c8c8083",
          8071 => x"0b87c094",
          8072 => x"940c9fba",
          8073 => x"0b81d394",
          8074 => x"0ca2bb0b",
          8075 => x"81d3980c",
          8076 => x"fee7b13f",
          8077 => x"feedd23f",
          8078 => x"81cfd851",
          8079 => x"fee4e13f",
          8080 => x"81cfe451",
          8081 => x"feeef23f",
          8082 => x"81a98051",
          8083 => x"feedb53f",
          8084 => x"8151ebed",
          8085 => x"3fefe23f",
          8086 => x"80040000",
          8087 => x"00ffffff",
          8088 => x"ff00ffff",
          8089 => x"ffff00ff",
          8090 => x"ffffff00",
          8091 => x"000014db",
          8092 => x"000014e1",
          8093 => x"000014e7",
          8094 => x"000014ed",
          8095 => x"000014f3",
          8096 => x"000051b1",
          8097 => x"00005135",
          8098 => x"0000513c",
          8099 => x"00005143",
          8100 => x"0000514a",
          8101 => x"00005151",
          8102 => x"00005158",
          8103 => x"0000515f",
          8104 => x"00005166",
          8105 => x"0000516d",
          8106 => x"00005174",
          8107 => x"0000517b",
          8108 => x"00005181",
          8109 => x"00005187",
          8110 => x"0000518d",
          8111 => x"00005193",
          8112 => x"00005199",
          8113 => x"0000519f",
          8114 => x"000051a5",
          8115 => x"000051ab",
          8116 => x"25642f25",
          8117 => x"642f2564",
          8118 => x"2025643a",
          8119 => x"25643a25",
          8120 => x"642e2564",
          8121 => x"25640a00",
          8122 => x"536f4320",
          8123 => x"436f6e66",
          8124 => x"69677572",
          8125 => x"6174696f",
          8126 => x"6e000000",
          8127 => x"20286672",
          8128 => x"6f6d2053",
          8129 => x"6f432063",
          8130 => x"6f6e6669",
          8131 => x"67290000",
          8132 => x"3a0a4465",
          8133 => x"76696365",
          8134 => x"7320696d",
          8135 => x"706c656d",
          8136 => x"656e7465",
          8137 => x"643a0a00",
          8138 => x"20202020",
          8139 => x"494e534e",
          8140 => x"20425241",
          8141 => x"4d202853",
          8142 => x"74617274",
          8143 => x"3d253038",
          8144 => x"582c2053",
          8145 => x"697a653d",
          8146 => x"25303858",
          8147 => x"292e0a00",
          8148 => x"20202020",
          8149 => x"4252414d",
          8150 => x"20285374",
          8151 => x"6172743d",
          8152 => x"25303858",
          8153 => x"2c205369",
          8154 => x"7a653d25",
          8155 => x"30385829",
          8156 => x"2e0a0000",
          8157 => x"20202020",
          8158 => x"52414d20",
          8159 => x"28537461",
          8160 => x"72743d25",
          8161 => x"3038582c",
          8162 => x"2053697a",
          8163 => x"653d2530",
          8164 => x"3858292e",
          8165 => x"0a000000",
          8166 => x"20202020",
          8167 => x"494f4354",
          8168 => x"4c0a0000",
          8169 => x"20202020",
          8170 => x"5053320a",
          8171 => x"00000000",
          8172 => x"20202020",
          8173 => x"5350490a",
          8174 => x"00000000",
          8175 => x"20202020",
          8176 => x"53442043",
          8177 => x"61726420",
          8178 => x"28446576",
          8179 => x"69636573",
          8180 => x"3d253032",
          8181 => x"58292e0a",
          8182 => x"00000000",
          8183 => x"20202020",
          8184 => x"494e5445",
          8185 => x"52525550",
          8186 => x"5420434f",
          8187 => x"4e54524f",
          8188 => x"4c4c4552",
          8189 => x"0a000000",
          8190 => x"20202020",
          8191 => x"54494d45",
          8192 => x"52312028",
          8193 => x"54696d65",
          8194 => x"72733d25",
          8195 => x"30315829",
          8196 => x"2e0a0000",
          8197 => x"41646472",
          8198 => x"65737365",
          8199 => x"733a0a00",
          8200 => x"20202020",
          8201 => x"43505520",
          8202 => x"52657365",
          8203 => x"74205665",
          8204 => x"63746f72",
          8205 => x"20416464",
          8206 => x"72657373",
          8207 => x"203d2025",
          8208 => x"3038580a",
          8209 => x"00000000",
          8210 => x"20202020",
          8211 => x"43505520",
          8212 => x"4d656d6f",
          8213 => x"72792053",
          8214 => x"74617274",
          8215 => x"20416464",
          8216 => x"72657373",
          8217 => x"203d2025",
          8218 => x"3038580a",
          8219 => x"00000000",
          8220 => x"20202020",
          8221 => x"53746163",
          8222 => x"6b205374",
          8223 => x"61727420",
          8224 => x"41646472",
          8225 => x"65737320",
          8226 => x"20202020",
          8227 => x"203d2025",
          8228 => x"3038580a",
          8229 => x"00000000",
          8230 => x"20202020",
          8231 => x"5a505520",
          8232 => x"49642020",
          8233 => x"20202020",
          8234 => x"20202020",
          8235 => x"20202020",
          8236 => x"20202020",
          8237 => x"203d2025",
          8238 => x"3038580a",
          8239 => x"00000000",
          8240 => x"20202020",
          8241 => x"53797374",
          8242 => x"656d2043",
          8243 => x"6c6f636b",
          8244 => x"20467265",
          8245 => x"71202020",
          8246 => x"20202020",
          8247 => x"203d2025",
          8248 => x"3038580a",
          8249 => x"00000000",
          8250 => x"536d616c",
          8251 => x"6c000000",
          8252 => x"4d656469",
          8253 => x"756d0000",
          8254 => x"466c6578",
          8255 => x"00000000",
          8256 => x"45564f00",
          8257 => x"45564f6d",
          8258 => x"696e0000",
          8259 => x"556e6b6e",
          8260 => x"6f776e00",
          8261 => x"53440000",
          8262 => x"222a2b2c",
          8263 => x"3a3b3c3d",
          8264 => x"3e3f5b5d",
          8265 => x"7c7f0000",
          8266 => x"46415400",
          8267 => x"46415433",
          8268 => x"32000000",
          8269 => x"ebfe904d",
          8270 => x"53444f53",
          8271 => x"352e3000",
          8272 => x"4e4f204e",
          8273 => x"414d4520",
          8274 => x"20202046",
          8275 => x"41543332",
          8276 => x"20202000",
          8277 => x"4e4f204e",
          8278 => x"414d4520",
          8279 => x"20202046",
          8280 => x"41542020",
          8281 => x"20202000",
          8282 => x"00006114",
          8283 => x"00000000",
          8284 => x"00000000",
          8285 => x"00000000",
          8286 => x"809a4541",
          8287 => x"8e418f80",
          8288 => x"45454549",
          8289 => x"49498e8f",
          8290 => x"9092924f",
          8291 => x"994f5555",
          8292 => x"59999a9b",
          8293 => x"9c9d9e9f",
          8294 => x"41494f55",
          8295 => x"a5a5a6a7",
          8296 => x"a8a9aaab",
          8297 => x"acadaeaf",
          8298 => x"b0b1b2b3",
          8299 => x"b4b5b6b7",
          8300 => x"b8b9babb",
          8301 => x"bcbdbebf",
          8302 => x"c0c1c2c3",
          8303 => x"c4c5c6c7",
          8304 => x"c8c9cacb",
          8305 => x"cccdcecf",
          8306 => x"d0d1d2d3",
          8307 => x"d4d5d6d7",
          8308 => x"d8d9dadb",
          8309 => x"dcdddedf",
          8310 => x"e0e1e2e3",
          8311 => x"e4e5e6e7",
          8312 => x"e8e9eaeb",
          8313 => x"ecedeeef",
          8314 => x"f0f1f2f3",
          8315 => x"f4f5f6f7",
          8316 => x"f8f9fafb",
          8317 => x"fcfdfeff",
          8318 => x"2b2e2c3b",
          8319 => x"3d5b5d2f",
          8320 => x"5c222a3a",
          8321 => x"3c3e3f7c",
          8322 => x"7f000000",
          8323 => x"00010004",
          8324 => x"00100040",
          8325 => x"01000200",
          8326 => x"00000000",
          8327 => x"00010002",
          8328 => x"00040008",
          8329 => x"00100020",
          8330 => x"00000000",
          8331 => x"64696e69",
          8332 => x"74000000",
          8333 => x"64696f63",
          8334 => x"746c0000",
          8335 => x"66696e69",
          8336 => x"74000000",
          8337 => x"666c6f61",
          8338 => x"64000000",
          8339 => x"66657865",
          8340 => x"63000000",
          8341 => x"6d636c65",
          8342 => x"61720000",
          8343 => x"6d64756d",
          8344 => x"70000000",
          8345 => x"6d656200",
          8346 => x"6d656800",
          8347 => x"6d657700",
          8348 => x"68696400",
          8349 => x"68696500",
          8350 => x"68666400",
          8351 => x"68666500",
          8352 => x"63616c6c",
          8353 => x"00000000",
          8354 => x"6a6d7000",
          8355 => x"72657374",
          8356 => x"61727400",
          8357 => x"72657365",
          8358 => x"74000000",
          8359 => x"696e666f",
          8360 => x"00000000",
          8361 => x"74657374",
          8362 => x"00000000",
          8363 => x"4469736b",
          8364 => x"20457272",
          8365 => x"6f720a00",
          8366 => x"496e7465",
          8367 => x"726e616c",
          8368 => x"20657272",
          8369 => x"6f722e0a",
          8370 => x"00000000",
          8371 => x"4469736b",
          8372 => x"206e6f74",
          8373 => x"20726561",
          8374 => x"64792e0a",
          8375 => x"00000000",
          8376 => x"4e6f2066",
          8377 => x"696c6520",
          8378 => x"666f756e",
          8379 => x"642e0a00",
          8380 => x"4e6f2070",
          8381 => x"61746820",
          8382 => x"666f756e",
          8383 => x"642e0a00",
          8384 => x"496e7661",
          8385 => x"6c696420",
          8386 => x"66696c65",
          8387 => x"6e616d65",
          8388 => x"2e0a0000",
          8389 => x"41636365",
          8390 => x"73732064",
          8391 => x"656e6965",
          8392 => x"642e0a00",
          8393 => x"46696c65",
          8394 => x"20616c72",
          8395 => x"65616479",
          8396 => x"20657869",
          8397 => x"7374732e",
          8398 => x"0a000000",
          8399 => x"46696c65",
          8400 => x"2068616e",
          8401 => x"646c6520",
          8402 => x"696e7661",
          8403 => x"6c69642e",
          8404 => x"0a000000",
          8405 => x"53442069",
          8406 => x"73207772",
          8407 => x"69746520",
          8408 => x"70726f74",
          8409 => x"65637465",
          8410 => x"642e0a00",
          8411 => x"44726976",
          8412 => x"65206e75",
          8413 => x"6d626572",
          8414 => x"20697320",
          8415 => x"696e7661",
          8416 => x"6c69642e",
          8417 => x"0a000000",
          8418 => x"4469736b",
          8419 => x"206e6f74",
          8420 => x"20656e61",
          8421 => x"626c6564",
          8422 => x"2e0a0000",
          8423 => x"4e6f2063",
          8424 => x"6f6d7061",
          8425 => x"7469626c",
          8426 => x"65206669",
          8427 => x"6c657379",
          8428 => x"7374656d",
          8429 => x"20666f75",
          8430 => x"6e64206f",
          8431 => x"6e206469",
          8432 => x"736b2e0a",
          8433 => x"00000000",
          8434 => x"466f726d",
          8435 => x"61742061",
          8436 => x"626f7274",
          8437 => x"65642e0a",
          8438 => x"00000000",
          8439 => x"54696d65",
          8440 => x"6f75742c",
          8441 => x"206f7065",
          8442 => x"72617469",
          8443 => x"6f6e2063",
          8444 => x"616e6365",
          8445 => x"6c6c6564",
          8446 => x"2e0a0000",
          8447 => x"46696c65",
          8448 => x"20697320",
          8449 => x"6c6f636b",
          8450 => x"65642e0a",
          8451 => x"00000000",
          8452 => x"496e7375",
          8453 => x"66666963",
          8454 => x"69656e74",
          8455 => x"206d656d",
          8456 => x"6f72792e",
          8457 => x"0a000000",
          8458 => x"546f6f20",
          8459 => x"6d616e79",
          8460 => x"206f7065",
          8461 => x"6e206669",
          8462 => x"6c65732e",
          8463 => x"0a000000",
          8464 => x"50617261",
          8465 => x"6d657465",
          8466 => x"72732069",
          8467 => x"6e636f72",
          8468 => x"72656374",
          8469 => x"2e0a0000",
          8470 => x"53756363",
          8471 => x"6573732e",
          8472 => x"0a000000",
          8473 => x"556e6b6e",
          8474 => x"6f776e20",
          8475 => x"6572726f",
          8476 => x"722e0a00",
          8477 => x"0a256c75",
          8478 => x"20627974",
          8479 => x"65732025",
          8480 => x"73206174",
          8481 => x"20256c75",
          8482 => x"20627974",
          8483 => x"65732f73",
          8484 => x"65632e0a",
          8485 => x"00000000",
          8486 => x"25303858",
          8487 => x"00000000",
          8488 => x"3a202000",
          8489 => x"25303458",
          8490 => x"00000000",
          8491 => x"20202020",
          8492 => x"20202020",
          8493 => x"00000000",
          8494 => x"25303258",
          8495 => x"00000000",
          8496 => x"20200000",
          8497 => x"207c0000",
          8498 => x"7c0d0a00",
          8499 => x"72656164",
          8500 => x"00000000",
          8501 => x"5a505554",
          8502 => x"41000000",
          8503 => x"0a2a2a20",
          8504 => x"25732028",
          8505 => x"00000000",
          8506 => x"31382f30",
          8507 => x"372f3230",
          8508 => x"31390000",
          8509 => x"76312e33",
          8510 => x"00000000",
          8511 => x"205a5055",
          8512 => x"2c207265",
          8513 => x"76202530",
          8514 => x"32782920",
          8515 => x"25732025",
          8516 => x"73202a2a",
          8517 => x"0a0a0000",
          8518 => x"5a505554",
          8519 => x"4120496e",
          8520 => x"74657272",
          8521 => x"75707420",
          8522 => x"48616e64",
          8523 => x"6c65720a",
          8524 => x"00000000",
          8525 => x"54696d65",
          8526 => x"7220696e",
          8527 => x"74657272",
          8528 => x"7570740a",
          8529 => x"00000000",
          8530 => x"50533220",
          8531 => x"696e7465",
          8532 => x"72727570",
          8533 => x"740a0000",
          8534 => x"494f4354",
          8535 => x"4c205244",
          8536 => x"20696e74",
          8537 => x"65727275",
          8538 => x"70740a00",
          8539 => x"494f4354",
          8540 => x"4c205752",
          8541 => x"20696e74",
          8542 => x"65727275",
          8543 => x"70740a00",
          8544 => x"55415254",
          8545 => x"30205258",
          8546 => x"20696e74",
          8547 => x"65727275",
          8548 => x"70740a00",
          8549 => x"55415254",
          8550 => x"30205458",
          8551 => x"20696e74",
          8552 => x"65727275",
          8553 => x"70740a00",
          8554 => x"55415254",
          8555 => x"31205258",
          8556 => x"20696e74",
          8557 => x"65727275",
          8558 => x"70740a00",
          8559 => x"55415254",
          8560 => x"31205458",
          8561 => x"20696e74",
          8562 => x"65727275",
          8563 => x"70740a00",
          8564 => x"53657474",
          8565 => x"696e6720",
          8566 => x"75702074",
          8567 => x"696d6572",
          8568 => x"2e2e2e0a",
          8569 => x"00000000",
          8570 => x"456e6162",
          8571 => x"6c696e67",
          8572 => x"2074696d",
          8573 => x"65722e2e",
          8574 => x"2e0a0000",
          8575 => x"303a0000",
          8576 => x"4661696c",
          8577 => x"65642074",
          8578 => x"6f20696e",
          8579 => x"69746961",
          8580 => x"6c697365",
          8581 => x"20736420",
          8582 => x"63617264",
          8583 => x"20302c20",
          8584 => x"706c6561",
          8585 => x"73652069",
          8586 => x"6e697420",
          8587 => x"6d616e75",
          8588 => x"616c6c79",
          8589 => x"2e0a0000",
          8590 => x"2a200000",
          8591 => x"42616420",
          8592 => x"6469736b",
          8593 => x"20696421",
          8594 => x"0a000000",
          8595 => x"496e6974",
          8596 => x"69616c69",
          8597 => x"7365642e",
          8598 => x"0a000000",
          8599 => x"4661696c",
          8600 => x"65642074",
          8601 => x"6f20696e",
          8602 => x"69746961",
          8603 => x"6c697365",
          8604 => x"2e0a0000",
          8605 => x"72633d25",
          8606 => x"640a0000",
          8607 => x"25753a00",
          8608 => x"436c6561",
          8609 => x"72696e67",
          8610 => x"2e2e2e00",
          8611 => x"44756d70",
          8612 => x"204d656d",
          8613 => x"6f72790a",
          8614 => x"00000000",
          8615 => x"0a436f6d",
          8616 => x"706c6574",
          8617 => x"652e0a00",
          8618 => x"25303858",
          8619 => x"20253032",
          8620 => x"582d0000",
          8621 => x"3f3f3f0a",
          8622 => x"00000000",
          8623 => x"25303858",
          8624 => x"20253034",
          8625 => x"582d0000",
          8626 => x"25303858",
          8627 => x"20253038",
          8628 => x"582d0000",
          8629 => x"44697361",
          8630 => x"626c696e",
          8631 => x"6720696e",
          8632 => x"74657272",
          8633 => x"75707473",
          8634 => x"0a000000",
          8635 => x"456e6162",
          8636 => x"6c696e67",
          8637 => x"20696e74",
          8638 => x"65727275",
          8639 => x"7074730a",
          8640 => x"00000000",
          8641 => x"44697361",
          8642 => x"626c6564",
          8643 => x"20756172",
          8644 => x"74206669",
          8645 => x"666f0a00",
          8646 => x"456e6162",
          8647 => x"6c696e67",
          8648 => x"20756172",
          8649 => x"74206669",
          8650 => x"666f0a00",
          8651 => x"45786563",
          8652 => x"7574696e",
          8653 => x"6720636f",
          8654 => x"64652040",
          8655 => x"20253038",
          8656 => x"78202e2e",
          8657 => x"2e0a0000",
          8658 => x"43616c6c",
          8659 => x"696e6720",
          8660 => x"636f6465",
          8661 => x"20402025",
          8662 => x"30387820",
          8663 => x"2e2e2e0a",
          8664 => x"00000000",
          8665 => x"43616c6c",
          8666 => x"20726574",
          8667 => x"75726e65",
          8668 => x"6420636f",
          8669 => x"64652028",
          8670 => x"2564292e",
          8671 => x"0a000000",
          8672 => x"52657374",
          8673 => x"61727469",
          8674 => x"6e672061",
          8675 => x"70706c69",
          8676 => x"63617469",
          8677 => x"6f6e2e2e",
          8678 => x"2e0a0000",
          8679 => x"436f6c64",
          8680 => x"20726562",
          8681 => x"6f6f7469",
          8682 => x"6e672e2e",
          8683 => x"2e0a0000",
          8684 => x"5a505500",
          8685 => x"62696e00",
          8686 => x"25643a5c",
          8687 => x"25735c25",
          8688 => x"732e2573",
          8689 => x"00000000",
          8690 => x"42616420",
          8691 => x"636f6d6d",
          8692 => x"616e642e",
          8693 => x"0a000000",
          8694 => x"52756e6e",
          8695 => x"696e672e",
          8696 => x"2e2e0a00",
          8697 => x"456e6162",
          8698 => x"6c696e67",
          8699 => x"20696e74",
          8700 => x"65727275",
          8701 => x"7074732e",
          8702 => x"2e2e0a00",
          8703 => x"00000000",
          8704 => x"00000000",
          8705 => x"00007fff",
          8706 => x"00000000",
          8707 => x"00007fff",
          8708 => x"00010000",
          8709 => x"00007fff",
          8710 => x"00000000",
          8711 => x"00000000",
          8712 => x"00007800",
          8713 => x"00000000",
          8714 => x"05f5e100",
          8715 => x"00010101",
          8716 => x"01010101",
          8717 => x"80010101",
          8718 => x"01000000",
          8719 => x"00000000",
          8720 => x"01000000",
          8721 => x"0000622c",
          8722 => x"01020100",
          8723 => x"00000000",
          8724 => x"00000000",
          8725 => x"00006234",
          8726 => x"01040100",
          8727 => x"00000000",
          8728 => x"00000000",
          8729 => x"0000623c",
          8730 => x"01140300",
          8731 => x"00000000",
          8732 => x"00000000",
          8733 => x"00006244",
          8734 => x"012b0300",
          8735 => x"00000000",
          8736 => x"00000000",
          8737 => x"0000624c",
          8738 => x"01300300",
          8739 => x"00000000",
          8740 => x"00000000",
          8741 => x"00006254",
          8742 => x"013c0400",
          8743 => x"00000000",
          8744 => x"00000000",
          8745 => x"0000625c",
          8746 => x"01400400",
          8747 => x"00000000",
          8748 => x"00000000",
          8749 => x"00006264",
          8750 => x"01410400",
          8751 => x"00000000",
          8752 => x"00000000",
          8753 => x"00006268",
          8754 => x"01420400",
          8755 => x"00000000",
          8756 => x"00000000",
          8757 => x"0000626c",
          8758 => x"01430400",
          8759 => x"00000000",
          8760 => x"00000000",
          8761 => x"00006270",
          8762 => x"01500500",
          8763 => x"00000000",
          8764 => x"00000000",
          8765 => x"00006274",
          8766 => x"01510500",
          8767 => x"00000000",
          8768 => x"00000000",
          8769 => x"00006278",
          8770 => x"01540500",
          8771 => x"00000000",
          8772 => x"00000000",
          8773 => x"0000627c",
          8774 => x"01550500",
          8775 => x"00000000",
          8776 => x"00000000",
          8777 => x"00006280",
          8778 => x"01790700",
          8779 => x"00000000",
          8780 => x"00000000",
          8781 => x"00006288",
          8782 => x"01780700",
          8783 => x"00000000",
          8784 => x"00000000",
          8785 => x"0000628c",
          8786 => x"01820800",
          8787 => x"00000000",
          8788 => x"00000000",
          8789 => x"00006294",
          8790 => x"01830800",
          8791 => x"00000000",
          8792 => x"00000000",
          8793 => x"0000629c",
          8794 => x"01850800",
          8795 => x"00000000",
          8796 => x"00000000",
          8797 => x"000062a4",
          8798 => x"01870800",
          8799 => x"00000000",
          8800 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;


end arch;

