-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBRAM;

architecture arch of SinglePortBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"a4",
             1 => x"0b",
             2 => x"04",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"a4",
             9 => x"0b",
            10 => x"04",
            11 => x"a4",
            12 => x"0b",
            13 => x"04",
            14 => x"a4",
            15 => x"0b",
            16 => x"04",
            17 => x"a4",
            18 => x"0b",
            19 => x"04",
            20 => x"a4",
            21 => x"0b",
            22 => x"04",
            23 => x"a5",
            24 => x"0b",
            25 => x"04",
            26 => x"a5",
            27 => x"0b",
            28 => x"04",
            29 => x"a5",
            30 => x"0b",
            31 => x"04",
            32 => x"a5",
            33 => x"0b",
            34 => x"04",
            35 => x"a6",
            36 => x"0b",
            37 => x"04",
            38 => x"a6",
            39 => x"0b",
            40 => x"04",
            41 => x"a6",
            42 => x"0b",
            43 => x"04",
            44 => x"a6",
            45 => x"0b",
            46 => x"04",
            47 => x"a7",
            48 => x"0b",
            49 => x"04",
            50 => x"a7",
            51 => x"0b",
            52 => x"04",
            53 => x"a7",
            54 => x"0b",
            55 => x"04",
            56 => x"a7",
            57 => x"0b",
            58 => x"04",
            59 => x"a8",
            60 => x"0b",
            61 => x"04",
            62 => x"a8",
            63 => x"0b",
            64 => x"04",
            65 => x"a8",
            66 => x"0b",
            67 => x"04",
            68 => x"a8",
            69 => x"0b",
            70 => x"04",
            71 => x"a9",
            72 => x"0b",
            73 => x"04",
            74 => x"a9",
            75 => x"0b",
            76 => x"04",
            77 => x"a9",
            78 => x"0b",
            79 => x"04",
            80 => x"a9",
            81 => x"0b",
            82 => x"04",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"04",
           129 => x"0c",
           130 => x"81",
           131 => x"83",
           132 => x"81",
           133 => x"80",
           134 => x"81",
           135 => x"83",
           136 => x"81",
           137 => x"80",
           138 => x"81",
           139 => x"83",
           140 => x"81",
           141 => x"80",
           142 => x"81",
           143 => x"83",
           144 => x"81",
           145 => x"80",
           146 => x"81",
           147 => x"83",
           148 => x"81",
           149 => x"80",
           150 => x"81",
           151 => x"83",
           152 => x"81",
           153 => x"80",
           154 => x"81",
           155 => x"83",
           156 => x"81",
           157 => x"80",
           158 => x"81",
           159 => x"83",
           160 => x"81",
           161 => x"80",
           162 => x"81",
           163 => x"83",
           164 => x"81",
           165 => x"80",
           166 => x"81",
           167 => x"83",
           168 => x"81",
           169 => x"80",
           170 => x"81",
           171 => x"83",
           172 => x"81",
           173 => x"80",
           174 => x"81",
           175 => x"83",
           176 => x"81",
           177 => x"b6",
           178 => x"ec",
           179 => x"80",
           180 => x"ec",
           181 => x"b1",
           182 => x"ec",
           183 => x"90",
           184 => x"ec",
           185 => x"2d",
           186 => x"08",
           187 => x"04",
           188 => x"0c",
           189 => x"81",
           190 => x"83",
           191 => x"81",
           192 => x"b2",
           193 => x"ec",
           194 => x"80",
           195 => x"ec",
           196 => x"fe",
           197 => x"ec",
           198 => x"80",
           199 => x"ec",
           200 => x"8b",
           201 => x"ec",
           202 => x"80",
           203 => x"ec",
           204 => x"83",
           205 => x"ec",
           206 => x"80",
           207 => x"ec",
           208 => x"86",
           209 => x"ec",
           210 => x"80",
           211 => x"ec",
           212 => x"90",
           213 => x"ec",
           214 => x"80",
           215 => x"ec",
           216 => x"99",
           217 => x"ec",
           218 => x"80",
           219 => x"ec",
           220 => x"89",
           221 => x"ec",
           222 => x"80",
           223 => x"ec",
           224 => x"93",
           225 => x"ec",
           226 => x"80",
           227 => x"ec",
           228 => x"94",
           229 => x"ec",
           230 => x"80",
           231 => x"ec",
           232 => x"95",
           233 => x"ec",
           234 => x"80",
           235 => x"ec",
           236 => x"9c",
           237 => x"ec",
           238 => x"80",
           239 => x"ec",
           240 => x"9a",
           241 => x"ec",
           242 => x"80",
           243 => x"ec",
           244 => x"9f",
           245 => x"ec",
           246 => x"80",
           247 => x"ec",
           248 => x"96",
           249 => x"ec",
           250 => x"80",
           251 => x"ec",
           252 => x"a2",
           253 => x"ec",
           254 => x"80",
           255 => x"ec",
           256 => x"a3",
           257 => x"ec",
           258 => x"80",
           259 => x"ec",
           260 => x"8b",
           261 => x"ec",
           262 => x"80",
           263 => x"ec",
           264 => x"8b",
           265 => x"ec",
           266 => x"80",
           267 => x"ec",
           268 => x"8c",
           269 => x"ec",
           270 => x"80",
           271 => x"ec",
           272 => x"96",
           273 => x"ec",
           274 => x"80",
           275 => x"ec",
           276 => x"a4",
           277 => x"ec",
           278 => x"80",
           279 => x"ec",
           280 => x"a6",
           281 => x"ec",
           282 => x"80",
           283 => x"ec",
           284 => x"a9",
           285 => x"ec",
           286 => x"80",
           287 => x"ec",
           288 => x"fd",
           289 => x"ec",
           290 => x"80",
           291 => x"ec",
           292 => x"ac",
           293 => x"ec",
           294 => x"80",
           295 => x"ec",
           296 => x"ce",
           297 => x"ec",
           298 => x"80",
           299 => x"ec",
           300 => x"d0",
           301 => x"ec",
           302 => x"80",
           303 => x"ec",
           304 => x"d2",
           305 => x"ec",
           306 => x"80",
           307 => x"ec",
           308 => x"f6",
           309 => x"ec",
           310 => x"90",
           311 => x"ec",
           312 => x"2d",
           313 => x"08",
           314 => x"04",
           315 => x"0c",
           316 => x"81",
           317 => x"83",
           318 => x"81",
           319 => x"81",
           320 => x"81",
           321 => x"83",
           322 => x"81",
           323 => x"82",
           324 => x"8e",
           325 => x"70",
           326 => x"0c",
           327 => x"aa",
           328 => x"80",
           329 => x"cc",
           330 => x"81",
           331 => x"02",
           332 => x"0c",
           333 => x"80",
           334 => x"ec",
           335 => x"08",
           336 => x"ec",
           337 => x"08",
           338 => x"3f",
           339 => x"08",
           340 => x"e0",
           341 => x"3d",
           342 => x"ec",
           343 => x"ec",
           344 => x"81",
           345 => x"fd",
           346 => x"53",
           347 => x"08",
           348 => x"52",
           349 => x"08",
           350 => x"51",
           351 => x"ec",
           352 => x"81",
           353 => x"54",
           354 => x"81",
           355 => x"04",
           356 => x"08",
           357 => x"ec",
           358 => x"0d",
           359 => x"ec",
           360 => x"05",
           361 => x"81",
           362 => x"f8",
           363 => x"ec",
           364 => x"05",
           365 => x"ec",
           366 => x"08",
           367 => x"81",
           368 => x"fc",
           369 => x"2e",
           370 => x"0b",
           371 => x"08",
           372 => x"24",
           373 => x"ec",
           374 => x"05",
           375 => x"ec",
           376 => x"05",
           377 => x"ec",
           378 => x"08",
           379 => x"ec",
           380 => x"0c",
           381 => x"81",
           382 => x"fc",
           383 => x"2e",
           384 => x"81",
           385 => x"8c",
           386 => x"ec",
           387 => x"05",
           388 => x"38",
           389 => x"08",
           390 => x"81",
           391 => x"8c",
           392 => x"81",
           393 => x"88",
           394 => x"ec",
           395 => x"05",
           396 => x"ec",
           397 => x"08",
           398 => x"ec",
           399 => x"0c",
           400 => x"08",
           401 => x"81",
           402 => x"ec",
           403 => x"0c",
           404 => x"08",
           405 => x"81",
           406 => x"ec",
           407 => x"0c",
           408 => x"81",
           409 => x"90",
           410 => x"2e",
           411 => x"ec",
           412 => x"05",
           413 => x"ec",
           414 => x"05",
           415 => x"39",
           416 => x"08",
           417 => x"70",
           418 => x"08",
           419 => x"51",
           420 => x"08",
           421 => x"81",
           422 => x"85",
           423 => x"ec",
           424 => x"fc",
           425 => x"79",
           426 => x"05",
           427 => x"57",
           428 => x"83",
           429 => x"38",
           430 => x"51",
           431 => x"a4",
           432 => x"52",
           433 => x"93",
           434 => x"70",
           435 => x"34",
           436 => x"71",
           437 => x"81",
           438 => x"74",
           439 => x"0c",
           440 => x"04",
           441 => x"2b",
           442 => x"71",
           443 => x"51",
           444 => x"72",
           445 => x"72",
           446 => x"05",
           447 => x"71",
           448 => x"53",
           449 => x"70",
           450 => x"0c",
           451 => x"84",
           452 => x"f0",
           453 => x"8f",
           454 => x"83",
           455 => x"38",
           456 => x"84",
           457 => x"fc",
           458 => x"83",
           459 => x"70",
           460 => x"39",
           461 => x"77",
           462 => x"07",
           463 => x"54",
           464 => x"38",
           465 => x"08",
           466 => x"71",
           467 => x"80",
           468 => x"75",
           469 => x"33",
           470 => x"06",
           471 => x"80",
           472 => x"72",
           473 => x"75",
           474 => x"06",
           475 => x"12",
           476 => x"33",
           477 => x"06",
           478 => x"52",
           479 => x"72",
           480 => x"81",
           481 => x"81",
           482 => x"71",
           483 => x"e0",
           484 => x"87",
           485 => x"71",
           486 => x"fb",
           487 => x"06",
           488 => x"82",
           489 => x"51",
           490 => x"97",
           491 => x"84",
           492 => x"54",
           493 => x"75",
           494 => x"38",
           495 => x"52",
           496 => x"80",
           497 => x"e0",
           498 => x"0d",
           499 => x"0d",
           500 => x"53",
           501 => x"52",
           502 => x"81",
           503 => x"81",
           504 => x"07",
           505 => x"52",
           506 => x"e8",
           507 => x"ec",
           508 => x"3d",
           509 => x"3d",
           510 => x"08",
           511 => x"56",
           512 => x"80",
           513 => x"33",
           514 => x"2e",
           515 => x"86",
           516 => x"52",
           517 => x"53",
           518 => x"13",
           519 => x"33",
           520 => x"06",
           521 => x"70",
           522 => x"38",
           523 => x"80",
           524 => x"74",
           525 => x"81",
           526 => x"70",
           527 => x"81",
           528 => x"80",
           529 => x"05",
           530 => x"76",
           531 => x"70",
           532 => x"0c",
           533 => x"04",
           534 => x"76",
           535 => x"80",
           536 => x"86",
           537 => x"52",
           538 => x"84",
           539 => x"e0",
           540 => x"80",
           541 => x"74",
           542 => x"ec",
           543 => x"3d",
           544 => x"3d",
           545 => x"11",
           546 => x"52",
           547 => x"70",
           548 => x"98",
           549 => x"33",
           550 => x"82",
           551 => x"26",
           552 => x"84",
           553 => x"83",
           554 => x"26",
           555 => x"85",
           556 => x"84",
           557 => x"26",
           558 => x"86",
           559 => x"85",
           560 => x"26",
           561 => x"88",
           562 => x"86",
           563 => x"e7",
           564 => x"38",
           565 => x"54",
           566 => x"87",
           567 => x"cc",
           568 => x"87",
           569 => x"0c",
           570 => x"c0",
           571 => x"82",
           572 => x"c0",
           573 => x"83",
           574 => x"c0",
           575 => x"84",
           576 => x"c0",
           577 => x"85",
           578 => x"c0",
           579 => x"86",
           580 => x"c0",
           581 => x"74",
           582 => x"a4",
           583 => x"c0",
           584 => x"80",
           585 => x"98",
           586 => x"52",
           587 => x"e0",
           588 => x"0d",
           589 => x"0d",
           590 => x"c0",
           591 => x"81",
           592 => x"c0",
           593 => x"5e",
           594 => x"87",
           595 => x"08",
           596 => x"1c",
           597 => x"98",
           598 => x"79",
           599 => x"87",
           600 => x"08",
           601 => x"1c",
           602 => x"98",
           603 => x"79",
           604 => x"87",
           605 => x"08",
           606 => x"1c",
           607 => x"98",
           608 => x"7b",
           609 => x"87",
           610 => x"08",
           611 => x"1c",
           612 => x"0c",
           613 => x"ff",
           614 => x"83",
           615 => x"58",
           616 => x"57",
           617 => x"56",
           618 => x"55",
           619 => x"54",
           620 => x"53",
           621 => x"ff",
           622 => x"d5",
           623 => x"c9",
           624 => x"0d",
           625 => x"0d",
           626 => x"33",
           627 => x"9f",
           628 => x"52",
           629 => x"81",
           630 => x"83",
           631 => x"fb",
           632 => x"0b",
           633 => x"88",
           634 => x"ff",
           635 => x"56",
           636 => x"84",
           637 => x"2e",
           638 => x"c0",
           639 => x"70",
           640 => x"2a",
           641 => x"53",
           642 => x"80",
           643 => x"71",
           644 => x"81",
           645 => x"70",
           646 => x"81",
           647 => x"06",
           648 => x"80",
           649 => x"71",
           650 => x"81",
           651 => x"70",
           652 => x"73",
           653 => x"51",
           654 => x"80",
           655 => x"2e",
           656 => x"c0",
           657 => x"75",
           658 => x"81",
           659 => x"87",
           660 => x"fb",
           661 => x"9f",
           662 => x"0b",
           663 => x"33",
           664 => x"06",
           665 => x"87",
           666 => x"51",
           667 => x"86",
           668 => x"94",
           669 => x"08",
           670 => x"70",
           671 => x"54",
           672 => x"2e",
           673 => x"91",
           674 => x"06",
           675 => x"d7",
           676 => x"32",
           677 => x"51",
           678 => x"2e",
           679 => x"93",
           680 => x"06",
           681 => x"ff",
           682 => x"81",
           683 => x"87",
           684 => x"52",
           685 => x"86",
           686 => x"94",
           687 => x"72",
           688 => x"0d",
           689 => x"0d",
           690 => x"74",
           691 => x"ff",
           692 => x"57",
           693 => x"80",
           694 => x"81",
           695 => x"15",
           696 => x"e9",
           697 => x"81",
           698 => x"57",
           699 => x"c0",
           700 => x"75",
           701 => x"38",
           702 => x"94",
           703 => x"70",
           704 => x"81",
           705 => x"52",
           706 => x"8c",
           707 => x"2a",
           708 => x"51",
           709 => x"38",
           710 => x"70",
           711 => x"51",
           712 => x"8d",
           713 => x"2a",
           714 => x"51",
           715 => x"be",
           716 => x"ff",
           717 => x"c0",
           718 => x"70",
           719 => x"38",
           720 => x"90",
           721 => x"0c",
           722 => x"33",
           723 => x"06",
           724 => x"70",
           725 => x"76",
           726 => x"0c",
           727 => x"04",
           728 => x"0b",
           729 => x"88",
           730 => x"ff",
           731 => x"87",
           732 => x"51",
           733 => x"86",
           734 => x"94",
           735 => x"08",
           736 => x"70",
           737 => x"51",
           738 => x"2e",
           739 => x"81",
           740 => x"87",
           741 => x"52",
           742 => x"86",
           743 => x"94",
           744 => x"08",
           745 => x"06",
           746 => x"0c",
           747 => x"0d",
           748 => x"0d",
           749 => x"e9",
           750 => x"81",
           751 => x"53",
           752 => x"84",
           753 => x"2e",
           754 => x"c0",
           755 => x"71",
           756 => x"2a",
           757 => x"51",
           758 => x"52",
           759 => x"a0",
           760 => x"ff",
           761 => x"c0",
           762 => x"70",
           763 => x"38",
           764 => x"90",
           765 => x"70",
           766 => x"98",
           767 => x"51",
           768 => x"e0",
           769 => x"0d",
           770 => x"0d",
           771 => x"80",
           772 => x"2a",
           773 => x"51",
           774 => x"84",
           775 => x"c0",
           776 => x"81",
           777 => x"87",
           778 => x"08",
           779 => x"0c",
           780 => x"94",
           781 => x"94",
           782 => x"9e",
           783 => x"e9",
           784 => x"c0",
           785 => x"81",
           786 => x"87",
           787 => x"08",
           788 => x"0c",
           789 => x"ac",
           790 => x"a4",
           791 => x"9e",
           792 => x"e9",
           793 => x"c0",
           794 => x"81",
           795 => x"87",
           796 => x"08",
           797 => x"0c",
           798 => x"bc",
           799 => x"b4",
           800 => x"9e",
           801 => x"e9",
           802 => x"c0",
           803 => x"81",
           804 => x"87",
           805 => x"08",
           806 => x"e9",
           807 => x"c0",
           808 => x"81",
           809 => x"87",
           810 => x"08",
           811 => x"0c",
           812 => x"8c",
           813 => x"cc",
           814 => x"81",
           815 => x"80",
           816 => x"9e",
           817 => x"84",
           818 => x"51",
           819 => x"80",
           820 => x"81",
           821 => x"e9",
           822 => x"0b",
           823 => x"90",
           824 => x"80",
           825 => x"52",
           826 => x"2e",
           827 => x"52",
           828 => x"d2",
           829 => x"87",
           830 => x"08",
           831 => x"0a",
           832 => x"52",
           833 => x"83",
           834 => x"71",
           835 => x"34",
           836 => x"c0",
           837 => x"70",
           838 => x"06",
           839 => x"70",
           840 => x"38",
           841 => x"81",
           842 => x"80",
           843 => x"9e",
           844 => x"a0",
           845 => x"51",
           846 => x"80",
           847 => x"81",
           848 => x"e9",
           849 => x"0b",
           850 => x"90",
           851 => x"80",
           852 => x"52",
           853 => x"2e",
           854 => x"52",
           855 => x"d6",
           856 => x"87",
           857 => x"08",
           858 => x"80",
           859 => x"52",
           860 => x"83",
           861 => x"71",
           862 => x"34",
           863 => x"c0",
           864 => x"70",
           865 => x"06",
           866 => x"70",
           867 => x"38",
           868 => x"81",
           869 => x"80",
           870 => x"9e",
           871 => x"81",
           872 => x"51",
           873 => x"80",
           874 => x"81",
           875 => x"e9",
           876 => x"0b",
           877 => x"90",
           878 => x"c0",
           879 => x"52",
           880 => x"2e",
           881 => x"52",
           882 => x"da",
           883 => x"87",
           884 => x"08",
           885 => x"06",
           886 => x"70",
           887 => x"38",
           888 => x"81",
           889 => x"87",
           890 => x"08",
           891 => x"06",
           892 => x"51",
           893 => x"81",
           894 => x"80",
           895 => x"9e",
           896 => x"84",
           897 => x"52",
           898 => x"2e",
           899 => x"52",
           900 => x"dd",
           901 => x"9e",
           902 => x"83",
           903 => x"84",
           904 => x"51",
           905 => x"de",
           906 => x"87",
           907 => x"08",
           908 => x"51",
           909 => x"80",
           910 => x"81",
           911 => x"e9",
           912 => x"c0",
           913 => x"70",
           914 => x"51",
           915 => x"e0",
           916 => x"0d",
           917 => x"0d",
           918 => x"51",
           919 => x"81",
           920 => x"54",
           921 => x"88",
           922 => x"8c",
           923 => x"3f",
           924 => x"51",
           925 => x"81",
           926 => x"54",
           927 => x"93",
           928 => x"ac",
           929 => x"b0",
           930 => x"52",
           931 => x"51",
           932 => x"81",
           933 => x"54",
           934 => x"93",
           935 => x"a4",
           936 => x"a8",
           937 => x"52",
           938 => x"51",
           939 => x"81",
           940 => x"54",
           941 => x"93",
           942 => x"8c",
           943 => x"90",
           944 => x"52",
           945 => x"51",
           946 => x"81",
           947 => x"54",
           948 => x"93",
           949 => x"94",
           950 => x"98",
           951 => x"52",
           952 => x"51",
           953 => x"81",
           954 => x"54",
           955 => x"93",
           956 => x"9c",
           957 => x"a0",
           958 => x"52",
           959 => x"51",
           960 => x"81",
           961 => x"54",
           962 => x"8d",
           963 => x"dc",
           964 => x"d7",
           965 => x"f1",
           966 => x"df",
           967 => x"80",
           968 => x"81",
           969 => x"52",
           970 => x"51",
           971 => x"81",
           972 => x"54",
           973 => x"8d",
           974 => x"de",
           975 => x"d8",
           976 => x"c5",
           977 => x"d1",
           978 => x"80",
           979 => x"81",
           980 => x"83",
           981 => x"e9",
           982 => x"73",
           983 => x"38",
           984 => x"51",
           985 => x"81",
           986 => x"54",
           987 => x"88",
           988 => x"c4",
           989 => x"3f",
           990 => x"33",
           991 => x"2e",
           992 => x"d8",
           993 => x"9d",
           994 => x"da",
           995 => x"80",
           996 => x"81",
           997 => x"83",
           998 => x"d8",
           999 => x"85",
          1000 => x"b4",
          1001 => x"d8",
          1002 => x"dd",
          1003 => x"b8",
          1004 => x"d9",
          1005 => x"d1",
          1006 => x"bc",
          1007 => x"d9",
          1008 => x"c5",
          1009 => x"ec",
          1010 => x"3f",
          1011 => x"22",
          1012 => x"f4",
          1013 => x"3f",
          1014 => x"08",
          1015 => x"c0",
          1016 => x"ea",
          1017 => x"ec",
          1018 => x"84",
          1019 => x"71",
          1020 => x"81",
          1021 => x"52",
          1022 => x"51",
          1023 => x"81",
          1024 => x"54",
          1025 => x"a8",
          1026 => x"c8",
          1027 => x"84",
          1028 => x"51",
          1029 => x"81",
          1030 => x"bd",
          1031 => x"76",
          1032 => x"54",
          1033 => x"08",
          1034 => x"c8",
          1035 => x"3f",
          1036 => x"33",
          1037 => x"2e",
          1038 => x"e9",
          1039 => x"bd",
          1040 => x"75",
          1041 => x"3f",
          1042 => x"08",
          1043 => x"29",
          1044 => x"54",
          1045 => x"e0",
          1046 => x"da",
          1047 => x"a9",
          1048 => x"d8",
          1049 => x"3f",
          1050 => x"04",
          1051 => x"02",
          1052 => x"ff",
          1053 => x"84",
          1054 => x"71",
          1055 => x"0b",
          1056 => x"05",
          1057 => x"04",
          1058 => x"51",
          1059 => x"db",
          1060 => x"39",
          1061 => x"51",
          1062 => x"db",
          1063 => x"39",
          1064 => x"51",
          1065 => x"db",
          1066 => x"f9",
          1067 => x"0d",
          1068 => x"80",
          1069 => x"0b",
          1070 => x"84",
          1071 => x"e9",
          1072 => x"c0",
          1073 => x"04",
          1074 => x"02",
          1075 => x"53",
          1076 => x"09",
          1077 => x"38",
          1078 => x"3f",
          1079 => x"08",
          1080 => x"2e",
          1081 => x"72",
          1082 => x"f8",
          1083 => x"81",
          1084 => x"8f",
          1085 => x"f0",
          1086 => x"80",
          1087 => x"72",
          1088 => x"84",
          1089 => x"fe",
          1090 => x"97",
          1091 => x"ec",
          1092 => x"81",
          1093 => x"54",
          1094 => x"3f",
          1095 => x"f0",
          1096 => x"0d",
          1097 => x"0d",
          1098 => x"33",
          1099 => x"06",
          1100 => x"80",
          1101 => x"72",
          1102 => x"51",
          1103 => x"ff",
          1104 => x"39",
          1105 => x"04",
          1106 => x"77",
          1107 => x"08",
          1108 => x"f0",
          1109 => x"73",
          1110 => x"ff",
          1111 => x"71",
          1112 => x"38",
          1113 => x"06",
          1114 => x"54",
          1115 => x"e7",
          1116 => x"ec",
          1117 => x"3d",
          1118 => x"3d",
          1119 => x"59",
          1120 => x"81",
          1121 => x"56",
          1122 => x"84",
          1123 => x"a5",
          1124 => x"06",
          1125 => x"80",
          1126 => x"81",
          1127 => x"58",
          1128 => x"b0",
          1129 => x"06",
          1130 => x"5a",
          1131 => x"ad",
          1132 => x"06",
          1133 => x"5a",
          1134 => x"05",
          1135 => x"75",
          1136 => x"81",
          1137 => x"77",
          1138 => x"08",
          1139 => x"05",
          1140 => x"5d",
          1141 => x"39",
          1142 => x"72",
          1143 => x"38",
          1144 => x"7b",
          1145 => x"05",
          1146 => x"70",
          1147 => x"33",
          1148 => x"39",
          1149 => x"32",
          1150 => x"72",
          1151 => x"78",
          1152 => x"70",
          1153 => x"07",
          1154 => x"07",
          1155 => x"51",
          1156 => x"80",
          1157 => x"79",
          1158 => x"70",
          1159 => x"33",
          1160 => x"80",
          1161 => x"38",
          1162 => x"e0",
          1163 => x"38",
          1164 => x"81",
          1165 => x"53",
          1166 => x"2e",
          1167 => x"73",
          1168 => x"a2",
          1169 => x"c3",
          1170 => x"38",
          1171 => x"24",
          1172 => x"80",
          1173 => x"8c",
          1174 => x"39",
          1175 => x"2e",
          1176 => x"81",
          1177 => x"80",
          1178 => x"80",
          1179 => x"d5",
          1180 => x"73",
          1181 => x"8e",
          1182 => x"39",
          1183 => x"2e",
          1184 => x"80",
          1185 => x"84",
          1186 => x"56",
          1187 => x"74",
          1188 => x"72",
          1189 => x"38",
          1190 => x"15",
          1191 => x"54",
          1192 => x"38",
          1193 => x"56",
          1194 => x"81",
          1195 => x"72",
          1196 => x"38",
          1197 => x"90",
          1198 => x"06",
          1199 => x"2e",
          1200 => x"51",
          1201 => x"74",
          1202 => x"53",
          1203 => x"fd",
          1204 => x"51",
          1205 => x"ef",
          1206 => x"19",
          1207 => x"53",
          1208 => x"39",
          1209 => x"39",
          1210 => x"39",
          1211 => x"39",
          1212 => x"39",
          1213 => x"d0",
          1214 => x"39",
          1215 => x"70",
          1216 => x"53",
          1217 => x"88",
          1218 => x"19",
          1219 => x"39",
          1220 => x"54",
          1221 => x"74",
          1222 => x"70",
          1223 => x"07",
          1224 => x"55",
          1225 => x"80",
          1226 => x"72",
          1227 => x"38",
          1228 => x"90",
          1229 => x"80",
          1230 => x"5e",
          1231 => x"74",
          1232 => x"3f",
          1233 => x"08",
          1234 => x"7c",
          1235 => x"54",
          1236 => x"81",
          1237 => x"55",
          1238 => x"92",
          1239 => x"53",
          1240 => x"2e",
          1241 => x"14",
          1242 => x"ff",
          1243 => x"14",
          1244 => x"70",
          1245 => x"34",
          1246 => x"30",
          1247 => x"9f",
          1248 => x"57",
          1249 => x"85",
          1250 => x"b1",
          1251 => x"2a",
          1252 => x"51",
          1253 => x"2e",
          1254 => x"3d",
          1255 => x"05",
          1256 => x"34",
          1257 => x"76",
          1258 => x"54",
          1259 => x"72",
          1260 => x"54",
          1261 => x"70",
          1262 => x"56",
          1263 => x"81",
          1264 => x"7b",
          1265 => x"73",
          1266 => x"3f",
          1267 => x"53",
          1268 => x"74",
          1269 => x"53",
          1270 => x"eb",
          1271 => x"77",
          1272 => x"53",
          1273 => x"14",
          1274 => x"54",
          1275 => x"3f",
          1276 => x"74",
          1277 => x"53",
          1278 => x"fb",
          1279 => x"51",
          1280 => x"ef",
          1281 => x"0d",
          1282 => x"0d",
          1283 => x"70",
          1284 => x"08",
          1285 => x"51",
          1286 => x"85",
          1287 => x"fe",
          1288 => x"81",
          1289 => x"85",
          1290 => x"52",
          1291 => x"ca",
          1292 => x"f8",
          1293 => x"73",
          1294 => x"81",
          1295 => x"84",
          1296 => x"fd",
          1297 => x"ec",
          1298 => x"81",
          1299 => x"87",
          1300 => x"53",
          1301 => x"fa",
          1302 => x"81",
          1303 => x"85",
          1304 => x"fb",
          1305 => x"79",
          1306 => x"08",
          1307 => x"57",
          1308 => x"71",
          1309 => x"e0",
          1310 => x"f4",
          1311 => x"2d",
          1312 => x"08",
          1313 => x"53",
          1314 => x"80",
          1315 => x"8d",
          1316 => x"72",
          1317 => x"30",
          1318 => x"51",
          1319 => x"80",
          1320 => x"71",
          1321 => x"38",
          1322 => x"97",
          1323 => x"25",
          1324 => x"16",
          1325 => x"25",
          1326 => x"14",
          1327 => x"34",
          1328 => x"72",
          1329 => x"3f",
          1330 => x"73",
          1331 => x"72",
          1332 => x"f7",
          1333 => x"53",
          1334 => x"e0",
          1335 => x"0d",
          1336 => x"0d",
          1337 => x"08",
          1338 => x"f4",
          1339 => x"76",
          1340 => x"ef",
          1341 => x"ec",
          1342 => x"3d",
          1343 => x"3d",
          1344 => x"5a",
          1345 => x"7a",
          1346 => x"08",
          1347 => x"53",
          1348 => x"09",
          1349 => x"38",
          1350 => x"0c",
          1351 => x"ad",
          1352 => x"06",
          1353 => x"76",
          1354 => x"0c",
          1355 => x"33",
          1356 => x"73",
          1357 => x"81",
          1358 => x"38",
          1359 => x"05",
          1360 => x"08",
          1361 => x"53",
          1362 => x"2e",
          1363 => x"57",
          1364 => x"2e",
          1365 => x"39",
          1366 => x"13",
          1367 => x"08",
          1368 => x"53",
          1369 => x"55",
          1370 => x"80",
          1371 => x"14",
          1372 => x"88",
          1373 => x"27",
          1374 => x"eb",
          1375 => x"53",
          1376 => x"89",
          1377 => x"38",
          1378 => x"55",
          1379 => x"8a",
          1380 => x"a0",
          1381 => x"c2",
          1382 => x"74",
          1383 => x"e0",
          1384 => x"ff",
          1385 => x"d0",
          1386 => x"ff",
          1387 => x"90",
          1388 => x"38",
          1389 => x"81",
          1390 => x"53",
          1391 => x"ca",
          1392 => x"27",
          1393 => x"77",
          1394 => x"08",
          1395 => x"0c",
          1396 => x"33",
          1397 => x"ff",
          1398 => x"80",
          1399 => x"74",
          1400 => x"79",
          1401 => x"74",
          1402 => x"0c",
          1403 => x"04",
          1404 => x"7a",
          1405 => x"80",
          1406 => x"58",
          1407 => x"33",
          1408 => x"a0",
          1409 => x"06",
          1410 => x"13",
          1411 => x"39",
          1412 => x"09",
          1413 => x"38",
          1414 => x"11",
          1415 => x"08",
          1416 => x"54",
          1417 => x"2e",
          1418 => x"80",
          1419 => x"08",
          1420 => x"0c",
          1421 => x"33",
          1422 => x"80",
          1423 => x"38",
          1424 => x"80",
          1425 => x"38",
          1426 => x"57",
          1427 => x"0c",
          1428 => x"33",
          1429 => x"39",
          1430 => x"74",
          1431 => x"38",
          1432 => x"80",
          1433 => x"89",
          1434 => x"38",
          1435 => x"d0",
          1436 => x"55",
          1437 => x"80",
          1438 => x"39",
          1439 => x"d9",
          1440 => x"80",
          1441 => x"27",
          1442 => x"80",
          1443 => x"89",
          1444 => x"70",
          1445 => x"55",
          1446 => x"70",
          1447 => x"55",
          1448 => x"27",
          1449 => x"14",
          1450 => x"06",
          1451 => x"74",
          1452 => x"73",
          1453 => x"38",
          1454 => x"14",
          1455 => x"05",
          1456 => x"08",
          1457 => x"54",
          1458 => x"39",
          1459 => x"84",
          1460 => x"55",
          1461 => x"81",
          1462 => x"ec",
          1463 => x"3d",
          1464 => x"3d",
          1465 => x"05",
          1466 => x"52",
          1467 => x"87",
          1468 => x"e8",
          1469 => x"71",
          1470 => x"0c",
          1471 => x"04",
          1472 => x"02",
          1473 => x"02",
          1474 => x"05",
          1475 => x"83",
          1476 => x"26",
          1477 => x"72",
          1478 => x"c0",
          1479 => x"53",
          1480 => x"74",
          1481 => x"38",
          1482 => x"73",
          1483 => x"c0",
          1484 => x"51",
          1485 => x"85",
          1486 => x"98",
          1487 => x"52",
          1488 => x"82",
          1489 => x"70",
          1490 => x"38",
          1491 => x"8c",
          1492 => x"ec",
          1493 => x"fc",
          1494 => x"52",
          1495 => x"87",
          1496 => x"08",
          1497 => x"2e",
          1498 => x"81",
          1499 => x"34",
          1500 => x"13",
          1501 => x"81",
          1502 => x"86",
          1503 => x"f3",
          1504 => x"62",
          1505 => x"05",
          1506 => x"57",
          1507 => x"83",
          1508 => x"fe",
          1509 => x"ec",
          1510 => x"06",
          1511 => x"71",
          1512 => x"71",
          1513 => x"2b",
          1514 => x"80",
          1515 => x"92",
          1516 => x"c0",
          1517 => x"41",
          1518 => x"5a",
          1519 => x"87",
          1520 => x"0c",
          1521 => x"84",
          1522 => x"08",
          1523 => x"70",
          1524 => x"53",
          1525 => x"2e",
          1526 => x"08",
          1527 => x"70",
          1528 => x"34",
          1529 => x"80",
          1530 => x"53",
          1531 => x"2e",
          1532 => x"53",
          1533 => x"26",
          1534 => x"80",
          1535 => x"87",
          1536 => x"08",
          1537 => x"38",
          1538 => x"8c",
          1539 => x"80",
          1540 => x"78",
          1541 => x"99",
          1542 => x"0c",
          1543 => x"8c",
          1544 => x"08",
          1545 => x"51",
          1546 => x"38",
          1547 => x"8d",
          1548 => x"17",
          1549 => x"81",
          1550 => x"53",
          1551 => x"2e",
          1552 => x"fc",
          1553 => x"52",
          1554 => x"7d",
          1555 => x"ed",
          1556 => x"80",
          1557 => x"71",
          1558 => x"38",
          1559 => x"53",
          1560 => x"e0",
          1561 => x"0d",
          1562 => x"0d",
          1563 => x"02",
          1564 => x"05",
          1565 => x"58",
          1566 => x"80",
          1567 => x"fc",
          1568 => x"ec",
          1569 => x"06",
          1570 => x"71",
          1571 => x"81",
          1572 => x"38",
          1573 => x"2b",
          1574 => x"80",
          1575 => x"92",
          1576 => x"c0",
          1577 => x"40",
          1578 => x"5a",
          1579 => x"c0",
          1580 => x"76",
          1581 => x"76",
          1582 => x"75",
          1583 => x"2a",
          1584 => x"51",
          1585 => x"80",
          1586 => x"7a",
          1587 => x"5c",
          1588 => x"81",
          1589 => x"81",
          1590 => x"06",
          1591 => x"80",
          1592 => x"87",
          1593 => x"08",
          1594 => x"38",
          1595 => x"8c",
          1596 => x"80",
          1597 => x"77",
          1598 => x"99",
          1599 => x"0c",
          1600 => x"8c",
          1601 => x"08",
          1602 => x"51",
          1603 => x"38",
          1604 => x"8d",
          1605 => x"70",
          1606 => x"84",
          1607 => x"5b",
          1608 => x"2e",
          1609 => x"fc",
          1610 => x"52",
          1611 => x"7d",
          1612 => x"f8",
          1613 => x"80",
          1614 => x"71",
          1615 => x"38",
          1616 => x"53",
          1617 => x"e0",
          1618 => x"0d",
          1619 => x"0d",
          1620 => x"05",
          1621 => x"02",
          1622 => x"05",
          1623 => x"54",
          1624 => x"fe",
          1625 => x"e0",
          1626 => x"53",
          1627 => x"80",
          1628 => x"0b",
          1629 => x"8c",
          1630 => x"71",
          1631 => x"dc",
          1632 => x"24",
          1633 => x"84",
          1634 => x"92",
          1635 => x"54",
          1636 => x"8d",
          1637 => x"39",
          1638 => x"80",
          1639 => x"cb",
          1640 => x"70",
          1641 => x"81",
          1642 => x"52",
          1643 => x"8a",
          1644 => x"98",
          1645 => x"71",
          1646 => x"c0",
          1647 => x"52",
          1648 => x"81",
          1649 => x"c0",
          1650 => x"53",
          1651 => x"82",
          1652 => x"71",
          1653 => x"39",
          1654 => x"39",
          1655 => x"77",
          1656 => x"81",
          1657 => x"72",
          1658 => x"84",
          1659 => x"73",
          1660 => x"0c",
          1661 => x"04",
          1662 => x"74",
          1663 => x"71",
          1664 => x"2b",
          1665 => x"e0",
          1666 => x"84",
          1667 => x"fd",
          1668 => x"83",
          1669 => x"12",
          1670 => x"2b",
          1671 => x"07",
          1672 => x"70",
          1673 => x"2b",
          1674 => x"07",
          1675 => x"0c",
          1676 => x"56",
          1677 => x"3d",
          1678 => x"3d",
          1679 => x"84",
          1680 => x"22",
          1681 => x"72",
          1682 => x"54",
          1683 => x"2a",
          1684 => x"34",
          1685 => x"04",
          1686 => x"73",
          1687 => x"70",
          1688 => x"05",
          1689 => x"88",
          1690 => x"72",
          1691 => x"54",
          1692 => x"2a",
          1693 => x"70",
          1694 => x"34",
          1695 => x"51",
          1696 => x"83",
          1697 => x"fe",
          1698 => x"75",
          1699 => x"51",
          1700 => x"92",
          1701 => x"81",
          1702 => x"73",
          1703 => x"55",
          1704 => x"51",
          1705 => x"3d",
          1706 => x"3d",
          1707 => x"76",
          1708 => x"72",
          1709 => x"05",
          1710 => x"11",
          1711 => x"38",
          1712 => x"04",
          1713 => x"78",
          1714 => x"56",
          1715 => x"81",
          1716 => x"74",
          1717 => x"56",
          1718 => x"31",
          1719 => x"52",
          1720 => x"80",
          1721 => x"71",
          1722 => x"38",
          1723 => x"e0",
          1724 => x"0d",
          1725 => x"0d",
          1726 => x"51",
          1727 => x"73",
          1728 => x"81",
          1729 => x"33",
          1730 => x"38",
          1731 => x"ec",
          1732 => x"3d",
          1733 => x"0b",
          1734 => x"0c",
          1735 => x"81",
          1736 => x"04",
          1737 => x"7b",
          1738 => x"83",
          1739 => x"5a",
          1740 => x"80",
          1741 => x"54",
          1742 => x"53",
          1743 => x"53",
          1744 => x"52",
          1745 => x"3f",
          1746 => x"08",
          1747 => x"81",
          1748 => x"81",
          1749 => x"83",
          1750 => x"16",
          1751 => x"18",
          1752 => x"18",
          1753 => x"58",
          1754 => x"9f",
          1755 => x"33",
          1756 => x"2e",
          1757 => x"93",
          1758 => x"76",
          1759 => x"52",
          1760 => x"51",
          1761 => x"83",
          1762 => x"79",
          1763 => x"0c",
          1764 => x"04",
          1765 => x"78",
          1766 => x"80",
          1767 => x"17",
          1768 => x"38",
          1769 => x"fc",
          1770 => x"e0",
          1771 => x"ec",
          1772 => x"38",
          1773 => x"53",
          1774 => x"81",
          1775 => x"f7",
          1776 => x"ec",
          1777 => x"2e",
          1778 => x"55",
          1779 => x"b0",
          1780 => x"81",
          1781 => x"88",
          1782 => x"f8",
          1783 => x"70",
          1784 => x"c0",
          1785 => x"e0",
          1786 => x"ec",
          1787 => x"91",
          1788 => x"55",
          1789 => x"09",
          1790 => x"f0",
          1791 => x"33",
          1792 => x"2e",
          1793 => x"80",
          1794 => x"80",
          1795 => x"e0",
          1796 => x"17",
          1797 => x"fd",
          1798 => x"d4",
          1799 => x"b2",
          1800 => x"96",
          1801 => x"85",
          1802 => x"75",
          1803 => x"3f",
          1804 => x"e4",
          1805 => x"98",
          1806 => x"9c",
          1807 => x"08",
          1808 => x"17",
          1809 => x"3f",
          1810 => x"52",
          1811 => x"51",
          1812 => x"a0",
          1813 => x"05",
          1814 => x"0c",
          1815 => x"75",
          1816 => x"33",
          1817 => x"3f",
          1818 => x"34",
          1819 => x"52",
          1820 => x"51",
          1821 => x"81",
          1822 => x"80",
          1823 => x"81",
          1824 => x"ec",
          1825 => x"3d",
          1826 => x"3d",
          1827 => x"1a",
          1828 => x"fe",
          1829 => x"54",
          1830 => x"73",
          1831 => x"8a",
          1832 => x"71",
          1833 => x"08",
          1834 => x"75",
          1835 => x"0c",
          1836 => x"04",
          1837 => x"7a",
          1838 => x"56",
          1839 => x"77",
          1840 => x"38",
          1841 => x"08",
          1842 => x"38",
          1843 => x"54",
          1844 => x"2e",
          1845 => x"72",
          1846 => x"38",
          1847 => x"8d",
          1848 => x"39",
          1849 => x"81",
          1850 => x"b6",
          1851 => x"2a",
          1852 => x"2a",
          1853 => x"05",
          1854 => x"55",
          1855 => x"81",
          1856 => x"81",
          1857 => x"83",
          1858 => x"b4",
          1859 => x"17",
          1860 => x"a4",
          1861 => x"55",
          1862 => x"57",
          1863 => x"3f",
          1864 => x"08",
          1865 => x"74",
          1866 => x"14",
          1867 => x"70",
          1868 => x"07",
          1869 => x"71",
          1870 => x"52",
          1871 => x"72",
          1872 => x"75",
          1873 => x"58",
          1874 => x"76",
          1875 => x"15",
          1876 => x"73",
          1877 => x"3f",
          1878 => x"08",
          1879 => x"76",
          1880 => x"06",
          1881 => x"05",
          1882 => x"3f",
          1883 => x"08",
          1884 => x"06",
          1885 => x"76",
          1886 => x"15",
          1887 => x"73",
          1888 => x"3f",
          1889 => x"08",
          1890 => x"82",
          1891 => x"06",
          1892 => x"05",
          1893 => x"3f",
          1894 => x"08",
          1895 => x"58",
          1896 => x"58",
          1897 => x"e0",
          1898 => x"0d",
          1899 => x"0d",
          1900 => x"5a",
          1901 => x"59",
          1902 => x"82",
          1903 => x"98",
          1904 => x"82",
          1905 => x"33",
          1906 => x"2e",
          1907 => x"72",
          1908 => x"38",
          1909 => x"8d",
          1910 => x"39",
          1911 => x"81",
          1912 => x"f7",
          1913 => x"2a",
          1914 => x"2a",
          1915 => x"05",
          1916 => x"55",
          1917 => x"81",
          1918 => x"59",
          1919 => x"08",
          1920 => x"74",
          1921 => x"16",
          1922 => x"16",
          1923 => x"59",
          1924 => x"53",
          1925 => x"8f",
          1926 => x"2b",
          1927 => x"74",
          1928 => x"71",
          1929 => x"72",
          1930 => x"0b",
          1931 => x"74",
          1932 => x"17",
          1933 => x"75",
          1934 => x"3f",
          1935 => x"08",
          1936 => x"e0",
          1937 => x"38",
          1938 => x"06",
          1939 => x"78",
          1940 => x"54",
          1941 => x"77",
          1942 => x"33",
          1943 => x"71",
          1944 => x"51",
          1945 => x"34",
          1946 => x"76",
          1947 => x"17",
          1948 => x"75",
          1949 => x"3f",
          1950 => x"08",
          1951 => x"e0",
          1952 => x"38",
          1953 => x"ff",
          1954 => x"10",
          1955 => x"76",
          1956 => x"51",
          1957 => x"be",
          1958 => x"2a",
          1959 => x"05",
          1960 => x"f9",
          1961 => x"ec",
          1962 => x"81",
          1963 => x"ab",
          1964 => x"0a",
          1965 => x"2b",
          1966 => x"70",
          1967 => x"70",
          1968 => x"54",
          1969 => x"81",
          1970 => x"8f",
          1971 => x"07",
          1972 => x"f7",
          1973 => x"0b",
          1974 => x"78",
          1975 => x"0c",
          1976 => x"04",
          1977 => x"7a",
          1978 => x"08",
          1979 => x"59",
          1980 => x"a4",
          1981 => x"17",
          1982 => x"38",
          1983 => x"aa",
          1984 => x"73",
          1985 => x"fd",
          1986 => x"ec",
          1987 => x"81",
          1988 => x"80",
          1989 => x"39",
          1990 => x"eb",
          1991 => x"80",
          1992 => x"ec",
          1993 => x"80",
          1994 => x"52",
          1995 => x"84",
          1996 => x"e0",
          1997 => x"ec",
          1998 => x"2e",
          1999 => x"81",
          2000 => x"81",
          2001 => x"81",
          2002 => x"ff",
          2003 => x"80",
          2004 => x"75",
          2005 => x"3f",
          2006 => x"08",
          2007 => x"16",
          2008 => x"90",
          2009 => x"55",
          2010 => x"27",
          2011 => x"15",
          2012 => x"84",
          2013 => x"07",
          2014 => x"17",
          2015 => x"76",
          2016 => x"a6",
          2017 => x"73",
          2018 => x"0c",
          2019 => x"04",
          2020 => x"7c",
          2021 => x"59",
          2022 => x"95",
          2023 => x"08",
          2024 => x"2e",
          2025 => x"17",
          2026 => x"b2",
          2027 => x"ae",
          2028 => x"7a",
          2029 => x"3f",
          2030 => x"81",
          2031 => x"27",
          2032 => x"81",
          2033 => x"55",
          2034 => x"08",
          2035 => x"d2",
          2036 => x"08",
          2037 => x"08",
          2038 => x"38",
          2039 => x"17",
          2040 => x"54",
          2041 => x"82",
          2042 => x"7a",
          2043 => x"06",
          2044 => x"81",
          2045 => x"17",
          2046 => x"83",
          2047 => x"75",
          2048 => x"f9",
          2049 => x"59",
          2050 => x"08",
          2051 => x"81",
          2052 => x"81",
          2053 => x"59",
          2054 => x"08",
          2055 => x"70",
          2056 => x"25",
          2057 => x"81",
          2058 => x"54",
          2059 => x"55",
          2060 => x"38",
          2061 => x"08",
          2062 => x"38",
          2063 => x"54",
          2064 => x"90",
          2065 => x"18",
          2066 => x"38",
          2067 => x"39",
          2068 => x"38",
          2069 => x"16",
          2070 => x"08",
          2071 => x"38",
          2072 => x"78",
          2073 => x"38",
          2074 => x"51",
          2075 => x"81",
          2076 => x"80",
          2077 => x"80",
          2078 => x"e0",
          2079 => x"09",
          2080 => x"38",
          2081 => x"08",
          2082 => x"e0",
          2083 => x"30",
          2084 => x"80",
          2085 => x"07",
          2086 => x"55",
          2087 => x"38",
          2088 => x"09",
          2089 => x"ae",
          2090 => x"80",
          2091 => x"53",
          2092 => x"51",
          2093 => x"81",
          2094 => x"81",
          2095 => x"30",
          2096 => x"e0",
          2097 => x"25",
          2098 => x"79",
          2099 => x"38",
          2100 => x"8f",
          2101 => x"79",
          2102 => x"f9",
          2103 => x"ec",
          2104 => x"74",
          2105 => x"8c",
          2106 => x"17",
          2107 => x"90",
          2108 => x"54",
          2109 => x"86",
          2110 => x"90",
          2111 => x"17",
          2112 => x"54",
          2113 => x"34",
          2114 => x"56",
          2115 => x"90",
          2116 => x"80",
          2117 => x"81",
          2118 => x"55",
          2119 => x"56",
          2120 => x"81",
          2121 => x"8c",
          2122 => x"f8",
          2123 => x"70",
          2124 => x"f0",
          2125 => x"e0",
          2126 => x"56",
          2127 => x"08",
          2128 => x"7b",
          2129 => x"f6",
          2130 => x"ec",
          2131 => x"ec",
          2132 => x"17",
          2133 => x"80",
          2134 => x"b4",
          2135 => x"57",
          2136 => x"77",
          2137 => x"81",
          2138 => x"15",
          2139 => x"78",
          2140 => x"81",
          2141 => x"53",
          2142 => x"15",
          2143 => x"e9",
          2144 => x"e0",
          2145 => x"df",
          2146 => x"22",
          2147 => x"30",
          2148 => x"70",
          2149 => x"51",
          2150 => x"81",
          2151 => x"8a",
          2152 => x"f8",
          2153 => x"7c",
          2154 => x"56",
          2155 => x"80",
          2156 => x"f1",
          2157 => x"06",
          2158 => x"e9",
          2159 => x"18",
          2160 => x"08",
          2161 => x"38",
          2162 => x"82",
          2163 => x"38",
          2164 => x"54",
          2165 => x"74",
          2166 => x"82",
          2167 => x"22",
          2168 => x"79",
          2169 => x"38",
          2170 => x"98",
          2171 => x"cd",
          2172 => x"22",
          2173 => x"54",
          2174 => x"26",
          2175 => x"52",
          2176 => x"b0",
          2177 => x"e0",
          2178 => x"ec",
          2179 => x"2e",
          2180 => x"0b",
          2181 => x"08",
          2182 => x"98",
          2183 => x"ec",
          2184 => x"85",
          2185 => x"bd",
          2186 => x"31",
          2187 => x"73",
          2188 => x"f4",
          2189 => x"ec",
          2190 => x"18",
          2191 => x"18",
          2192 => x"08",
          2193 => x"72",
          2194 => x"38",
          2195 => x"58",
          2196 => x"89",
          2197 => x"18",
          2198 => x"ff",
          2199 => x"05",
          2200 => x"80",
          2201 => x"ec",
          2202 => x"3d",
          2203 => x"3d",
          2204 => x"08",
          2205 => x"a0",
          2206 => x"54",
          2207 => x"77",
          2208 => x"80",
          2209 => x"0c",
          2210 => x"53",
          2211 => x"80",
          2212 => x"38",
          2213 => x"06",
          2214 => x"b5",
          2215 => x"98",
          2216 => x"14",
          2217 => x"92",
          2218 => x"2a",
          2219 => x"56",
          2220 => x"26",
          2221 => x"80",
          2222 => x"16",
          2223 => x"77",
          2224 => x"53",
          2225 => x"38",
          2226 => x"51",
          2227 => x"81",
          2228 => x"53",
          2229 => x"0b",
          2230 => x"08",
          2231 => x"38",
          2232 => x"ec",
          2233 => x"2e",
          2234 => x"98",
          2235 => x"ec",
          2236 => x"80",
          2237 => x"8a",
          2238 => x"15",
          2239 => x"80",
          2240 => x"14",
          2241 => x"51",
          2242 => x"81",
          2243 => x"53",
          2244 => x"ec",
          2245 => x"2e",
          2246 => x"82",
          2247 => x"e0",
          2248 => x"ba",
          2249 => x"81",
          2250 => x"ff",
          2251 => x"81",
          2252 => x"52",
          2253 => x"f3",
          2254 => x"e0",
          2255 => x"72",
          2256 => x"72",
          2257 => x"f2",
          2258 => x"ec",
          2259 => x"15",
          2260 => x"15",
          2261 => x"b4",
          2262 => x"0c",
          2263 => x"81",
          2264 => x"8a",
          2265 => x"f7",
          2266 => x"7d",
          2267 => x"5b",
          2268 => x"76",
          2269 => x"3f",
          2270 => x"08",
          2271 => x"e0",
          2272 => x"38",
          2273 => x"08",
          2274 => x"08",
          2275 => x"f0",
          2276 => x"ec",
          2277 => x"81",
          2278 => x"80",
          2279 => x"ec",
          2280 => x"18",
          2281 => x"51",
          2282 => x"81",
          2283 => x"81",
          2284 => x"81",
          2285 => x"e0",
          2286 => x"83",
          2287 => x"77",
          2288 => x"72",
          2289 => x"38",
          2290 => x"75",
          2291 => x"81",
          2292 => x"a5",
          2293 => x"e0",
          2294 => x"52",
          2295 => x"8e",
          2296 => x"e0",
          2297 => x"ec",
          2298 => x"2e",
          2299 => x"73",
          2300 => x"81",
          2301 => x"87",
          2302 => x"ec",
          2303 => x"3d",
          2304 => x"3d",
          2305 => x"11",
          2306 => x"ec",
          2307 => x"e0",
          2308 => x"ff",
          2309 => x"33",
          2310 => x"71",
          2311 => x"81",
          2312 => x"94",
          2313 => x"d0",
          2314 => x"e0",
          2315 => x"73",
          2316 => x"81",
          2317 => x"85",
          2318 => x"fc",
          2319 => x"79",
          2320 => x"ff",
          2321 => x"12",
          2322 => x"eb",
          2323 => x"70",
          2324 => x"72",
          2325 => x"81",
          2326 => x"73",
          2327 => x"94",
          2328 => x"d6",
          2329 => x"0d",
          2330 => x"0d",
          2331 => x"55",
          2332 => x"5a",
          2333 => x"08",
          2334 => x"8a",
          2335 => x"08",
          2336 => x"ee",
          2337 => x"ec",
          2338 => x"81",
          2339 => x"80",
          2340 => x"15",
          2341 => x"55",
          2342 => x"38",
          2343 => x"e6",
          2344 => x"33",
          2345 => x"70",
          2346 => x"58",
          2347 => x"86",
          2348 => x"ec",
          2349 => x"73",
          2350 => x"83",
          2351 => x"73",
          2352 => x"38",
          2353 => x"06",
          2354 => x"80",
          2355 => x"75",
          2356 => x"38",
          2357 => x"08",
          2358 => x"54",
          2359 => x"2e",
          2360 => x"83",
          2361 => x"73",
          2362 => x"38",
          2363 => x"51",
          2364 => x"81",
          2365 => x"58",
          2366 => x"08",
          2367 => x"15",
          2368 => x"38",
          2369 => x"0b",
          2370 => x"77",
          2371 => x"0c",
          2372 => x"04",
          2373 => x"77",
          2374 => x"54",
          2375 => x"51",
          2376 => x"81",
          2377 => x"55",
          2378 => x"08",
          2379 => x"14",
          2380 => x"51",
          2381 => x"81",
          2382 => x"55",
          2383 => x"08",
          2384 => x"53",
          2385 => x"08",
          2386 => x"08",
          2387 => x"3f",
          2388 => x"14",
          2389 => x"08",
          2390 => x"3f",
          2391 => x"17",
          2392 => x"ec",
          2393 => x"3d",
          2394 => x"3d",
          2395 => x"08",
          2396 => x"54",
          2397 => x"53",
          2398 => x"81",
          2399 => x"8d",
          2400 => x"08",
          2401 => x"34",
          2402 => x"15",
          2403 => x"0d",
          2404 => x"0d",
          2405 => x"57",
          2406 => x"17",
          2407 => x"08",
          2408 => x"82",
          2409 => x"89",
          2410 => x"55",
          2411 => x"14",
          2412 => x"16",
          2413 => x"71",
          2414 => x"38",
          2415 => x"09",
          2416 => x"38",
          2417 => x"73",
          2418 => x"81",
          2419 => x"ae",
          2420 => x"05",
          2421 => x"15",
          2422 => x"70",
          2423 => x"34",
          2424 => x"8a",
          2425 => x"38",
          2426 => x"05",
          2427 => x"81",
          2428 => x"17",
          2429 => x"12",
          2430 => x"34",
          2431 => x"9c",
          2432 => x"e8",
          2433 => x"ec",
          2434 => x"0c",
          2435 => x"e7",
          2436 => x"ec",
          2437 => x"17",
          2438 => x"51",
          2439 => x"81",
          2440 => x"84",
          2441 => x"3d",
          2442 => x"3d",
          2443 => x"08",
          2444 => x"61",
          2445 => x"55",
          2446 => x"2e",
          2447 => x"55",
          2448 => x"2e",
          2449 => x"80",
          2450 => x"94",
          2451 => x"1c",
          2452 => x"81",
          2453 => x"61",
          2454 => x"56",
          2455 => x"2e",
          2456 => x"83",
          2457 => x"73",
          2458 => x"70",
          2459 => x"25",
          2460 => x"51",
          2461 => x"38",
          2462 => x"0c",
          2463 => x"51",
          2464 => x"26",
          2465 => x"80",
          2466 => x"34",
          2467 => x"51",
          2468 => x"81",
          2469 => x"55",
          2470 => x"91",
          2471 => x"1d",
          2472 => x"8b",
          2473 => x"79",
          2474 => x"3f",
          2475 => x"57",
          2476 => x"55",
          2477 => x"2e",
          2478 => x"80",
          2479 => x"18",
          2480 => x"1a",
          2481 => x"70",
          2482 => x"2a",
          2483 => x"07",
          2484 => x"5a",
          2485 => x"8c",
          2486 => x"54",
          2487 => x"81",
          2488 => x"39",
          2489 => x"70",
          2490 => x"2a",
          2491 => x"75",
          2492 => x"8c",
          2493 => x"2e",
          2494 => x"a0",
          2495 => x"38",
          2496 => x"0c",
          2497 => x"76",
          2498 => x"38",
          2499 => x"b8",
          2500 => x"70",
          2501 => x"5a",
          2502 => x"76",
          2503 => x"38",
          2504 => x"70",
          2505 => x"dc",
          2506 => x"72",
          2507 => x"80",
          2508 => x"51",
          2509 => x"73",
          2510 => x"38",
          2511 => x"18",
          2512 => x"1a",
          2513 => x"55",
          2514 => x"2e",
          2515 => x"83",
          2516 => x"73",
          2517 => x"70",
          2518 => x"25",
          2519 => x"51",
          2520 => x"38",
          2521 => x"75",
          2522 => x"81",
          2523 => x"81",
          2524 => x"27",
          2525 => x"73",
          2526 => x"38",
          2527 => x"70",
          2528 => x"32",
          2529 => x"80",
          2530 => x"2a",
          2531 => x"56",
          2532 => x"81",
          2533 => x"57",
          2534 => x"f5",
          2535 => x"2b",
          2536 => x"25",
          2537 => x"80",
          2538 => x"dc",
          2539 => x"57",
          2540 => x"e6",
          2541 => x"ec",
          2542 => x"2e",
          2543 => x"18",
          2544 => x"1a",
          2545 => x"56",
          2546 => x"3f",
          2547 => x"08",
          2548 => x"e8",
          2549 => x"54",
          2550 => x"80",
          2551 => x"17",
          2552 => x"34",
          2553 => x"11",
          2554 => x"74",
          2555 => x"75",
          2556 => x"d0",
          2557 => x"3f",
          2558 => x"08",
          2559 => x"9f",
          2560 => x"99",
          2561 => x"e0",
          2562 => x"ff",
          2563 => x"79",
          2564 => x"74",
          2565 => x"57",
          2566 => x"77",
          2567 => x"76",
          2568 => x"38",
          2569 => x"73",
          2570 => x"09",
          2571 => x"38",
          2572 => x"84",
          2573 => x"27",
          2574 => x"39",
          2575 => x"f2",
          2576 => x"80",
          2577 => x"54",
          2578 => x"34",
          2579 => x"58",
          2580 => x"f2",
          2581 => x"ec",
          2582 => x"81",
          2583 => x"80",
          2584 => x"1b",
          2585 => x"51",
          2586 => x"81",
          2587 => x"56",
          2588 => x"08",
          2589 => x"9c",
          2590 => x"33",
          2591 => x"80",
          2592 => x"38",
          2593 => x"bf",
          2594 => x"86",
          2595 => x"15",
          2596 => x"2a",
          2597 => x"51",
          2598 => x"92",
          2599 => x"79",
          2600 => x"e4",
          2601 => x"ec",
          2602 => x"2e",
          2603 => x"52",
          2604 => x"ba",
          2605 => x"39",
          2606 => x"33",
          2607 => x"80",
          2608 => x"74",
          2609 => x"81",
          2610 => x"38",
          2611 => x"70",
          2612 => x"82",
          2613 => x"54",
          2614 => x"96",
          2615 => x"06",
          2616 => x"2e",
          2617 => x"ff",
          2618 => x"1c",
          2619 => x"80",
          2620 => x"81",
          2621 => x"ba",
          2622 => x"b6",
          2623 => x"2a",
          2624 => x"51",
          2625 => x"38",
          2626 => x"70",
          2627 => x"81",
          2628 => x"55",
          2629 => x"e1",
          2630 => x"08",
          2631 => x"1d",
          2632 => x"7c",
          2633 => x"3f",
          2634 => x"08",
          2635 => x"fa",
          2636 => x"81",
          2637 => x"8f",
          2638 => x"f6",
          2639 => x"5b",
          2640 => x"70",
          2641 => x"59",
          2642 => x"73",
          2643 => x"c6",
          2644 => x"81",
          2645 => x"70",
          2646 => x"52",
          2647 => x"8d",
          2648 => x"38",
          2649 => x"09",
          2650 => x"a5",
          2651 => x"d0",
          2652 => x"ff",
          2653 => x"53",
          2654 => x"91",
          2655 => x"73",
          2656 => x"d0",
          2657 => x"71",
          2658 => x"f7",
          2659 => x"81",
          2660 => x"55",
          2661 => x"55",
          2662 => x"81",
          2663 => x"74",
          2664 => x"56",
          2665 => x"12",
          2666 => x"70",
          2667 => x"38",
          2668 => x"81",
          2669 => x"51",
          2670 => x"51",
          2671 => x"89",
          2672 => x"70",
          2673 => x"53",
          2674 => x"70",
          2675 => x"51",
          2676 => x"09",
          2677 => x"38",
          2678 => x"38",
          2679 => x"77",
          2680 => x"70",
          2681 => x"2a",
          2682 => x"07",
          2683 => x"51",
          2684 => x"8f",
          2685 => x"84",
          2686 => x"83",
          2687 => x"94",
          2688 => x"74",
          2689 => x"38",
          2690 => x"0c",
          2691 => x"86",
          2692 => x"90",
          2693 => x"81",
          2694 => x"8c",
          2695 => x"fa",
          2696 => x"56",
          2697 => x"17",
          2698 => x"b0",
          2699 => x"52",
          2700 => x"e0",
          2701 => x"81",
          2702 => x"81",
          2703 => x"b2",
          2704 => x"b4",
          2705 => x"e0",
          2706 => x"ff",
          2707 => x"55",
          2708 => x"d5",
          2709 => x"06",
          2710 => x"80",
          2711 => x"33",
          2712 => x"81",
          2713 => x"81",
          2714 => x"81",
          2715 => x"eb",
          2716 => x"70",
          2717 => x"07",
          2718 => x"73",
          2719 => x"81",
          2720 => x"81",
          2721 => x"83",
          2722 => x"e0",
          2723 => x"16",
          2724 => x"3f",
          2725 => x"08",
          2726 => x"e0",
          2727 => x"9d",
          2728 => x"81",
          2729 => x"81",
          2730 => x"e0",
          2731 => x"ec",
          2732 => x"81",
          2733 => x"80",
          2734 => x"82",
          2735 => x"ec",
          2736 => x"3d",
          2737 => x"3d",
          2738 => x"84",
          2739 => x"05",
          2740 => x"80",
          2741 => x"51",
          2742 => x"81",
          2743 => x"58",
          2744 => x"0b",
          2745 => x"08",
          2746 => x"38",
          2747 => x"08",
          2748 => x"ec",
          2749 => x"08",
          2750 => x"56",
          2751 => x"86",
          2752 => x"75",
          2753 => x"fe",
          2754 => x"54",
          2755 => x"2e",
          2756 => x"14",
          2757 => x"ca",
          2758 => x"e0",
          2759 => x"06",
          2760 => x"54",
          2761 => x"38",
          2762 => x"86",
          2763 => x"82",
          2764 => x"06",
          2765 => x"56",
          2766 => x"38",
          2767 => x"80",
          2768 => x"81",
          2769 => x"52",
          2770 => x"51",
          2771 => x"81",
          2772 => x"81",
          2773 => x"81",
          2774 => x"83",
          2775 => x"87",
          2776 => x"2e",
          2777 => x"82",
          2778 => x"06",
          2779 => x"56",
          2780 => x"38",
          2781 => x"74",
          2782 => x"a3",
          2783 => x"e0",
          2784 => x"06",
          2785 => x"2e",
          2786 => x"80",
          2787 => x"3d",
          2788 => x"83",
          2789 => x"15",
          2790 => x"53",
          2791 => x"8d",
          2792 => x"15",
          2793 => x"3f",
          2794 => x"08",
          2795 => x"70",
          2796 => x"0c",
          2797 => x"16",
          2798 => x"80",
          2799 => x"80",
          2800 => x"54",
          2801 => x"84",
          2802 => x"5b",
          2803 => x"80",
          2804 => x"7a",
          2805 => x"fc",
          2806 => x"ec",
          2807 => x"ff",
          2808 => x"77",
          2809 => x"81",
          2810 => x"76",
          2811 => x"81",
          2812 => x"2e",
          2813 => x"8d",
          2814 => x"26",
          2815 => x"bf",
          2816 => x"f4",
          2817 => x"e0",
          2818 => x"ff",
          2819 => x"84",
          2820 => x"81",
          2821 => x"38",
          2822 => x"51",
          2823 => x"81",
          2824 => x"83",
          2825 => x"58",
          2826 => x"80",
          2827 => x"db",
          2828 => x"ec",
          2829 => x"77",
          2830 => x"80",
          2831 => x"82",
          2832 => x"c4",
          2833 => x"11",
          2834 => x"06",
          2835 => x"8d",
          2836 => x"26",
          2837 => x"74",
          2838 => x"78",
          2839 => x"c1",
          2840 => x"59",
          2841 => x"15",
          2842 => x"2e",
          2843 => x"13",
          2844 => x"72",
          2845 => x"38",
          2846 => x"eb",
          2847 => x"14",
          2848 => x"3f",
          2849 => x"08",
          2850 => x"e0",
          2851 => x"23",
          2852 => x"57",
          2853 => x"83",
          2854 => x"c7",
          2855 => x"d8",
          2856 => x"e0",
          2857 => x"ff",
          2858 => x"8d",
          2859 => x"14",
          2860 => x"3f",
          2861 => x"08",
          2862 => x"14",
          2863 => x"3f",
          2864 => x"08",
          2865 => x"06",
          2866 => x"72",
          2867 => x"97",
          2868 => x"22",
          2869 => x"84",
          2870 => x"5a",
          2871 => x"83",
          2872 => x"14",
          2873 => x"79",
          2874 => x"b0",
          2875 => x"ec",
          2876 => x"81",
          2877 => x"80",
          2878 => x"38",
          2879 => x"08",
          2880 => x"ff",
          2881 => x"38",
          2882 => x"83",
          2883 => x"83",
          2884 => x"74",
          2885 => x"85",
          2886 => x"89",
          2887 => x"76",
          2888 => x"c3",
          2889 => x"70",
          2890 => x"7b",
          2891 => x"73",
          2892 => x"17",
          2893 => x"ac",
          2894 => x"55",
          2895 => x"09",
          2896 => x"38",
          2897 => x"51",
          2898 => x"81",
          2899 => x"83",
          2900 => x"53",
          2901 => x"82",
          2902 => x"82",
          2903 => x"e0",
          2904 => x"ab",
          2905 => x"e0",
          2906 => x"0c",
          2907 => x"53",
          2908 => x"56",
          2909 => x"81",
          2910 => x"13",
          2911 => x"74",
          2912 => x"82",
          2913 => x"74",
          2914 => x"81",
          2915 => x"06",
          2916 => x"83",
          2917 => x"2a",
          2918 => x"72",
          2919 => x"26",
          2920 => x"ff",
          2921 => x"0c",
          2922 => x"15",
          2923 => x"0b",
          2924 => x"76",
          2925 => x"81",
          2926 => x"38",
          2927 => x"51",
          2928 => x"81",
          2929 => x"83",
          2930 => x"53",
          2931 => x"09",
          2932 => x"f9",
          2933 => x"52",
          2934 => x"b8",
          2935 => x"e0",
          2936 => x"38",
          2937 => x"08",
          2938 => x"84",
          2939 => x"d8",
          2940 => x"ec",
          2941 => x"ff",
          2942 => x"72",
          2943 => x"2e",
          2944 => x"80",
          2945 => x"14",
          2946 => x"3f",
          2947 => x"08",
          2948 => x"a4",
          2949 => x"81",
          2950 => x"84",
          2951 => x"d7",
          2952 => x"ec",
          2953 => x"8a",
          2954 => x"2e",
          2955 => x"9d",
          2956 => x"14",
          2957 => x"3f",
          2958 => x"08",
          2959 => x"84",
          2960 => x"d7",
          2961 => x"ec",
          2962 => x"15",
          2963 => x"34",
          2964 => x"22",
          2965 => x"72",
          2966 => x"23",
          2967 => x"23",
          2968 => x"15",
          2969 => x"75",
          2970 => x"0c",
          2971 => x"04",
          2972 => x"77",
          2973 => x"73",
          2974 => x"38",
          2975 => x"72",
          2976 => x"38",
          2977 => x"71",
          2978 => x"38",
          2979 => x"84",
          2980 => x"52",
          2981 => x"09",
          2982 => x"38",
          2983 => x"51",
          2984 => x"81",
          2985 => x"81",
          2986 => x"88",
          2987 => x"08",
          2988 => x"39",
          2989 => x"73",
          2990 => x"74",
          2991 => x"0c",
          2992 => x"04",
          2993 => x"02",
          2994 => x"7a",
          2995 => x"fc",
          2996 => x"f4",
          2997 => x"54",
          2998 => x"ec",
          2999 => x"bc",
          3000 => x"e0",
          3001 => x"81",
          3002 => x"70",
          3003 => x"73",
          3004 => x"38",
          3005 => x"78",
          3006 => x"2e",
          3007 => x"74",
          3008 => x"0c",
          3009 => x"80",
          3010 => x"80",
          3011 => x"70",
          3012 => x"51",
          3013 => x"81",
          3014 => x"54",
          3015 => x"e0",
          3016 => x"0d",
          3017 => x"0d",
          3018 => x"05",
          3019 => x"33",
          3020 => x"54",
          3021 => x"84",
          3022 => x"bf",
          3023 => x"98",
          3024 => x"53",
          3025 => x"05",
          3026 => x"fa",
          3027 => x"e0",
          3028 => x"ec",
          3029 => x"a4",
          3030 => x"68",
          3031 => x"70",
          3032 => x"c6",
          3033 => x"e0",
          3034 => x"ec",
          3035 => x"38",
          3036 => x"05",
          3037 => x"2b",
          3038 => x"80",
          3039 => x"86",
          3040 => x"06",
          3041 => x"2e",
          3042 => x"74",
          3043 => x"38",
          3044 => x"09",
          3045 => x"38",
          3046 => x"f8",
          3047 => x"e0",
          3048 => x"39",
          3049 => x"33",
          3050 => x"73",
          3051 => x"77",
          3052 => x"81",
          3053 => x"73",
          3054 => x"38",
          3055 => x"bc",
          3056 => x"07",
          3057 => x"b4",
          3058 => x"2a",
          3059 => x"51",
          3060 => x"2e",
          3061 => x"62",
          3062 => x"e8",
          3063 => x"ec",
          3064 => x"82",
          3065 => x"52",
          3066 => x"51",
          3067 => x"62",
          3068 => x"8b",
          3069 => x"53",
          3070 => x"51",
          3071 => x"80",
          3072 => x"05",
          3073 => x"3f",
          3074 => x"0b",
          3075 => x"75",
          3076 => x"f1",
          3077 => x"11",
          3078 => x"80",
          3079 => x"97",
          3080 => x"51",
          3081 => x"81",
          3082 => x"55",
          3083 => x"08",
          3084 => x"b7",
          3085 => x"c4",
          3086 => x"05",
          3087 => x"2a",
          3088 => x"51",
          3089 => x"80",
          3090 => x"84",
          3091 => x"39",
          3092 => x"70",
          3093 => x"54",
          3094 => x"a9",
          3095 => x"06",
          3096 => x"2e",
          3097 => x"55",
          3098 => x"73",
          3099 => x"d6",
          3100 => x"ec",
          3101 => x"ff",
          3102 => x"0c",
          3103 => x"ec",
          3104 => x"f8",
          3105 => x"2a",
          3106 => x"51",
          3107 => x"2e",
          3108 => x"80",
          3109 => x"7a",
          3110 => x"a0",
          3111 => x"a4",
          3112 => x"53",
          3113 => x"e6",
          3114 => x"ec",
          3115 => x"ec",
          3116 => x"1b",
          3117 => x"05",
          3118 => x"d3",
          3119 => x"e0",
          3120 => x"e0",
          3121 => x"0c",
          3122 => x"56",
          3123 => x"84",
          3124 => x"90",
          3125 => x"0b",
          3126 => x"80",
          3127 => x"0c",
          3128 => x"1a",
          3129 => x"2a",
          3130 => x"51",
          3131 => x"2e",
          3132 => x"81",
          3133 => x"80",
          3134 => x"38",
          3135 => x"08",
          3136 => x"8a",
          3137 => x"89",
          3138 => x"59",
          3139 => x"76",
          3140 => x"d7",
          3141 => x"ec",
          3142 => x"81",
          3143 => x"81",
          3144 => x"82",
          3145 => x"e0",
          3146 => x"09",
          3147 => x"38",
          3148 => x"78",
          3149 => x"30",
          3150 => x"80",
          3151 => x"77",
          3152 => x"38",
          3153 => x"06",
          3154 => x"c3",
          3155 => x"1a",
          3156 => x"38",
          3157 => x"06",
          3158 => x"2e",
          3159 => x"52",
          3160 => x"a6",
          3161 => x"e0",
          3162 => x"82",
          3163 => x"75",
          3164 => x"ec",
          3165 => x"9c",
          3166 => x"39",
          3167 => x"74",
          3168 => x"ec",
          3169 => x"3d",
          3170 => x"3d",
          3171 => x"65",
          3172 => x"5d",
          3173 => x"0c",
          3174 => x"05",
          3175 => x"f9",
          3176 => x"ec",
          3177 => x"81",
          3178 => x"8a",
          3179 => x"33",
          3180 => x"2e",
          3181 => x"56",
          3182 => x"90",
          3183 => x"06",
          3184 => x"74",
          3185 => x"b6",
          3186 => x"82",
          3187 => x"34",
          3188 => x"aa",
          3189 => x"91",
          3190 => x"56",
          3191 => x"8c",
          3192 => x"1a",
          3193 => x"74",
          3194 => x"38",
          3195 => x"80",
          3196 => x"38",
          3197 => x"70",
          3198 => x"56",
          3199 => x"b2",
          3200 => x"11",
          3201 => x"77",
          3202 => x"5b",
          3203 => x"38",
          3204 => x"88",
          3205 => x"8f",
          3206 => x"08",
          3207 => x"d5",
          3208 => x"ec",
          3209 => x"81",
          3210 => x"9f",
          3211 => x"2e",
          3212 => x"74",
          3213 => x"98",
          3214 => x"7e",
          3215 => x"3f",
          3216 => x"08",
          3217 => x"83",
          3218 => x"e0",
          3219 => x"89",
          3220 => x"77",
          3221 => x"d6",
          3222 => x"7f",
          3223 => x"58",
          3224 => x"75",
          3225 => x"75",
          3226 => x"77",
          3227 => x"7c",
          3228 => x"33",
          3229 => x"3f",
          3230 => x"08",
          3231 => x"7e",
          3232 => x"56",
          3233 => x"2e",
          3234 => x"16",
          3235 => x"55",
          3236 => x"94",
          3237 => x"53",
          3238 => x"b0",
          3239 => x"31",
          3240 => x"05",
          3241 => x"3f",
          3242 => x"56",
          3243 => x"9c",
          3244 => x"19",
          3245 => x"06",
          3246 => x"31",
          3247 => x"76",
          3248 => x"7b",
          3249 => x"08",
          3250 => x"d1",
          3251 => x"ec",
          3252 => x"81",
          3253 => x"94",
          3254 => x"ff",
          3255 => x"05",
          3256 => x"cf",
          3257 => x"76",
          3258 => x"17",
          3259 => x"1e",
          3260 => x"18",
          3261 => x"5e",
          3262 => x"39",
          3263 => x"81",
          3264 => x"90",
          3265 => x"f2",
          3266 => x"63",
          3267 => x"40",
          3268 => x"7e",
          3269 => x"fc",
          3270 => x"51",
          3271 => x"81",
          3272 => x"55",
          3273 => x"08",
          3274 => x"18",
          3275 => x"80",
          3276 => x"74",
          3277 => x"39",
          3278 => x"70",
          3279 => x"81",
          3280 => x"56",
          3281 => x"80",
          3282 => x"38",
          3283 => x"0b",
          3284 => x"82",
          3285 => x"39",
          3286 => x"19",
          3287 => x"83",
          3288 => x"18",
          3289 => x"56",
          3290 => x"27",
          3291 => x"09",
          3292 => x"2e",
          3293 => x"94",
          3294 => x"83",
          3295 => x"56",
          3296 => x"38",
          3297 => x"22",
          3298 => x"89",
          3299 => x"55",
          3300 => x"75",
          3301 => x"18",
          3302 => x"9c",
          3303 => x"85",
          3304 => x"08",
          3305 => x"d7",
          3306 => x"ec",
          3307 => x"81",
          3308 => x"80",
          3309 => x"38",
          3310 => x"ff",
          3311 => x"ff",
          3312 => x"38",
          3313 => x"0c",
          3314 => x"85",
          3315 => x"19",
          3316 => x"b0",
          3317 => x"19",
          3318 => x"81",
          3319 => x"74",
          3320 => x"3f",
          3321 => x"08",
          3322 => x"98",
          3323 => x"7e",
          3324 => x"3f",
          3325 => x"08",
          3326 => x"d2",
          3327 => x"e0",
          3328 => x"89",
          3329 => x"78",
          3330 => x"d5",
          3331 => x"7f",
          3332 => x"58",
          3333 => x"75",
          3334 => x"75",
          3335 => x"78",
          3336 => x"7c",
          3337 => x"33",
          3338 => x"3f",
          3339 => x"08",
          3340 => x"7e",
          3341 => x"78",
          3342 => x"74",
          3343 => x"38",
          3344 => x"b0",
          3345 => x"31",
          3346 => x"05",
          3347 => x"51",
          3348 => x"7e",
          3349 => x"83",
          3350 => x"89",
          3351 => x"db",
          3352 => x"08",
          3353 => x"26",
          3354 => x"51",
          3355 => x"81",
          3356 => x"fd",
          3357 => x"77",
          3358 => x"55",
          3359 => x"0c",
          3360 => x"83",
          3361 => x"80",
          3362 => x"55",
          3363 => x"83",
          3364 => x"9c",
          3365 => x"7e",
          3366 => x"3f",
          3367 => x"08",
          3368 => x"75",
          3369 => x"94",
          3370 => x"ff",
          3371 => x"05",
          3372 => x"3f",
          3373 => x"0b",
          3374 => x"7b",
          3375 => x"08",
          3376 => x"76",
          3377 => x"08",
          3378 => x"1c",
          3379 => x"08",
          3380 => x"5c",
          3381 => x"83",
          3382 => x"74",
          3383 => x"fd",
          3384 => x"18",
          3385 => x"07",
          3386 => x"19",
          3387 => x"75",
          3388 => x"0c",
          3389 => x"04",
          3390 => x"7a",
          3391 => x"05",
          3392 => x"56",
          3393 => x"81",
          3394 => x"57",
          3395 => x"08",
          3396 => x"90",
          3397 => x"86",
          3398 => x"06",
          3399 => x"73",
          3400 => x"e9",
          3401 => x"08",
          3402 => x"cc",
          3403 => x"ec",
          3404 => x"81",
          3405 => x"80",
          3406 => x"16",
          3407 => x"33",
          3408 => x"55",
          3409 => x"34",
          3410 => x"53",
          3411 => x"08",
          3412 => x"3f",
          3413 => x"52",
          3414 => x"c9",
          3415 => x"88",
          3416 => x"96",
          3417 => x"f0",
          3418 => x"92",
          3419 => x"ca",
          3420 => x"81",
          3421 => x"34",
          3422 => x"df",
          3423 => x"e0",
          3424 => x"33",
          3425 => x"55",
          3426 => x"17",
          3427 => x"ec",
          3428 => x"3d",
          3429 => x"3d",
          3430 => x"52",
          3431 => x"3f",
          3432 => x"08",
          3433 => x"e0",
          3434 => x"86",
          3435 => x"52",
          3436 => x"bc",
          3437 => x"e0",
          3438 => x"ec",
          3439 => x"38",
          3440 => x"08",
          3441 => x"81",
          3442 => x"86",
          3443 => x"ff",
          3444 => x"3d",
          3445 => x"3f",
          3446 => x"0b",
          3447 => x"08",
          3448 => x"81",
          3449 => x"81",
          3450 => x"80",
          3451 => x"ec",
          3452 => x"3d",
          3453 => x"3d",
          3454 => x"93",
          3455 => x"52",
          3456 => x"e9",
          3457 => x"ec",
          3458 => x"81",
          3459 => x"80",
          3460 => x"58",
          3461 => x"3d",
          3462 => x"e0",
          3463 => x"ec",
          3464 => x"81",
          3465 => x"bc",
          3466 => x"c7",
          3467 => x"98",
          3468 => x"73",
          3469 => x"38",
          3470 => x"12",
          3471 => x"39",
          3472 => x"33",
          3473 => x"70",
          3474 => x"55",
          3475 => x"2e",
          3476 => x"7f",
          3477 => x"54",
          3478 => x"81",
          3479 => x"94",
          3480 => x"39",
          3481 => x"08",
          3482 => x"81",
          3483 => x"85",
          3484 => x"ec",
          3485 => x"3d",
          3486 => x"3d",
          3487 => x"5b",
          3488 => x"34",
          3489 => x"3d",
          3490 => x"52",
          3491 => x"e8",
          3492 => x"ec",
          3493 => x"81",
          3494 => x"82",
          3495 => x"43",
          3496 => x"11",
          3497 => x"58",
          3498 => x"80",
          3499 => x"38",
          3500 => x"3d",
          3501 => x"d5",
          3502 => x"ec",
          3503 => x"81",
          3504 => x"82",
          3505 => x"52",
          3506 => x"c8",
          3507 => x"e0",
          3508 => x"ec",
          3509 => x"c1",
          3510 => x"7b",
          3511 => x"3f",
          3512 => x"08",
          3513 => x"74",
          3514 => x"3f",
          3515 => x"08",
          3516 => x"e0",
          3517 => x"38",
          3518 => x"51",
          3519 => x"81",
          3520 => x"57",
          3521 => x"08",
          3522 => x"52",
          3523 => x"f2",
          3524 => x"ec",
          3525 => x"a6",
          3526 => x"74",
          3527 => x"3f",
          3528 => x"08",
          3529 => x"e0",
          3530 => x"cc",
          3531 => x"2e",
          3532 => x"86",
          3533 => x"81",
          3534 => x"81",
          3535 => x"3d",
          3536 => x"52",
          3537 => x"c9",
          3538 => x"3d",
          3539 => x"11",
          3540 => x"5a",
          3541 => x"2e",
          3542 => x"b9",
          3543 => x"16",
          3544 => x"33",
          3545 => x"73",
          3546 => x"16",
          3547 => x"26",
          3548 => x"75",
          3549 => x"38",
          3550 => x"05",
          3551 => x"6f",
          3552 => x"ff",
          3553 => x"55",
          3554 => x"74",
          3555 => x"38",
          3556 => x"11",
          3557 => x"74",
          3558 => x"39",
          3559 => x"09",
          3560 => x"38",
          3561 => x"11",
          3562 => x"74",
          3563 => x"81",
          3564 => x"70",
          3565 => x"dc",
          3566 => x"08",
          3567 => x"5c",
          3568 => x"73",
          3569 => x"38",
          3570 => x"1a",
          3571 => x"55",
          3572 => x"38",
          3573 => x"73",
          3574 => x"38",
          3575 => x"76",
          3576 => x"74",
          3577 => x"33",
          3578 => x"05",
          3579 => x"15",
          3580 => x"ba",
          3581 => x"05",
          3582 => x"ff",
          3583 => x"06",
          3584 => x"57",
          3585 => x"18",
          3586 => x"54",
          3587 => x"70",
          3588 => x"34",
          3589 => x"ee",
          3590 => x"34",
          3591 => x"e0",
          3592 => x"0d",
          3593 => x"0d",
          3594 => x"3d",
          3595 => x"71",
          3596 => x"ec",
          3597 => x"ec",
          3598 => x"81",
          3599 => x"82",
          3600 => x"15",
          3601 => x"82",
          3602 => x"15",
          3603 => x"76",
          3604 => x"90",
          3605 => x"81",
          3606 => x"06",
          3607 => x"72",
          3608 => x"56",
          3609 => x"54",
          3610 => x"17",
          3611 => x"78",
          3612 => x"38",
          3613 => x"22",
          3614 => x"59",
          3615 => x"78",
          3616 => x"76",
          3617 => x"51",
          3618 => x"3f",
          3619 => x"08",
          3620 => x"54",
          3621 => x"53",
          3622 => x"3f",
          3623 => x"08",
          3624 => x"38",
          3625 => x"75",
          3626 => x"18",
          3627 => x"31",
          3628 => x"57",
          3629 => x"b1",
          3630 => x"08",
          3631 => x"38",
          3632 => x"51",
          3633 => x"81",
          3634 => x"54",
          3635 => x"08",
          3636 => x"9a",
          3637 => x"e0",
          3638 => x"81",
          3639 => x"ec",
          3640 => x"16",
          3641 => x"16",
          3642 => x"2e",
          3643 => x"76",
          3644 => x"dc",
          3645 => x"31",
          3646 => x"18",
          3647 => x"90",
          3648 => x"81",
          3649 => x"06",
          3650 => x"56",
          3651 => x"9a",
          3652 => x"74",
          3653 => x"3f",
          3654 => x"08",
          3655 => x"e0",
          3656 => x"81",
          3657 => x"56",
          3658 => x"52",
          3659 => x"84",
          3660 => x"e0",
          3661 => x"ff",
          3662 => x"81",
          3663 => x"38",
          3664 => x"98",
          3665 => x"a6",
          3666 => x"16",
          3667 => x"39",
          3668 => x"16",
          3669 => x"75",
          3670 => x"53",
          3671 => x"aa",
          3672 => x"79",
          3673 => x"3f",
          3674 => x"08",
          3675 => x"0b",
          3676 => x"82",
          3677 => x"39",
          3678 => x"16",
          3679 => x"bb",
          3680 => x"2a",
          3681 => x"08",
          3682 => x"15",
          3683 => x"15",
          3684 => x"90",
          3685 => x"16",
          3686 => x"33",
          3687 => x"53",
          3688 => x"34",
          3689 => x"06",
          3690 => x"2e",
          3691 => x"9c",
          3692 => x"85",
          3693 => x"16",
          3694 => x"72",
          3695 => x"0c",
          3696 => x"04",
          3697 => x"79",
          3698 => x"75",
          3699 => x"8a",
          3700 => x"89",
          3701 => x"52",
          3702 => x"05",
          3703 => x"3f",
          3704 => x"08",
          3705 => x"e0",
          3706 => x"38",
          3707 => x"7a",
          3708 => x"d8",
          3709 => x"ec",
          3710 => x"81",
          3711 => x"80",
          3712 => x"16",
          3713 => x"2b",
          3714 => x"74",
          3715 => x"86",
          3716 => x"84",
          3717 => x"06",
          3718 => x"73",
          3719 => x"38",
          3720 => x"52",
          3721 => x"da",
          3722 => x"e0",
          3723 => x"0c",
          3724 => x"14",
          3725 => x"23",
          3726 => x"51",
          3727 => x"81",
          3728 => x"55",
          3729 => x"09",
          3730 => x"38",
          3731 => x"39",
          3732 => x"84",
          3733 => x"0c",
          3734 => x"81",
          3735 => x"89",
          3736 => x"fc",
          3737 => x"87",
          3738 => x"53",
          3739 => x"e7",
          3740 => x"ec",
          3741 => x"38",
          3742 => x"08",
          3743 => x"3d",
          3744 => x"3d",
          3745 => x"89",
          3746 => x"54",
          3747 => x"54",
          3748 => x"81",
          3749 => x"53",
          3750 => x"08",
          3751 => x"74",
          3752 => x"ec",
          3753 => x"73",
          3754 => x"3f",
          3755 => x"08",
          3756 => x"39",
          3757 => x"08",
          3758 => x"d3",
          3759 => x"ec",
          3760 => x"81",
          3761 => x"84",
          3762 => x"06",
          3763 => x"53",
          3764 => x"ec",
          3765 => x"38",
          3766 => x"51",
          3767 => x"72",
          3768 => x"cf",
          3769 => x"ec",
          3770 => x"32",
          3771 => x"72",
          3772 => x"70",
          3773 => x"08",
          3774 => x"54",
          3775 => x"ec",
          3776 => x"3d",
          3777 => x"3d",
          3778 => x"80",
          3779 => x"70",
          3780 => x"52",
          3781 => x"3f",
          3782 => x"08",
          3783 => x"e0",
          3784 => x"64",
          3785 => x"d6",
          3786 => x"ec",
          3787 => x"81",
          3788 => x"a0",
          3789 => x"cb",
          3790 => x"98",
          3791 => x"73",
          3792 => x"38",
          3793 => x"39",
          3794 => x"88",
          3795 => x"75",
          3796 => x"3f",
          3797 => x"e0",
          3798 => x"0d",
          3799 => x"0d",
          3800 => x"5c",
          3801 => x"3d",
          3802 => x"93",
          3803 => x"d6",
          3804 => x"e0",
          3805 => x"ec",
          3806 => x"80",
          3807 => x"0c",
          3808 => x"11",
          3809 => x"90",
          3810 => x"56",
          3811 => x"74",
          3812 => x"75",
          3813 => x"e4",
          3814 => x"81",
          3815 => x"5b",
          3816 => x"81",
          3817 => x"75",
          3818 => x"73",
          3819 => x"81",
          3820 => x"82",
          3821 => x"76",
          3822 => x"f0",
          3823 => x"f4",
          3824 => x"e0",
          3825 => x"d1",
          3826 => x"e0",
          3827 => x"ce",
          3828 => x"e0",
          3829 => x"81",
          3830 => x"07",
          3831 => x"05",
          3832 => x"53",
          3833 => x"98",
          3834 => x"26",
          3835 => x"f9",
          3836 => x"08",
          3837 => x"08",
          3838 => x"98",
          3839 => x"81",
          3840 => x"58",
          3841 => x"3f",
          3842 => x"08",
          3843 => x"e0",
          3844 => x"38",
          3845 => x"77",
          3846 => x"5d",
          3847 => x"74",
          3848 => x"81",
          3849 => x"b4",
          3850 => x"bb",
          3851 => x"ec",
          3852 => x"ff",
          3853 => x"30",
          3854 => x"1b",
          3855 => x"5b",
          3856 => x"39",
          3857 => x"ff",
          3858 => x"81",
          3859 => x"f0",
          3860 => x"30",
          3861 => x"1b",
          3862 => x"5b",
          3863 => x"83",
          3864 => x"58",
          3865 => x"92",
          3866 => x"0c",
          3867 => x"12",
          3868 => x"33",
          3869 => x"54",
          3870 => x"34",
          3871 => x"e0",
          3872 => x"0d",
          3873 => x"0d",
          3874 => x"fc",
          3875 => x"52",
          3876 => x"3f",
          3877 => x"08",
          3878 => x"e0",
          3879 => x"38",
          3880 => x"56",
          3881 => x"38",
          3882 => x"70",
          3883 => x"81",
          3884 => x"55",
          3885 => x"80",
          3886 => x"38",
          3887 => x"54",
          3888 => x"08",
          3889 => x"38",
          3890 => x"81",
          3891 => x"53",
          3892 => x"52",
          3893 => x"8c",
          3894 => x"e0",
          3895 => x"19",
          3896 => x"c9",
          3897 => x"08",
          3898 => x"ff",
          3899 => x"81",
          3900 => x"ff",
          3901 => x"06",
          3902 => x"56",
          3903 => x"08",
          3904 => x"81",
          3905 => x"82",
          3906 => x"75",
          3907 => x"54",
          3908 => x"08",
          3909 => x"27",
          3910 => x"17",
          3911 => x"ec",
          3912 => x"76",
          3913 => x"3f",
          3914 => x"08",
          3915 => x"08",
          3916 => x"90",
          3917 => x"c0",
          3918 => x"90",
          3919 => x"80",
          3920 => x"75",
          3921 => x"75",
          3922 => x"ec",
          3923 => x"3d",
          3924 => x"3d",
          3925 => x"a0",
          3926 => x"05",
          3927 => x"51",
          3928 => x"81",
          3929 => x"55",
          3930 => x"08",
          3931 => x"78",
          3932 => x"08",
          3933 => x"70",
          3934 => x"ae",
          3935 => x"e0",
          3936 => x"ec",
          3937 => x"db",
          3938 => x"fb",
          3939 => x"85",
          3940 => x"06",
          3941 => x"86",
          3942 => x"c7",
          3943 => x"2b",
          3944 => x"24",
          3945 => x"02",
          3946 => x"33",
          3947 => x"58",
          3948 => x"76",
          3949 => x"6b",
          3950 => x"cc",
          3951 => x"ec",
          3952 => x"84",
          3953 => x"06",
          3954 => x"73",
          3955 => x"d4",
          3956 => x"81",
          3957 => x"94",
          3958 => x"81",
          3959 => x"5a",
          3960 => x"08",
          3961 => x"8a",
          3962 => x"54",
          3963 => x"81",
          3964 => x"55",
          3965 => x"08",
          3966 => x"81",
          3967 => x"52",
          3968 => x"e5",
          3969 => x"e0",
          3970 => x"ec",
          3971 => x"38",
          3972 => x"cf",
          3973 => x"e0",
          3974 => x"88",
          3975 => x"e0",
          3976 => x"38",
          3977 => x"c2",
          3978 => x"e0",
          3979 => x"e0",
          3980 => x"81",
          3981 => x"07",
          3982 => x"55",
          3983 => x"2e",
          3984 => x"80",
          3985 => x"80",
          3986 => x"77",
          3987 => x"3f",
          3988 => x"08",
          3989 => x"38",
          3990 => x"ba",
          3991 => x"ec",
          3992 => x"74",
          3993 => x"0c",
          3994 => x"04",
          3995 => x"82",
          3996 => x"c0",
          3997 => x"3d",
          3998 => x"3f",
          3999 => x"08",
          4000 => x"e0",
          4001 => x"38",
          4002 => x"52",
          4003 => x"52",
          4004 => x"3f",
          4005 => x"08",
          4006 => x"e0",
          4007 => x"88",
          4008 => x"39",
          4009 => x"08",
          4010 => x"81",
          4011 => x"38",
          4012 => x"05",
          4013 => x"2a",
          4014 => x"55",
          4015 => x"81",
          4016 => x"5a",
          4017 => x"3d",
          4018 => x"c1",
          4019 => x"ec",
          4020 => x"55",
          4021 => x"e0",
          4022 => x"87",
          4023 => x"e0",
          4024 => x"09",
          4025 => x"38",
          4026 => x"ec",
          4027 => x"2e",
          4028 => x"86",
          4029 => x"81",
          4030 => x"81",
          4031 => x"ec",
          4032 => x"78",
          4033 => x"3f",
          4034 => x"08",
          4035 => x"e0",
          4036 => x"38",
          4037 => x"52",
          4038 => x"ff",
          4039 => x"78",
          4040 => x"b4",
          4041 => x"54",
          4042 => x"15",
          4043 => x"b2",
          4044 => x"ca",
          4045 => x"b6",
          4046 => x"53",
          4047 => x"53",
          4048 => x"3f",
          4049 => x"b4",
          4050 => x"d4",
          4051 => x"b6",
          4052 => x"54",
          4053 => x"d5",
          4054 => x"53",
          4055 => x"11",
          4056 => x"d7",
          4057 => x"81",
          4058 => x"34",
          4059 => x"a4",
          4060 => x"e0",
          4061 => x"ec",
          4062 => x"38",
          4063 => x"0a",
          4064 => x"05",
          4065 => x"d0",
          4066 => x"64",
          4067 => x"c9",
          4068 => x"54",
          4069 => x"15",
          4070 => x"81",
          4071 => x"34",
          4072 => x"b8",
          4073 => x"ec",
          4074 => x"8b",
          4075 => x"75",
          4076 => x"ff",
          4077 => x"73",
          4078 => x"0c",
          4079 => x"04",
          4080 => x"a9",
          4081 => x"51",
          4082 => x"82",
          4083 => x"ff",
          4084 => x"a9",
          4085 => x"ee",
          4086 => x"e0",
          4087 => x"ec",
          4088 => x"d3",
          4089 => x"a9",
          4090 => x"9d",
          4091 => x"58",
          4092 => x"81",
          4093 => x"55",
          4094 => x"08",
          4095 => x"02",
          4096 => x"33",
          4097 => x"54",
          4098 => x"82",
          4099 => x"53",
          4100 => x"52",
          4101 => x"88",
          4102 => x"b4",
          4103 => x"53",
          4104 => x"3d",
          4105 => x"ff",
          4106 => x"aa",
          4107 => x"73",
          4108 => x"3f",
          4109 => x"08",
          4110 => x"e0",
          4111 => x"63",
          4112 => x"81",
          4113 => x"65",
          4114 => x"2e",
          4115 => x"55",
          4116 => x"81",
          4117 => x"84",
          4118 => x"06",
          4119 => x"73",
          4120 => x"3f",
          4121 => x"08",
          4122 => x"e0",
          4123 => x"38",
          4124 => x"53",
          4125 => x"95",
          4126 => x"16",
          4127 => x"87",
          4128 => x"05",
          4129 => x"34",
          4130 => x"70",
          4131 => x"81",
          4132 => x"55",
          4133 => x"74",
          4134 => x"73",
          4135 => x"78",
          4136 => x"83",
          4137 => x"16",
          4138 => x"2a",
          4139 => x"51",
          4140 => x"80",
          4141 => x"38",
          4142 => x"80",
          4143 => x"52",
          4144 => x"be",
          4145 => x"e0",
          4146 => x"51",
          4147 => x"3f",
          4148 => x"ec",
          4149 => x"2e",
          4150 => x"81",
          4151 => x"52",
          4152 => x"b5",
          4153 => x"ec",
          4154 => x"80",
          4155 => x"58",
          4156 => x"e0",
          4157 => x"38",
          4158 => x"54",
          4159 => x"09",
          4160 => x"38",
          4161 => x"52",
          4162 => x"af",
          4163 => x"81",
          4164 => x"34",
          4165 => x"ec",
          4166 => x"38",
          4167 => x"ca",
          4168 => x"e0",
          4169 => x"ec",
          4170 => x"38",
          4171 => x"b5",
          4172 => x"ec",
          4173 => x"74",
          4174 => x"0c",
          4175 => x"04",
          4176 => x"02",
          4177 => x"33",
          4178 => x"80",
          4179 => x"57",
          4180 => x"95",
          4181 => x"52",
          4182 => x"d2",
          4183 => x"ec",
          4184 => x"81",
          4185 => x"80",
          4186 => x"5a",
          4187 => x"3d",
          4188 => x"c9",
          4189 => x"ec",
          4190 => x"81",
          4191 => x"b8",
          4192 => x"cf",
          4193 => x"a0",
          4194 => x"55",
          4195 => x"75",
          4196 => x"71",
          4197 => x"33",
          4198 => x"74",
          4199 => x"57",
          4200 => x"8b",
          4201 => x"54",
          4202 => x"15",
          4203 => x"ff",
          4204 => x"81",
          4205 => x"55",
          4206 => x"e0",
          4207 => x"0d",
          4208 => x"0d",
          4209 => x"53",
          4210 => x"05",
          4211 => x"51",
          4212 => x"81",
          4213 => x"55",
          4214 => x"08",
          4215 => x"76",
          4216 => x"93",
          4217 => x"51",
          4218 => x"81",
          4219 => x"55",
          4220 => x"08",
          4221 => x"80",
          4222 => x"81",
          4223 => x"86",
          4224 => x"38",
          4225 => x"86",
          4226 => x"90",
          4227 => x"54",
          4228 => x"ff",
          4229 => x"76",
          4230 => x"83",
          4231 => x"51",
          4232 => x"3f",
          4233 => x"08",
          4234 => x"ec",
          4235 => x"3d",
          4236 => x"3d",
          4237 => x"5c",
          4238 => x"98",
          4239 => x"52",
          4240 => x"d1",
          4241 => x"ec",
          4242 => x"ec",
          4243 => x"70",
          4244 => x"08",
          4245 => x"51",
          4246 => x"80",
          4247 => x"38",
          4248 => x"06",
          4249 => x"80",
          4250 => x"38",
          4251 => x"5f",
          4252 => x"3d",
          4253 => x"ff",
          4254 => x"81",
          4255 => x"57",
          4256 => x"08",
          4257 => x"74",
          4258 => x"c3",
          4259 => x"ec",
          4260 => x"81",
          4261 => x"bf",
          4262 => x"e0",
          4263 => x"e0",
          4264 => x"59",
          4265 => x"81",
          4266 => x"56",
          4267 => x"33",
          4268 => x"16",
          4269 => x"27",
          4270 => x"56",
          4271 => x"80",
          4272 => x"80",
          4273 => x"ff",
          4274 => x"70",
          4275 => x"56",
          4276 => x"e8",
          4277 => x"76",
          4278 => x"81",
          4279 => x"80",
          4280 => x"57",
          4281 => x"78",
          4282 => x"51",
          4283 => x"2e",
          4284 => x"73",
          4285 => x"38",
          4286 => x"08",
          4287 => x"b1",
          4288 => x"ec",
          4289 => x"81",
          4290 => x"a7",
          4291 => x"33",
          4292 => x"c3",
          4293 => x"2e",
          4294 => x"e4",
          4295 => x"2e",
          4296 => x"56",
          4297 => x"05",
          4298 => x"e3",
          4299 => x"e0",
          4300 => x"76",
          4301 => x"0c",
          4302 => x"04",
          4303 => x"82",
          4304 => x"ff",
          4305 => x"9d",
          4306 => x"fa",
          4307 => x"e0",
          4308 => x"e0",
          4309 => x"81",
          4310 => x"83",
          4311 => x"53",
          4312 => x"3d",
          4313 => x"ff",
          4314 => x"73",
          4315 => x"70",
          4316 => x"52",
          4317 => x"9f",
          4318 => x"bc",
          4319 => x"74",
          4320 => x"6d",
          4321 => x"70",
          4322 => x"af",
          4323 => x"ec",
          4324 => x"2e",
          4325 => x"70",
          4326 => x"57",
          4327 => x"fd",
          4328 => x"e0",
          4329 => x"8d",
          4330 => x"2b",
          4331 => x"81",
          4332 => x"86",
          4333 => x"e0",
          4334 => x"9f",
          4335 => x"ff",
          4336 => x"54",
          4337 => x"8a",
          4338 => x"70",
          4339 => x"06",
          4340 => x"ff",
          4341 => x"38",
          4342 => x"15",
          4343 => x"80",
          4344 => x"74",
          4345 => x"b0",
          4346 => x"89",
          4347 => x"e0",
          4348 => x"81",
          4349 => x"88",
          4350 => x"26",
          4351 => x"39",
          4352 => x"86",
          4353 => x"81",
          4354 => x"ff",
          4355 => x"38",
          4356 => x"54",
          4357 => x"81",
          4358 => x"81",
          4359 => x"78",
          4360 => x"5a",
          4361 => x"6d",
          4362 => x"81",
          4363 => x"57",
          4364 => x"9f",
          4365 => x"38",
          4366 => x"54",
          4367 => x"81",
          4368 => x"b1",
          4369 => x"2e",
          4370 => x"a7",
          4371 => x"15",
          4372 => x"54",
          4373 => x"09",
          4374 => x"38",
          4375 => x"76",
          4376 => x"41",
          4377 => x"52",
          4378 => x"52",
          4379 => x"b3",
          4380 => x"e0",
          4381 => x"ec",
          4382 => x"f7",
          4383 => x"74",
          4384 => x"e5",
          4385 => x"e0",
          4386 => x"ec",
          4387 => x"38",
          4388 => x"38",
          4389 => x"74",
          4390 => x"39",
          4391 => x"08",
          4392 => x"81",
          4393 => x"38",
          4394 => x"74",
          4395 => x"38",
          4396 => x"51",
          4397 => x"3f",
          4398 => x"08",
          4399 => x"e0",
          4400 => x"a0",
          4401 => x"e0",
          4402 => x"51",
          4403 => x"3f",
          4404 => x"0b",
          4405 => x"8b",
          4406 => x"67",
          4407 => x"a7",
          4408 => x"81",
          4409 => x"34",
          4410 => x"ad",
          4411 => x"ec",
          4412 => x"73",
          4413 => x"ec",
          4414 => x"3d",
          4415 => x"3d",
          4416 => x"02",
          4417 => x"cb",
          4418 => x"3d",
          4419 => x"72",
          4420 => x"5a",
          4421 => x"81",
          4422 => x"58",
          4423 => x"08",
          4424 => x"91",
          4425 => x"77",
          4426 => x"7c",
          4427 => x"38",
          4428 => x"59",
          4429 => x"90",
          4430 => x"81",
          4431 => x"06",
          4432 => x"73",
          4433 => x"54",
          4434 => x"82",
          4435 => x"39",
          4436 => x"8b",
          4437 => x"11",
          4438 => x"2b",
          4439 => x"54",
          4440 => x"fe",
          4441 => x"ff",
          4442 => x"70",
          4443 => x"07",
          4444 => x"ec",
          4445 => x"8c",
          4446 => x"40",
          4447 => x"55",
          4448 => x"88",
          4449 => x"08",
          4450 => x"38",
          4451 => x"77",
          4452 => x"56",
          4453 => x"51",
          4454 => x"3f",
          4455 => x"55",
          4456 => x"08",
          4457 => x"38",
          4458 => x"ec",
          4459 => x"2e",
          4460 => x"81",
          4461 => x"ff",
          4462 => x"38",
          4463 => x"08",
          4464 => x"16",
          4465 => x"2e",
          4466 => x"87",
          4467 => x"74",
          4468 => x"74",
          4469 => x"81",
          4470 => x"38",
          4471 => x"ff",
          4472 => x"2e",
          4473 => x"7b",
          4474 => x"80",
          4475 => x"81",
          4476 => x"81",
          4477 => x"06",
          4478 => x"56",
          4479 => x"52",
          4480 => x"af",
          4481 => x"ec",
          4482 => x"81",
          4483 => x"80",
          4484 => x"81",
          4485 => x"56",
          4486 => x"d3",
          4487 => x"ff",
          4488 => x"7c",
          4489 => x"55",
          4490 => x"b3",
          4491 => x"1b",
          4492 => x"1b",
          4493 => x"33",
          4494 => x"54",
          4495 => x"34",
          4496 => x"fe",
          4497 => x"08",
          4498 => x"74",
          4499 => x"75",
          4500 => x"16",
          4501 => x"33",
          4502 => x"73",
          4503 => x"77",
          4504 => x"ec",
          4505 => x"3d",
          4506 => x"3d",
          4507 => x"02",
          4508 => x"eb",
          4509 => x"3d",
          4510 => x"59",
          4511 => x"8b",
          4512 => x"81",
          4513 => x"24",
          4514 => x"81",
          4515 => x"84",
          4516 => x"fc",
          4517 => x"51",
          4518 => x"2e",
          4519 => x"75",
          4520 => x"e0",
          4521 => x"06",
          4522 => x"7e",
          4523 => x"d0",
          4524 => x"e0",
          4525 => x"06",
          4526 => x"56",
          4527 => x"74",
          4528 => x"76",
          4529 => x"81",
          4530 => x"8a",
          4531 => x"b2",
          4532 => x"fc",
          4533 => x"52",
          4534 => x"a4",
          4535 => x"ec",
          4536 => x"38",
          4537 => x"80",
          4538 => x"74",
          4539 => x"26",
          4540 => x"15",
          4541 => x"74",
          4542 => x"38",
          4543 => x"80",
          4544 => x"84",
          4545 => x"92",
          4546 => x"80",
          4547 => x"38",
          4548 => x"06",
          4549 => x"2e",
          4550 => x"56",
          4551 => x"78",
          4552 => x"89",
          4553 => x"2b",
          4554 => x"43",
          4555 => x"38",
          4556 => x"30",
          4557 => x"77",
          4558 => x"91",
          4559 => x"c2",
          4560 => x"f8",
          4561 => x"52",
          4562 => x"a4",
          4563 => x"56",
          4564 => x"08",
          4565 => x"77",
          4566 => x"77",
          4567 => x"e0",
          4568 => x"45",
          4569 => x"bf",
          4570 => x"8e",
          4571 => x"26",
          4572 => x"74",
          4573 => x"48",
          4574 => x"75",
          4575 => x"38",
          4576 => x"81",
          4577 => x"fa",
          4578 => x"2a",
          4579 => x"56",
          4580 => x"2e",
          4581 => x"87",
          4582 => x"82",
          4583 => x"38",
          4584 => x"55",
          4585 => x"83",
          4586 => x"81",
          4587 => x"56",
          4588 => x"80",
          4589 => x"38",
          4590 => x"83",
          4591 => x"06",
          4592 => x"78",
          4593 => x"91",
          4594 => x"0b",
          4595 => x"22",
          4596 => x"80",
          4597 => x"74",
          4598 => x"38",
          4599 => x"56",
          4600 => x"17",
          4601 => x"57",
          4602 => x"2e",
          4603 => x"75",
          4604 => x"79",
          4605 => x"fe",
          4606 => x"81",
          4607 => x"84",
          4608 => x"05",
          4609 => x"5e",
          4610 => x"80",
          4611 => x"e0",
          4612 => x"8a",
          4613 => x"fd",
          4614 => x"75",
          4615 => x"38",
          4616 => x"78",
          4617 => x"8c",
          4618 => x"0b",
          4619 => x"22",
          4620 => x"80",
          4621 => x"74",
          4622 => x"38",
          4623 => x"56",
          4624 => x"17",
          4625 => x"57",
          4626 => x"2e",
          4627 => x"75",
          4628 => x"79",
          4629 => x"fe",
          4630 => x"81",
          4631 => x"10",
          4632 => x"81",
          4633 => x"9f",
          4634 => x"38",
          4635 => x"ec",
          4636 => x"81",
          4637 => x"05",
          4638 => x"2a",
          4639 => x"56",
          4640 => x"17",
          4641 => x"81",
          4642 => x"60",
          4643 => x"65",
          4644 => x"12",
          4645 => x"30",
          4646 => x"74",
          4647 => x"59",
          4648 => x"7d",
          4649 => x"81",
          4650 => x"76",
          4651 => x"41",
          4652 => x"76",
          4653 => x"90",
          4654 => x"62",
          4655 => x"51",
          4656 => x"26",
          4657 => x"75",
          4658 => x"31",
          4659 => x"65",
          4660 => x"fe",
          4661 => x"81",
          4662 => x"58",
          4663 => x"09",
          4664 => x"38",
          4665 => x"08",
          4666 => x"26",
          4667 => x"78",
          4668 => x"79",
          4669 => x"78",
          4670 => x"86",
          4671 => x"82",
          4672 => x"06",
          4673 => x"83",
          4674 => x"81",
          4675 => x"27",
          4676 => x"8f",
          4677 => x"55",
          4678 => x"26",
          4679 => x"59",
          4680 => x"62",
          4681 => x"74",
          4682 => x"38",
          4683 => x"88",
          4684 => x"e0",
          4685 => x"26",
          4686 => x"86",
          4687 => x"1a",
          4688 => x"79",
          4689 => x"38",
          4690 => x"80",
          4691 => x"2e",
          4692 => x"83",
          4693 => x"9f",
          4694 => x"8b",
          4695 => x"06",
          4696 => x"74",
          4697 => x"84",
          4698 => x"52",
          4699 => x"a2",
          4700 => x"53",
          4701 => x"52",
          4702 => x"a2",
          4703 => x"80",
          4704 => x"51",
          4705 => x"3f",
          4706 => x"34",
          4707 => x"ff",
          4708 => x"1b",
          4709 => x"a2",
          4710 => x"90",
          4711 => x"83",
          4712 => x"70",
          4713 => x"80",
          4714 => x"55",
          4715 => x"ff",
          4716 => x"66",
          4717 => x"ff",
          4718 => x"38",
          4719 => x"ff",
          4720 => x"1b",
          4721 => x"f2",
          4722 => x"74",
          4723 => x"51",
          4724 => x"3f",
          4725 => x"1c",
          4726 => x"98",
          4727 => x"a0",
          4728 => x"ff",
          4729 => x"51",
          4730 => x"3f",
          4731 => x"1b",
          4732 => x"e4",
          4733 => x"2e",
          4734 => x"80",
          4735 => x"88",
          4736 => x"80",
          4737 => x"ff",
          4738 => x"7c",
          4739 => x"51",
          4740 => x"3f",
          4741 => x"1b",
          4742 => x"bc",
          4743 => x"b0",
          4744 => x"a0",
          4745 => x"52",
          4746 => x"ff",
          4747 => x"ff",
          4748 => x"c0",
          4749 => x"0b",
          4750 => x"34",
          4751 => x"db",
          4752 => x"c7",
          4753 => x"39",
          4754 => x"0a",
          4755 => x"51",
          4756 => x"3f",
          4757 => x"ff",
          4758 => x"1b",
          4759 => x"da",
          4760 => x"0b",
          4761 => x"a9",
          4762 => x"34",
          4763 => x"dc",
          4764 => x"1b",
          4765 => x"8f",
          4766 => x"d5",
          4767 => x"1b",
          4768 => x"ff",
          4769 => x"81",
          4770 => x"7a",
          4771 => x"ff",
          4772 => x"81",
          4773 => x"e0",
          4774 => x"38",
          4775 => x"09",
          4776 => x"ee",
          4777 => x"60",
          4778 => x"7a",
          4779 => x"ff",
          4780 => x"84",
          4781 => x"52",
          4782 => x"9f",
          4783 => x"8b",
          4784 => x"52",
          4785 => x"9f",
          4786 => x"8a",
          4787 => x"52",
          4788 => x"51",
          4789 => x"3f",
          4790 => x"83",
          4791 => x"ff",
          4792 => x"82",
          4793 => x"1b",
          4794 => x"ec",
          4795 => x"d5",
          4796 => x"ff",
          4797 => x"75",
          4798 => x"05",
          4799 => x"7e",
          4800 => x"e5",
          4801 => x"60",
          4802 => x"52",
          4803 => x"9a",
          4804 => x"53",
          4805 => x"51",
          4806 => x"3f",
          4807 => x"58",
          4808 => x"09",
          4809 => x"38",
          4810 => x"51",
          4811 => x"3f",
          4812 => x"1b",
          4813 => x"a0",
          4814 => x"52",
          4815 => x"91",
          4816 => x"ff",
          4817 => x"81",
          4818 => x"f8",
          4819 => x"7a",
          4820 => x"84",
          4821 => x"61",
          4822 => x"26",
          4823 => x"57",
          4824 => x"53",
          4825 => x"51",
          4826 => x"3f",
          4827 => x"08",
          4828 => x"84",
          4829 => x"ec",
          4830 => x"7a",
          4831 => x"aa",
          4832 => x"75",
          4833 => x"56",
          4834 => x"81",
          4835 => x"80",
          4836 => x"38",
          4837 => x"83",
          4838 => x"63",
          4839 => x"74",
          4840 => x"38",
          4841 => x"54",
          4842 => x"52",
          4843 => x"99",
          4844 => x"ec",
          4845 => x"c1",
          4846 => x"75",
          4847 => x"56",
          4848 => x"8c",
          4849 => x"2e",
          4850 => x"56",
          4851 => x"ff",
          4852 => x"84",
          4853 => x"2e",
          4854 => x"56",
          4855 => x"58",
          4856 => x"38",
          4857 => x"77",
          4858 => x"ff",
          4859 => x"82",
          4860 => x"78",
          4861 => x"c2",
          4862 => x"1b",
          4863 => x"34",
          4864 => x"16",
          4865 => x"82",
          4866 => x"83",
          4867 => x"84",
          4868 => x"67",
          4869 => x"fd",
          4870 => x"51",
          4871 => x"3f",
          4872 => x"16",
          4873 => x"e0",
          4874 => x"bf",
          4875 => x"86",
          4876 => x"ec",
          4877 => x"16",
          4878 => x"83",
          4879 => x"ff",
          4880 => x"66",
          4881 => x"1b",
          4882 => x"8c",
          4883 => x"77",
          4884 => x"7e",
          4885 => x"91",
          4886 => x"81",
          4887 => x"a2",
          4888 => x"80",
          4889 => x"ff",
          4890 => x"81",
          4891 => x"e0",
          4892 => x"89",
          4893 => x"8a",
          4894 => x"86",
          4895 => x"e0",
          4896 => x"81",
          4897 => x"99",
          4898 => x"f5",
          4899 => x"60",
          4900 => x"79",
          4901 => x"5a",
          4902 => x"78",
          4903 => x"8d",
          4904 => x"55",
          4905 => x"fc",
          4906 => x"51",
          4907 => x"7a",
          4908 => x"81",
          4909 => x"8c",
          4910 => x"74",
          4911 => x"38",
          4912 => x"81",
          4913 => x"81",
          4914 => x"8a",
          4915 => x"06",
          4916 => x"76",
          4917 => x"76",
          4918 => x"55",
          4919 => x"e0",
          4920 => x"0d",
          4921 => x"0d",
          4922 => x"70",
          4923 => x"74",
          4924 => x"ea",
          4925 => x"74",
          4926 => x"14",
          4927 => x"de",
          4928 => x"55",
          4929 => x"55",
          4930 => x"2e",
          4931 => x"56",
          4932 => x"9f",
          4933 => x"51",
          4934 => x"38",
          4935 => x"09",
          4936 => x"38",
          4937 => x"81",
          4938 => x"72",
          4939 => x"29",
          4940 => x"05",
          4941 => x"70",
          4942 => x"fe",
          4943 => x"81",
          4944 => x"8b",
          4945 => x"33",
          4946 => x"2e",
          4947 => x"81",
          4948 => x"ff",
          4949 => x"96",
          4950 => x"38",
          4951 => x"81",
          4952 => x"88",
          4953 => x"ff",
          4954 => x"52",
          4955 => x"81",
          4956 => x"84",
          4957 => x"90",
          4958 => x"08",
          4959 => x"fc",
          4960 => x"39",
          4961 => x"51",
          4962 => x"81",
          4963 => x"80",
          4964 => x"df",
          4965 => x"eb",
          4966 => x"c0",
          4967 => x"39",
          4968 => x"51",
          4969 => x"81",
          4970 => x"80",
          4971 => x"df",
          4972 => x"cf",
          4973 => x"8c",
          4974 => x"39",
          4975 => x"51",
          4976 => x"81",
          4977 => x"bb",
          4978 => x"d8",
          4979 => x"81",
          4980 => x"af",
          4981 => x"98",
          4982 => x"81",
          4983 => x"a3",
          4984 => x"cc",
          4985 => x"81",
          4986 => x"97",
          4987 => x"f8",
          4988 => x"81",
          4989 => x"8b",
          4990 => x"a8",
          4991 => x"81",
          4992 => x"ff",
          4993 => x"83",
          4994 => x"fb",
          4995 => x"79",
          4996 => x"87",
          4997 => x"38",
          4998 => x"87",
          4999 => x"91",
          5000 => x"52",
          5001 => x"ee",
          5002 => x"ec",
          5003 => x"75",
          5004 => x"f7",
          5005 => x"e0",
          5006 => x"53",
          5007 => x"e2",
          5008 => x"8b",
          5009 => x"3d",
          5010 => x"3d",
          5011 => x"84",
          5012 => x"05",
          5013 => x"80",
          5014 => x"70",
          5015 => x"25",
          5016 => x"59",
          5017 => x"87",
          5018 => x"38",
          5019 => x"76",
          5020 => x"ff",
          5021 => x"93",
          5022 => x"ff",
          5023 => x"76",
          5024 => x"70",
          5025 => x"9d",
          5026 => x"e0",
          5027 => x"ec",
          5028 => x"38",
          5029 => x"08",
          5030 => x"88",
          5031 => x"e0",
          5032 => x"3d",
          5033 => x"84",
          5034 => x"52",
          5035 => x"da",
          5036 => x"e0",
          5037 => x"ec",
          5038 => x"38",
          5039 => x"80",
          5040 => x"74",
          5041 => x"59",
          5042 => x"96",
          5043 => x"51",
          5044 => x"76",
          5045 => x"07",
          5046 => x"30",
          5047 => x"72",
          5048 => x"51",
          5049 => x"2e",
          5050 => x"e2",
          5051 => x"c0",
          5052 => x"52",
          5053 => x"93",
          5054 => x"75",
          5055 => x"0c",
          5056 => x"04",
          5057 => x"7b",
          5058 => x"b3",
          5059 => x"58",
          5060 => x"53",
          5061 => x"51",
          5062 => x"81",
          5063 => x"a4",
          5064 => x"2e",
          5065 => x"81",
          5066 => x"98",
          5067 => x"7f",
          5068 => x"e0",
          5069 => x"7d",
          5070 => x"81",
          5071 => x"57",
          5072 => x"04",
          5073 => x"e0",
          5074 => x"0d",
          5075 => x"0d",
          5076 => x"02",
          5077 => x"cf",
          5078 => x"73",
          5079 => x"5f",
          5080 => x"5e",
          5081 => x"81",
          5082 => x"ff",
          5083 => x"81",
          5084 => x"ff",
          5085 => x"80",
          5086 => x"27",
          5087 => x"7b",
          5088 => x"38",
          5089 => x"a7",
          5090 => x"39",
          5091 => x"72",
          5092 => x"38",
          5093 => x"81",
          5094 => x"ff",
          5095 => x"89",
          5096 => x"88",
          5097 => x"fd",
          5098 => x"55",
          5099 => x"74",
          5100 => x"7a",
          5101 => x"72",
          5102 => x"e2",
          5103 => x"88",
          5104 => x"39",
          5105 => x"51",
          5106 => x"3f",
          5107 => x"a1",
          5108 => x"53",
          5109 => x"8e",
          5110 => x"52",
          5111 => x"51",
          5112 => x"3f",
          5113 => x"e3",
          5114 => x"82",
          5115 => x"15",
          5116 => x"ff",
          5117 => x"ff",
          5118 => x"e3",
          5119 => x"82",
          5120 => x"55",
          5121 => x"bc",
          5122 => x"70",
          5123 => x"80",
          5124 => x"27",
          5125 => x"56",
          5126 => x"74",
          5127 => x"81",
          5128 => x"06",
          5129 => x"06",
          5130 => x"80",
          5131 => x"73",
          5132 => x"85",
          5133 => x"83",
          5134 => x"ff",
          5135 => x"81",
          5136 => x"39",
          5137 => x"51",
          5138 => x"3f",
          5139 => x"1c",
          5140 => x"f6",
          5141 => x"ec",
          5142 => x"2b",
          5143 => x"51",
          5144 => x"2e",
          5145 => x"ab",
          5146 => x"c5",
          5147 => x"e0",
          5148 => x"70",
          5149 => x"a0",
          5150 => x"72",
          5151 => x"30",
          5152 => x"73",
          5153 => x"51",
          5154 => x"57",
          5155 => x"73",
          5156 => x"76",
          5157 => x"81",
          5158 => x"80",
          5159 => x"7c",
          5160 => x"78",
          5161 => x"38",
          5162 => x"81",
          5163 => x"8f",
          5164 => x"fc",
          5165 => x"9b",
          5166 => x"e3",
          5167 => x"e3",
          5168 => x"ff",
          5169 => x"81",
          5170 => x"51",
          5171 => x"3f",
          5172 => x"54",
          5173 => x"53",
          5174 => x"33",
          5175 => x"c8",
          5176 => x"a5",
          5177 => x"2e",
          5178 => x"fa",
          5179 => x"3d",
          5180 => x"3d",
          5181 => x"96",
          5182 => x"fe",
          5183 => x"81",
          5184 => x"c1",
          5185 => x"e4",
          5186 => x"b9",
          5187 => x"fe",
          5188 => x"72",
          5189 => x"81",
          5190 => x"71",
          5191 => x"38",
          5192 => x"f1",
          5193 => x"e3",
          5194 => x"f3",
          5195 => x"51",
          5196 => x"3f",
          5197 => x"70",
          5198 => x"52",
          5199 => x"95",
          5200 => x"fe",
          5201 => x"81",
          5202 => x"fe",
          5203 => x"80",
          5204 => x"f1",
          5205 => x"2a",
          5206 => x"51",
          5207 => x"2e",
          5208 => x"51",
          5209 => x"3f",
          5210 => x"51",
          5211 => x"3f",
          5212 => x"f0",
          5213 => x"84",
          5214 => x"06",
          5215 => x"80",
          5216 => x"81",
          5217 => x"bd",
          5218 => x"b4",
          5219 => x"b5",
          5220 => x"fe",
          5221 => x"72",
          5222 => x"81",
          5223 => x"71",
          5224 => x"38",
          5225 => x"f0",
          5226 => x"e4",
          5227 => x"f2",
          5228 => x"51",
          5229 => x"3f",
          5230 => x"70",
          5231 => x"52",
          5232 => x"95",
          5233 => x"fe",
          5234 => x"81",
          5235 => x"fe",
          5236 => x"80",
          5237 => x"ed",
          5238 => x"2a",
          5239 => x"51",
          5240 => x"2e",
          5241 => x"51",
          5242 => x"3f",
          5243 => x"51",
          5244 => x"3f",
          5245 => x"ef",
          5246 => x"88",
          5247 => x"06",
          5248 => x"80",
          5249 => x"81",
          5250 => x"b9",
          5251 => x"84",
          5252 => x"b1",
          5253 => x"fe",
          5254 => x"fe",
          5255 => x"84",
          5256 => x"fb",
          5257 => x"79",
          5258 => x"56",
          5259 => x"51",
          5260 => x"3f",
          5261 => x"33",
          5262 => x"38",
          5263 => x"e5",
          5264 => x"83",
          5265 => x"b9",
          5266 => x"ec",
          5267 => x"70",
          5268 => x"08",
          5269 => x"82",
          5270 => x"51",
          5271 => x"e9",
          5272 => x"e9",
          5273 => x"73",
          5274 => x"81",
          5275 => x"82",
          5276 => x"74",
          5277 => x"f4",
          5278 => x"ec",
          5279 => x"2e",
          5280 => x"ec",
          5281 => x"fe",
          5282 => x"8e",
          5283 => x"e4",
          5284 => x"3f",
          5285 => x"e9",
          5286 => x"e9",
          5287 => x"73",
          5288 => x"81",
          5289 => x"74",
          5290 => x"ff",
          5291 => x"80",
          5292 => x"e0",
          5293 => x"0d",
          5294 => x"0d",
          5295 => x"82",
          5296 => x"5f",
          5297 => x"7c",
          5298 => x"b4",
          5299 => x"e0",
          5300 => x"06",
          5301 => x"2e",
          5302 => x"a2",
          5303 => x"d4",
          5304 => x"70",
          5305 => x"82",
          5306 => x"53",
          5307 => x"ee",
          5308 => x"b7",
          5309 => x"ec",
          5310 => x"2e",
          5311 => x"e5",
          5312 => x"c1",
          5313 => x"5f",
          5314 => x"90",
          5315 => x"95",
          5316 => x"70",
          5317 => x"f8",
          5318 => x"fe",
          5319 => x"3d",
          5320 => x"51",
          5321 => x"81",
          5322 => x"90",
          5323 => x"2c",
          5324 => x"80",
          5325 => x"b3",
          5326 => x"c2",
          5327 => x"78",
          5328 => x"d5",
          5329 => x"24",
          5330 => x"80",
          5331 => x"38",
          5332 => x"80",
          5333 => x"e9",
          5334 => x"c0",
          5335 => x"38",
          5336 => x"24",
          5337 => x"78",
          5338 => x"92",
          5339 => x"39",
          5340 => x"2e",
          5341 => x"78",
          5342 => x"92",
          5343 => x"c3",
          5344 => x"38",
          5345 => x"2e",
          5346 => x"8a",
          5347 => x"81",
          5348 => x"99",
          5349 => x"83",
          5350 => x"78",
          5351 => x"89",
          5352 => x"9d",
          5353 => x"85",
          5354 => x"38",
          5355 => x"b4",
          5356 => x"11",
          5357 => x"05",
          5358 => x"c2",
          5359 => x"e0",
          5360 => x"fe",
          5361 => x"3d",
          5362 => x"53",
          5363 => x"51",
          5364 => x"3f",
          5365 => x"08",
          5366 => x"ad",
          5367 => x"fe",
          5368 => x"ff",
          5369 => x"ff",
          5370 => x"81",
          5371 => x"86",
          5372 => x"e0",
          5373 => x"e6",
          5374 => x"fa",
          5375 => x"63",
          5376 => x"7b",
          5377 => x"38",
          5378 => x"7a",
          5379 => x"5c",
          5380 => x"26",
          5381 => x"e1",
          5382 => x"ff",
          5383 => x"ff",
          5384 => x"ff",
          5385 => x"81",
          5386 => x"80",
          5387 => x"38",
          5388 => x"fc",
          5389 => x"84",
          5390 => x"81",
          5391 => x"ec",
          5392 => x"2e",
          5393 => x"b4",
          5394 => x"11",
          5395 => x"05",
          5396 => x"aa",
          5397 => x"e0",
          5398 => x"fd",
          5399 => x"e6",
          5400 => x"f9",
          5401 => x"5a",
          5402 => x"81",
          5403 => x"59",
          5404 => x"05",
          5405 => x"34",
          5406 => x"42",
          5407 => x"3d",
          5408 => x"53",
          5409 => x"51",
          5410 => x"3f",
          5411 => x"08",
          5412 => x"f5",
          5413 => x"fe",
          5414 => x"ff",
          5415 => x"ff",
          5416 => x"81",
          5417 => x"80",
          5418 => x"38",
          5419 => x"f8",
          5420 => x"84",
          5421 => x"80",
          5422 => x"ec",
          5423 => x"2e",
          5424 => x"81",
          5425 => x"fe",
          5426 => x"63",
          5427 => x"27",
          5428 => x"70",
          5429 => x"5e",
          5430 => x"7c",
          5431 => x"78",
          5432 => x"79",
          5433 => x"52",
          5434 => x"51",
          5435 => x"3f",
          5436 => x"81",
          5437 => x"d5",
          5438 => x"d8",
          5439 => x"39",
          5440 => x"80",
          5441 => x"84",
          5442 => x"ff",
          5443 => x"ec",
          5444 => x"df",
          5445 => x"d4",
          5446 => x"80",
          5447 => x"81",
          5448 => x"44",
          5449 => x"81",
          5450 => x"59",
          5451 => x"88",
          5452 => x"94",
          5453 => x"39",
          5454 => x"33",
          5455 => x"2e",
          5456 => x"e9",
          5457 => x"ab",
          5458 => x"d7",
          5459 => x"80",
          5460 => x"81",
          5461 => x"44",
          5462 => x"e9",
          5463 => x"78",
          5464 => x"38",
          5465 => x"08",
          5466 => x"81",
          5467 => x"fc",
          5468 => x"b4",
          5469 => x"11",
          5470 => x"05",
          5471 => x"fe",
          5472 => x"e0",
          5473 => x"38",
          5474 => x"33",
          5475 => x"2e",
          5476 => x"e9",
          5477 => x"80",
          5478 => x"e9",
          5479 => x"78",
          5480 => x"38",
          5481 => x"08",
          5482 => x"81",
          5483 => x"59",
          5484 => x"88",
          5485 => x"a0",
          5486 => x"39",
          5487 => x"33",
          5488 => x"2e",
          5489 => x"e9",
          5490 => x"99",
          5491 => x"d2",
          5492 => x"80",
          5493 => x"81",
          5494 => x"43",
          5495 => x"e9",
          5496 => x"05",
          5497 => x"fe",
          5498 => x"ff",
          5499 => x"fe",
          5500 => x"81",
          5501 => x"80",
          5502 => x"80",
          5503 => x"7a",
          5504 => x"38",
          5505 => x"90",
          5506 => x"70",
          5507 => x"2a",
          5508 => x"51",
          5509 => x"78",
          5510 => x"38",
          5511 => x"83",
          5512 => x"81",
          5513 => x"fe",
          5514 => x"a0",
          5515 => x"61",
          5516 => x"63",
          5517 => x"3f",
          5518 => x"51",
          5519 => x"3f",
          5520 => x"b4",
          5521 => x"11",
          5522 => x"05",
          5523 => x"ae",
          5524 => x"e0",
          5525 => x"f9",
          5526 => x"3d",
          5527 => x"53",
          5528 => x"51",
          5529 => x"3f",
          5530 => x"08",
          5531 => x"38",
          5532 => x"80",
          5533 => x"79",
          5534 => x"05",
          5535 => x"fe",
          5536 => x"ff",
          5537 => x"fe",
          5538 => x"81",
          5539 => x"e0",
          5540 => x"39",
          5541 => x"54",
          5542 => x"f8",
          5543 => x"e9",
          5544 => x"52",
          5545 => x"fb",
          5546 => x"45",
          5547 => x"78",
          5548 => x"d5",
          5549 => x"27",
          5550 => x"3d",
          5551 => x"53",
          5552 => x"51",
          5553 => x"3f",
          5554 => x"08",
          5555 => x"38",
          5556 => x"80",
          5557 => x"79",
          5558 => x"05",
          5559 => x"39",
          5560 => x"51",
          5561 => x"3f",
          5562 => x"b4",
          5563 => x"11",
          5564 => x"05",
          5565 => x"f8",
          5566 => x"e0",
          5567 => x"f8",
          5568 => x"3d",
          5569 => x"53",
          5570 => x"51",
          5571 => x"3f",
          5572 => x"08",
          5573 => x"38",
          5574 => x"be",
          5575 => x"70",
          5576 => x"23",
          5577 => x"3d",
          5578 => x"53",
          5579 => x"51",
          5580 => x"3f",
          5581 => x"08",
          5582 => x"cd",
          5583 => x"22",
          5584 => x"e7",
          5585 => x"f9",
          5586 => x"f8",
          5587 => x"fe",
          5588 => x"79",
          5589 => x"59",
          5590 => x"f7",
          5591 => x"9f",
          5592 => x"60",
          5593 => x"d5",
          5594 => x"fe",
          5595 => x"ff",
          5596 => x"fe",
          5597 => x"81",
          5598 => x"80",
          5599 => x"60",
          5600 => x"05",
          5601 => x"82",
          5602 => x"78",
          5603 => x"39",
          5604 => x"51",
          5605 => x"3f",
          5606 => x"b4",
          5607 => x"11",
          5608 => x"05",
          5609 => x"c8",
          5610 => x"e0",
          5611 => x"f6",
          5612 => x"3d",
          5613 => x"53",
          5614 => x"51",
          5615 => x"3f",
          5616 => x"08",
          5617 => x"38",
          5618 => x"0c",
          5619 => x"05",
          5620 => x"fe",
          5621 => x"ff",
          5622 => x"fe",
          5623 => x"81",
          5624 => x"e4",
          5625 => x"39",
          5626 => x"54",
          5627 => x"98",
          5628 => x"95",
          5629 => x"52",
          5630 => x"f8",
          5631 => x"45",
          5632 => x"78",
          5633 => x"81",
          5634 => x"27",
          5635 => x"3d",
          5636 => x"53",
          5637 => x"51",
          5638 => x"3f",
          5639 => x"08",
          5640 => x"38",
          5641 => x"0c",
          5642 => x"05",
          5643 => x"39",
          5644 => x"51",
          5645 => x"3f",
          5646 => x"b4",
          5647 => x"11",
          5648 => x"05",
          5649 => x"b6",
          5650 => x"e0",
          5651 => x"f5",
          5652 => x"52",
          5653 => x"51",
          5654 => x"3f",
          5655 => x"04",
          5656 => x"80",
          5657 => x"84",
          5658 => x"f9",
          5659 => x"ec",
          5660 => x"2e",
          5661 => x"63",
          5662 => x"c0",
          5663 => x"89",
          5664 => x"78",
          5665 => x"e0",
          5666 => x"f4",
          5667 => x"ec",
          5668 => x"81",
          5669 => x"fe",
          5670 => x"f4",
          5671 => x"e7",
          5672 => x"f1",
          5673 => x"d8",
          5674 => x"dd",
          5675 => x"94",
          5676 => x"f1",
          5677 => x"ff",
          5678 => x"eb",
          5679 => x"c9",
          5680 => x"33",
          5681 => x"80",
          5682 => x"38",
          5683 => x"59",
          5684 => x"81",
          5685 => x"3d",
          5686 => x"51",
          5687 => x"3f",
          5688 => x"08",
          5689 => x"7a",
          5690 => x"38",
          5691 => x"89",
          5692 => x"2e",
          5693 => x"cd",
          5694 => x"2e",
          5695 => x"c5",
          5696 => x"a8",
          5697 => x"81",
          5698 => x"80",
          5699 => x"b0",
          5700 => x"ff",
          5701 => x"fe",
          5702 => x"bb",
          5703 => x"d0",
          5704 => x"ff",
          5705 => x"fe",
          5706 => x"ab",
          5707 => x"81",
          5708 => x"80",
          5709 => x"c0",
          5710 => x"ff",
          5711 => x"fe",
          5712 => x"93",
          5713 => x"80",
          5714 => x"cc",
          5715 => x"ff",
          5716 => x"fe",
          5717 => x"81",
          5718 => x"81",
          5719 => x"80",
          5720 => x"11",
          5721 => x"55",
          5722 => x"80",
          5723 => x"80",
          5724 => x"3d",
          5725 => x"51",
          5726 => x"81",
          5727 => x"81",
          5728 => x"09",
          5729 => x"72",
          5730 => x"51",
          5731 => x"80",
          5732 => x"26",
          5733 => x"5a",
          5734 => x"59",
          5735 => x"8d",
          5736 => x"70",
          5737 => x"5c",
          5738 => x"bb",
          5739 => x"32",
          5740 => x"07",
          5741 => x"38",
          5742 => x"09",
          5743 => x"c9",
          5744 => x"d4",
          5745 => x"c1",
          5746 => x"39",
          5747 => x"80",
          5748 => x"94",
          5749 => x"94",
          5750 => x"54",
          5751 => x"80",
          5752 => x"fe",
          5753 => x"81",
          5754 => x"90",
          5755 => x"55",
          5756 => x"80",
          5757 => x"fe",
          5758 => x"72",
          5759 => x"08",
          5760 => x"87",
          5761 => x"70",
          5762 => x"87",
          5763 => x"72",
          5764 => x"97",
          5765 => x"e0",
          5766 => x"75",
          5767 => x"87",
          5768 => x"73",
          5769 => x"83",
          5770 => x"ec",
          5771 => x"75",
          5772 => x"83",
          5773 => x"94",
          5774 => x"80",
          5775 => x"c0",
          5776 => x"b3",
          5777 => x"ec",
          5778 => x"e0",
          5779 => x"f4",
          5780 => x"b5",
          5781 => x"de",
          5782 => x"e4",
          5783 => x"c5",
          5784 => x"f0",
          5785 => x"bd",
          5786 => x"f2",
          5787 => x"c1",
          5788 => x"ec",
          5789 => x"c1",
          5790 => x"00",
          5791 => x"88",
          5792 => x"8e",
          5793 => x"94",
          5794 => x"9a",
          5795 => x"a0",
          5796 => x"f9",
          5797 => x"7d",
          5798 => x"84",
          5799 => x"8b",
          5800 => x"92",
          5801 => x"99",
          5802 => x"a0",
          5803 => x"a7",
          5804 => x"ae",
          5805 => x"b5",
          5806 => x"bc",
          5807 => x"c3",
          5808 => x"c9",
          5809 => x"cf",
          5810 => x"d5",
          5811 => x"db",
          5812 => x"e1",
          5813 => x"e7",
          5814 => x"ed",
          5815 => x"f3",
          5816 => x"25",
          5817 => x"64",
          5818 => x"3a",
          5819 => x"25",
          5820 => x"64",
          5821 => x"00",
          5822 => x"20",
          5823 => x"66",
          5824 => x"72",
          5825 => x"6f",
          5826 => x"00",
          5827 => x"72",
          5828 => x"53",
          5829 => x"63",
          5830 => x"69",
          5831 => x"00",
          5832 => x"65",
          5833 => x"65",
          5834 => x"6d",
          5835 => x"6d",
          5836 => x"65",
          5837 => x"00",
          5838 => x"20",
          5839 => x"53",
          5840 => x"4d",
          5841 => x"25",
          5842 => x"3a",
          5843 => x"58",
          5844 => x"00",
          5845 => x"20",
          5846 => x"41",
          5847 => x"20",
          5848 => x"25",
          5849 => x"3a",
          5850 => x"58",
          5851 => x"00",
          5852 => x"20",
          5853 => x"4e",
          5854 => x"41",
          5855 => x"25",
          5856 => x"3a",
          5857 => x"58",
          5858 => x"00",
          5859 => x"20",
          5860 => x"4d",
          5861 => x"20",
          5862 => x"25",
          5863 => x"3a",
          5864 => x"58",
          5865 => x"00",
          5866 => x"20",
          5867 => x"20",
          5868 => x"20",
          5869 => x"25",
          5870 => x"3a",
          5871 => x"58",
          5872 => x"00",
          5873 => x"20",
          5874 => x"43",
          5875 => x"20",
          5876 => x"44",
          5877 => x"63",
          5878 => x"3d",
          5879 => x"64",
          5880 => x"00",
          5881 => x"20",
          5882 => x"45",
          5883 => x"20",
          5884 => x"54",
          5885 => x"72",
          5886 => x"3d",
          5887 => x"64",
          5888 => x"00",
          5889 => x"20",
          5890 => x"52",
          5891 => x"52",
          5892 => x"43",
          5893 => x"6e",
          5894 => x"3d",
          5895 => x"64",
          5896 => x"00",
          5897 => x"20",
          5898 => x"48",
          5899 => x"45",
          5900 => x"53",
          5901 => x"00",
          5902 => x"20",
          5903 => x"49",
          5904 => x"00",
          5905 => x"20",
          5906 => x"54",
          5907 => x"00",
          5908 => x"20",
          5909 => x"0a",
          5910 => x"00",
          5911 => x"20",
          5912 => x"0a",
          5913 => x"00",
          5914 => x"72",
          5915 => x"65",
          5916 => x"00",
          5917 => x"20",
          5918 => x"20",
          5919 => x"65",
          5920 => x"65",
          5921 => x"72",
          5922 => x"64",
          5923 => x"73",
          5924 => x"25",
          5925 => x"0a",
          5926 => x"00",
          5927 => x"20",
          5928 => x"20",
          5929 => x"6f",
          5930 => x"53",
          5931 => x"74",
          5932 => x"64",
          5933 => x"73",
          5934 => x"25",
          5935 => x"0a",
          5936 => x"00",
          5937 => x"20",
          5938 => x"63",
          5939 => x"74",
          5940 => x"20",
          5941 => x"72",
          5942 => x"20",
          5943 => x"20",
          5944 => x"25",
          5945 => x"0a",
          5946 => x"00",
          5947 => x"63",
          5948 => x"00",
          5949 => x"20",
          5950 => x"20",
          5951 => x"20",
          5952 => x"20",
          5953 => x"20",
          5954 => x"20",
          5955 => x"20",
          5956 => x"25",
          5957 => x"0a",
          5958 => x"00",
          5959 => x"20",
          5960 => x"74",
          5961 => x"43",
          5962 => x"6b",
          5963 => x"65",
          5964 => x"20",
          5965 => x"20",
          5966 => x"25",
          5967 => x"30",
          5968 => x"48",
          5969 => x"00",
          5970 => x"20",
          5971 => x"41",
          5972 => x"6c",
          5973 => x"20",
          5974 => x"71",
          5975 => x"20",
          5976 => x"20",
          5977 => x"25",
          5978 => x"30",
          5979 => x"48",
          5980 => x"00",
          5981 => x"20",
          5982 => x"68",
          5983 => x"65",
          5984 => x"52",
          5985 => x"43",
          5986 => x"6b",
          5987 => x"65",
          5988 => x"25",
          5989 => x"30",
          5990 => x"48",
          5991 => x"00",
          5992 => x"6c",
          5993 => x"00",
          5994 => x"69",
          5995 => x"00",
          5996 => x"78",
          5997 => x"00",
          5998 => x"00",
          5999 => x"6d",
          6000 => x"00",
          6001 => x"6e",
          6002 => x"00",
          6003 => x"00",
          6004 => x"2c",
          6005 => x"3d",
          6006 => x"5d",
          6007 => x"00",
          6008 => x"00",
          6009 => x"33",
          6010 => x"00",
          6011 => x"4d",
          6012 => x"53",
          6013 => x"00",
          6014 => x"4e",
          6015 => x"20",
          6016 => x"46",
          6017 => x"32",
          6018 => x"00",
          6019 => x"4e",
          6020 => x"20",
          6021 => x"46",
          6022 => x"20",
          6023 => x"00",
          6024 => x"cc",
          6025 => x"00",
          6026 => x"00",
          6027 => x"00",
          6028 => x"41",
          6029 => x"80",
          6030 => x"49",
          6031 => x"8f",
          6032 => x"4f",
          6033 => x"55",
          6034 => x"9b",
          6035 => x"9f",
          6036 => x"55",
          6037 => x"a7",
          6038 => x"ab",
          6039 => x"af",
          6040 => x"b3",
          6041 => x"b7",
          6042 => x"bb",
          6043 => x"bf",
          6044 => x"c3",
          6045 => x"c7",
          6046 => x"cb",
          6047 => x"cf",
          6048 => x"d3",
          6049 => x"d7",
          6050 => x"db",
          6051 => x"df",
          6052 => x"e3",
          6053 => x"e7",
          6054 => x"eb",
          6055 => x"ef",
          6056 => x"f3",
          6057 => x"f7",
          6058 => x"fb",
          6059 => x"ff",
          6060 => x"3b",
          6061 => x"2f",
          6062 => x"3a",
          6063 => x"7c",
          6064 => x"00",
          6065 => x"04",
          6066 => x"40",
          6067 => x"00",
          6068 => x"00",
          6069 => x"02",
          6070 => x"08",
          6071 => x"20",
          6072 => x"00",
          6073 => x"69",
          6074 => x"00",
          6075 => x"63",
          6076 => x"00",
          6077 => x"69",
          6078 => x"00",
          6079 => x"61",
          6080 => x"00",
          6081 => x"65",
          6082 => x"00",
          6083 => x"65",
          6084 => x"00",
          6085 => x"70",
          6086 => x"00",
          6087 => x"66",
          6088 => x"00",
          6089 => x"6d",
          6090 => x"00",
          6091 => x"00",
          6092 => x"00",
          6093 => x"00",
          6094 => x"00",
          6095 => x"00",
          6096 => x"00",
          6097 => x"00",
          6098 => x"6c",
          6099 => x"00",
          6100 => x"00",
          6101 => x"74",
          6102 => x"00",
          6103 => x"65",
          6104 => x"00",
          6105 => x"6f",
          6106 => x"00",
          6107 => x"74",
          6108 => x"00",
          6109 => x"73",
          6110 => x"00",
          6111 => x"6b",
          6112 => x"72",
          6113 => x"00",
          6114 => x"65",
          6115 => x"6c",
          6116 => x"72",
          6117 => x"0a",
          6118 => x"00",
          6119 => x"6b",
          6120 => x"74",
          6121 => x"61",
          6122 => x"0a",
          6123 => x"00",
          6124 => x"66",
          6125 => x"20",
          6126 => x"6e",
          6127 => x"00",
          6128 => x"70",
          6129 => x"20",
          6130 => x"6e",
          6131 => x"00",
          6132 => x"61",
          6133 => x"20",
          6134 => x"65",
          6135 => x"65",
          6136 => x"00",
          6137 => x"65",
          6138 => x"64",
          6139 => x"65",
          6140 => x"00",
          6141 => x"65",
          6142 => x"72",
          6143 => x"79",
          6144 => x"69",
          6145 => x"2e",
          6146 => x"00",
          6147 => x"65",
          6148 => x"6e",
          6149 => x"20",
          6150 => x"61",
          6151 => x"2e",
          6152 => x"00",
          6153 => x"69",
          6154 => x"72",
          6155 => x"20",
          6156 => x"74",
          6157 => x"65",
          6158 => x"00",
          6159 => x"76",
          6160 => x"75",
          6161 => x"72",
          6162 => x"20",
          6163 => x"61",
          6164 => x"2e",
          6165 => x"00",
          6166 => x"6b",
          6167 => x"74",
          6168 => x"61",
          6169 => x"64",
          6170 => x"00",
          6171 => x"63",
          6172 => x"61",
          6173 => x"6c",
          6174 => x"69",
          6175 => x"79",
          6176 => x"6d",
          6177 => x"75",
          6178 => x"6f",
          6179 => x"69",
          6180 => x"0a",
          6181 => x"00",
          6182 => x"6d",
          6183 => x"61",
          6184 => x"74",
          6185 => x"0a",
          6186 => x"00",
          6187 => x"65",
          6188 => x"2c",
          6189 => x"65",
          6190 => x"69",
          6191 => x"63",
          6192 => x"65",
          6193 => x"64",
          6194 => x"00",
          6195 => x"65",
          6196 => x"20",
          6197 => x"6b",
          6198 => x"0a",
          6199 => x"00",
          6200 => x"75",
          6201 => x"63",
          6202 => x"74",
          6203 => x"6d",
          6204 => x"2e",
          6205 => x"00",
          6206 => x"20",
          6207 => x"79",
          6208 => x"65",
          6209 => x"69",
          6210 => x"2e",
          6211 => x"00",
          6212 => x"61",
          6213 => x"65",
          6214 => x"69",
          6215 => x"72",
          6216 => x"74",
          6217 => x"00",
          6218 => x"63",
          6219 => x"2e",
          6220 => x"00",
          6221 => x"6e",
          6222 => x"20",
          6223 => x"6f",
          6224 => x"00",
          6225 => x"75",
          6226 => x"74",
          6227 => x"25",
          6228 => x"74",
          6229 => x"75",
          6230 => x"74",
          6231 => x"73",
          6232 => x"0a",
          6233 => x"00",
          6234 => x"64",
          6235 => x"00",
          6236 => x"58",
          6237 => x"00",
          6238 => x"00",
          6239 => x"58",
          6240 => x"00",
          6241 => x"20",
          6242 => x"20",
          6243 => x"00",
          6244 => x"58",
          6245 => x"00",
          6246 => x"00",
          6247 => x"00",
          6248 => x"00",
          6249 => x"00",
          6250 => x"20",
          6251 => x"28",
          6252 => x"00",
          6253 => x"30",
          6254 => x"30",
          6255 => x"00",
          6256 => x"30",
          6257 => x"00",
          6258 => x"55",
          6259 => x"65",
          6260 => x"30",
          6261 => x"20",
          6262 => x"25",
          6263 => x"2a",
          6264 => x"00",
          6265 => x"20",
          6266 => x"65",
          6267 => x"70",
          6268 => x"61",
          6269 => x"65",
          6270 => x"00",
          6271 => x"65",
          6272 => x"6e",
          6273 => x"72",
          6274 => x"0a",
          6275 => x"00",
          6276 => x"20",
          6277 => x"65",
          6278 => x"70",
          6279 => x"00",
          6280 => x"54",
          6281 => x"44",
          6282 => x"74",
          6283 => x"75",
          6284 => x"00",
          6285 => x"54",
          6286 => x"52",
          6287 => x"74",
          6288 => x"75",
          6289 => x"00",
          6290 => x"54",
          6291 => x"58",
          6292 => x"74",
          6293 => x"75",
          6294 => x"00",
          6295 => x"54",
          6296 => x"58",
          6297 => x"74",
          6298 => x"75",
          6299 => x"00",
          6300 => x"54",
          6301 => x"58",
          6302 => x"74",
          6303 => x"75",
          6304 => x"00",
          6305 => x"54",
          6306 => x"58",
          6307 => x"74",
          6308 => x"75",
          6309 => x"00",
          6310 => x"74",
          6311 => x"20",
          6312 => x"74",
          6313 => x"72",
          6314 => x"0a",
          6315 => x"00",
          6316 => x"62",
          6317 => x"67",
          6318 => x"6d",
          6319 => x"2e",
          6320 => x"00",
          6321 => x"6f",
          6322 => x"63",
          6323 => x"74",
          6324 => x"00",
          6325 => x"00",
          6326 => x"6c",
          6327 => x"74",
          6328 => x"6e",
          6329 => x"61",
          6330 => x"65",
          6331 => x"20",
          6332 => x"64",
          6333 => x"20",
          6334 => x"61",
          6335 => x"69",
          6336 => x"20",
          6337 => x"75",
          6338 => x"79",
          6339 => x"00",
          6340 => x"00",
          6341 => x"61",
          6342 => x"67",
          6343 => x"2e",
          6344 => x"00",
          6345 => x"79",
          6346 => x"2e",
          6347 => x"00",
          6348 => x"70",
          6349 => x"6e",
          6350 => x"2e",
          6351 => x"00",
          6352 => x"6c",
          6353 => x"30",
          6354 => x"2d",
          6355 => x"38",
          6356 => x"25",
          6357 => x"29",
          6358 => x"00",
          6359 => x"70",
          6360 => x"6d",
          6361 => x"0a",
          6362 => x"00",
          6363 => x"6d",
          6364 => x"74",
          6365 => x"00",
          6366 => x"58",
          6367 => x"32",
          6368 => x"00",
          6369 => x"0a",
          6370 => x"00",
          6371 => x"58",
          6372 => x"34",
          6373 => x"00",
          6374 => x"58",
          6375 => x"38",
          6376 => x"00",
          6377 => x"63",
          6378 => x"6e",
          6379 => x"6f",
          6380 => x"40",
          6381 => x"38",
          6382 => x"2e",
          6383 => x"00",
          6384 => x"6c",
          6385 => x"20",
          6386 => x"65",
          6387 => x"25",
          6388 => x"20",
          6389 => x"0a",
          6390 => x"00",
          6391 => x"6c",
          6392 => x"74",
          6393 => x"65",
          6394 => x"6f",
          6395 => x"28",
          6396 => x"2e",
          6397 => x"00",
          6398 => x"74",
          6399 => x"69",
          6400 => x"61",
          6401 => x"69",
          6402 => x"69",
          6403 => x"2e",
          6404 => x"00",
          6405 => x"64",
          6406 => x"62",
          6407 => x"69",
          6408 => x"2e",
          6409 => x"00",
          6410 => x"00",
          6411 => x"00",
          6412 => x"5c",
          6413 => x"25",
          6414 => x"73",
          6415 => x"00",
          6416 => x"5c",
          6417 => x"25",
          6418 => x"00",
          6419 => x"5c",
          6420 => x"00",
          6421 => x"20",
          6422 => x"6d",
          6423 => x"2e",
          6424 => x"00",
          6425 => x"6e",
          6426 => x"2e",
          6427 => x"00",
          6428 => x"62",
          6429 => x"67",
          6430 => x"74",
          6431 => x"75",
          6432 => x"2e",
          6433 => x"00",
          6434 => x"00",
          6435 => x"00",
          6436 => x"ff",
          6437 => x"00",
          6438 => x"ff",
          6439 => x"00",
          6440 => x"ff",
          6441 => x"00",
          6442 => x"00",
          6443 => x"00",
          6444 => x"ff",
          6445 => x"00",
          6446 => x"00",
          6447 => x"00",
          6448 => x"00",
          6449 => x"00",
          6450 => x"00",
          6451 => x"00",
          6452 => x"00",
          6453 => x"01",
          6454 => x"01",
          6455 => x"01",
          6456 => x"00",
          6457 => x"00",
          6458 => x"00",
          6459 => x"00",
          6460 => x"e4",
          6461 => x"00",
          6462 => x"00",
          6463 => x"00",
          6464 => x"ec",
          6465 => x"00",
          6466 => x"00",
          6467 => x"00",
          6468 => x"f4",
          6469 => x"00",
          6470 => x"00",
          6471 => x"00",
          6472 => x"fc",
          6473 => x"00",
          6474 => x"00",
          6475 => x"00",
          6476 => x"04",
          6477 => x"00",
          6478 => x"00",
          6479 => x"00",
          6480 => x"0c",
          6481 => x"00",
          6482 => x"00",
          6483 => x"00",
          6484 => x"14",
          6485 => x"00",
          6486 => x"00",
          6487 => x"00",
          6488 => x"1c",
          6489 => x"00",
          6490 => x"00",
          6491 => x"00",
          6492 => x"24",
          6493 => x"00",
          6494 => x"00",
          6495 => x"00",
          6496 => x"2c",
          6497 => x"00",
          6498 => x"00",
          6499 => x"00",
          6500 => x"30",
          6501 => x"00",
          6502 => x"00",
          6503 => x"00",
          6504 => x"34",
          6505 => x"00",
          6506 => x"00",
          6507 => x"00",
          6508 => x"38",
          6509 => x"00",
          6510 => x"00",
          6511 => x"00",
          6512 => x"3c",
          6513 => x"00",
          6514 => x"00",
          6515 => x"00",
          6516 => x"40",
          6517 => x"00",
          6518 => x"00",
          6519 => x"00",
          6520 => x"44",
          6521 => x"00",
          6522 => x"00",
          6523 => x"00",
          6524 => x"48",
          6525 => x"00",
          6526 => x"00",
          6527 => x"00",
          6528 => x"50",
          6529 => x"00",
          6530 => x"00",
          6531 => x"00",
          6532 => x"54",
          6533 => x"00",
          6534 => x"00",
          6535 => x"00",
          6536 => x"5c",
          6537 => x"00",
          6538 => x"00",
          6539 => x"00",
          6540 => x"64",
          6541 => x"00",
          6542 => x"00",
          6543 => x"00",
          6544 => x"6c",
          6545 => x"00",
          6546 => x"00",
          6547 => x"00",
          6548 => x"74",
          6549 => x"00",
          6550 => x"00",
          6551 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"8b",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"0b",
            10 => x"84",
            11 => x"0b",
            12 => x"0b",
            13 => x"a3",
            14 => x"0b",
            15 => x"0b",
            16 => x"c3",
            17 => x"0b",
            18 => x"0b",
            19 => x"e3",
            20 => x"0b",
            21 => x"0b",
            22 => x"83",
            23 => x"0b",
            24 => x"0b",
            25 => x"a3",
            26 => x"0b",
            27 => x"0b",
            28 => x"c3",
            29 => x"0b",
            30 => x"0b",
            31 => x"e1",
            32 => x"0b",
            33 => x"0b",
            34 => x"ff",
            35 => x"0b",
            36 => x"0b",
            37 => x"9e",
            38 => x"0b",
            39 => x"0b",
            40 => x"be",
            41 => x"0b",
            42 => x"0b",
            43 => x"de",
            44 => x"0b",
            45 => x"0b",
            46 => x"fe",
            47 => x"0b",
            48 => x"0b",
            49 => x"9e",
            50 => x"0b",
            51 => x"0b",
            52 => x"be",
            53 => x"0b",
            54 => x"0b",
            55 => x"de",
            56 => x"0b",
            57 => x"0b",
            58 => x"fe",
            59 => x"0b",
            60 => x"0b",
            61 => x"9e",
            62 => x"0b",
            63 => x"0b",
            64 => x"be",
            65 => x"0b",
            66 => x"0b",
            67 => x"de",
            68 => x"0b",
            69 => x"0b",
            70 => x"fe",
            71 => x"0b",
            72 => x"0b",
            73 => x"9e",
            74 => x"0b",
            75 => x"0b",
            76 => x"be",
            77 => x"0b",
            78 => x"0b",
            79 => x"dd",
            80 => x"0b",
            81 => x"0b",
            82 => x"fb",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"80",
           129 => x"ec",
           130 => x"2d",
           131 => x"08",
           132 => x"04",
           133 => x"0c",
           134 => x"2d",
           135 => x"08",
           136 => x"04",
           137 => x"0c",
           138 => x"2d",
           139 => x"08",
           140 => x"04",
           141 => x"0c",
           142 => x"2d",
           143 => x"08",
           144 => x"04",
           145 => x"0c",
           146 => x"2d",
           147 => x"08",
           148 => x"04",
           149 => x"0c",
           150 => x"2d",
           151 => x"08",
           152 => x"04",
           153 => x"0c",
           154 => x"2d",
           155 => x"08",
           156 => x"04",
           157 => x"0c",
           158 => x"2d",
           159 => x"08",
           160 => x"04",
           161 => x"0c",
           162 => x"2d",
           163 => x"08",
           164 => x"04",
           165 => x"0c",
           166 => x"2d",
           167 => x"08",
           168 => x"04",
           169 => x"0c",
           170 => x"2d",
           171 => x"08",
           172 => x"04",
           173 => x"0c",
           174 => x"2d",
           175 => x"08",
           176 => x"04",
           177 => x"0c",
           178 => x"81",
           179 => x"83",
           180 => x"81",
           181 => x"b7",
           182 => x"ec",
           183 => x"80",
           184 => x"ec",
           185 => x"cd",
           186 => x"ec",
           187 => x"90",
           188 => x"ec",
           189 => x"2d",
           190 => x"08",
           191 => x"04",
           192 => x"0c",
           193 => x"81",
           194 => x"83",
           195 => x"81",
           196 => x"80",
           197 => x"81",
           198 => x"83",
           199 => x"81",
           200 => x"81",
           201 => x"81",
           202 => x"83",
           203 => x"81",
           204 => x"81",
           205 => x"81",
           206 => x"83",
           207 => x"81",
           208 => x"81",
           209 => x"81",
           210 => x"83",
           211 => x"81",
           212 => x"81",
           213 => x"81",
           214 => x"83",
           215 => x"81",
           216 => x"81",
           217 => x"81",
           218 => x"83",
           219 => x"81",
           220 => x"81",
           221 => x"81",
           222 => x"83",
           223 => x"81",
           224 => x"81",
           225 => x"81",
           226 => x"83",
           227 => x"81",
           228 => x"81",
           229 => x"81",
           230 => x"83",
           231 => x"81",
           232 => x"81",
           233 => x"81",
           234 => x"83",
           235 => x"81",
           236 => x"81",
           237 => x"81",
           238 => x"83",
           239 => x"81",
           240 => x"81",
           241 => x"81",
           242 => x"83",
           243 => x"81",
           244 => x"81",
           245 => x"81",
           246 => x"83",
           247 => x"81",
           248 => x"81",
           249 => x"81",
           250 => x"83",
           251 => x"81",
           252 => x"81",
           253 => x"81",
           254 => x"83",
           255 => x"81",
           256 => x"81",
           257 => x"81",
           258 => x"83",
           259 => x"81",
           260 => x"81",
           261 => x"81",
           262 => x"83",
           263 => x"81",
           264 => x"81",
           265 => x"81",
           266 => x"83",
           267 => x"81",
           268 => x"81",
           269 => x"81",
           270 => x"83",
           271 => x"81",
           272 => x"81",
           273 => x"81",
           274 => x"83",
           275 => x"81",
           276 => x"81",
           277 => x"81",
           278 => x"83",
           279 => x"81",
           280 => x"81",
           281 => x"81",
           282 => x"83",
           283 => x"81",
           284 => x"81",
           285 => x"81",
           286 => x"83",
           287 => x"81",
           288 => x"80",
           289 => x"81",
           290 => x"83",
           291 => x"81",
           292 => x"81",
           293 => x"81",
           294 => x"83",
           295 => x"81",
           296 => x"80",
           297 => x"81",
           298 => x"83",
           299 => x"81",
           300 => x"80",
           301 => x"81",
           302 => x"83",
           303 => x"81",
           304 => x"80",
           305 => x"81",
           306 => x"83",
           307 => x"81",
           308 => x"af",
           309 => x"ec",
           310 => x"80",
           311 => x"ec",
           312 => x"d8",
           313 => x"ec",
           314 => x"90",
           315 => x"ec",
           316 => x"2d",
           317 => x"08",
           318 => x"04",
           319 => x"0c",
           320 => x"2d",
           321 => x"08",
           322 => x"04",
           323 => x"70",
           324 => x"27",
           325 => x"71",
           326 => x"53",
           327 => x"0b",
           328 => x"a4",
           329 => x"d3",
           330 => x"04",
           331 => x"08",
           332 => x"ec",
           333 => x"0d",
           334 => x"ec",
           335 => x"05",
           336 => x"ec",
           337 => x"05",
           338 => x"c5",
           339 => x"e0",
           340 => x"ec",
           341 => x"85",
           342 => x"ec",
           343 => x"81",
           344 => x"02",
           345 => x"0c",
           346 => x"81",
           347 => x"ec",
           348 => x"08",
           349 => x"ec",
           350 => x"08",
           351 => x"81",
           352 => x"70",
           353 => x"0c",
           354 => x"0d",
           355 => x"0c",
           356 => x"ec",
           357 => x"ec",
           358 => x"3d",
           359 => x"81",
           360 => x"fc",
           361 => x"0b",
           362 => x"08",
           363 => x"81",
           364 => x"8c",
           365 => x"ec",
           366 => x"05",
           367 => x"38",
           368 => x"08",
           369 => x"80",
           370 => x"80",
           371 => x"ec",
           372 => x"08",
           373 => x"81",
           374 => x"8c",
           375 => x"81",
           376 => x"8c",
           377 => x"ec",
           378 => x"05",
           379 => x"ec",
           380 => x"05",
           381 => x"39",
           382 => x"08",
           383 => x"80",
           384 => x"38",
           385 => x"08",
           386 => x"81",
           387 => x"88",
           388 => x"ad",
           389 => x"ec",
           390 => x"08",
           391 => x"08",
           392 => x"31",
           393 => x"08",
           394 => x"81",
           395 => x"f8",
           396 => x"ec",
           397 => x"05",
           398 => x"ec",
           399 => x"05",
           400 => x"ec",
           401 => x"08",
           402 => x"ec",
           403 => x"05",
           404 => x"ec",
           405 => x"08",
           406 => x"ec",
           407 => x"05",
           408 => x"39",
           409 => x"08",
           410 => x"80",
           411 => x"81",
           412 => x"88",
           413 => x"81",
           414 => x"f4",
           415 => x"91",
           416 => x"ec",
           417 => x"08",
           418 => x"ec",
           419 => x"0c",
           420 => x"ec",
           421 => x"08",
           422 => x"0c",
           423 => x"81",
           424 => x"04",
           425 => x"76",
           426 => x"8c",
           427 => x"33",
           428 => x"55",
           429 => x"8a",
           430 => x"06",
           431 => x"2e",
           432 => x"12",
           433 => x"2e",
           434 => x"73",
           435 => x"55",
           436 => x"52",
           437 => x"09",
           438 => x"38",
           439 => x"e0",
           440 => x"0d",
           441 => x"88",
           442 => x"70",
           443 => x"07",
           444 => x"8f",
           445 => x"38",
           446 => x"84",
           447 => x"72",
           448 => x"05",
           449 => x"71",
           450 => x"53",
           451 => x"70",
           452 => x"0c",
           453 => x"71",
           454 => x"38",
           455 => x"90",
           456 => x"70",
           457 => x"0c",
           458 => x"71",
           459 => x"38",
           460 => x"8e",
           461 => x"0d",
           462 => x"72",
           463 => x"53",
           464 => x"93",
           465 => x"73",
           466 => x"54",
           467 => x"2e",
           468 => x"73",
           469 => x"71",
           470 => x"ff",
           471 => x"70",
           472 => x"38",
           473 => x"70",
           474 => x"81",
           475 => x"81",
           476 => x"71",
           477 => x"ff",
           478 => x"54",
           479 => x"38",
           480 => x"73",
           481 => x"75",
           482 => x"71",
           483 => x"ec",
           484 => x"52",
           485 => x"04",
           486 => x"f7",
           487 => x"14",
           488 => x"84",
           489 => x"06",
           490 => x"70",
           491 => x"14",
           492 => x"08",
           493 => x"71",
           494 => x"dc",
           495 => x"54",
           496 => x"39",
           497 => x"ec",
           498 => x"3d",
           499 => x"3d",
           500 => x"83",
           501 => x"2b",
           502 => x"3f",
           503 => x"08",
           504 => x"72",
           505 => x"54",
           506 => x"25",
           507 => x"81",
           508 => x"84",
           509 => x"fb",
           510 => x"70",
           511 => x"53",
           512 => x"2e",
           513 => x"71",
           514 => x"a0",
           515 => x"06",
           516 => x"12",
           517 => x"71",
           518 => x"81",
           519 => x"73",
           520 => x"ff",
           521 => x"55",
           522 => x"83",
           523 => x"70",
           524 => x"38",
           525 => x"73",
           526 => x"51",
           527 => x"09",
           528 => x"38",
           529 => x"81",
           530 => x"72",
           531 => x"51",
           532 => x"e0",
           533 => x"0d",
           534 => x"0d",
           535 => x"08",
           536 => x"38",
           537 => x"05",
           538 => x"9b",
           539 => x"ec",
           540 => x"38",
           541 => x"39",
           542 => x"81",
           543 => x"86",
           544 => x"fc",
           545 => x"82",
           546 => x"05",
           547 => x"52",
           548 => x"81",
           549 => x"13",
           550 => x"51",
           551 => x"9e",
           552 => x"38",
           553 => x"51",
           554 => x"97",
           555 => x"38",
           556 => x"51",
           557 => x"bb",
           558 => x"38",
           559 => x"51",
           560 => x"bb",
           561 => x"38",
           562 => x"55",
           563 => x"87",
           564 => x"d9",
           565 => x"22",
           566 => x"73",
           567 => x"80",
           568 => x"0b",
           569 => x"9c",
           570 => x"87",
           571 => x"0c",
           572 => x"87",
           573 => x"0c",
           574 => x"87",
           575 => x"0c",
           576 => x"87",
           577 => x"0c",
           578 => x"87",
           579 => x"0c",
           580 => x"87",
           581 => x"0c",
           582 => x"98",
           583 => x"87",
           584 => x"0c",
           585 => x"c0",
           586 => x"80",
           587 => x"ec",
           588 => x"3d",
           589 => x"3d",
           590 => x"87",
           591 => x"5d",
           592 => x"87",
           593 => x"08",
           594 => x"23",
           595 => x"b8",
           596 => x"82",
           597 => x"c0",
           598 => x"5a",
           599 => x"34",
           600 => x"b0",
           601 => x"84",
           602 => x"c0",
           603 => x"5a",
           604 => x"34",
           605 => x"a8",
           606 => x"86",
           607 => x"c0",
           608 => x"5c",
           609 => x"23",
           610 => x"a0",
           611 => x"8a",
           612 => x"7d",
           613 => x"ff",
           614 => x"7b",
           615 => x"06",
           616 => x"33",
           617 => x"33",
           618 => x"33",
           619 => x"33",
           620 => x"33",
           621 => x"ff",
           622 => x"81",
           623 => x"94",
           624 => x"3d",
           625 => x"3d",
           626 => x"05",
           627 => x"70",
           628 => x"52",
           629 => x"0b",
           630 => x"34",
           631 => x"04",
           632 => x"77",
           633 => x"e9",
           634 => x"81",
           635 => x"55",
           636 => x"94",
           637 => x"80",
           638 => x"87",
           639 => x"51",
           640 => x"96",
           641 => x"06",
           642 => x"70",
           643 => x"38",
           644 => x"70",
           645 => x"51",
           646 => x"72",
           647 => x"81",
           648 => x"70",
           649 => x"38",
           650 => x"70",
           651 => x"51",
           652 => x"38",
           653 => x"06",
           654 => x"94",
           655 => x"80",
           656 => x"87",
           657 => x"52",
           658 => x"75",
           659 => x"0c",
           660 => x"04",
           661 => x"02",
           662 => x"0b",
           663 => x"88",
           664 => x"ff",
           665 => x"56",
           666 => x"84",
           667 => x"2e",
           668 => x"c0",
           669 => x"70",
           670 => x"2a",
           671 => x"53",
           672 => x"80",
           673 => x"71",
           674 => x"81",
           675 => x"70",
           676 => x"81",
           677 => x"06",
           678 => x"80",
           679 => x"71",
           680 => x"81",
           681 => x"70",
           682 => x"73",
           683 => x"51",
           684 => x"80",
           685 => x"2e",
           686 => x"c0",
           687 => x"75",
           688 => x"3d",
           689 => x"3d",
           690 => x"80",
           691 => x"81",
           692 => x"53",
           693 => x"2e",
           694 => x"71",
           695 => x"81",
           696 => x"81",
           697 => x"70",
           698 => x"59",
           699 => x"87",
           700 => x"51",
           701 => x"86",
           702 => x"94",
           703 => x"08",
           704 => x"70",
           705 => x"54",
           706 => x"2e",
           707 => x"91",
           708 => x"06",
           709 => x"d7",
           710 => x"32",
           711 => x"51",
           712 => x"2e",
           713 => x"93",
           714 => x"06",
           715 => x"ff",
           716 => x"81",
           717 => x"87",
           718 => x"52",
           719 => x"86",
           720 => x"94",
           721 => x"72",
           722 => x"74",
           723 => x"ff",
           724 => x"57",
           725 => x"38",
           726 => x"e0",
           727 => x"0d",
           728 => x"0d",
           729 => x"e9",
           730 => x"81",
           731 => x"52",
           732 => x"84",
           733 => x"2e",
           734 => x"c0",
           735 => x"70",
           736 => x"2a",
           737 => x"51",
           738 => x"80",
           739 => x"71",
           740 => x"51",
           741 => x"80",
           742 => x"2e",
           743 => x"c0",
           744 => x"71",
           745 => x"ff",
           746 => x"e0",
           747 => x"3d",
           748 => x"3d",
           749 => x"81",
           750 => x"70",
           751 => x"52",
           752 => x"94",
           753 => x"80",
           754 => x"87",
           755 => x"52",
           756 => x"82",
           757 => x"06",
           758 => x"ff",
           759 => x"2e",
           760 => x"81",
           761 => x"87",
           762 => x"52",
           763 => x"86",
           764 => x"94",
           765 => x"08",
           766 => x"70",
           767 => x"53",
           768 => x"ec",
           769 => x"3d",
           770 => x"3d",
           771 => x"9e",
           772 => x"9c",
           773 => x"51",
           774 => x"2e",
           775 => x"87",
           776 => x"08",
           777 => x"0c",
           778 => x"a8",
           779 => x"90",
           780 => x"9e",
           781 => x"e9",
           782 => x"c0",
           783 => x"81",
           784 => x"87",
           785 => x"08",
           786 => x"0c",
           787 => x"a0",
           788 => x"a0",
           789 => x"9e",
           790 => x"e9",
           791 => x"c0",
           792 => x"81",
           793 => x"87",
           794 => x"08",
           795 => x"0c",
           796 => x"b8",
           797 => x"b0",
           798 => x"9e",
           799 => x"e9",
           800 => x"c0",
           801 => x"81",
           802 => x"87",
           803 => x"08",
           804 => x"0c",
           805 => x"80",
           806 => x"81",
           807 => x"87",
           808 => x"08",
           809 => x"0c",
           810 => x"88",
           811 => x"c8",
           812 => x"9e",
           813 => x"e9",
           814 => x"0b",
           815 => x"34",
           816 => x"c0",
           817 => x"70",
           818 => x"06",
           819 => x"70",
           820 => x"38",
           821 => x"81",
           822 => x"80",
           823 => x"9e",
           824 => x"88",
           825 => x"51",
           826 => x"80",
           827 => x"81",
           828 => x"e9",
           829 => x"0b",
           830 => x"90",
           831 => x"80",
           832 => x"52",
           833 => x"2e",
           834 => x"52",
           835 => x"d3",
           836 => x"87",
           837 => x"08",
           838 => x"80",
           839 => x"52",
           840 => x"83",
           841 => x"71",
           842 => x"34",
           843 => x"c0",
           844 => x"70",
           845 => x"06",
           846 => x"70",
           847 => x"38",
           848 => x"81",
           849 => x"80",
           850 => x"9e",
           851 => x"90",
           852 => x"51",
           853 => x"80",
           854 => x"81",
           855 => x"e9",
           856 => x"0b",
           857 => x"90",
           858 => x"80",
           859 => x"52",
           860 => x"2e",
           861 => x"52",
           862 => x"d7",
           863 => x"87",
           864 => x"08",
           865 => x"80",
           866 => x"52",
           867 => x"83",
           868 => x"71",
           869 => x"34",
           870 => x"c0",
           871 => x"70",
           872 => x"06",
           873 => x"70",
           874 => x"38",
           875 => x"81",
           876 => x"80",
           877 => x"9e",
           878 => x"80",
           879 => x"51",
           880 => x"80",
           881 => x"81",
           882 => x"e9",
           883 => x"0b",
           884 => x"90",
           885 => x"80",
           886 => x"52",
           887 => x"83",
           888 => x"71",
           889 => x"34",
           890 => x"90",
           891 => x"80",
           892 => x"2a",
           893 => x"70",
           894 => x"34",
           895 => x"c0",
           896 => x"70",
           897 => x"51",
           898 => x"80",
           899 => x"81",
           900 => x"e9",
           901 => x"c0",
           902 => x"70",
           903 => x"70",
           904 => x"51",
           905 => x"e9",
           906 => x"0b",
           907 => x"90",
           908 => x"06",
           909 => x"70",
           910 => x"38",
           911 => x"81",
           912 => x"87",
           913 => x"08",
           914 => x"51",
           915 => x"e9",
           916 => x"3d",
           917 => x"3d",
           918 => x"f8",
           919 => x"3f",
           920 => x"33",
           921 => x"2e",
           922 => x"d6",
           923 => x"b6",
           924 => x"a0",
           925 => x"3f",
           926 => x"33",
           927 => x"2e",
           928 => x"e9",
           929 => x"e9",
           930 => x"54",
           931 => x"b8",
           932 => x"3f",
           933 => x"33",
           934 => x"2e",
           935 => x"e9",
           936 => x"e9",
           937 => x"54",
           938 => x"d4",
           939 => x"3f",
           940 => x"33",
           941 => x"2e",
           942 => x"e9",
           943 => x"e9",
           944 => x"54",
           945 => x"f0",
           946 => x"3f",
           947 => x"33",
           948 => x"2e",
           949 => x"e9",
           950 => x"e9",
           951 => x"54",
           952 => x"8c",
           953 => x"3f",
           954 => x"33",
           955 => x"2e",
           956 => x"e9",
           957 => x"e9",
           958 => x"54",
           959 => x"a8",
           960 => x"3f",
           961 => x"33",
           962 => x"2e",
           963 => x"e9",
           964 => x"81",
           965 => x"89",
           966 => x"e9",
           967 => x"73",
           968 => x"38",
           969 => x"33",
           970 => x"e4",
           971 => x"3f",
           972 => x"33",
           973 => x"2e",
           974 => x"e9",
           975 => x"81",
           976 => x"89",
           977 => x"e9",
           978 => x"73",
           979 => x"38",
           980 => x"51",
           981 => x"81",
           982 => x"54",
           983 => x"88",
           984 => x"b8",
           985 => x"3f",
           986 => x"33",
           987 => x"2e",
           988 => x"d8",
           989 => x"ae",
           990 => x"d9",
           991 => x"80",
           992 => x"81",
           993 => x"83",
           994 => x"e9",
           995 => x"73",
           996 => x"38",
           997 => x"51",
           998 => x"81",
           999 => x"83",
          1000 => x"e9",
          1001 => x"81",
          1002 => x"88",
          1003 => x"e9",
          1004 => x"81",
          1005 => x"88",
          1006 => x"e9",
          1007 => x"81",
          1008 => x"88",
          1009 => x"d9",
          1010 => x"da",
          1011 => x"c0",
          1012 => x"d9",
          1013 => x"b2",
          1014 => x"c4",
          1015 => x"84",
          1016 => x"51",
          1017 => x"81",
          1018 => x"bd",
          1019 => x"76",
          1020 => x"54",
          1021 => x"08",
          1022 => x"9c",
          1023 => x"3f",
          1024 => x"33",
          1025 => x"2e",
          1026 => x"e9",
          1027 => x"bd",
          1028 => x"75",
          1029 => x"3f",
          1030 => x"08",
          1031 => x"29",
          1032 => x"54",
          1033 => x"e0",
          1034 => x"da",
          1035 => x"da",
          1036 => x"d2",
          1037 => x"80",
          1038 => x"81",
          1039 => x"56",
          1040 => x"52",
          1041 => x"e4",
          1042 => x"e0",
          1043 => x"c0",
          1044 => x"31",
          1045 => x"ec",
          1046 => x"81",
          1047 => x"87",
          1048 => x"e6",
          1049 => x"be",
          1050 => x"0d",
          1051 => x"0d",
          1052 => x"33",
          1053 => x"71",
          1054 => x"38",
          1055 => x"0b",
          1056 => x"fc",
          1057 => x"08",
          1058 => x"a0",
          1059 => x"81",
          1060 => x"97",
          1061 => x"b0",
          1062 => x"81",
          1063 => x"8b",
          1064 => x"bc",
          1065 => x"81",
          1066 => x"80",
          1067 => x"3d",
          1068 => x"88",
          1069 => x"80",
          1070 => x"96",
          1071 => x"81",
          1072 => x"87",
          1073 => x"0c",
          1074 => x"0d",
          1075 => x"33",
          1076 => x"2e",
          1077 => x"85",
          1078 => x"ed",
          1079 => x"f8",
          1080 => x"80",
          1081 => x"72",
          1082 => x"ec",
          1083 => x"05",
          1084 => x"0c",
          1085 => x"ec",
          1086 => x"71",
          1087 => x"38",
          1088 => x"2d",
          1089 => x"04",
          1090 => x"02",
          1091 => x"81",
          1092 => x"76",
          1093 => x"0c",
          1094 => x"ad",
          1095 => x"ec",
          1096 => x"3d",
          1097 => x"3d",
          1098 => x"73",
          1099 => x"ff",
          1100 => x"71",
          1101 => x"38",
          1102 => x"06",
          1103 => x"54",
          1104 => x"e7",
          1105 => x"0d",
          1106 => x"0d",
          1107 => x"f0",
          1108 => x"ec",
          1109 => x"54",
          1110 => x"81",
          1111 => x"53",
          1112 => x"8e",
          1113 => x"ff",
          1114 => x"14",
          1115 => x"3f",
          1116 => x"81",
          1117 => x"86",
          1118 => x"ec",
          1119 => x"68",
          1120 => x"70",
          1121 => x"33",
          1122 => x"2e",
          1123 => x"75",
          1124 => x"81",
          1125 => x"38",
          1126 => x"70",
          1127 => x"33",
          1128 => x"75",
          1129 => x"81",
          1130 => x"81",
          1131 => x"75",
          1132 => x"81",
          1133 => x"82",
          1134 => x"81",
          1135 => x"56",
          1136 => x"09",
          1137 => x"38",
          1138 => x"71",
          1139 => x"81",
          1140 => x"59",
          1141 => x"9d",
          1142 => x"53",
          1143 => x"95",
          1144 => x"29",
          1145 => x"76",
          1146 => x"79",
          1147 => x"5b",
          1148 => x"e5",
          1149 => x"ec",
          1150 => x"70",
          1151 => x"25",
          1152 => x"32",
          1153 => x"72",
          1154 => x"73",
          1155 => x"58",
          1156 => x"73",
          1157 => x"38",
          1158 => x"79",
          1159 => x"5b",
          1160 => x"75",
          1161 => x"de",
          1162 => x"80",
          1163 => x"89",
          1164 => x"70",
          1165 => x"55",
          1166 => x"cf",
          1167 => x"38",
          1168 => x"24",
          1169 => x"80",
          1170 => x"8e",
          1171 => x"c3",
          1172 => x"73",
          1173 => x"81",
          1174 => x"99",
          1175 => x"c4",
          1176 => x"38",
          1177 => x"73",
          1178 => x"81",
          1179 => x"80",
          1180 => x"38",
          1181 => x"2e",
          1182 => x"f9",
          1183 => x"d8",
          1184 => x"38",
          1185 => x"77",
          1186 => x"08",
          1187 => x"80",
          1188 => x"55",
          1189 => x"8d",
          1190 => x"70",
          1191 => x"51",
          1192 => x"f5",
          1193 => x"2a",
          1194 => x"74",
          1195 => x"53",
          1196 => x"8f",
          1197 => x"fc",
          1198 => x"81",
          1199 => x"80",
          1200 => x"73",
          1201 => x"3f",
          1202 => x"56",
          1203 => x"27",
          1204 => x"a0",
          1205 => x"3f",
          1206 => x"84",
          1207 => x"33",
          1208 => x"93",
          1209 => x"95",
          1210 => x"91",
          1211 => x"8d",
          1212 => x"89",
          1213 => x"fb",
          1214 => x"86",
          1215 => x"2a",
          1216 => x"51",
          1217 => x"2e",
          1218 => x"84",
          1219 => x"86",
          1220 => x"78",
          1221 => x"08",
          1222 => x"32",
          1223 => x"72",
          1224 => x"51",
          1225 => x"74",
          1226 => x"38",
          1227 => x"88",
          1228 => x"7a",
          1229 => x"55",
          1230 => x"3d",
          1231 => x"52",
          1232 => x"9b",
          1233 => x"e0",
          1234 => x"06",
          1235 => x"52",
          1236 => x"3f",
          1237 => x"08",
          1238 => x"27",
          1239 => x"14",
          1240 => x"f8",
          1241 => x"87",
          1242 => x"81",
          1243 => x"b0",
          1244 => x"7d",
          1245 => x"5f",
          1246 => x"75",
          1247 => x"07",
          1248 => x"54",
          1249 => x"26",
          1250 => x"ff",
          1251 => x"84",
          1252 => x"06",
          1253 => x"80",
          1254 => x"96",
          1255 => x"e0",
          1256 => x"73",
          1257 => x"57",
          1258 => x"06",
          1259 => x"54",
          1260 => x"a0",
          1261 => x"2a",
          1262 => x"54",
          1263 => x"38",
          1264 => x"76",
          1265 => x"38",
          1266 => x"fd",
          1267 => x"06",
          1268 => x"38",
          1269 => x"56",
          1270 => x"26",
          1271 => x"3d",
          1272 => x"05",
          1273 => x"ff",
          1274 => x"53",
          1275 => x"d9",
          1276 => x"38",
          1277 => x"56",
          1278 => x"27",
          1279 => x"a0",
          1280 => x"3f",
          1281 => x"3d",
          1282 => x"3d",
          1283 => x"70",
          1284 => x"52",
          1285 => x"73",
          1286 => x"3f",
          1287 => x"04",
          1288 => x"74",
          1289 => x"0c",
          1290 => x"05",
          1291 => x"fa",
          1292 => x"ec",
          1293 => x"80",
          1294 => x"0b",
          1295 => x"0c",
          1296 => x"04",
          1297 => x"81",
          1298 => x"76",
          1299 => x"0c",
          1300 => x"05",
          1301 => x"53",
          1302 => x"72",
          1303 => x"0c",
          1304 => x"04",
          1305 => x"77",
          1306 => x"f4",
          1307 => x"54",
          1308 => x"54",
          1309 => x"80",
          1310 => x"ec",
          1311 => x"71",
          1312 => x"e0",
          1313 => x"06",
          1314 => x"2e",
          1315 => x"72",
          1316 => x"38",
          1317 => x"70",
          1318 => x"25",
          1319 => x"73",
          1320 => x"38",
          1321 => x"86",
          1322 => x"54",
          1323 => x"73",
          1324 => x"ff",
          1325 => x"72",
          1326 => x"74",
          1327 => x"72",
          1328 => x"54",
          1329 => x"81",
          1330 => x"39",
          1331 => x"80",
          1332 => x"51",
          1333 => x"81",
          1334 => x"ec",
          1335 => x"3d",
          1336 => x"3d",
          1337 => x"f4",
          1338 => x"ec",
          1339 => x"53",
          1340 => x"fe",
          1341 => x"81",
          1342 => x"84",
          1343 => x"f8",
          1344 => x"7c",
          1345 => x"70",
          1346 => x"75",
          1347 => x"55",
          1348 => x"2e",
          1349 => x"87",
          1350 => x"76",
          1351 => x"73",
          1352 => x"81",
          1353 => x"81",
          1354 => x"77",
          1355 => x"70",
          1356 => x"58",
          1357 => x"09",
          1358 => x"c2",
          1359 => x"81",
          1360 => x"75",
          1361 => x"55",
          1362 => x"e2",
          1363 => x"90",
          1364 => x"f8",
          1365 => x"8f",
          1366 => x"81",
          1367 => x"75",
          1368 => x"55",
          1369 => x"81",
          1370 => x"27",
          1371 => x"d0",
          1372 => x"55",
          1373 => x"73",
          1374 => x"80",
          1375 => x"14",
          1376 => x"72",
          1377 => x"e0",
          1378 => x"80",
          1379 => x"39",
          1380 => x"55",
          1381 => x"80",
          1382 => x"e0",
          1383 => x"38",
          1384 => x"81",
          1385 => x"53",
          1386 => x"81",
          1387 => x"53",
          1388 => x"8e",
          1389 => x"70",
          1390 => x"55",
          1391 => x"27",
          1392 => x"77",
          1393 => x"74",
          1394 => x"76",
          1395 => x"77",
          1396 => x"70",
          1397 => x"55",
          1398 => x"77",
          1399 => x"38",
          1400 => x"74",
          1401 => x"55",
          1402 => x"e0",
          1403 => x"0d",
          1404 => x"0d",
          1405 => x"56",
          1406 => x"0c",
          1407 => x"70",
          1408 => x"73",
          1409 => x"81",
          1410 => x"81",
          1411 => x"ed",
          1412 => x"2e",
          1413 => x"8e",
          1414 => x"08",
          1415 => x"76",
          1416 => x"56",
          1417 => x"b0",
          1418 => x"06",
          1419 => x"75",
          1420 => x"76",
          1421 => x"70",
          1422 => x"73",
          1423 => x"8b",
          1424 => x"73",
          1425 => x"85",
          1426 => x"82",
          1427 => x"76",
          1428 => x"70",
          1429 => x"ac",
          1430 => x"a0",
          1431 => x"fa",
          1432 => x"53",
          1433 => x"57",
          1434 => x"98",
          1435 => x"39",
          1436 => x"80",
          1437 => x"26",
          1438 => x"86",
          1439 => x"80",
          1440 => x"57",
          1441 => x"74",
          1442 => x"38",
          1443 => x"27",
          1444 => x"14",
          1445 => x"06",
          1446 => x"14",
          1447 => x"06",
          1448 => x"74",
          1449 => x"f9",
          1450 => x"ff",
          1451 => x"89",
          1452 => x"38",
          1453 => x"c5",
          1454 => x"29",
          1455 => x"81",
          1456 => x"76",
          1457 => x"56",
          1458 => x"ba",
          1459 => x"2e",
          1460 => x"30",
          1461 => x"0c",
          1462 => x"81",
          1463 => x"8a",
          1464 => x"ff",
          1465 => x"8f",
          1466 => x"81",
          1467 => x"26",
          1468 => x"e9",
          1469 => x"52",
          1470 => x"e0",
          1471 => x"0d",
          1472 => x"0d",
          1473 => x"33",
          1474 => x"9f",
          1475 => x"53",
          1476 => x"81",
          1477 => x"38",
          1478 => x"87",
          1479 => x"11",
          1480 => x"54",
          1481 => x"84",
          1482 => x"54",
          1483 => x"87",
          1484 => x"11",
          1485 => x"0c",
          1486 => x"c0",
          1487 => x"70",
          1488 => x"70",
          1489 => x"51",
          1490 => x"8a",
          1491 => x"98",
          1492 => x"70",
          1493 => x"08",
          1494 => x"06",
          1495 => x"38",
          1496 => x"8c",
          1497 => x"80",
          1498 => x"71",
          1499 => x"14",
          1500 => x"e8",
          1501 => x"70",
          1502 => x"0c",
          1503 => x"04",
          1504 => x"60",
          1505 => x"8c",
          1506 => x"33",
          1507 => x"5b",
          1508 => x"5a",
          1509 => x"81",
          1510 => x"81",
          1511 => x"52",
          1512 => x"38",
          1513 => x"84",
          1514 => x"92",
          1515 => x"c0",
          1516 => x"87",
          1517 => x"13",
          1518 => x"57",
          1519 => x"0b",
          1520 => x"8c",
          1521 => x"0c",
          1522 => x"75",
          1523 => x"2a",
          1524 => x"51",
          1525 => x"80",
          1526 => x"7b",
          1527 => x"7b",
          1528 => x"5d",
          1529 => x"59",
          1530 => x"06",
          1531 => x"73",
          1532 => x"81",
          1533 => x"ff",
          1534 => x"72",
          1535 => x"38",
          1536 => x"8c",
          1537 => x"c3",
          1538 => x"98",
          1539 => x"71",
          1540 => x"38",
          1541 => x"2e",
          1542 => x"76",
          1543 => x"92",
          1544 => x"72",
          1545 => x"06",
          1546 => x"f7",
          1547 => x"5a",
          1548 => x"80",
          1549 => x"70",
          1550 => x"5a",
          1551 => x"80",
          1552 => x"73",
          1553 => x"06",
          1554 => x"38",
          1555 => x"fe",
          1556 => x"fc",
          1557 => x"52",
          1558 => x"83",
          1559 => x"71",
          1560 => x"ec",
          1561 => x"3d",
          1562 => x"3d",
          1563 => x"64",
          1564 => x"bf",
          1565 => x"40",
          1566 => x"59",
          1567 => x"58",
          1568 => x"81",
          1569 => x"81",
          1570 => x"52",
          1571 => x"09",
          1572 => x"b1",
          1573 => x"84",
          1574 => x"92",
          1575 => x"c0",
          1576 => x"87",
          1577 => x"13",
          1578 => x"56",
          1579 => x"87",
          1580 => x"0c",
          1581 => x"82",
          1582 => x"58",
          1583 => x"84",
          1584 => x"06",
          1585 => x"71",
          1586 => x"38",
          1587 => x"05",
          1588 => x"0c",
          1589 => x"73",
          1590 => x"81",
          1591 => x"71",
          1592 => x"38",
          1593 => x"8c",
          1594 => x"d0",
          1595 => x"98",
          1596 => x"71",
          1597 => x"38",
          1598 => x"2e",
          1599 => x"76",
          1600 => x"92",
          1601 => x"72",
          1602 => x"06",
          1603 => x"f7",
          1604 => x"59",
          1605 => x"1a",
          1606 => x"06",
          1607 => x"59",
          1608 => x"80",
          1609 => x"73",
          1610 => x"06",
          1611 => x"38",
          1612 => x"fe",
          1613 => x"fc",
          1614 => x"52",
          1615 => x"83",
          1616 => x"71",
          1617 => x"ec",
          1618 => x"3d",
          1619 => x"3d",
          1620 => x"84",
          1621 => x"33",
          1622 => x"a7",
          1623 => x"54",
          1624 => x"fa",
          1625 => x"ec",
          1626 => x"06",
          1627 => x"72",
          1628 => x"85",
          1629 => x"98",
          1630 => x"56",
          1631 => x"80",
          1632 => x"76",
          1633 => x"74",
          1634 => x"c0",
          1635 => x"54",
          1636 => x"2e",
          1637 => x"d4",
          1638 => x"2e",
          1639 => x"80",
          1640 => x"08",
          1641 => x"70",
          1642 => x"51",
          1643 => x"2e",
          1644 => x"c0",
          1645 => x"52",
          1646 => x"87",
          1647 => x"08",
          1648 => x"38",
          1649 => x"87",
          1650 => x"14",
          1651 => x"70",
          1652 => x"52",
          1653 => x"96",
          1654 => x"92",
          1655 => x"0a",
          1656 => x"39",
          1657 => x"0c",
          1658 => x"39",
          1659 => x"54",
          1660 => x"e0",
          1661 => x"0d",
          1662 => x"0d",
          1663 => x"33",
          1664 => x"88",
          1665 => x"ec",
          1666 => x"51",
          1667 => x"04",
          1668 => x"75",
          1669 => x"82",
          1670 => x"90",
          1671 => x"2b",
          1672 => x"33",
          1673 => x"88",
          1674 => x"71",
          1675 => x"e0",
          1676 => x"54",
          1677 => x"85",
          1678 => x"ff",
          1679 => x"02",
          1680 => x"05",
          1681 => x"70",
          1682 => x"05",
          1683 => x"88",
          1684 => x"72",
          1685 => x"0d",
          1686 => x"0d",
          1687 => x"52",
          1688 => x"81",
          1689 => x"70",
          1690 => x"70",
          1691 => x"05",
          1692 => x"88",
          1693 => x"72",
          1694 => x"54",
          1695 => x"2a",
          1696 => x"34",
          1697 => x"04",
          1698 => x"76",
          1699 => x"54",
          1700 => x"2e",
          1701 => x"70",
          1702 => x"33",
          1703 => x"05",
          1704 => x"11",
          1705 => x"84",
          1706 => x"fe",
          1707 => x"77",
          1708 => x"53",
          1709 => x"81",
          1710 => x"ff",
          1711 => x"f4",
          1712 => x"0d",
          1713 => x"0d",
          1714 => x"56",
          1715 => x"70",
          1716 => x"33",
          1717 => x"05",
          1718 => x"71",
          1719 => x"56",
          1720 => x"72",
          1721 => x"38",
          1722 => x"e2",
          1723 => x"ec",
          1724 => x"3d",
          1725 => x"3d",
          1726 => x"54",
          1727 => x"71",
          1728 => x"38",
          1729 => x"70",
          1730 => x"f3",
          1731 => x"81",
          1732 => x"84",
          1733 => x"80",
          1734 => x"e0",
          1735 => x"0b",
          1736 => x"0c",
          1737 => x"0d",
          1738 => x"0b",
          1739 => x"56",
          1740 => x"2e",
          1741 => x"81",
          1742 => x"08",
          1743 => x"70",
          1744 => x"33",
          1745 => x"a2",
          1746 => x"e0",
          1747 => x"09",
          1748 => x"38",
          1749 => x"08",
          1750 => x"b0",
          1751 => x"a4",
          1752 => x"9c",
          1753 => x"56",
          1754 => x"27",
          1755 => x"16",
          1756 => x"82",
          1757 => x"06",
          1758 => x"54",
          1759 => x"78",
          1760 => x"33",
          1761 => x"3f",
          1762 => x"5a",
          1763 => x"e0",
          1764 => x"0d",
          1765 => x"0d",
          1766 => x"56",
          1767 => x"b0",
          1768 => x"af",
          1769 => x"fe",
          1770 => x"ec",
          1771 => x"81",
          1772 => x"9f",
          1773 => x"74",
          1774 => x"52",
          1775 => x"51",
          1776 => x"81",
          1777 => x"80",
          1778 => x"ff",
          1779 => x"74",
          1780 => x"76",
          1781 => x"0c",
          1782 => x"04",
          1783 => x"7a",
          1784 => x"fe",
          1785 => x"ec",
          1786 => x"81",
          1787 => x"81",
          1788 => x"33",
          1789 => x"2e",
          1790 => x"80",
          1791 => x"17",
          1792 => x"81",
          1793 => x"06",
          1794 => x"84",
          1795 => x"ec",
          1796 => x"b4",
          1797 => x"56",
          1798 => x"82",
          1799 => x"84",
          1800 => x"fc",
          1801 => x"8b",
          1802 => x"52",
          1803 => x"a9",
          1804 => x"85",
          1805 => x"84",
          1806 => x"fc",
          1807 => x"17",
          1808 => x"9c",
          1809 => x"91",
          1810 => x"08",
          1811 => x"17",
          1812 => x"3f",
          1813 => x"81",
          1814 => x"19",
          1815 => x"53",
          1816 => x"17",
          1817 => x"82",
          1818 => x"18",
          1819 => x"80",
          1820 => x"33",
          1821 => x"3f",
          1822 => x"08",
          1823 => x"38",
          1824 => x"81",
          1825 => x"8a",
          1826 => x"fb",
          1827 => x"fe",
          1828 => x"08",
          1829 => x"56",
          1830 => x"74",
          1831 => x"38",
          1832 => x"75",
          1833 => x"16",
          1834 => x"53",
          1835 => x"e0",
          1836 => x"0d",
          1837 => x"0d",
          1838 => x"08",
          1839 => x"81",
          1840 => x"df",
          1841 => x"15",
          1842 => x"d7",
          1843 => x"33",
          1844 => x"82",
          1845 => x"38",
          1846 => x"89",
          1847 => x"2e",
          1848 => x"bf",
          1849 => x"2e",
          1850 => x"81",
          1851 => x"81",
          1852 => x"89",
          1853 => x"08",
          1854 => x"52",
          1855 => x"3f",
          1856 => x"08",
          1857 => x"74",
          1858 => x"14",
          1859 => x"81",
          1860 => x"2a",
          1861 => x"05",
          1862 => x"57",
          1863 => x"f5",
          1864 => x"e0",
          1865 => x"38",
          1866 => x"06",
          1867 => x"33",
          1868 => x"78",
          1869 => x"06",
          1870 => x"5c",
          1871 => x"53",
          1872 => x"38",
          1873 => x"06",
          1874 => x"39",
          1875 => x"a4",
          1876 => x"52",
          1877 => x"bd",
          1878 => x"e0",
          1879 => x"38",
          1880 => x"fe",
          1881 => x"b4",
          1882 => x"8d",
          1883 => x"e0",
          1884 => x"ff",
          1885 => x"39",
          1886 => x"a4",
          1887 => x"52",
          1888 => x"91",
          1889 => x"e0",
          1890 => x"76",
          1891 => x"fc",
          1892 => x"b4",
          1893 => x"f8",
          1894 => x"e0",
          1895 => x"06",
          1896 => x"81",
          1897 => x"ec",
          1898 => x"3d",
          1899 => x"3d",
          1900 => x"7e",
          1901 => x"82",
          1902 => x"27",
          1903 => x"76",
          1904 => x"27",
          1905 => x"75",
          1906 => x"79",
          1907 => x"38",
          1908 => x"89",
          1909 => x"2e",
          1910 => x"80",
          1911 => x"2e",
          1912 => x"81",
          1913 => x"81",
          1914 => x"89",
          1915 => x"08",
          1916 => x"52",
          1917 => x"3f",
          1918 => x"08",
          1919 => x"e0",
          1920 => x"38",
          1921 => x"06",
          1922 => x"81",
          1923 => x"06",
          1924 => x"77",
          1925 => x"2e",
          1926 => x"84",
          1927 => x"06",
          1928 => x"06",
          1929 => x"53",
          1930 => x"81",
          1931 => x"34",
          1932 => x"a4",
          1933 => x"52",
          1934 => x"d9",
          1935 => x"e0",
          1936 => x"ec",
          1937 => x"94",
          1938 => x"ff",
          1939 => x"05",
          1940 => x"54",
          1941 => x"38",
          1942 => x"74",
          1943 => x"06",
          1944 => x"07",
          1945 => x"74",
          1946 => x"39",
          1947 => x"a4",
          1948 => x"52",
          1949 => x"9d",
          1950 => x"e0",
          1951 => x"ec",
          1952 => x"d8",
          1953 => x"ff",
          1954 => x"76",
          1955 => x"06",
          1956 => x"05",
          1957 => x"3f",
          1958 => x"87",
          1959 => x"08",
          1960 => x"51",
          1961 => x"81",
          1962 => x"59",
          1963 => x"08",
          1964 => x"f0",
          1965 => x"82",
          1966 => x"06",
          1967 => x"05",
          1968 => x"54",
          1969 => x"3f",
          1970 => x"08",
          1971 => x"74",
          1972 => x"51",
          1973 => x"81",
          1974 => x"34",
          1975 => x"e0",
          1976 => x"0d",
          1977 => x"0d",
          1978 => x"72",
          1979 => x"56",
          1980 => x"27",
          1981 => x"98",
          1982 => x"9d",
          1983 => x"2e",
          1984 => x"53",
          1985 => x"51",
          1986 => x"81",
          1987 => x"54",
          1988 => x"08",
          1989 => x"93",
          1990 => x"80",
          1991 => x"54",
          1992 => x"81",
          1993 => x"54",
          1994 => x"74",
          1995 => x"fb",
          1996 => x"ec",
          1997 => x"81",
          1998 => x"80",
          1999 => x"38",
          2000 => x"08",
          2001 => x"38",
          2002 => x"08",
          2003 => x"38",
          2004 => x"52",
          2005 => x"d6",
          2006 => x"e0",
          2007 => x"98",
          2008 => x"11",
          2009 => x"57",
          2010 => x"74",
          2011 => x"81",
          2012 => x"0c",
          2013 => x"81",
          2014 => x"84",
          2015 => x"55",
          2016 => x"ff",
          2017 => x"54",
          2018 => x"e0",
          2019 => x"0d",
          2020 => x"0d",
          2021 => x"08",
          2022 => x"79",
          2023 => x"17",
          2024 => x"80",
          2025 => x"98",
          2026 => x"26",
          2027 => x"58",
          2028 => x"52",
          2029 => x"fd",
          2030 => x"74",
          2031 => x"08",
          2032 => x"38",
          2033 => x"08",
          2034 => x"e0",
          2035 => x"82",
          2036 => x"17",
          2037 => x"e0",
          2038 => x"c7",
          2039 => x"90",
          2040 => x"56",
          2041 => x"2e",
          2042 => x"77",
          2043 => x"81",
          2044 => x"38",
          2045 => x"98",
          2046 => x"26",
          2047 => x"56",
          2048 => x"51",
          2049 => x"80",
          2050 => x"e0",
          2051 => x"09",
          2052 => x"38",
          2053 => x"08",
          2054 => x"e0",
          2055 => x"30",
          2056 => x"80",
          2057 => x"07",
          2058 => x"08",
          2059 => x"55",
          2060 => x"ef",
          2061 => x"e0",
          2062 => x"95",
          2063 => x"08",
          2064 => x"27",
          2065 => x"98",
          2066 => x"89",
          2067 => x"85",
          2068 => x"db",
          2069 => x"81",
          2070 => x"17",
          2071 => x"89",
          2072 => x"75",
          2073 => x"ac",
          2074 => x"7a",
          2075 => x"3f",
          2076 => x"08",
          2077 => x"38",
          2078 => x"ec",
          2079 => x"2e",
          2080 => x"86",
          2081 => x"e0",
          2082 => x"ec",
          2083 => x"70",
          2084 => x"07",
          2085 => x"7c",
          2086 => x"55",
          2087 => x"f8",
          2088 => x"2e",
          2089 => x"ff",
          2090 => x"55",
          2091 => x"ff",
          2092 => x"76",
          2093 => x"3f",
          2094 => x"08",
          2095 => x"08",
          2096 => x"ec",
          2097 => x"80",
          2098 => x"55",
          2099 => x"94",
          2100 => x"2e",
          2101 => x"53",
          2102 => x"51",
          2103 => x"81",
          2104 => x"55",
          2105 => x"75",
          2106 => x"98",
          2107 => x"05",
          2108 => x"56",
          2109 => x"26",
          2110 => x"15",
          2111 => x"84",
          2112 => x"07",
          2113 => x"18",
          2114 => x"ff",
          2115 => x"2e",
          2116 => x"39",
          2117 => x"39",
          2118 => x"08",
          2119 => x"81",
          2120 => x"74",
          2121 => x"0c",
          2122 => x"04",
          2123 => x"7a",
          2124 => x"f3",
          2125 => x"ec",
          2126 => x"81",
          2127 => x"e0",
          2128 => x"38",
          2129 => x"51",
          2130 => x"81",
          2131 => x"81",
          2132 => x"b0",
          2133 => x"84",
          2134 => x"52",
          2135 => x"52",
          2136 => x"3f",
          2137 => x"39",
          2138 => x"8a",
          2139 => x"75",
          2140 => x"38",
          2141 => x"19",
          2142 => x"81",
          2143 => x"ed",
          2144 => x"ec",
          2145 => x"2e",
          2146 => x"15",
          2147 => x"70",
          2148 => x"07",
          2149 => x"53",
          2150 => x"75",
          2151 => x"0c",
          2152 => x"04",
          2153 => x"7a",
          2154 => x"58",
          2155 => x"f0",
          2156 => x"80",
          2157 => x"9f",
          2158 => x"80",
          2159 => x"90",
          2160 => x"17",
          2161 => x"aa",
          2162 => x"53",
          2163 => x"88",
          2164 => x"08",
          2165 => x"38",
          2166 => x"53",
          2167 => x"17",
          2168 => x"72",
          2169 => x"fe",
          2170 => x"08",
          2171 => x"80",
          2172 => x"16",
          2173 => x"2b",
          2174 => x"75",
          2175 => x"73",
          2176 => x"f5",
          2177 => x"ec",
          2178 => x"81",
          2179 => x"ff",
          2180 => x"81",
          2181 => x"e0",
          2182 => x"38",
          2183 => x"81",
          2184 => x"26",
          2185 => x"58",
          2186 => x"73",
          2187 => x"39",
          2188 => x"51",
          2189 => x"81",
          2190 => x"98",
          2191 => x"94",
          2192 => x"17",
          2193 => x"58",
          2194 => x"9a",
          2195 => x"81",
          2196 => x"74",
          2197 => x"98",
          2198 => x"83",
          2199 => x"b4",
          2200 => x"0c",
          2201 => x"81",
          2202 => x"8a",
          2203 => x"f8",
          2204 => x"70",
          2205 => x"08",
          2206 => x"57",
          2207 => x"0a",
          2208 => x"38",
          2209 => x"15",
          2210 => x"08",
          2211 => x"72",
          2212 => x"cb",
          2213 => x"ff",
          2214 => x"81",
          2215 => x"13",
          2216 => x"94",
          2217 => x"74",
          2218 => x"85",
          2219 => x"22",
          2220 => x"73",
          2221 => x"38",
          2222 => x"8a",
          2223 => x"05",
          2224 => x"06",
          2225 => x"8a",
          2226 => x"73",
          2227 => x"3f",
          2228 => x"08",
          2229 => x"81",
          2230 => x"e0",
          2231 => x"ff",
          2232 => x"81",
          2233 => x"ff",
          2234 => x"38",
          2235 => x"81",
          2236 => x"26",
          2237 => x"7b",
          2238 => x"98",
          2239 => x"55",
          2240 => x"94",
          2241 => x"73",
          2242 => x"3f",
          2243 => x"08",
          2244 => x"81",
          2245 => x"80",
          2246 => x"38",
          2247 => x"ec",
          2248 => x"2e",
          2249 => x"55",
          2250 => x"08",
          2251 => x"38",
          2252 => x"08",
          2253 => x"fb",
          2254 => x"ec",
          2255 => x"38",
          2256 => x"0c",
          2257 => x"51",
          2258 => x"81",
          2259 => x"98",
          2260 => x"90",
          2261 => x"16",
          2262 => x"15",
          2263 => x"74",
          2264 => x"0c",
          2265 => x"04",
          2266 => x"7b",
          2267 => x"5b",
          2268 => x"52",
          2269 => x"ac",
          2270 => x"e0",
          2271 => x"ec",
          2272 => x"ec",
          2273 => x"e0",
          2274 => x"17",
          2275 => x"51",
          2276 => x"81",
          2277 => x"54",
          2278 => x"08",
          2279 => x"81",
          2280 => x"9c",
          2281 => x"33",
          2282 => x"72",
          2283 => x"09",
          2284 => x"38",
          2285 => x"ec",
          2286 => x"72",
          2287 => x"55",
          2288 => x"53",
          2289 => x"8e",
          2290 => x"56",
          2291 => x"09",
          2292 => x"38",
          2293 => x"ec",
          2294 => x"81",
          2295 => x"fd",
          2296 => x"ec",
          2297 => x"81",
          2298 => x"80",
          2299 => x"38",
          2300 => x"09",
          2301 => x"38",
          2302 => x"81",
          2303 => x"8b",
          2304 => x"fd",
          2305 => x"9a",
          2306 => x"eb",
          2307 => x"ec",
          2308 => x"ff",
          2309 => x"70",
          2310 => x"53",
          2311 => x"09",
          2312 => x"38",
          2313 => x"eb",
          2314 => x"ec",
          2315 => x"2b",
          2316 => x"72",
          2317 => x"0c",
          2318 => x"04",
          2319 => x"77",
          2320 => x"ff",
          2321 => x"9a",
          2322 => x"55",
          2323 => x"76",
          2324 => x"53",
          2325 => x"09",
          2326 => x"38",
          2327 => x"52",
          2328 => x"eb",
          2329 => x"3d",
          2330 => x"3d",
          2331 => x"5b",
          2332 => x"08",
          2333 => x"15",
          2334 => x"81",
          2335 => x"15",
          2336 => x"51",
          2337 => x"81",
          2338 => x"58",
          2339 => x"08",
          2340 => x"9c",
          2341 => x"33",
          2342 => x"86",
          2343 => x"80",
          2344 => x"13",
          2345 => x"06",
          2346 => x"06",
          2347 => x"72",
          2348 => x"81",
          2349 => x"53",
          2350 => x"2e",
          2351 => x"53",
          2352 => x"a9",
          2353 => x"74",
          2354 => x"72",
          2355 => x"38",
          2356 => x"99",
          2357 => x"e0",
          2358 => x"06",
          2359 => x"88",
          2360 => x"06",
          2361 => x"54",
          2362 => x"a0",
          2363 => x"74",
          2364 => x"3f",
          2365 => x"08",
          2366 => x"e0",
          2367 => x"98",
          2368 => x"fa",
          2369 => x"80",
          2370 => x"0c",
          2371 => x"e0",
          2372 => x"0d",
          2373 => x"0d",
          2374 => x"57",
          2375 => x"73",
          2376 => x"3f",
          2377 => x"08",
          2378 => x"e0",
          2379 => x"98",
          2380 => x"75",
          2381 => x"3f",
          2382 => x"08",
          2383 => x"e0",
          2384 => x"a0",
          2385 => x"e0",
          2386 => x"14",
          2387 => x"db",
          2388 => x"a0",
          2389 => x"14",
          2390 => x"ac",
          2391 => x"83",
          2392 => x"81",
          2393 => x"87",
          2394 => x"fd",
          2395 => x"70",
          2396 => x"08",
          2397 => x"55",
          2398 => x"3f",
          2399 => x"08",
          2400 => x"13",
          2401 => x"73",
          2402 => x"83",
          2403 => x"3d",
          2404 => x"3d",
          2405 => x"57",
          2406 => x"89",
          2407 => x"17",
          2408 => x"81",
          2409 => x"70",
          2410 => x"55",
          2411 => x"08",
          2412 => x"81",
          2413 => x"52",
          2414 => x"a8",
          2415 => x"2e",
          2416 => x"84",
          2417 => x"52",
          2418 => x"09",
          2419 => x"38",
          2420 => x"81",
          2421 => x"81",
          2422 => x"73",
          2423 => x"55",
          2424 => x"55",
          2425 => x"c5",
          2426 => x"88",
          2427 => x"0b",
          2428 => x"9c",
          2429 => x"8b",
          2430 => x"17",
          2431 => x"08",
          2432 => x"52",
          2433 => x"81",
          2434 => x"76",
          2435 => x"51",
          2436 => x"81",
          2437 => x"86",
          2438 => x"12",
          2439 => x"3f",
          2440 => x"08",
          2441 => x"88",
          2442 => x"f3",
          2443 => x"70",
          2444 => x"80",
          2445 => x"51",
          2446 => x"af",
          2447 => x"81",
          2448 => x"dc",
          2449 => x"74",
          2450 => x"38",
          2451 => x"88",
          2452 => x"39",
          2453 => x"80",
          2454 => x"56",
          2455 => x"af",
          2456 => x"06",
          2457 => x"56",
          2458 => x"32",
          2459 => x"80",
          2460 => x"51",
          2461 => x"dc",
          2462 => x"1c",
          2463 => x"33",
          2464 => x"9f",
          2465 => x"ff",
          2466 => x"1c",
          2467 => x"7a",
          2468 => x"3f",
          2469 => x"08",
          2470 => x"39",
          2471 => x"a0",
          2472 => x"5e",
          2473 => x"52",
          2474 => x"ff",
          2475 => x"59",
          2476 => x"33",
          2477 => x"ae",
          2478 => x"06",
          2479 => x"78",
          2480 => x"81",
          2481 => x"32",
          2482 => x"9f",
          2483 => x"26",
          2484 => x"53",
          2485 => x"73",
          2486 => x"17",
          2487 => x"34",
          2488 => x"db",
          2489 => x"32",
          2490 => x"9f",
          2491 => x"54",
          2492 => x"2e",
          2493 => x"80",
          2494 => x"75",
          2495 => x"bd",
          2496 => x"7e",
          2497 => x"a0",
          2498 => x"bd",
          2499 => x"82",
          2500 => x"18",
          2501 => x"1a",
          2502 => x"a0",
          2503 => x"fc",
          2504 => x"32",
          2505 => x"80",
          2506 => x"30",
          2507 => x"71",
          2508 => x"51",
          2509 => x"55",
          2510 => x"ac",
          2511 => x"81",
          2512 => x"78",
          2513 => x"51",
          2514 => x"af",
          2515 => x"06",
          2516 => x"55",
          2517 => x"32",
          2518 => x"80",
          2519 => x"51",
          2520 => x"db",
          2521 => x"39",
          2522 => x"09",
          2523 => x"38",
          2524 => x"7c",
          2525 => x"54",
          2526 => x"a2",
          2527 => x"32",
          2528 => x"ae",
          2529 => x"72",
          2530 => x"9f",
          2531 => x"51",
          2532 => x"74",
          2533 => x"88",
          2534 => x"fe",
          2535 => x"98",
          2536 => x"80",
          2537 => x"75",
          2538 => x"81",
          2539 => x"33",
          2540 => x"51",
          2541 => x"81",
          2542 => x"80",
          2543 => x"78",
          2544 => x"81",
          2545 => x"5a",
          2546 => x"d2",
          2547 => x"e0",
          2548 => x"80",
          2549 => x"1c",
          2550 => x"27",
          2551 => x"79",
          2552 => x"74",
          2553 => x"7a",
          2554 => x"74",
          2555 => x"39",
          2556 => x"db",
          2557 => x"fe",
          2558 => x"e0",
          2559 => x"ff",
          2560 => x"73",
          2561 => x"38",
          2562 => x"81",
          2563 => x"54",
          2564 => x"75",
          2565 => x"17",
          2566 => x"39",
          2567 => x"0c",
          2568 => x"99",
          2569 => x"54",
          2570 => x"2e",
          2571 => x"84",
          2572 => x"34",
          2573 => x"76",
          2574 => x"8b",
          2575 => x"81",
          2576 => x"56",
          2577 => x"80",
          2578 => x"1b",
          2579 => x"08",
          2580 => x"51",
          2581 => x"81",
          2582 => x"56",
          2583 => x"08",
          2584 => x"98",
          2585 => x"76",
          2586 => x"3f",
          2587 => x"08",
          2588 => x"e0",
          2589 => x"38",
          2590 => x"70",
          2591 => x"73",
          2592 => x"be",
          2593 => x"33",
          2594 => x"73",
          2595 => x"8b",
          2596 => x"83",
          2597 => x"06",
          2598 => x"73",
          2599 => x"53",
          2600 => x"51",
          2601 => x"81",
          2602 => x"80",
          2603 => x"75",
          2604 => x"f3",
          2605 => x"9f",
          2606 => x"1c",
          2607 => x"74",
          2608 => x"38",
          2609 => x"09",
          2610 => x"e7",
          2611 => x"2a",
          2612 => x"77",
          2613 => x"51",
          2614 => x"2e",
          2615 => x"81",
          2616 => x"80",
          2617 => x"38",
          2618 => x"ab",
          2619 => x"55",
          2620 => x"75",
          2621 => x"73",
          2622 => x"55",
          2623 => x"82",
          2624 => x"06",
          2625 => x"ab",
          2626 => x"33",
          2627 => x"70",
          2628 => x"55",
          2629 => x"2e",
          2630 => x"1b",
          2631 => x"06",
          2632 => x"52",
          2633 => x"db",
          2634 => x"e0",
          2635 => x"0c",
          2636 => x"74",
          2637 => x"0c",
          2638 => x"04",
          2639 => x"7c",
          2640 => x"08",
          2641 => x"55",
          2642 => x"59",
          2643 => x"81",
          2644 => x"70",
          2645 => x"33",
          2646 => x"52",
          2647 => x"2e",
          2648 => x"ee",
          2649 => x"2e",
          2650 => x"81",
          2651 => x"33",
          2652 => x"81",
          2653 => x"52",
          2654 => x"26",
          2655 => x"14",
          2656 => x"06",
          2657 => x"52",
          2658 => x"80",
          2659 => x"0b",
          2660 => x"59",
          2661 => x"7a",
          2662 => x"70",
          2663 => x"33",
          2664 => x"05",
          2665 => x"9f",
          2666 => x"53",
          2667 => x"89",
          2668 => x"70",
          2669 => x"54",
          2670 => x"12",
          2671 => x"26",
          2672 => x"12",
          2673 => x"06",
          2674 => x"30",
          2675 => x"51",
          2676 => x"2e",
          2677 => x"85",
          2678 => x"be",
          2679 => x"74",
          2680 => x"30",
          2681 => x"9f",
          2682 => x"2a",
          2683 => x"54",
          2684 => x"2e",
          2685 => x"15",
          2686 => x"55",
          2687 => x"ff",
          2688 => x"39",
          2689 => x"86",
          2690 => x"7c",
          2691 => x"51",
          2692 => x"ed",
          2693 => x"70",
          2694 => x"0c",
          2695 => x"04",
          2696 => x"78",
          2697 => x"83",
          2698 => x"0b",
          2699 => x"79",
          2700 => x"e2",
          2701 => x"55",
          2702 => x"08",
          2703 => x"84",
          2704 => x"df",
          2705 => x"ec",
          2706 => x"ff",
          2707 => x"83",
          2708 => x"d4",
          2709 => x"81",
          2710 => x"38",
          2711 => x"17",
          2712 => x"74",
          2713 => x"09",
          2714 => x"38",
          2715 => x"81",
          2716 => x"30",
          2717 => x"79",
          2718 => x"54",
          2719 => x"74",
          2720 => x"09",
          2721 => x"38",
          2722 => x"db",
          2723 => x"ea",
          2724 => x"b1",
          2725 => x"e0",
          2726 => x"ec",
          2727 => x"2e",
          2728 => x"53",
          2729 => x"52",
          2730 => x"51",
          2731 => x"81",
          2732 => x"55",
          2733 => x"08",
          2734 => x"38",
          2735 => x"81",
          2736 => x"88",
          2737 => x"f2",
          2738 => x"02",
          2739 => x"cb",
          2740 => x"55",
          2741 => x"60",
          2742 => x"3f",
          2743 => x"08",
          2744 => x"80",
          2745 => x"e0",
          2746 => x"fc",
          2747 => x"e0",
          2748 => x"81",
          2749 => x"70",
          2750 => x"8c",
          2751 => x"2e",
          2752 => x"73",
          2753 => x"81",
          2754 => x"33",
          2755 => x"80",
          2756 => x"81",
          2757 => x"d7",
          2758 => x"ec",
          2759 => x"ff",
          2760 => x"06",
          2761 => x"98",
          2762 => x"2e",
          2763 => x"74",
          2764 => x"81",
          2765 => x"8a",
          2766 => x"ac",
          2767 => x"39",
          2768 => x"77",
          2769 => x"81",
          2770 => x"33",
          2771 => x"3f",
          2772 => x"08",
          2773 => x"70",
          2774 => x"55",
          2775 => x"86",
          2776 => x"80",
          2777 => x"74",
          2778 => x"81",
          2779 => x"8a",
          2780 => x"f4",
          2781 => x"53",
          2782 => x"fd",
          2783 => x"ec",
          2784 => x"ff",
          2785 => x"82",
          2786 => x"06",
          2787 => x"8c",
          2788 => x"58",
          2789 => x"f6",
          2790 => x"58",
          2791 => x"2e",
          2792 => x"fa",
          2793 => x"e8",
          2794 => x"e0",
          2795 => x"78",
          2796 => x"5a",
          2797 => x"90",
          2798 => x"75",
          2799 => x"38",
          2800 => x"3d",
          2801 => x"70",
          2802 => x"08",
          2803 => x"7a",
          2804 => x"38",
          2805 => x"51",
          2806 => x"81",
          2807 => x"81",
          2808 => x"81",
          2809 => x"38",
          2810 => x"83",
          2811 => x"38",
          2812 => x"84",
          2813 => x"38",
          2814 => x"81",
          2815 => x"38",
          2816 => x"db",
          2817 => x"ec",
          2818 => x"ff",
          2819 => x"72",
          2820 => x"09",
          2821 => x"d0",
          2822 => x"14",
          2823 => x"3f",
          2824 => x"08",
          2825 => x"06",
          2826 => x"38",
          2827 => x"51",
          2828 => x"81",
          2829 => x"58",
          2830 => x"0c",
          2831 => x"33",
          2832 => x"80",
          2833 => x"ff",
          2834 => x"ff",
          2835 => x"55",
          2836 => x"81",
          2837 => x"38",
          2838 => x"06",
          2839 => x"80",
          2840 => x"52",
          2841 => x"8a",
          2842 => x"80",
          2843 => x"ff",
          2844 => x"53",
          2845 => x"86",
          2846 => x"83",
          2847 => x"c5",
          2848 => x"f5",
          2849 => x"e0",
          2850 => x"ec",
          2851 => x"15",
          2852 => x"06",
          2853 => x"76",
          2854 => x"80",
          2855 => x"da",
          2856 => x"ec",
          2857 => x"ff",
          2858 => x"74",
          2859 => x"d4",
          2860 => x"dc",
          2861 => x"e0",
          2862 => x"c2",
          2863 => x"b9",
          2864 => x"e0",
          2865 => x"ff",
          2866 => x"56",
          2867 => x"83",
          2868 => x"14",
          2869 => x"71",
          2870 => x"5a",
          2871 => x"26",
          2872 => x"8a",
          2873 => x"74",
          2874 => x"ff",
          2875 => x"81",
          2876 => x"55",
          2877 => x"08",
          2878 => x"ec",
          2879 => x"e0",
          2880 => x"ff",
          2881 => x"83",
          2882 => x"74",
          2883 => x"26",
          2884 => x"57",
          2885 => x"26",
          2886 => x"57",
          2887 => x"56",
          2888 => x"82",
          2889 => x"15",
          2890 => x"0c",
          2891 => x"0c",
          2892 => x"a4",
          2893 => x"1d",
          2894 => x"54",
          2895 => x"2e",
          2896 => x"af",
          2897 => x"14",
          2898 => x"3f",
          2899 => x"08",
          2900 => x"06",
          2901 => x"72",
          2902 => x"79",
          2903 => x"80",
          2904 => x"d9",
          2905 => x"ec",
          2906 => x"15",
          2907 => x"2b",
          2908 => x"8d",
          2909 => x"2e",
          2910 => x"77",
          2911 => x"0c",
          2912 => x"76",
          2913 => x"38",
          2914 => x"70",
          2915 => x"81",
          2916 => x"53",
          2917 => x"89",
          2918 => x"56",
          2919 => x"08",
          2920 => x"38",
          2921 => x"15",
          2922 => x"8c",
          2923 => x"80",
          2924 => x"34",
          2925 => x"09",
          2926 => x"92",
          2927 => x"14",
          2928 => x"3f",
          2929 => x"08",
          2930 => x"06",
          2931 => x"2e",
          2932 => x"80",
          2933 => x"1b",
          2934 => x"db",
          2935 => x"ec",
          2936 => x"ea",
          2937 => x"e0",
          2938 => x"34",
          2939 => x"51",
          2940 => x"81",
          2941 => x"83",
          2942 => x"53",
          2943 => x"d5",
          2944 => x"06",
          2945 => x"b4",
          2946 => x"84",
          2947 => x"e0",
          2948 => x"85",
          2949 => x"09",
          2950 => x"38",
          2951 => x"51",
          2952 => x"81",
          2953 => x"86",
          2954 => x"f2",
          2955 => x"06",
          2956 => x"9c",
          2957 => x"d8",
          2958 => x"e0",
          2959 => x"0c",
          2960 => x"51",
          2961 => x"81",
          2962 => x"8c",
          2963 => x"74",
          2964 => x"8c",
          2965 => x"53",
          2966 => x"8c",
          2967 => x"15",
          2968 => x"94",
          2969 => x"56",
          2970 => x"e0",
          2971 => x"0d",
          2972 => x"0d",
          2973 => x"55",
          2974 => x"b9",
          2975 => x"53",
          2976 => x"b1",
          2977 => x"52",
          2978 => x"a9",
          2979 => x"22",
          2980 => x"57",
          2981 => x"2e",
          2982 => x"99",
          2983 => x"33",
          2984 => x"3f",
          2985 => x"08",
          2986 => x"71",
          2987 => x"74",
          2988 => x"83",
          2989 => x"78",
          2990 => x"52",
          2991 => x"e0",
          2992 => x"0d",
          2993 => x"0d",
          2994 => x"33",
          2995 => x"3d",
          2996 => x"56",
          2997 => x"8b",
          2998 => x"81",
          2999 => x"24",
          3000 => x"ec",
          3001 => x"29",
          3002 => x"05",
          3003 => x"55",
          3004 => x"84",
          3005 => x"34",
          3006 => x"80",
          3007 => x"80",
          3008 => x"75",
          3009 => x"75",
          3010 => x"38",
          3011 => x"3d",
          3012 => x"05",
          3013 => x"3f",
          3014 => x"08",
          3015 => x"ec",
          3016 => x"3d",
          3017 => x"3d",
          3018 => x"84",
          3019 => x"05",
          3020 => x"89",
          3021 => x"2e",
          3022 => x"77",
          3023 => x"54",
          3024 => x"05",
          3025 => x"84",
          3026 => x"f6",
          3027 => x"ec",
          3028 => x"81",
          3029 => x"84",
          3030 => x"5c",
          3031 => x"3d",
          3032 => x"ed",
          3033 => x"ec",
          3034 => x"81",
          3035 => x"92",
          3036 => x"d7",
          3037 => x"98",
          3038 => x"73",
          3039 => x"38",
          3040 => x"9c",
          3041 => x"80",
          3042 => x"38",
          3043 => x"95",
          3044 => x"2e",
          3045 => x"aa",
          3046 => x"ea",
          3047 => x"ec",
          3048 => x"9e",
          3049 => x"05",
          3050 => x"54",
          3051 => x"38",
          3052 => x"70",
          3053 => x"54",
          3054 => x"8e",
          3055 => x"83",
          3056 => x"88",
          3057 => x"83",
          3058 => x"83",
          3059 => x"06",
          3060 => x"80",
          3061 => x"38",
          3062 => x"51",
          3063 => x"81",
          3064 => x"56",
          3065 => x"0a",
          3066 => x"05",
          3067 => x"3f",
          3068 => x"0b",
          3069 => x"80",
          3070 => x"7a",
          3071 => x"3f",
          3072 => x"9c",
          3073 => x"d1",
          3074 => x"81",
          3075 => x"34",
          3076 => x"80",
          3077 => x"b0",
          3078 => x"54",
          3079 => x"52",
          3080 => x"05",
          3081 => x"3f",
          3082 => x"08",
          3083 => x"e0",
          3084 => x"38",
          3085 => x"82",
          3086 => x"b2",
          3087 => x"84",
          3088 => x"06",
          3089 => x"73",
          3090 => x"38",
          3091 => x"ad",
          3092 => x"2a",
          3093 => x"51",
          3094 => x"2e",
          3095 => x"81",
          3096 => x"80",
          3097 => x"87",
          3098 => x"39",
          3099 => x"51",
          3100 => x"81",
          3101 => x"7b",
          3102 => x"12",
          3103 => x"81",
          3104 => x"81",
          3105 => x"83",
          3106 => x"06",
          3107 => x"80",
          3108 => x"77",
          3109 => x"58",
          3110 => x"08",
          3111 => x"63",
          3112 => x"63",
          3113 => x"57",
          3114 => x"81",
          3115 => x"81",
          3116 => x"88",
          3117 => x"9c",
          3118 => x"d2",
          3119 => x"ec",
          3120 => x"ec",
          3121 => x"1b",
          3122 => x"0c",
          3123 => x"22",
          3124 => x"77",
          3125 => x"80",
          3126 => x"34",
          3127 => x"1a",
          3128 => x"94",
          3129 => x"85",
          3130 => x"06",
          3131 => x"80",
          3132 => x"38",
          3133 => x"08",
          3134 => x"84",
          3135 => x"e0",
          3136 => x"0c",
          3137 => x"70",
          3138 => x"52",
          3139 => x"39",
          3140 => x"51",
          3141 => x"81",
          3142 => x"57",
          3143 => x"08",
          3144 => x"38",
          3145 => x"ec",
          3146 => x"2e",
          3147 => x"83",
          3148 => x"75",
          3149 => x"74",
          3150 => x"07",
          3151 => x"54",
          3152 => x"8a",
          3153 => x"75",
          3154 => x"73",
          3155 => x"98",
          3156 => x"a9",
          3157 => x"ff",
          3158 => x"80",
          3159 => x"76",
          3160 => x"d6",
          3161 => x"ec",
          3162 => x"38",
          3163 => x"39",
          3164 => x"81",
          3165 => x"05",
          3166 => x"84",
          3167 => x"0c",
          3168 => x"81",
          3169 => x"97",
          3170 => x"f2",
          3171 => x"63",
          3172 => x"40",
          3173 => x"7e",
          3174 => x"fc",
          3175 => x"51",
          3176 => x"81",
          3177 => x"55",
          3178 => x"08",
          3179 => x"19",
          3180 => x"80",
          3181 => x"74",
          3182 => x"39",
          3183 => x"81",
          3184 => x"56",
          3185 => x"82",
          3186 => x"39",
          3187 => x"1a",
          3188 => x"82",
          3189 => x"0b",
          3190 => x"81",
          3191 => x"39",
          3192 => x"94",
          3193 => x"55",
          3194 => x"83",
          3195 => x"7b",
          3196 => x"89",
          3197 => x"08",
          3198 => x"06",
          3199 => x"81",
          3200 => x"8a",
          3201 => x"05",
          3202 => x"06",
          3203 => x"a8",
          3204 => x"38",
          3205 => x"55",
          3206 => x"19",
          3207 => x"51",
          3208 => x"81",
          3209 => x"55",
          3210 => x"ff",
          3211 => x"ff",
          3212 => x"38",
          3213 => x"0c",
          3214 => x"52",
          3215 => x"cb",
          3216 => x"e0",
          3217 => x"ff",
          3218 => x"ec",
          3219 => x"7c",
          3220 => x"57",
          3221 => x"80",
          3222 => x"1a",
          3223 => x"22",
          3224 => x"75",
          3225 => x"38",
          3226 => x"58",
          3227 => x"53",
          3228 => x"1b",
          3229 => x"88",
          3230 => x"e0",
          3231 => x"38",
          3232 => x"33",
          3233 => x"80",
          3234 => x"b0",
          3235 => x"31",
          3236 => x"27",
          3237 => x"80",
          3238 => x"52",
          3239 => x"77",
          3240 => x"7d",
          3241 => x"e0",
          3242 => x"2b",
          3243 => x"76",
          3244 => x"94",
          3245 => x"ff",
          3246 => x"71",
          3247 => x"7b",
          3248 => x"38",
          3249 => x"19",
          3250 => x"51",
          3251 => x"81",
          3252 => x"fe",
          3253 => x"53",
          3254 => x"83",
          3255 => x"b4",
          3256 => x"51",
          3257 => x"7b",
          3258 => x"08",
          3259 => x"76",
          3260 => x"08",
          3261 => x"0c",
          3262 => x"f3",
          3263 => x"75",
          3264 => x"0c",
          3265 => x"04",
          3266 => x"60",
          3267 => x"40",
          3268 => x"80",
          3269 => x"3d",
          3270 => x"77",
          3271 => x"3f",
          3272 => x"08",
          3273 => x"e0",
          3274 => x"91",
          3275 => x"74",
          3276 => x"38",
          3277 => x"b8",
          3278 => x"33",
          3279 => x"70",
          3280 => x"56",
          3281 => x"74",
          3282 => x"a4",
          3283 => x"82",
          3284 => x"34",
          3285 => x"98",
          3286 => x"91",
          3287 => x"56",
          3288 => x"94",
          3289 => x"11",
          3290 => x"76",
          3291 => x"75",
          3292 => x"80",
          3293 => x"38",
          3294 => x"70",
          3295 => x"56",
          3296 => x"fd",
          3297 => x"11",
          3298 => x"77",
          3299 => x"5c",
          3300 => x"38",
          3301 => x"88",
          3302 => x"74",
          3303 => x"52",
          3304 => x"18",
          3305 => x"51",
          3306 => x"81",
          3307 => x"55",
          3308 => x"08",
          3309 => x"ab",
          3310 => x"2e",
          3311 => x"74",
          3312 => x"95",
          3313 => x"19",
          3314 => x"08",
          3315 => x"88",
          3316 => x"55",
          3317 => x"9c",
          3318 => x"09",
          3319 => x"38",
          3320 => x"c1",
          3321 => x"e0",
          3322 => x"38",
          3323 => x"52",
          3324 => x"97",
          3325 => x"e0",
          3326 => x"fe",
          3327 => x"ec",
          3328 => x"7c",
          3329 => x"57",
          3330 => x"80",
          3331 => x"1b",
          3332 => x"22",
          3333 => x"75",
          3334 => x"38",
          3335 => x"59",
          3336 => x"53",
          3337 => x"1a",
          3338 => x"be",
          3339 => x"e0",
          3340 => x"38",
          3341 => x"08",
          3342 => x"56",
          3343 => x"9b",
          3344 => x"53",
          3345 => x"77",
          3346 => x"7d",
          3347 => x"16",
          3348 => x"3f",
          3349 => x"0b",
          3350 => x"78",
          3351 => x"80",
          3352 => x"18",
          3353 => x"08",
          3354 => x"7e",
          3355 => x"3f",
          3356 => x"08",
          3357 => x"7e",
          3358 => x"0c",
          3359 => x"19",
          3360 => x"08",
          3361 => x"84",
          3362 => x"57",
          3363 => x"27",
          3364 => x"56",
          3365 => x"52",
          3366 => x"f9",
          3367 => x"e0",
          3368 => x"38",
          3369 => x"52",
          3370 => x"83",
          3371 => x"b4",
          3372 => x"d4",
          3373 => x"81",
          3374 => x"34",
          3375 => x"7e",
          3376 => x"0c",
          3377 => x"1a",
          3378 => x"94",
          3379 => x"1b",
          3380 => x"5e",
          3381 => x"27",
          3382 => x"55",
          3383 => x"0c",
          3384 => x"90",
          3385 => x"c0",
          3386 => x"90",
          3387 => x"56",
          3388 => x"e0",
          3389 => x"0d",
          3390 => x"0d",
          3391 => x"fc",
          3392 => x"52",
          3393 => x"3f",
          3394 => x"08",
          3395 => x"e0",
          3396 => x"38",
          3397 => x"70",
          3398 => x"81",
          3399 => x"55",
          3400 => x"80",
          3401 => x"16",
          3402 => x"51",
          3403 => x"81",
          3404 => x"57",
          3405 => x"08",
          3406 => x"a4",
          3407 => x"11",
          3408 => x"55",
          3409 => x"16",
          3410 => x"08",
          3411 => x"75",
          3412 => x"e8",
          3413 => x"08",
          3414 => x"51",
          3415 => x"82",
          3416 => x"52",
          3417 => x"c9",
          3418 => x"52",
          3419 => x"c9",
          3420 => x"54",
          3421 => x"15",
          3422 => x"cc",
          3423 => x"ec",
          3424 => x"17",
          3425 => x"06",
          3426 => x"90",
          3427 => x"81",
          3428 => x"8a",
          3429 => x"fc",
          3430 => x"70",
          3431 => x"d9",
          3432 => x"e0",
          3433 => x"ec",
          3434 => x"38",
          3435 => x"05",
          3436 => x"f1",
          3437 => x"ec",
          3438 => x"81",
          3439 => x"87",
          3440 => x"e0",
          3441 => x"72",
          3442 => x"0c",
          3443 => x"04",
          3444 => x"84",
          3445 => x"e4",
          3446 => x"80",
          3447 => x"e0",
          3448 => x"38",
          3449 => x"08",
          3450 => x"34",
          3451 => x"81",
          3452 => x"83",
          3453 => x"ef",
          3454 => x"53",
          3455 => x"05",
          3456 => x"51",
          3457 => x"81",
          3458 => x"55",
          3459 => x"08",
          3460 => x"76",
          3461 => x"93",
          3462 => x"51",
          3463 => x"81",
          3464 => x"55",
          3465 => x"08",
          3466 => x"80",
          3467 => x"70",
          3468 => x"56",
          3469 => x"89",
          3470 => x"94",
          3471 => x"b2",
          3472 => x"05",
          3473 => x"2a",
          3474 => x"51",
          3475 => x"80",
          3476 => x"76",
          3477 => x"52",
          3478 => x"3f",
          3479 => x"08",
          3480 => x"8e",
          3481 => x"e0",
          3482 => x"09",
          3483 => x"38",
          3484 => x"81",
          3485 => x"93",
          3486 => x"e4",
          3487 => x"6f",
          3488 => x"7a",
          3489 => x"9e",
          3490 => x"05",
          3491 => x"51",
          3492 => x"81",
          3493 => x"57",
          3494 => x"08",
          3495 => x"7b",
          3496 => x"94",
          3497 => x"55",
          3498 => x"73",
          3499 => x"ed",
          3500 => x"93",
          3501 => x"55",
          3502 => x"81",
          3503 => x"57",
          3504 => x"08",
          3505 => x"68",
          3506 => x"c9",
          3507 => x"ec",
          3508 => x"81",
          3509 => x"82",
          3510 => x"52",
          3511 => x"a3",
          3512 => x"e0",
          3513 => x"52",
          3514 => x"b8",
          3515 => x"e0",
          3516 => x"ec",
          3517 => x"a2",
          3518 => x"74",
          3519 => x"3f",
          3520 => x"08",
          3521 => x"e0",
          3522 => x"69",
          3523 => x"d9",
          3524 => x"81",
          3525 => x"2e",
          3526 => x"52",
          3527 => x"cf",
          3528 => x"e0",
          3529 => x"ec",
          3530 => x"2e",
          3531 => x"84",
          3532 => x"06",
          3533 => x"57",
          3534 => x"76",
          3535 => x"9e",
          3536 => x"05",
          3537 => x"dc",
          3538 => x"90",
          3539 => x"81",
          3540 => x"56",
          3541 => x"80",
          3542 => x"02",
          3543 => x"81",
          3544 => x"70",
          3545 => x"56",
          3546 => x"81",
          3547 => x"78",
          3548 => x"38",
          3549 => x"99",
          3550 => x"81",
          3551 => x"18",
          3552 => x"18",
          3553 => x"58",
          3554 => x"33",
          3555 => x"ee",
          3556 => x"6f",
          3557 => x"af",
          3558 => x"8d",
          3559 => x"2e",
          3560 => x"8a",
          3561 => x"6f",
          3562 => x"af",
          3563 => x"0b",
          3564 => x"33",
          3565 => x"81",
          3566 => x"70",
          3567 => x"52",
          3568 => x"56",
          3569 => x"8d",
          3570 => x"70",
          3571 => x"51",
          3572 => x"f5",
          3573 => x"54",
          3574 => x"a7",
          3575 => x"74",
          3576 => x"38",
          3577 => x"73",
          3578 => x"81",
          3579 => x"81",
          3580 => x"39",
          3581 => x"81",
          3582 => x"74",
          3583 => x"81",
          3584 => x"91",
          3585 => x"6e",
          3586 => x"59",
          3587 => x"7a",
          3588 => x"5c",
          3589 => x"26",
          3590 => x"7a",
          3591 => x"ec",
          3592 => x"3d",
          3593 => x"3d",
          3594 => x"8d",
          3595 => x"54",
          3596 => x"55",
          3597 => x"81",
          3598 => x"53",
          3599 => x"08",
          3600 => x"91",
          3601 => x"72",
          3602 => x"8c",
          3603 => x"73",
          3604 => x"38",
          3605 => x"70",
          3606 => x"81",
          3607 => x"57",
          3608 => x"73",
          3609 => x"08",
          3610 => x"94",
          3611 => x"75",
          3612 => x"97",
          3613 => x"11",
          3614 => x"2b",
          3615 => x"73",
          3616 => x"38",
          3617 => x"16",
          3618 => x"a0",
          3619 => x"e0",
          3620 => x"78",
          3621 => x"55",
          3622 => x"90",
          3623 => x"e0",
          3624 => x"96",
          3625 => x"70",
          3626 => x"94",
          3627 => x"71",
          3628 => x"08",
          3629 => x"53",
          3630 => x"15",
          3631 => x"a6",
          3632 => x"74",
          3633 => x"3f",
          3634 => x"08",
          3635 => x"e0",
          3636 => x"81",
          3637 => x"ec",
          3638 => x"2e",
          3639 => x"81",
          3640 => x"88",
          3641 => x"98",
          3642 => x"80",
          3643 => x"38",
          3644 => x"80",
          3645 => x"77",
          3646 => x"08",
          3647 => x"0c",
          3648 => x"70",
          3649 => x"81",
          3650 => x"5a",
          3651 => x"2e",
          3652 => x"52",
          3653 => x"f9",
          3654 => x"e0",
          3655 => x"ec",
          3656 => x"38",
          3657 => x"08",
          3658 => x"73",
          3659 => x"c7",
          3660 => x"ec",
          3661 => x"73",
          3662 => x"38",
          3663 => x"af",
          3664 => x"73",
          3665 => x"27",
          3666 => x"98",
          3667 => x"a0",
          3668 => x"08",
          3669 => x"0c",
          3670 => x"06",
          3671 => x"2e",
          3672 => x"52",
          3673 => x"a3",
          3674 => x"e0",
          3675 => x"82",
          3676 => x"34",
          3677 => x"c4",
          3678 => x"91",
          3679 => x"53",
          3680 => x"89",
          3681 => x"e0",
          3682 => x"94",
          3683 => x"8c",
          3684 => x"27",
          3685 => x"8c",
          3686 => x"15",
          3687 => x"07",
          3688 => x"16",
          3689 => x"ff",
          3690 => x"80",
          3691 => x"77",
          3692 => x"2e",
          3693 => x"9c",
          3694 => x"53",
          3695 => x"e0",
          3696 => x"0d",
          3697 => x"0d",
          3698 => x"54",
          3699 => x"81",
          3700 => x"53",
          3701 => x"05",
          3702 => x"84",
          3703 => x"e7",
          3704 => x"e0",
          3705 => x"ec",
          3706 => x"ea",
          3707 => x"0c",
          3708 => x"51",
          3709 => x"81",
          3710 => x"55",
          3711 => x"08",
          3712 => x"ab",
          3713 => x"98",
          3714 => x"80",
          3715 => x"38",
          3716 => x"70",
          3717 => x"81",
          3718 => x"57",
          3719 => x"ad",
          3720 => x"08",
          3721 => x"d3",
          3722 => x"ec",
          3723 => x"17",
          3724 => x"86",
          3725 => x"17",
          3726 => x"75",
          3727 => x"3f",
          3728 => x"08",
          3729 => x"2e",
          3730 => x"85",
          3731 => x"86",
          3732 => x"2e",
          3733 => x"76",
          3734 => x"73",
          3735 => x"0c",
          3736 => x"04",
          3737 => x"76",
          3738 => x"05",
          3739 => x"53",
          3740 => x"81",
          3741 => x"87",
          3742 => x"e0",
          3743 => x"86",
          3744 => x"fb",
          3745 => x"79",
          3746 => x"05",
          3747 => x"56",
          3748 => x"3f",
          3749 => x"08",
          3750 => x"e0",
          3751 => x"38",
          3752 => x"81",
          3753 => x"52",
          3754 => x"f8",
          3755 => x"e0",
          3756 => x"ca",
          3757 => x"e0",
          3758 => x"51",
          3759 => x"81",
          3760 => x"53",
          3761 => x"08",
          3762 => x"81",
          3763 => x"80",
          3764 => x"81",
          3765 => x"a6",
          3766 => x"73",
          3767 => x"3f",
          3768 => x"51",
          3769 => x"81",
          3770 => x"84",
          3771 => x"70",
          3772 => x"2c",
          3773 => x"e0",
          3774 => x"51",
          3775 => x"81",
          3776 => x"87",
          3777 => x"ee",
          3778 => x"57",
          3779 => x"3d",
          3780 => x"3d",
          3781 => x"af",
          3782 => x"e0",
          3783 => x"ec",
          3784 => x"38",
          3785 => x"51",
          3786 => x"81",
          3787 => x"55",
          3788 => x"08",
          3789 => x"80",
          3790 => x"70",
          3791 => x"58",
          3792 => x"85",
          3793 => x"8d",
          3794 => x"2e",
          3795 => x"52",
          3796 => x"be",
          3797 => x"ec",
          3798 => x"3d",
          3799 => x"3d",
          3800 => x"55",
          3801 => x"92",
          3802 => x"52",
          3803 => x"de",
          3804 => x"ec",
          3805 => x"81",
          3806 => x"82",
          3807 => x"74",
          3808 => x"98",
          3809 => x"11",
          3810 => x"59",
          3811 => x"75",
          3812 => x"38",
          3813 => x"81",
          3814 => x"5b",
          3815 => x"82",
          3816 => x"39",
          3817 => x"08",
          3818 => x"59",
          3819 => x"09",
          3820 => x"38",
          3821 => x"57",
          3822 => x"3d",
          3823 => x"c1",
          3824 => x"ec",
          3825 => x"2e",
          3826 => x"ec",
          3827 => x"2e",
          3828 => x"ec",
          3829 => x"70",
          3830 => x"08",
          3831 => x"7a",
          3832 => x"7f",
          3833 => x"54",
          3834 => x"77",
          3835 => x"80",
          3836 => x"15",
          3837 => x"e0",
          3838 => x"75",
          3839 => x"52",
          3840 => x"52",
          3841 => x"8d",
          3842 => x"e0",
          3843 => x"ec",
          3844 => x"d6",
          3845 => x"33",
          3846 => x"1a",
          3847 => x"54",
          3848 => x"09",
          3849 => x"38",
          3850 => x"ff",
          3851 => x"81",
          3852 => x"83",
          3853 => x"70",
          3854 => x"25",
          3855 => x"59",
          3856 => x"9b",
          3857 => x"51",
          3858 => x"3f",
          3859 => x"08",
          3860 => x"70",
          3861 => x"25",
          3862 => x"59",
          3863 => x"75",
          3864 => x"7a",
          3865 => x"ff",
          3866 => x"7c",
          3867 => x"90",
          3868 => x"11",
          3869 => x"56",
          3870 => x"15",
          3871 => x"ec",
          3872 => x"3d",
          3873 => x"3d",
          3874 => x"3d",
          3875 => x"70",
          3876 => x"dd",
          3877 => x"e0",
          3878 => x"ec",
          3879 => x"a8",
          3880 => x"33",
          3881 => x"a0",
          3882 => x"33",
          3883 => x"70",
          3884 => x"55",
          3885 => x"73",
          3886 => x"8e",
          3887 => x"08",
          3888 => x"18",
          3889 => x"80",
          3890 => x"38",
          3891 => x"08",
          3892 => x"08",
          3893 => x"c4",
          3894 => x"ec",
          3895 => x"88",
          3896 => x"80",
          3897 => x"17",
          3898 => x"51",
          3899 => x"3f",
          3900 => x"08",
          3901 => x"81",
          3902 => x"81",
          3903 => x"e0",
          3904 => x"09",
          3905 => x"38",
          3906 => x"39",
          3907 => x"77",
          3908 => x"e0",
          3909 => x"08",
          3910 => x"98",
          3911 => x"81",
          3912 => x"52",
          3913 => x"bd",
          3914 => x"e0",
          3915 => x"17",
          3916 => x"0c",
          3917 => x"80",
          3918 => x"73",
          3919 => x"75",
          3920 => x"38",
          3921 => x"34",
          3922 => x"81",
          3923 => x"89",
          3924 => x"e2",
          3925 => x"53",
          3926 => x"a4",
          3927 => x"3d",
          3928 => x"3f",
          3929 => x"08",
          3930 => x"e0",
          3931 => x"38",
          3932 => x"3d",
          3933 => x"3d",
          3934 => x"d1",
          3935 => x"ec",
          3936 => x"81",
          3937 => x"81",
          3938 => x"80",
          3939 => x"70",
          3940 => x"81",
          3941 => x"56",
          3942 => x"81",
          3943 => x"98",
          3944 => x"74",
          3945 => x"38",
          3946 => x"05",
          3947 => x"06",
          3948 => x"55",
          3949 => x"38",
          3950 => x"51",
          3951 => x"81",
          3952 => x"74",
          3953 => x"81",
          3954 => x"56",
          3955 => x"80",
          3956 => x"54",
          3957 => x"08",
          3958 => x"2e",
          3959 => x"73",
          3960 => x"e0",
          3961 => x"52",
          3962 => x"52",
          3963 => x"3f",
          3964 => x"08",
          3965 => x"e0",
          3966 => x"38",
          3967 => x"08",
          3968 => x"cc",
          3969 => x"ec",
          3970 => x"81",
          3971 => x"86",
          3972 => x"80",
          3973 => x"ec",
          3974 => x"2e",
          3975 => x"ec",
          3976 => x"c0",
          3977 => x"ce",
          3978 => x"ec",
          3979 => x"ec",
          3980 => x"70",
          3981 => x"08",
          3982 => x"51",
          3983 => x"80",
          3984 => x"73",
          3985 => x"38",
          3986 => x"52",
          3987 => x"95",
          3988 => x"e0",
          3989 => x"8c",
          3990 => x"ff",
          3991 => x"81",
          3992 => x"55",
          3993 => x"e0",
          3994 => x"0d",
          3995 => x"0d",
          3996 => x"3d",
          3997 => x"9a",
          3998 => x"cb",
          3999 => x"e0",
          4000 => x"ec",
          4001 => x"b0",
          4002 => x"69",
          4003 => x"70",
          4004 => x"97",
          4005 => x"e0",
          4006 => x"ec",
          4007 => x"38",
          4008 => x"94",
          4009 => x"e0",
          4010 => x"09",
          4011 => x"88",
          4012 => x"df",
          4013 => x"85",
          4014 => x"51",
          4015 => x"74",
          4016 => x"78",
          4017 => x"8a",
          4018 => x"57",
          4019 => x"81",
          4020 => x"75",
          4021 => x"ec",
          4022 => x"38",
          4023 => x"ec",
          4024 => x"2e",
          4025 => x"83",
          4026 => x"81",
          4027 => x"ff",
          4028 => x"06",
          4029 => x"54",
          4030 => x"73",
          4031 => x"81",
          4032 => x"52",
          4033 => x"a4",
          4034 => x"e0",
          4035 => x"ec",
          4036 => x"9a",
          4037 => x"a0",
          4038 => x"51",
          4039 => x"3f",
          4040 => x"0b",
          4041 => x"78",
          4042 => x"bf",
          4043 => x"88",
          4044 => x"80",
          4045 => x"ff",
          4046 => x"75",
          4047 => x"11",
          4048 => x"f8",
          4049 => x"78",
          4050 => x"80",
          4051 => x"ff",
          4052 => x"78",
          4053 => x"80",
          4054 => x"7f",
          4055 => x"d4",
          4056 => x"c9",
          4057 => x"54",
          4058 => x"15",
          4059 => x"cb",
          4060 => x"ec",
          4061 => x"81",
          4062 => x"b2",
          4063 => x"b2",
          4064 => x"96",
          4065 => x"b5",
          4066 => x"53",
          4067 => x"51",
          4068 => x"64",
          4069 => x"8b",
          4070 => x"54",
          4071 => x"15",
          4072 => x"ff",
          4073 => x"81",
          4074 => x"54",
          4075 => x"53",
          4076 => x"51",
          4077 => x"3f",
          4078 => x"e0",
          4079 => x"0d",
          4080 => x"0d",
          4081 => x"05",
          4082 => x"3f",
          4083 => x"3d",
          4084 => x"52",
          4085 => x"d5",
          4086 => x"ec",
          4087 => x"81",
          4088 => x"82",
          4089 => x"4d",
          4090 => x"52",
          4091 => x"52",
          4092 => x"3f",
          4093 => x"08",
          4094 => x"e0",
          4095 => x"38",
          4096 => x"05",
          4097 => x"06",
          4098 => x"73",
          4099 => x"a0",
          4100 => x"08",
          4101 => x"ff",
          4102 => x"ff",
          4103 => x"ac",
          4104 => x"92",
          4105 => x"54",
          4106 => x"3f",
          4107 => x"52",
          4108 => x"f7",
          4109 => x"e0",
          4110 => x"ec",
          4111 => x"38",
          4112 => x"09",
          4113 => x"38",
          4114 => x"08",
          4115 => x"88",
          4116 => x"39",
          4117 => x"08",
          4118 => x"81",
          4119 => x"38",
          4120 => x"b1",
          4121 => x"e0",
          4122 => x"ec",
          4123 => x"c8",
          4124 => x"93",
          4125 => x"ff",
          4126 => x"8d",
          4127 => x"b4",
          4128 => x"af",
          4129 => x"17",
          4130 => x"33",
          4131 => x"70",
          4132 => x"55",
          4133 => x"38",
          4134 => x"54",
          4135 => x"34",
          4136 => x"0b",
          4137 => x"8b",
          4138 => x"84",
          4139 => x"06",
          4140 => x"73",
          4141 => x"e5",
          4142 => x"2e",
          4143 => x"75",
          4144 => x"c6",
          4145 => x"ec",
          4146 => x"78",
          4147 => x"bb",
          4148 => x"81",
          4149 => x"80",
          4150 => x"38",
          4151 => x"08",
          4152 => x"ff",
          4153 => x"81",
          4154 => x"79",
          4155 => x"58",
          4156 => x"ec",
          4157 => x"c0",
          4158 => x"33",
          4159 => x"2e",
          4160 => x"99",
          4161 => x"75",
          4162 => x"c6",
          4163 => x"54",
          4164 => x"15",
          4165 => x"81",
          4166 => x"9c",
          4167 => x"c8",
          4168 => x"ec",
          4169 => x"81",
          4170 => x"8c",
          4171 => x"ff",
          4172 => x"81",
          4173 => x"55",
          4174 => x"e0",
          4175 => x"0d",
          4176 => x"0d",
          4177 => x"05",
          4178 => x"05",
          4179 => x"33",
          4180 => x"53",
          4181 => x"05",
          4182 => x"51",
          4183 => x"81",
          4184 => x"55",
          4185 => x"08",
          4186 => x"78",
          4187 => x"95",
          4188 => x"51",
          4189 => x"81",
          4190 => x"55",
          4191 => x"08",
          4192 => x"80",
          4193 => x"81",
          4194 => x"86",
          4195 => x"38",
          4196 => x"61",
          4197 => x"12",
          4198 => x"7a",
          4199 => x"51",
          4200 => x"74",
          4201 => x"78",
          4202 => x"83",
          4203 => x"51",
          4204 => x"3f",
          4205 => x"08",
          4206 => x"ec",
          4207 => x"3d",
          4208 => x"3d",
          4209 => x"82",
          4210 => x"d0",
          4211 => x"3d",
          4212 => x"3f",
          4213 => x"08",
          4214 => x"e0",
          4215 => x"38",
          4216 => x"52",
          4217 => x"05",
          4218 => x"3f",
          4219 => x"08",
          4220 => x"e0",
          4221 => x"02",
          4222 => x"33",
          4223 => x"54",
          4224 => x"a6",
          4225 => x"22",
          4226 => x"71",
          4227 => x"53",
          4228 => x"51",
          4229 => x"3f",
          4230 => x"0b",
          4231 => x"76",
          4232 => x"b8",
          4233 => x"e0",
          4234 => x"81",
          4235 => x"93",
          4236 => x"ea",
          4237 => x"6b",
          4238 => x"53",
          4239 => x"05",
          4240 => x"51",
          4241 => x"81",
          4242 => x"81",
          4243 => x"30",
          4244 => x"e0",
          4245 => x"25",
          4246 => x"79",
          4247 => x"85",
          4248 => x"75",
          4249 => x"73",
          4250 => x"f9",
          4251 => x"80",
          4252 => x"8d",
          4253 => x"54",
          4254 => x"3f",
          4255 => x"08",
          4256 => x"e0",
          4257 => x"38",
          4258 => x"51",
          4259 => x"81",
          4260 => x"57",
          4261 => x"08",
          4262 => x"ec",
          4263 => x"ec",
          4264 => x"5b",
          4265 => x"18",
          4266 => x"18",
          4267 => x"74",
          4268 => x"81",
          4269 => x"78",
          4270 => x"8b",
          4271 => x"54",
          4272 => x"75",
          4273 => x"38",
          4274 => x"1b",
          4275 => x"55",
          4276 => x"2e",
          4277 => x"39",
          4278 => x"09",
          4279 => x"38",
          4280 => x"80",
          4281 => x"70",
          4282 => x"25",
          4283 => x"80",
          4284 => x"38",
          4285 => x"bc",
          4286 => x"11",
          4287 => x"ff",
          4288 => x"81",
          4289 => x"57",
          4290 => x"08",
          4291 => x"70",
          4292 => x"80",
          4293 => x"83",
          4294 => x"80",
          4295 => x"84",
          4296 => x"a7",
          4297 => x"b4",
          4298 => x"ad",
          4299 => x"ec",
          4300 => x"0c",
          4301 => x"e0",
          4302 => x"0d",
          4303 => x"0d",
          4304 => x"3d",
          4305 => x"52",
          4306 => x"ce",
          4307 => x"ec",
          4308 => x"ec",
          4309 => x"54",
          4310 => x"08",
          4311 => x"8b",
          4312 => x"8b",
          4313 => x"59",
          4314 => x"3f",
          4315 => x"33",
          4316 => x"06",
          4317 => x"57",
          4318 => x"81",
          4319 => x"58",
          4320 => x"06",
          4321 => x"4e",
          4322 => x"ff",
          4323 => x"81",
          4324 => x"80",
          4325 => x"6c",
          4326 => x"53",
          4327 => x"ae",
          4328 => x"ec",
          4329 => x"2e",
          4330 => x"88",
          4331 => x"6d",
          4332 => x"55",
          4333 => x"ec",
          4334 => x"ff",
          4335 => x"83",
          4336 => x"51",
          4337 => x"26",
          4338 => x"15",
          4339 => x"ff",
          4340 => x"80",
          4341 => x"87",
          4342 => x"b0",
          4343 => x"74",
          4344 => x"38",
          4345 => x"dd",
          4346 => x"ae",
          4347 => x"ec",
          4348 => x"38",
          4349 => x"27",
          4350 => x"89",
          4351 => x"8b",
          4352 => x"27",
          4353 => x"55",
          4354 => x"81",
          4355 => x"8f",
          4356 => x"2a",
          4357 => x"70",
          4358 => x"34",
          4359 => x"74",
          4360 => x"05",
          4361 => x"17",
          4362 => x"70",
          4363 => x"52",
          4364 => x"73",
          4365 => x"c8",
          4366 => x"33",
          4367 => x"73",
          4368 => x"81",
          4369 => x"80",
          4370 => x"02",
          4371 => x"76",
          4372 => x"51",
          4373 => x"2e",
          4374 => x"87",
          4375 => x"57",
          4376 => x"79",
          4377 => x"80",
          4378 => x"70",
          4379 => x"ba",
          4380 => x"ec",
          4381 => x"81",
          4382 => x"80",
          4383 => x"52",
          4384 => x"bf",
          4385 => x"ec",
          4386 => x"81",
          4387 => x"8d",
          4388 => x"c4",
          4389 => x"e5",
          4390 => x"c6",
          4391 => x"e0",
          4392 => x"09",
          4393 => x"cc",
          4394 => x"76",
          4395 => x"c4",
          4396 => x"74",
          4397 => x"b0",
          4398 => x"e0",
          4399 => x"ec",
          4400 => x"38",
          4401 => x"ec",
          4402 => x"67",
          4403 => x"db",
          4404 => x"88",
          4405 => x"34",
          4406 => x"52",
          4407 => x"ab",
          4408 => x"54",
          4409 => x"15",
          4410 => x"ff",
          4411 => x"81",
          4412 => x"54",
          4413 => x"81",
          4414 => x"9c",
          4415 => x"f2",
          4416 => x"62",
          4417 => x"80",
          4418 => x"93",
          4419 => x"55",
          4420 => x"5e",
          4421 => x"3f",
          4422 => x"08",
          4423 => x"e0",
          4424 => x"38",
          4425 => x"58",
          4426 => x"38",
          4427 => x"97",
          4428 => x"08",
          4429 => x"38",
          4430 => x"70",
          4431 => x"81",
          4432 => x"55",
          4433 => x"87",
          4434 => x"39",
          4435 => x"90",
          4436 => x"82",
          4437 => x"8a",
          4438 => x"89",
          4439 => x"7f",
          4440 => x"56",
          4441 => x"3f",
          4442 => x"06",
          4443 => x"72",
          4444 => x"81",
          4445 => x"05",
          4446 => x"7c",
          4447 => x"55",
          4448 => x"27",
          4449 => x"16",
          4450 => x"83",
          4451 => x"76",
          4452 => x"80",
          4453 => x"79",
          4454 => x"99",
          4455 => x"7f",
          4456 => x"14",
          4457 => x"83",
          4458 => x"81",
          4459 => x"81",
          4460 => x"38",
          4461 => x"08",
          4462 => x"95",
          4463 => x"e0",
          4464 => x"81",
          4465 => x"7b",
          4466 => x"06",
          4467 => x"39",
          4468 => x"56",
          4469 => x"09",
          4470 => x"b9",
          4471 => x"80",
          4472 => x"80",
          4473 => x"78",
          4474 => x"7a",
          4475 => x"38",
          4476 => x"73",
          4477 => x"81",
          4478 => x"ff",
          4479 => x"74",
          4480 => x"ff",
          4481 => x"81",
          4482 => x"58",
          4483 => x"08",
          4484 => x"74",
          4485 => x"16",
          4486 => x"73",
          4487 => x"39",
          4488 => x"7e",
          4489 => x"0c",
          4490 => x"2e",
          4491 => x"88",
          4492 => x"8c",
          4493 => x"1a",
          4494 => x"07",
          4495 => x"1b",
          4496 => x"08",
          4497 => x"16",
          4498 => x"75",
          4499 => x"38",
          4500 => x"90",
          4501 => x"15",
          4502 => x"54",
          4503 => x"34",
          4504 => x"81",
          4505 => x"90",
          4506 => x"e9",
          4507 => x"6d",
          4508 => x"80",
          4509 => x"9d",
          4510 => x"5c",
          4511 => x"3f",
          4512 => x"0b",
          4513 => x"08",
          4514 => x"38",
          4515 => x"08",
          4516 => x"ec",
          4517 => x"08",
          4518 => x"80",
          4519 => x"80",
          4520 => x"ec",
          4521 => x"ff",
          4522 => x"52",
          4523 => x"a0",
          4524 => x"ec",
          4525 => x"ff",
          4526 => x"06",
          4527 => x"56",
          4528 => x"38",
          4529 => x"70",
          4530 => x"55",
          4531 => x"8b",
          4532 => x"3d",
          4533 => x"83",
          4534 => x"ff",
          4535 => x"81",
          4536 => x"99",
          4537 => x"74",
          4538 => x"38",
          4539 => x"80",
          4540 => x"ff",
          4541 => x"55",
          4542 => x"83",
          4543 => x"78",
          4544 => x"38",
          4545 => x"26",
          4546 => x"81",
          4547 => x"8b",
          4548 => x"79",
          4549 => x"80",
          4550 => x"93",
          4551 => x"39",
          4552 => x"6e",
          4553 => x"89",
          4554 => x"48",
          4555 => x"83",
          4556 => x"61",
          4557 => x"25",
          4558 => x"55",
          4559 => x"8a",
          4560 => x"3d",
          4561 => x"81",
          4562 => x"ff",
          4563 => x"81",
          4564 => x"e0",
          4565 => x"38",
          4566 => x"70",
          4567 => x"ec",
          4568 => x"56",
          4569 => x"38",
          4570 => x"55",
          4571 => x"75",
          4572 => x"38",
          4573 => x"70",
          4574 => x"ff",
          4575 => x"83",
          4576 => x"78",
          4577 => x"89",
          4578 => x"81",
          4579 => x"06",
          4580 => x"80",
          4581 => x"77",
          4582 => x"74",
          4583 => x"8d",
          4584 => x"06",
          4585 => x"2e",
          4586 => x"77",
          4587 => x"93",
          4588 => x"74",
          4589 => x"cb",
          4590 => x"7d",
          4591 => x"81",
          4592 => x"38",
          4593 => x"66",
          4594 => x"81",
          4595 => x"d4",
          4596 => x"74",
          4597 => x"38",
          4598 => x"98",
          4599 => x"d4",
          4600 => x"82",
          4601 => x"57",
          4602 => x"80",
          4603 => x"76",
          4604 => x"38",
          4605 => x"51",
          4606 => x"3f",
          4607 => x"08",
          4608 => x"87",
          4609 => x"2a",
          4610 => x"5c",
          4611 => x"ec",
          4612 => x"80",
          4613 => x"44",
          4614 => x"0a",
          4615 => x"ec",
          4616 => x"39",
          4617 => x"66",
          4618 => x"81",
          4619 => x"c4",
          4620 => x"74",
          4621 => x"38",
          4622 => x"98",
          4623 => x"c4",
          4624 => x"82",
          4625 => x"57",
          4626 => x"80",
          4627 => x"76",
          4628 => x"38",
          4629 => x"51",
          4630 => x"3f",
          4631 => x"08",
          4632 => x"57",
          4633 => x"08",
          4634 => x"96",
          4635 => x"81",
          4636 => x"10",
          4637 => x"08",
          4638 => x"72",
          4639 => x"59",
          4640 => x"ff",
          4641 => x"5d",
          4642 => x"44",
          4643 => x"11",
          4644 => x"70",
          4645 => x"71",
          4646 => x"06",
          4647 => x"52",
          4648 => x"40",
          4649 => x"09",
          4650 => x"38",
          4651 => x"18",
          4652 => x"39",
          4653 => x"79",
          4654 => x"70",
          4655 => x"58",
          4656 => x"76",
          4657 => x"38",
          4658 => x"7d",
          4659 => x"70",
          4660 => x"55",
          4661 => x"3f",
          4662 => x"08",
          4663 => x"2e",
          4664 => x"9b",
          4665 => x"e0",
          4666 => x"f5",
          4667 => x"38",
          4668 => x"38",
          4669 => x"59",
          4670 => x"38",
          4671 => x"7d",
          4672 => x"81",
          4673 => x"38",
          4674 => x"0b",
          4675 => x"08",
          4676 => x"78",
          4677 => x"1a",
          4678 => x"c0",
          4679 => x"74",
          4680 => x"39",
          4681 => x"55",
          4682 => x"8f",
          4683 => x"fd",
          4684 => x"ec",
          4685 => x"f5",
          4686 => x"78",
          4687 => x"79",
          4688 => x"80",
          4689 => x"f1",
          4690 => x"39",
          4691 => x"81",
          4692 => x"06",
          4693 => x"55",
          4694 => x"27",
          4695 => x"81",
          4696 => x"56",
          4697 => x"38",
          4698 => x"80",
          4699 => x"ff",
          4700 => x"8b",
          4701 => x"ec",
          4702 => x"ff",
          4703 => x"84",
          4704 => x"1b",
          4705 => x"b3",
          4706 => x"1c",
          4707 => x"ff",
          4708 => x"8e",
          4709 => x"a1",
          4710 => x"0b",
          4711 => x"7d",
          4712 => x"30",
          4713 => x"84",
          4714 => x"51",
          4715 => x"51",
          4716 => x"3f",
          4717 => x"83",
          4718 => x"90",
          4719 => x"ff",
          4720 => x"93",
          4721 => x"a0",
          4722 => x"39",
          4723 => x"1b",
          4724 => x"85",
          4725 => x"95",
          4726 => x"52",
          4727 => x"ff",
          4728 => x"81",
          4729 => x"1b",
          4730 => x"cf",
          4731 => x"9c",
          4732 => x"a0",
          4733 => x"83",
          4734 => x"06",
          4735 => x"82",
          4736 => x"52",
          4737 => x"51",
          4738 => x"3f",
          4739 => x"1b",
          4740 => x"c5",
          4741 => x"ac",
          4742 => x"a0",
          4743 => x"52",
          4744 => x"ff",
          4745 => x"86",
          4746 => x"51",
          4747 => x"3f",
          4748 => x"80",
          4749 => x"a9",
          4750 => x"1c",
          4751 => x"81",
          4752 => x"80",
          4753 => x"ae",
          4754 => x"b2",
          4755 => x"1b",
          4756 => x"85",
          4757 => x"ff",
          4758 => x"96",
          4759 => x"9f",
          4760 => x"80",
          4761 => x"34",
          4762 => x"1c",
          4763 => x"81",
          4764 => x"ab",
          4765 => x"a0",
          4766 => x"d4",
          4767 => x"fe",
          4768 => x"59",
          4769 => x"3f",
          4770 => x"53",
          4771 => x"51",
          4772 => x"3f",
          4773 => x"ec",
          4774 => x"e7",
          4775 => x"2e",
          4776 => x"80",
          4777 => x"54",
          4778 => x"53",
          4779 => x"51",
          4780 => x"3f",
          4781 => x"80",
          4782 => x"ff",
          4783 => x"84",
          4784 => x"d2",
          4785 => x"ff",
          4786 => x"86",
          4787 => x"f2",
          4788 => x"1b",
          4789 => x"81",
          4790 => x"52",
          4791 => x"51",
          4792 => x"3f",
          4793 => x"ec",
          4794 => x"9e",
          4795 => x"d4",
          4796 => x"51",
          4797 => x"3f",
          4798 => x"87",
          4799 => x"52",
          4800 => x"9a",
          4801 => x"54",
          4802 => x"7a",
          4803 => x"ff",
          4804 => x"65",
          4805 => x"7a",
          4806 => x"8f",
          4807 => x"80",
          4808 => x"2e",
          4809 => x"9a",
          4810 => x"7a",
          4811 => x"a9",
          4812 => x"84",
          4813 => x"9e",
          4814 => x"0a",
          4815 => x"51",
          4816 => x"ff",
          4817 => x"7d",
          4818 => x"38",
          4819 => x"52",
          4820 => x"9e",
          4821 => x"55",
          4822 => x"62",
          4823 => x"74",
          4824 => x"75",
          4825 => x"7e",
          4826 => x"fe",
          4827 => x"e0",
          4828 => x"38",
          4829 => x"81",
          4830 => x"52",
          4831 => x"9e",
          4832 => x"16",
          4833 => x"56",
          4834 => x"38",
          4835 => x"77",
          4836 => x"8d",
          4837 => x"7d",
          4838 => x"38",
          4839 => x"57",
          4840 => x"83",
          4841 => x"76",
          4842 => x"7a",
          4843 => x"ff",
          4844 => x"81",
          4845 => x"81",
          4846 => x"16",
          4847 => x"56",
          4848 => x"38",
          4849 => x"83",
          4850 => x"86",
          4851 => x"ff",
          4852 => x"38",
          4853 => x"82",
          4854 => x"81",
          4855 => x"06",
          4856 => x"fe",
          4857 => x"53",
          4858 => x"51",
          4859 => x"3f",
          4860 => x"52",
          4861 => x"9c",
          4862 => x"be",
          4863 => x"75",
          4864 => x"81",
          4865 => x"0b",
          4866 => x"77",
          4867 => x"75",
          4868 => x"60",
          4869 => x"80",
          4870 => x"75",
          4871 => x"8c",
          4872 => x"85",
          4873 => x"ec",
          4874 => x"2a",
          4875 => x"75",
          4876 => x"81",
          4877 => x"87",
          4878 => x"52",
          4879 => x"51",
          4880 => x"3f",
          4881 => x"ca",
          4882 => x"9c",
          4883 => x"54",
          4884 => x"52",
          4885 => x"98",
          4886 => x"56",
          4887 => x"08",
          4888 => x"53",
          4889 => x"51",
          4890 => x"3f",
          4891 => x"ec",
          4892 => x"38",
          4893 => x"56",
          4894 => x"56",
          4895 => x"ec",
          4896 => x"75",
          4897 => x"0c",
          4898 => x"04",
          4899 => x"7d",
          4900 => x"80",
          4901 => x"05",
          4902 => x"76",
          4903 => x"38",
          4904 => x"11",
          4905 => x"53",
          4906 => x"79",
          4907 => x"3f",
          4908 => x"09",
          4909 => x"38",
          4910 => x"55",
          4911 => x"db",
          4912 => x"70",
          4913 => x"34",
          4914 => x"74",
          4915 => x"81",
          4916 => x"80",
          4917 => x"55",
          4918 => x"76",
          4919 => x"ec",
          4920 => x"3d",
          4921 => x"3d",
          4922 => x"08",
          4923 => x"57",
          4924 => x"80",
          4925 => x"39",
          4926 => x"85",
          4927 => x"80",
          4928 => x"15",
          4929 => x"33",
          4930 => x"a0",
          4931 => x"81",
          4932 => x"70",
          4933 => x"06",
          4934 => x"e6",
          4935 => x"2e",
          4936 => x"88",
          4937 => x"70",
          4938 => x"34",
          4939 => x"90",
          4940 => x"f0",
          4941 => x"53",
          4942 => x"54",
          4943 => x"3f",
          4944 => x"08",
          4945 => x"14",
          4946 => x"81",
          4947 => x"38",
          4948 => x"81",
          4949 => x"53",
          4950 => x"d2",
          4951 => x"72",
          4952 => x"0c",
          4953 => x"04",
          4954 => x"73",
          4955 => x"26",
          4956 => x"71",
          4957 => x"d5",
          4958 => x"71",
          4959 => x"de",
          4960 => x"80",
          4961 => x"88",
          4962 => x"39",
          4963 => x"51",
          4964 => x"81",
          4965 => x"80",
          4966 => x"df",
          4967 => x"e4",
          4968 => x"d0",
          4969 => x"39",
          4970 => x"51",
          4971 => x"81",
          4972 => x"80",
          4973 => x"e0",
          4974 => x"c8",
          4975 => x"a4",
          4976 => x"39",
          4977 => x"51",
          4978 => x"e0",
          4979 => x"39",
          4980 => x"51",
          4981 => x"e1",
          4982 => x"39",
          4983 => x"51",
          4984 => x"e1",
          4985 => x"39",
          4986 => x"51",
          4987 => x"e1",
          4988 => x"39",
          4989 => x"51",
          4990 => x"e2",
          4991 => x"39",
          4992 => x"51",
          4993 => x"3f",
          4994 => x"04",
          4995 => x"77",
          4996 => x"74",
          4997 => x"8a",
          4998 => x"75",
          4999 => x"51",
          5000 => x"e8",
          5001 => x"fe",
          5002 => x"81",
          5003 => x"52",
          5004 => x"ed",
          5005 => x"ec",
          5006 => x"79",
          5007 => x"81",
          5008 => x"ff",
          5009 => x"87",
          5010 => x"ec",
          5011 => x"02",
          5012 => x"e3",
          5013 => x"57",
          5014 => x"30",
          5015 => x"73",
          5016 => x"59",
          5017 => x"77",
          5018 => x"83",
          5019 => x"74",
          5020 => x"81",
          5021 => x"55",
          5022 => x"80",
          5023 => x"53",
          5024 => x"3d",
          5025 => x"c1",
          5026 => x"ec",
          5027 => x"81",
          5028 => x"b8",
          5029 => x"e0",
          5030 => x"98",
          5031 => x"ec",
          5032 => x"96",
          5033 => x"54",
          5034 => x"77",
          5035 => x"c5",
          5036 => x"ec",
          5037 => x"81",
          5038 => x"90",
          5039 => x"74",
          5040 => x"38",
          5041 => x"19",
          5042 => x"39",
          5043 => x"05",
          5044 => x"3f",
          5045 => x"78",
          5046 => x"7b",
          5047 => x"2a",
          5048 => x"57",
          5049 => x"80",
          5050 => x"81",
          5051 => x"87",
          5052 => x"08",
          5053 => x"fe",
          5054 => x"56",
          5055 => x"e0",
          5056 => x"0d",
          5057 => x"0d",
          5058 => x"05",
          5059 => x"57",
          5060 => x"80",
          5061 => x"79",
          5062 => x"3f",
          5063 => x"08",
          5064 => x"80",
          5065 => x"75",
          5066 => x"38",
          5067 => x"55",
          5068 => x"ec",
          5069 => x"52",
          5070 => x"2d",
          5071 => x"08",
          5072 => x"77",
          5073 => x"ec",
          5074 => x"3d",
          5075 => x"3d",
          5076 => x"63",
          5077 => x"80",
          5078 => x"73",
          5079 => x"41",
          5080 => x"5e",
          5081 => x"52",
          5082 => x"51",
          5083 => x"3f",
          5084 => x"51",
          5085 => x"3f",
          5086 => x"79",
          5087 => x"38",
          5088 => x"89",
          5089 => x"2e",
          5090 => x"c6",
          5091 => x"53",
          5092 => x"8e",
          5093 => x"52",
          5094 => x"51",
          5095 => x"3f",
          5096 => x"e3",
          5097 => x"82",
          5098 => x"15",
          5099 => x"39",
          5100 => x"72",
          5101 => x"38",
          5102 => x"81",
          5103 => x"ff",
          5104 => x"89",
          5105 => x"84",
          5106 => x"da",
          5107 => x"55",
          5108 => x"18",
          5109 => x"27",
          5110 => x"33",
          5111 => x"90",
          5112 => x"a6",
          5113 => x"81",
          5114 => x"ff",
          5115 => x"81",
          5116 => x"51",
          5117 => x"3f",
          5118 => x"81",
          5119 => x"ff",
          5120 => x"80",
          5121 => x"27",
          5122 => x"18",
          5123 => x"53",
          5124 => x"7a",
          5125 => x"81",
          5126 => x"9f",
          5127 => x"38",
          5128 => x"73",
          5129 => x"ff",
          5130 => x"72",
          5131 => x"38",
          5132 => x"26",
          5133 => x"51",
          5134 => x"51",
          5135 => x"3f",
          5136 => x"c1",
          5137 => x"a0",
          5138 => x"da",
          5139 => x"79",
          5140 => x"fe",
          5141 => x"81",
          5142 => x"98",
          5143 => x"2c",
          5144 => x"a0",
          5145 => x"06",
          5146 => x"f6",
          5147 => x"ec",
          5148 => x"2b",
          5149 => x"70",
          5150 => x"30",
          5151 => x"70",
          5152 => x"07",
          5153 => x"06",
          5154 => x"59",
          5155 => x"80",
          5156 => x"38",
          5157 => x"09",
          5158 => x"38",
          5159 => x"39",
          5160 => x"72",
          5161 => x"be",
          5162 => x"72",
          5163 => x"0c",
          5164 => x"04",
          5165 => x"02",
          5166 => x"81",
          5167 => x"81",
          5168 => x"55",
          5169 => x"3f",
          5170 => x"22",
          5171 => x"9d",
          5172 => x"b4",
          5173 => x"c0",
          5174 => x"c1",
          5175 => x"e3",
          5176 => x"86",
          5177 => x"80",
          5178 => x"fe",
          5179 => x"86",
          5180 => x"fe",
          5181 => x"c0",
          5182 => x"53",
          5183 => x"3f",
          5184 => x"f1",
          5185 => x"e3",
          5186 => x"f3",
          5187 => x"51",
          5188 => x"3f",
          5189 => x"70",
          5190 => x"52",
          5191 => x"95",
          5192 => x"fe",
          5193 => x"81",
          5194 => x"fe",
          5195 => x"80",
          5196 => x"92",
          5197 => x"2a",
          5198 => x"51",
          5199 => x"2e",
          5200 => x"51",
          5201 => x"3f",
          5202 => x"51",
          5203 => x"3f",
          5204 => x"f0",
          5205 => x"83",
          5206 => x"06",
          5207 => x"80",
          5208 => x"81",
          5209 => x"de",
          5210 => x"a0",
          5211 => x"d6",
          5212 => x"fe",
          5213 => x"72",
          5214 => x"81",
          5215 => x"71",
          5216 => x"38",
          5217 => x"f0",
          5218 => x"e4",
          5219 => x"f2",
          5220 => x"51",
          5221 => x"3f",
          5222 => x"70",
          5223 => x"52",
          5224 => x"95",
          5225 => x"fe",
          5226 => x"81",
          5227 => x"fe",
          5228 => x"80",
          5229 => x"8e",
          5230 => x"2a",
          5231 => x"51",
          5232 => x"2e",
          5233 => x"51",
          5234 => x"3f",
          5235 => x"51",
          5236 => x"3f",
          5237 => x"ef",
          5238 => x"87",
          5239 => x"06",
          5240 => x"80",
          5241 => x"81",
          5242 => x"da",
          5243 => x"f0",
          5244 => x"d2",
          5245 => x"fe",
          5246 => x"72",
          5247 => x"81",
          5248 => x"71",
          5249 => x"38",
          5250 => x"ef",
          5251 => x"e5",
          5252 => x"f1",
          5253 => x"51",
          5254 => x"3f",
          5255 => x"3f",
          5256 => x"04",
          5257 => x"77",
          5258 => x"56",
          5259 => x"75",
          5260 => x"f0",
          5261 => x"ec",
          5262 => x"a7",
          5263 => x"81",
          5264 => x"82",
          5265 => x"ff",
          5266 => x"81",
          5267 => x"30",
          5268 => x"e0",
          5269 => x"25",
          5270 => x"51",
          5271 => x"81",
          5272 => x"81",
          5273 => x"54",
          5274 => x"09",
          5275 => x"38",
          5276 => x"53",
          5277 => x"51",
          5278 => x"81",
          5279 => x"80",
          5280 => x"81",
          5281 => x"51",
          5282 => x"3f",
          5283 => x"83",
          5284 => x"83",
          5285 => x"81",
          5286 => x"81",
          5287 => x"54",
          5288 => x"09",
          5289 => x"38",
          5290 => x"51",
          5291 => x"3f",
          5292 => x"ec",
          5293 => x"3d",
          5294 => x"3d",
          5295 => x"71",
          5296 => x"0c",
          5297 => x"52",
          5298 => x"88",
          5299 => x"ec",
          5300 => x"ff",
          5301 => x"7d",
          5302 => x"06",
          5303 => x"e5",
          5304 => x"3d",
          5305 => x"ff",
          5306 => x"7c",
          5307 => x"81",
          5308 => x"ff",
          5309 => x"81",
          5310 => x"7d",
          5311 => x"81",
          5312 => x"8d",
          5313 => x"70",
          5314 => x"e6",
          5315 => x"fc",
          5316 => x"3d",
          5317 => x"80",
          5318 => x"51",
          5319 => x"b4",
          5320 => x"05",
          5321 => x"3f",
          5322 => x"08",
          5323 => x"90",
          5324 => x"78",
          5325 => x"87",
          5326 => x"80",
          5327 => x"38",
          5328 => x"81",
          5329 => x"bd",
          5330 => x"78",
          5331 => x"ba",
          5332 => x"2e",
          5333 => x"8a",
          5334 => x"80",
          5335 => x"a1",
          5336 => x"c0",
          5337 => x"38",
          5338 => x"82",
          5339 => x"d2",
          5340 => x"f9",
          5341 => x"38",
          5342 => x"24",
          5343 => x"80",
          5344 => x"98",
          5345 => x"f8",
          5346 => x"38",
          5347 => x"78",
          5348 => x"8a",
          5349 => x"81",
          5350 => x"38",
          5351 => x"2e",
          5352 => x"8a",
          5353 => x"81",
          5354 => x"8f",
          5355 => x"39",
          5356 => x"80",
          5357 => x"84",
          5358 => x"82",
          5359 => x"ec",
          5360 => x"2e",
          5361 => x"b4",
          5362 => x"11",
          5363 => x"05",
          5364 => x"ab",
          5365 => x"e0",
          5366 => x"fe",
          5367 => x"3d",
          5368 => x"53",
          5369 => x"51",
          5370 => x"3f",
          5371 => x"08",
          5372 => x"ec",
          5373 => x"81",
          5374 => x"fe",
          5375 => x"63",
          5376 => x"79",
          5377 => x"f2",
          5378 => x"78",
          5379 => x"05",
          5380 => x"7a",
          5381 => x"81",
          5382 => x"3d",
          5383 => x"53",
          5384 => x"51",
          5385 => x"3f",
          5386 => x"08",
          5387 => x"da",
          5388 => x"fe",
          5389 => x"ff",
          5390 => x"ff",
          5391 => x"81",
          5392 => x"80",
          5393 => x"38",
          5394 => x"f8",
          5395 => x"84",
          5396 => x"81",
          5397 => x"ec",
          5398 => x"2e",
          5399 => x"81",
          5400 => x"fe",
          5401 => x"63",
          5402 => x"27",
          5403 => x"61",
          5404 => x"81",
          5405 => x"79",
          5406 => x"05",
          5407 => x"b4",
          5408 => x"11",
          5409 => x"05",
          5410 => x"f3",
          5411 => x"e0",
          5412 => x"fc",
          5413 => x"3d",
          5414 => x"53",
          5415 => x"51",
          5416 => x"3f",
          5417 => x"08",
          5418 => x"de",
          5419 => x"fe",
          5420 => x"ff",
          5421 => x"ff",
          5422 => x"81",
          5423 => x"80",
          5424 => x"38",
          5425 => x"51",
          5426 => x"3f",
          5427 => x"63",
          5428 => x"61",
          5429 => x"33",
          5430 => x"78",
          5431 => x"38",
          5432 => x"54",
          5433 => x"79",
          5434 => x"c0",
          5435 => x"9a",
          5436 => x"62",
          5437 => x"5a",
          5438 => x"e6",
          5439 => x"bd",
          5440 => x"ff",
          5441 => x"ff",
          5442 => x"fe",
          5443 => x"81",
          5444 => x"80",
          5445 => x"e9",
          5446 => x"78",
          5447 => x"38",
          5448 => x"08",
          5449 => x"39",
          5450 => x"33",
          5451 => x"2e",
          5452 => x"e9",
          5453 => x"bc",
          5454 => x"d6",
          5455 => x"80",
          5456 => x"81",
          5457 => x"44",
          5458 => x"e9",
          5459 => x"78",
          5460 => x"38",
          5461 => x"08",
          5462 => x"81",
          5463 => x"59",
          5464 => x"88",
          5465 => x"ac",
          5466 => x"39",
          5467 => x"08",
          5468 => x"44",
          5469 => x"fc",
          5470 => x"84",
          5471 => x"fe",
          5472 => x"ec",
          5473 => x"de",
          5474 => x"d4",
          5475 => x"80",
          5476 => x"81",
          5477 => x"43",
          5478 => x"81",
          5479 => x"59",
          5480 => x"88",
          5481 => x"98",
          5482 => x"39",
          5483 => x"33",
          5484 => x"2e",
          5485 => x"e9",
          5486 => x"aa",
          5487 => x"d7",
          5488 => x"80",
          5489 => x"81",
          5490 => x"43",
          5491 => x"e9",
          5492 => x"78",
          5493 => x"38",
          5494 => x"08",
          5495 => x"81",
          5496 => x"88",
          5497 => x"3d",
          5498 => x"53",
          5499 => x"51",
          5500 => x"3f",
          5501 => x"08",
          5502 => x"38",
          5503 => x"5c",
          5504 => x"83",
          5505 => x"7a",
          5506 => x"30",
          5507 => x"9f",
          5508 => x"06",
          5509 => x"5a",
          5510 => x"88",
          5511 => x"2e",
          5512 => x"42",
          5513 => x"51",
          5514 => x"3f",
          5515 => x"54",
          5516 => x"52",
          5517 => x"96",
          5518 => x"ec",
          5519 => x"e6",
          5520 => x"39",
          5521 => x"80",
          5522 => x"84",
          5523 => x"fd",
          5524 => x"ec",
          5525 => x"2e",
          5526 => x"b4",
          5527 => x"11",
          5528 => x"05",
          5529 => x"97",
          5530 => x"e0",
          5531 => x"a5",
          5532 => x"02",
          5533 => x"33",
          5534 => x"81",
          5535 => x"3d",
          5536 => x"53",
          5537 => x"51",
          5538 => x"3f",
          5539 => x"08",
          5540 => x"f6",
          5541 => x"33",
          5542 => x"e6",
          5543 => x"fa",
          5544 => x"f8",
          5545 => x"fe",
          5546 => x"79",
          5547 => x"59",
          5548 => x"f8",
          5549 => x"79",
          5550 => x"b4",
          5551 => x"11",
          5552 => x"05",
          5553 => x"b7",
          5554 => x"e0",
          5555 => x"91",
          5556 => x"02",
          5557 => x"33",
          5558 => x"81",
          5559 => x"b5",
          5560 => x"84",
          5561 => x"be",
          5562 => x"39",
          5563 => x"f4",
          5564 => x"84",
          5565 => x"fd",
          5566 => x"ec",
          5567 => x"2e",
          5568 => x"b4",
          5569 => x"11",
          5570 => x"05",
          5571 => x"e1",
          5572 => x"e0",
          5573 => x"a6",
          5574 => x"02",
          5575 => x"79",
          5576 => x"5b",
          5577 => x"b4",
          5578 => x"11",
          5579 => x"05",
          5580 => x"bd",
          5581 => x"e0",
          5582 => x"f7",
          5583 => x"70",
          5584 => x"81",
          5585 => x"fe",
          5586 => x"80",
          5587 => x"51",
          5588 => x"3f",
          5589 => x"33",
          5590 => x"2e",
          5591 => x"78",
          5592 => x"38",
          5593 => x"41",
          5594 => x"3d",
          5595 => x"53",
          5596 => x"51",
          5597 => x"3f",
          5598 => x"08",
          5599 => x"38",
          5600 => x"be",
          5601 => x"70",
          5602 => x"23",
          5603 => x"ae",
          5604 => x"84",
          5605 => x"8e",
          5606 => x"39",
          5607 => x"f4",
          5608 => x"84",
          5609 => x"fc",
          5610 => x"ec",
          5611 => x"2e",
          5612 => x"b4",
          5613 => x"11",
          5614 => x"05",
          5615 => x"b1",
          5616 => x"e0",
          5617 => x"a1",
          5618 => x"71",
          5619 => x"84",
          5620 => x"3d",
          5621 => x"53",
          5622 => x"51",
          5623 => x"3f",
          5624 => x"08",
          5625 => x"a2",
          5626 => x"08",
          5627 => x"e7",
          5628 => x"f8",
          5629 => x"f8",
          5630 => x"fe",
          5631 => x"79",
          5632 => x"59",
          5633 => x"f6",
          5634 => x"79",
          5635 => x"b4",
          5636 => x"11",
          5637 => x"05",
          5638 => x"d5",
          5639 => x"e0",
          5640 => x"8d",
          5641 => x"71",
          5642 => x"84",
          5643 => x"b9",
          5644 => x"84",
          5645 => x"ee",
          5646 => x"39",
          5647 => x"80",
          5648 => x"84",
          5649 => x"f9",
          5650 => x"ec",
          5651 => x"2e",
          5652 => x"63",
          5653 => x"a4",
          5654 => x"ae",
          5655 => x"78",
          5656 => x"ff",
          5657 => x"ff",
          5658 => x"fe",
          5659 => x"81",
          5660 => x"80",
          5661 => x"38",
          5662 => x"e7",
          5663 => x"f7",
          5664 => x"59",
          5665 => x"ec",
          5666 => x"2e",
          5667 => x"81",
          5668 => x"52",
          5669 => x"51",
          5670 => x"3f",
          5671 => x"81",
          5672 => x"fe",
          5673 => x"fe",
          5674 => x"f4",
          5675 => x"e8",
          5676 => x"f0",
          5677 => x"59",
          5678 => x"fe",
          5679 => x"f4",
          5680 => x"70",
          5681 => x"78",
          5682 => x"be",
          5683 => x"06",
          5684 => x"2e",
          5685 => x"b4",
          5686 => x"05",
          5687 => x"97",
          5688 => x"e0",
          5689 => x"5b",
          5690 => x"b2",
          5691 => x"24",
          5692 => x"81",
          5693 => x"80",
          5694 => x"83",
          5695 => x"80",
          5696 => x"e8",
          5697 => x"55",
          5698 => x"54",
          5699 => x"e8",
          5700 => x"3d",
          5701 => x"51",
          5702 => x"3f",
          5703 => x"e8",
          5704 => x"3d",
          5705 => x"51",
          5706 => x"3f",
          5707 => x"55",
          5708 => x"54",
          5709 => x"e8",
          5710 => x"3d",
          5711 => x"51",
          5712 => x"3f",
          5713 => x"54",
          5714 => x"e8",
          5715 => x"3d",
          5716 => x"51",
          5717 => x"3f",
          5718 => x"58",
          5719 => x"57",
          5720 => x"81",
          5721 => x"05",
          5722 => x"83",
          5723 => x"83",
          5724 => x"b4",
          5725 => x"05",
          5726 => x"3f",
          5727 => x"08",
          5728 => x"08",
          5729 => x"70",
          5730 => x"25",
          5731 => x"5f",
          5732 => x"83",
          5733 => x"81",
          5734 => x"06",
          5735 => x"2e",
          5736 => x"1b",
          5737 => x"06",
          5738 => x"fe",
          5739 => x"81",
          5740 => x"32",
          5741 => x"8a",
          5742 => x"2e",
          5743 => x"f2",
          5744 => x"e8",
          5745 => x"f4",
          5746 => x"be",
          5747 => x"0d",
          5748 => x"ed",
          5749 => x"c0",
          5750 => x"08",
          5751 => x"84",
          5752 => x"51",
          5753 => x"3f",
          5754 => x"08",
          5755 => x"08",
          5756 => x"84",
          5757 => x"51",
          5758 => x"3f",
          5759 => x"e0",
          5760 => x"0c",
          5761 => x"9c",
          5762 => x"55",
          5763 => x"52",
          5764 => x"d6",
          5765 => x"ec",
          5766 => x"2b",
          5767 => x"53",
          5768 => x"52",
          5769 => x"d6",
          5770 => x"81",
          5771 => x"07",
          5772 => x"80",
          5773 => x"c0",
          5774 => x"8c",
          5775 => x"87",
          5776 => x"0c",
          5777 => x"81",
          5778 => x"b6",
          5779 => x"ec",
          5780 => x"e3",
          5781 => x"ec",
          5782 => x"e8",
          5783 => x"ed",
          5784 => x"e8",
          5785 => x"ed",
          5786 => x"c1",
          5787 => x"ec",
          5788 => x"51",
          5789 => x"f0",
          5790 => x"04",
          5791 => x"20",
          5792 => x"20",
          5793 => x"20",
          5794 => x"20",
          5795 => x"20",
          5796 => x"5d",
          5797 => x"5d",
          5798 => x"5d",
          5799 => x"5d",
          5800 => x"5d",
          5801 => x"5d",
          5802 => x"5d",
          5803 => x"5d",
          5804 => x"5d",
          5805 => x"5d",
          5806 => x"5d",
          5807 => x"5d",
          5808 => x"5d",
          5809 => x"5d",
          5810 => x"5d",
          5811 => x"5d",
          5812 => x"5d",
          5813 => x"5d",
          5814 => x"5d",
          5815 => x"5d",
          5816 => x"2f",
          5817 => x"25",
          5818 => x"64",
          5819 => x"3a",
          5820 => x"25",
          5821 => x"0a",
          5822 => x"43",
          5823 => x"6e",
          5824 => x"75",
          5825 => x"69",
          5826 => x"00",
          5827 => x"66",
          5828 => x"20",
          5829 => x"20",
          5830 => x"66",
          5831 => x"00",
          5832 => x"44",
          5833 => x"63",
          5834 => x"69",
          5835 => x"65",
          5836 => x"74",
          5837 => x"0a",
          5838 => x"20",
          5839 => x"20",
          5840 => x"41",
          5841 => x"28",
          5842 => x"58",
          5843 => x"38",
          5844 => x"0a",
          5845 => x"20",
          5846 => x"52",
          5847 => x"20",
          5848 => x"28",
          5849 => x"58",
          5850 => x"38",
          5851 => x"0a",
          5852 => x"20",
          5853 => x"53",
          5854 => x"52",
          5855 => x"28",
          5856 => x"58",
          5857 => x"38",
          5858 => x"0a",
          5859 => x"20",
          5860 => x"41",
          5861 => x"20",
          5862 => x"28",
          5863 => x"58",
          5864 => x"38",
          5865 => x"0a",
          5866 => x"20",
          5867 => x"4d",
          5868 => x"20",
          5869 => x"28",
          5870 => x"58",
          5871 => x"38",
          5872 => x"0a",
          5873 => x"20",
          5874 => x"20",
          5875 => x"44",
          5876 => x"28",
          5877 => x"69",
          5878 => x"20",
          5879 => x"32",
          5880 => x"0a",
          5881 => x"20",
          5882 => x"4d",
          5883 => x"20",
          5884 => x"28",
          5885 => x"65",
          5886 => x"20",
          5887 => x"32",
          5888 => x"0a",
          5889 => x"20",
          5890 => x"54",
          5891 => x"54",
          5892 => x"28",
          5893 => x"6e",
          5894 => x"73",
          5895 => x"32",
          5896 => x"0a",
          5897 => x"20",
          5898 => x"53",
          5899 => x"4e",
          5900 => x"55",
          5901 => x"00",
          5902 => x"20",
          5903 => x"20",
          5904 => x"0a",
          5905 => x"20",
          5906 => x"43",
          5907 => x"00",
          5908 => x"20",
          5909 => x"32",
          5910 => x"00",
          5911 => x"20",
          5912 => x"49",
          5913 => x"00",
          5914 => x"64",
          5915 => x"73",
          5916 => x"0a",
          5917 => x"20",
          5918 => x"55",
          5919 => x"73",
          5920 => x"56",
          5921 => x"6f",
          5922 => x"64",
          5923 => x"73",
          5924 => x"20",
          5925 => x"58",
          5926 => x"00",
          5927 => x"20",
          5928 => x"55",
          5929 => x"6d",
          5930 => x"20",
          5931 => x"72",
          5932 => x"64",
          5933 => x"73",
          5934 => x"20",
          5935 => x"58",
          5936 => x"00",
          5937 => x"20",
          5938 => x"61",
          5939 => x"53",
          5940 => x"74",
          5941 => x"64",
          5942 => x"73",
          5943 => x"20",
          5944 => x"20",
          5945 => x"58",
          5946 => x"00",
          5947 => x"73",
          5948 => x"00",
          5949 => x"20",
          5950 => x"55",
          5951 => x"20",
          5952 => x"20",
          5953 => x"20",
          5954 => x"20",
          5955 => x"20",
          5956 => x"20",
          5957 => x"58",
          5958 => x"00",
          5959 => x"20",
          5960 => x"73",
          5961 => x"20",
          5962 => x"63",
          5963 => x"72",
          5964 => x"20",
          5965 => x"20",
          5966 => x"20",
          5967 => x"25",
          5968 => x"4d",
          5969 => x"00",
          5970 => x"20",
          5971 => x"52",
          5972 => x"43",
          5973 => x"6b",
          5974 => x"65",
          5975 => x"20",
          5976 => x"20",
          5977 => x"20",
          5978 => x"25",
          5979 => x"4d",
          5980 => x"00",
          5981 => x"20",
          5982 => x"73",
          5983 => x"6e",
          5984 => x"44",
          5985 => x"20",
          5986 => x"63",
          5987 => x"72",
          5988 => x"20",
          5989 => x"25",
          5990 => x"4d",
          5991 => x"00",
          5992 => x"61",
          5993 => x"00",
          5994 => x"64",
          5995 => x"00",
          5996 => x"65",
          5997 => x"00",
          5998 => x"4f",
          5999 => x"4f",
          6000 => x"00",
          6001 => x"6b",
          6002 => x"6e",
          6003 => x"00",
          6004 => x"2b",
          6005 => x"3c",
          6006 => x"5b",
          6007 => x"00",
          6008 => x"54",
          6009 => x"54",
          6010 => x"00",
          6011 => x"90",
          6012 => x"4f",
          6013 => x"30",
          6014 => x"20",
          6015 => x"45",
          6016 => x"20",
          6017 => x"33",
          6018 => x"20",
          6019 => x"20",
          6020 => x"45",
          6021 => x"20",
          6022 => x"20",
          6023 => x"20",
          6024 => x"6d",
          6025 => x"00",
          6026 => x"00",
          6027 => x"00",
          6028 => x"45",
          6029 => x"8f",
          6030 => x"45",
          6031 => x"8e",
          6032 => x"92",
          6033 => x"55",
          6034 => x"9a",
          6035 => x"9e",
          6036 => x"4f",
          6037 => x"a6",
          6038 => x"aa",
          6039 => x"ae",
          6040 => x"b2",
          6041 => x"b6",
          6042 => x"ba",
          6043 => x"be",
          6044 => x"c2",
          6045 => x"c6",
          6046 => x"ca",
          6047 => x"ce",
          6048 => x"d2",
          6049 => x"d6",
          6050 => x"da",
          6051 => x"de",
          6052 => x"e2",
          6053 => x"e6",
          6054 => x"ea",
          6055 => x"ee",
          6056 => x"f2",
          6057 => x"f6",
          6058 => x"fa",
          6059 => x"fe",
          6060 => x"2c",
          6061 => x"5d",
          6062 => x"2a",
          6063 => x"3f",
          6064 => x"00",
          6065 => x"00",
          6066 => x"00",
          6067 => x"02",
          6068 => x"00",
          6069 => x"00",
          6070 => x"00",
          6071 => x"00",
          6072 => x"00",
          6073 => x"6e",
          6074 => x"00",
          6075 => x"6f",
          6076 => x"00",
          6077 => x"6e",
          6078 => x"00",
          6079 => x"6f",
          6080 => x"00",
          6081 => x"78",
          6082 => x"00",
          6083 => x"6c",
          6084 => x"00",
          6085 => x"6f",
          6086 => x"00",
          6087 => x"69",
          6088 => x"00",
          6089 => x"75",
          6090 => x"00",
          6091 => x"62",
          6092 => x"68",
          6093 => x"77",
          6094 => x"64",
          6095 => x"65",
          6096 => x"64",
          6097 => x"65",
          6098 => x"6c",
          6099 => x"00",
          6100 => x"70",
          6101 => x"73",
          6102 => x"74",
          6103 => x"73",
          6104 => x"00",
          6105 => x"66",
          6106 => x"00",
          6107 => x"73",
          6108 => x"00",
          6109 => x"61",
          6110 => x"00",
          6111 => x"73",
          6112 => x"72",
          6113 => x"0a",
          6114 => x"74",
          6115 => x"61",
          6116 => x"72",
          6117 => x"2e",
          6118 => x"00",
          6119 => x"73",
          6120 => x"6f",
          6121 => x"65",
          6122 => x"2e",
          6123 => x"00",
          6124 => x"20",
          6125 => x"65",
          6126 => x"75",
          6127 => x"0a",
          6128 => x"20",
          6129 => x"68",
          6130 => x"75",
          6131 => x"0a",
          6132 => x"76",
          6133 => x"64",
          6134 => x"6c",
          6135 => x"6d",
          6136 => x"00",
          6137 => x"63",
          6138 => x"20",
          6139 => x"69",
          6140 => x"0a",
          6141 => x"6c",
          6142 => x"6c",
          6143 => x"64",
          6144 => x"78",
          6145 => x"73",
          6146 => x"00",
          6147 => x"6c",
          6148 => x"61",
          6149 => x"65",
          6150 => x"76",
          6151 => x"64",
          6152 => x"00",
          6153 => x"20",
          6154 => x"77",
          6155 => x"65",
          6156 => x"6f",
          6157 => x"74",
          6158 => x"0a",
          6159 => x"69",
          6160 => x"6e",
          6161 => x"65",
          6162 => x"73",
          6163 => x"76",
          6164 => x"64",
          6165 => x"00",
          6166 => x"73",
          6167 => x"6f",
          6168 => x"6e",
          6169 => x"65",
          6170 => x"00",
          6171 => x"20",
          6172 => x"70",
          6173 => x"62",
          6174 => x"66",
          6175 => x"73",
          6176 => x"65",
          6177 => x"6f",
          6178 => x"20",
          6179 => x"64",
          6180 => x"2e",
          6181 => x"00",
          6182 => x"72",
          6183 => x"20",
          6184 => x"72",
          6185 => x"2e",
          6186 => x"00",
          6187 => x"6d",
          6188 => x"74",
          6189 => x"70",
          6190 => x"74",
          6191 => x"20",
          6192 => x"63",
          6193 => x"65",
          6194 => x"00",
          6195 => x"6c",
          6196 => x"73",
          6197 => x"63",
          6198 => x"2e",
          6199 => x"00",
          6200 => x"73",
          6201 => x"69",
          6202 => x"6e",
          6203 => x"65",
          6204 => x"79",
          6205 => x"00",
          6206 => x"6f",
          6207 => x"6e",
          6208 => x"70",
          6209 => x"66",
          6210 => x"73",
          6211 => x"00",
          6212 => x"72",
          6213 => x"74",
          6214 => x"20",
          6215 => x"6f",
          6216 => x"63",
          6217 => x"00",
          6218 => x"63",
          6219 => x"73",
          6220 => x"00",
          6221 => x"6b",
          6222 => x"6e",
          6223 => x"72",
          6224 => x"0a",
          6225 => x"6c",
          6226 => x"79",
          6227 => x"20",
          6228 => x"61",
          6229 => x"6c",
          6230 => x"79",
          6231 => x"2f",
          6232 => x"2e",
          6233 => x"00",
          6234 => x"61",
          6235 => x"00",
          6236 => x"38",
          6237 => x"00",
          6238 => x"20",
          6239 => x"34",
          6240 => x"00",
          6241 => x"20",
          6242 => x"20",
          6243 => x"00",
          6244 => x"32",
          6245 => x"00",
          6246 => x"00",
          6247 => x"00",
          6248 => x"0a",
          6249 => x"53",
          6250 => x"2a",
          6251 => x"20",
          6252 => x"00",
          6253 => x"2f",
          6254 => x"32",
          6255 => x"00",
          6256 => x"2e",
          6257 => x"00",
          6258 => x"50",
          6259 => x"72",
          6260 => x"25",
          6261 => x"29",
          6262 => x"20",
          6263 => x"2a",
          6264 => x"00",
          6265 => x"55",
          6266 => x"74",
          6267 => x"75",
          6268 => x"48",
          6269 => x"6c",
          6270 => x"00",
          6271 => x"6d",
          6272 => x"69",
          6273 => x"72",
          6274 => x"74",
          6275 => x"00",
          6276 => x"32",
          6277 => x"74",
          6278 => x"75",
          6279 => x"00",
          6280 => x"43",
          6281 => x"52",
          6282 => x"6e",
          6283 => x"72",
          6284 => x"0a",
          6285 => x"43",
          6286 => x"57",
          6287 => x"6e",
          6288 => x"72",
          6289 => x"0a",
          6290 => x"52",
          6291 => x"52",
          6292 => x"6e",
          6293 => x"72",
          6294 => x"0a",
          6295 => x"52",
          6296 => x"54",
          6297 => x"6e",
          6298 => x"72",
          6299 => x"0a",
          6300 => x"52",
          6301 => x"52",
          6302 => x"6e",
          6303 => x"72",
          6304 => x"0a",
          6305 => x"52",
          6306 => x"54",
          6307 => x"6e",
          6308 => x"72",
          6309 => x"0a",
          6310 => x"74",
          6311 => x"67",
          6312 => x"20",
          6313 => x"65",
          6314 => x"2e",
          6315 => x"00",
          6316 => x"61",
          6317 => x"6e",
          6318 => x"69",
          6319 => x"2e",
          6320 => x"00",
          6321 => x"74",
          6322 => x"65",
          6323 => x"61",
          6324 => x"00",
          6325 => x"00",
          6326 => x"69",
          6327 => x"20",
          6328 => x"69",
          6329 => x"69",
          6330 => x"73",
          6331 => x"64",
          6332 => x"72",
          6333 => x"2c",
          6334 => x"65",
          6335 => x"20",
          6336 => x"74",
          6337 => x"6e",
          6338 => x"6c",
          6339 => x"00",
          6340 => x"00",
          6341 => x"65",
          6342 => x"6e",
          6343 => x"2e",
          6344 => x"00",
          6345 => x"70",
          6346 => x"67",
          6347 => x"00",
          6348 => x"6d",
          6349 => x"69",
          6350 => x"2e",
          6351 => x"00",
          6352 => x"38",
          6353 => x"25",
          6354 => x"29",
          6355 => x"30",
          6356 => x"28",
          6357 => x"78",
          6358 => x"00",
          6359 => x"6d",
          6360 => x"65",
          6361 => x"79",
          6362 => x"00",
          6363 => x"6f",
          6364 => x"65",
          6365 => x"0a",
          6366 => x"38",
          6367 => x"30",
          6368 => x"00",
          6369 => x"3f",
          6370 => x"00",
          6371 => x"38",
          6372 => x"30",
          6373 => x"00",
          6374 => x"38",
          6375 => x"30",
          6376 => x"00",
          6377 => x"65",
          6378 => x"69",
          6379 => x"63",
          6380 => x"20",
          6381 => x"30",
          6382 => x"2e",
          6383 => x"00",
          6384 => x"6c",
          6385 => x"67",
          6386 => x"64",
          6387 => x"20",
          6388 => x"78",
          6389 => x"2e",
          6390 => x"00",
          6391 => x"6c",
          6392 => x"65",
          6393 => x"6e",
          6394 => x"63",
          6395 => x"20",
          6396 => x"29",
          6397 => x"00",
          6398 => x"73",
          6399 => x"74",
          6400 => x"20",
          6401 => x"6c",
          6402 => x"74",
          6403 => x"2e",
          6404 => x"00",
          6405 => x"6c",
          6406 => x"65",
          6407 => x"74",
          6408 => x"2e",
          6409 => x"00",
          6410 => x"55",
          6411 => x"6e",
          6412 => x"3a",
          6413 => x"5c",
          6414 => x"25",
          6415 => x"00",
          6416 => x"3a",
          6417 => x"5c",
          6418 => x"00",
          6419 => x"3a",
          6420 => x"00",
          6421 => x"64",
          6422 => x"6d",
          6423 => x"64",
          6424 => x"00",
          6425 => x"6e",
          6426 => x"67",
          6427 => x"0a",
          6428 => x"61",
          6429 => x"6e",
          6430 => x"6e",
          6431 => x"72",
          6432 => x"73",
          6433 => x"0a",
          6434 => x"00",
          6435 => x"00",
          6436 => x"7f",
          6437 => x"00",
          6438 => x"7f",
          6439 => x"00",
          6440 => x"7f",
          6441 => x"00",
          6442 => x"00",
          6443 => x"00",
          6444 => x"ff",
          6445 => x"00",
          6446 => x"00",
          6447 => x"78",
          6448 => x"00",
          6449 => x"e1",
          6450 => x"e1",
          6451 => x"e1",
          6452 => x"00",
          6453 => x"01",
          6454 => x"01",
          6455 => x"10",
          6456 => x"00",
          6457 => x"00",
          6458 => x"00",
          6459 => x"00",
          6460 => x"6e",
          6461 => x"01",
          6462 => x"00",
          6463 => x"00",
          6464 => x"6e",
          6465 => x"01",
          6466 => x"00",
          6467 => x"00",
          6468 => x"6e",
          6469 => x"03",
          6470 => x"00",
          6471 => x"00",
          6472 => x"6e",
          6473 => x"03",
          6474 => x"00",
          6475 => x"00",
          6476 => x"6f",
          6477 => x"03",
          6478 => x"00",
          6479 => x"00",
          6480 => x"6f",
          6481 => x"04",
          6482 => x"00",
          6483 => x"00",
          6484 => x"6f",
          6485 => x"04",
          6486 => x"00",
          6487 => x"00",
          6488 => x"6f",
          6489 => x"04",
          6490 => x"00",
          6491 => x"00",
          6492 => x"6f",
          6493 => x"04",
          6494 => x"00",
          6495 => x"00",
          6496 => x"6f",
          6497 => x"04",
          6498 => x"00",
          6499 => x"00",
          6500 => x"6f",
          6501 => x"04",
          6502 => x"00",
          6503 => x"00",
          6504 => x"6f",
          6505 => x"04",
          6506 => x"00",
          6507 => x"00",
          6508 => x"6f",
          6509 => x"05",
          6510 => x"00",
          6511 => x"00",
          6512 => x"6f",
          6513 => x"05",
          6514 => x"00",
          6515 => x"00",
          6516 => x"6f",
          6517 => x"05",
          6518 => x"00",
          6519 => x"00",
          6520 => x"6f",
          6521 => x"05",
          6522 => x"00",
          6523 => x"00",
          6524 => x"6f",
          6525 => x"07",
          6526 => x"00",
          6527 => x"00",
          6528 => x"6f",
          6529 => x"07",
          6530 => x"00",
          6531 => x"00",
          6532 => x"6f",
          6533 => x"08",
          6534 => x"00",
          6535 => x"00",
          6536 => x"6f",
          6537 => x"08",
          6538 => x"00",
          6539 => x"00",
          6540 => x"6f",
          6541 => x"08",
          6542 => x"00",
          6543 => x"00",
          6544 => x"6f",
          6545 => x"08",
          6546 => x"00",
          6547 => x"00",
          6548 => x"6f",
          6549 => x"09",
          6550 => x"00",
          6551 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"aa",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"04",
            10 => x"a4",
            11 => x"0b",
            12 => x"04",
            13 => x"a4",
            14 => x"0b",
            15 => x"04",
            16 => x"a4",
            17 => x"0b",
            18 => x"04",
            19 => x"a4",
            20 => x"0b",
            21 => x"04",
            22 => x"a5",
            23 => x"0b",
            24 => x"04",
            25 => x"a5",
            26 => x"0b",
            27 => x"04",
            28 => x"a5",
            29 => x"0b",
            30 => x"04",
            31 => x"a5",
            32 => x"0b",
            33 => x"04",
            34 => x"a5",
            35 => x"0b",
            36 => x"04",
            37 => x"a6",
            38 => x"0b",
            39 => x"04",
            40 => x"a6",
            41 => x"0b",
            42 => x"04",
            43 => x"a6",
            44 => x"0b",
            45 => x"04",
            46 => x"a6",
            47 => x"0b",
            48 => x"04",
            49 => x"a7",
            50 => x"0b",
            51 => x"04",
            52 => x"a7",
            53 => x"0b",
            54 => x"04",
            55 => x"a7",
            56 => x"0b",
            57 => x"04",
            58 => x"a7",
            59 => x"0b",
            60 => x"04",
            61 => x"a8",
            62 => x"0b",
            63 => x"04",
            64 => x"a8",
            65 => x"0b",
            66 => x"04",
            67 => x"a8",
            68 => x"0b",
            69 => x"04",
            70 => x"a8",
            71 => x"0b",
            72 => x"04",
            73 => x"a9",
            74 => x"0b",
            75 => x"04",
            76 => x"a9",
            77 => x"0b",
            78 => x"04",
            79 => x"a9",
            80 => x"0b",
            81 => x"04",
            82 => x"a9",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"a4",
           129 => x"ec",
           130 => x"d3",
           131 => x"ec",
           132 => x"90",
           133 => x"ec",
           134 => x"c8",
           135 => x"ec",
           136 => x"90",
           137 => x"ec",
           138 => x"87",
           139 => x"ec",
           140 => x"90",
           141 => x"ec",
           142 => x"a5",
           143 => x"ec",
           144 => x"90",
           145 => x"ec",
           146 => x"e3",
           147 => x"ec",
           148 => x"90",
           149 => x"ec",
           150 => x"e1",
           151 => x"ec",
           152 => x"90",
           153 => x"ec",
           154 => x"c8",
           155 => x"ec",
           156 => x"90",
           157 => x"ec",
           158 => x"fe",
           159 => x"ec",
           160 => x"90",
           161 => x"ec",
           162 => x"f0",
           163 => x"ec",
           164 => x"90",
           165 => x"ec",
           166 => x"89",
           167 => x"ec",
           168 => x"90",
           169 => x"ec",
           170 => x"9f",
           171 => x"ec",
           172 => x"90",
           173 => x"ec",
           174 => x"c3",
           175 => x"ec",
           176 => x"90",
           177 => x"ec",
           178 => x"2d",
           179 => x"08",
           180 => x"04",
           181 => x"0c",
           182 => x"81",
           183 => x"83",
           184 => x"81",
           185 => x"af",
           186 => x"ec",
           187 => x"80",
           188 => x"ec",
           189 => x"82",
           190 => x"ec",
           191 => x"90",
           192 => x"ec",
           193 => x"2d",
           194 => x"08",
           195 => x"04",
           196 => x"0c",
           197 => x"2d",
           198 => x"08",
           199 => x"04",
           200 => x"0c",
           201 => x"2d",
           202 => x"08",
           203 => x"04",
           204 => x"0c",
           205 => x"2d",
           206 => x"08",
           207 => x"04",
           208 => x"0c",
           209 => x"2d",
           210 => x"08",
           211 => x"04",
           212 => x"0c",
           213 => x"2d",
           214 => x"08",
           215 => x"04",
           216 => x"0c",
           217 => x"2d",
           218 => x"08",
           219 => x"04",
           220 => x"0c",
           221 => x"2d",
           222 => x"08",
           223 => x"04",
           224 => x"0c",
           225 => x"2d",
           226 => x"08",
           227 => x"04",
           228 => x"0c",
           229 => x"2d",
           230 => x"08",
           231 => x"04",
           232 => x"0c",
           233 => x"2d",
           234 => x"08",
           235 => x"04",
           236 => x"0c",
           237 => x"2d",
           238 => x"08",
           239 => x"04",
           240 => x"0c",
           241 => x"2d",
           242 => x"08",
           243 => x"04",
           244 => x"0c",
           245 => x"2d",
           246 => x"08",
           247 => x"04",
           248 => x"0c",
           249 => x"2d",
           250 => x"08",
           251 => x"04",
           252 => x"0c",
           253 => x"2d",
           254 => x"08",
           255 => x"04",
           256 => x"0c",
           257 => x"2d",
           258 => x"08",
           259 => x"04",
           260 => x"0c",
           261 => x"2d",
           262 => x"08",
           263 => x"04",
           264 => x"0c",
           265 => x"2d",
           266 => x"08",
           267 => x"04",
           268 => x"0c",
           269 => x"2d",
           270 => x"08",
           271 => x"04",
           272 => x"0c",
           273 => x"2d",
           274 => x"08",
           275 => x"04",
           276 => x"0c",
           277 => x"2d",
           278 => x"08",
           279 => x"04",
           280 => x"0c",
           281 => x"2d",
           282 => x"08",
           283 => x"04",
           284 => x"0c",
           285 => x"2d",
           286 => x"08",
           287 => x"04",
           288 => x"0c",
           289 => x"2d",
           290 => x"08",
           291 => x"04",
           292 => x"0c",
           293 => x"2d",
           294 => x"08",
           295 => x"04",
           296 => x"0c",
           297 => x"2d",
           298 => x"08",
           299 => x"04",
           300 => x"0c",
           301 => x"2d",
           302 => x"08",
           303 => x"04",
           304 => x"0c",
           305 => x"2d",
           306 => x"08",
           307 => x"04",
           308 => x"0c",
           309 => x"81",
           310 => x"83",
           311 => x"81",
           312 => x"b0",
           313 => x"ec",
           314 => x"80",
           315 => x"ec",
           316 => x"c5",
           317 => x"ec",
           318 => x"90",
           319 => x"ec",
           320 => x"e7",
           321 => x"ec",
           322 => x"90",
           323 => x"e0",
           324 => x"8c",
           325 => x"80",
           326 => x"05",
           327 => x"0b",
           328 => x"04",
           329 => x"81",
           330 => x"3c",
           331 => x"ec",
           332 => x"ec",
           333 => x"3d",
           334 => x"81",
           335 => x"8c",
           336 => x"81",
           337 => x"88",
           338 => x"80",
           339 => x"ec",
           340 => x"81",
           341 => x"54",
           342 => x"81",
           343 => x"04",
           344 => x"08",
           345 => x"ec",
           346 => x"0d",
           347 => x"ec",
           348 => x"05",
           349 => x"ec",
           350 => x"05",
           351 => x"3f",
           352 => x"08",
           353 => x"e0",
           354 => x"3d",
           355 => x"ec",
           356 => x"ec",
           357 => x"81",
           358 => x"fd",
           359 => x"0b",
           360 => x"08",
           361 => x"80",
           362 => x"ec",
           363 => x"0c",
           364 => x"08",
           365 => x"81",
           366 => x"88",
           367 => x"b9",
           368 => x"ec",
           369 => x"08",
           370 => x"38",
           371 => x"ec",
           372 => x"05",
           373 => x"38",
           374 => x"08",
           375 => x"10",
           376 => x"08",
           377 => x"81",
           378 => x"fc",
           379 => x"81",
           380 => x"fc",
           381 => x"b8",
           382 => x"ec",
           383 => x"08",
           384 => x"e1",
           385 => x"ec",
           386 => x"08",
           387 => x"08",
           388 => x"26",
           389 => x"ec",
           390 => x"05",
           391 => x"ec",
           392 => x"08",
           393 => x"ec",
           394 => x"0c",
           395 => x"08",
           396 => x"81",
           397 => x"fc",
           398 => x"81",
           399 => x"f8",
           400 => x"ec",
           401 => x"05",
           402 => x"81",
           403 => x"fc",
           404 => x"ec",
           405 => x"05",
           406 => x"81",
           407 => x"8c",
           408 => x"95",
           409 => x"ec",
           410 => x"08",
           411 => x"38",
           412 => x"08",
           413 => x"70",
           414 => x"08",
           415 => x"51",
           416 => x"ec",
           417 => x"05",
           418 => x"ec",
           419 => x"05",
           420 => x"ec",
           421 => x"05",
           422 => x"e0",
           423 => x"0d",
           424 => x"0c",
           425 => x"0d",
           426 => x"02",
           427 => x"05",
           428 => x"53",
           429 => x"27",
           430 => x"83",
           431 => x"80",
           432 => x"ff",
           433 => x"ff",
           434 => x"73",
           435 => x"05",
           436 => x"12",
           437 => x"2e",
           438 => x"ef",
           439 => x"ec",
           440 => x"3d",
           441 => x"74",
           442 => x"07",
           443 => x"2b",
           444 => x"51",
           445 => x"a5",
           446 => x"70",
           447 => x"0c",
           448 => x"84",
           449 => x"72",
           450 => x"05",
           451 => x"71",
           452 => x"53",
           453 => x"52",
           454 => x"dd",
           455 => x"27",
           456 => x"71",
           457 => x"53",
           458 => x"52",
           459 => x"f2",
           460 => x"ff",
           461 => x"3d",
           462 => x"70",
           463 => x"06",
           464 => x"70",
           465 => x"73",
           466 => x"56",
           467 => x"08",
           468 => x"38",
           469 => x"52",
           470 => x"81",
           471 => x"54",
           472 => x"9d",
           473 => x"55",
           474 => x"09",
           475 => x"38",
           476 => x"14",
           477 => x"81",
           478 => x"56",
           479 => x"e5",
           480 => x"55",
           481 => x"06",
           482 => x"06",
           483 => x"81",
           484 => x"52",
           485 => x"0d",
           486 => x"70",
           487 => x"ff",
           488 => x"f8",
           489 => x"80",
           490 => x"51",
           491 => x"84",
           492 => x"71",
           493 => x"54",
           494 => x"2e",
           495 => x"75",
           496 => x"94",
           497 => x"81",
           498 => x"87",
           499 => x"fe",
           500 => x"52",
           501 => x"88",
           502 => x"86",
           503 => x"e0",
           504 => x"06",
           505 => x"14",
           506 => x"80",
           507 => x"71",
           508 => x"0c",
           509 => x"04",
           510 => x"77",
           511 => x"53",
           512 => x"80",
           513 => x"38",
           514 => x"70",
           515 => x"81",
           516 => x"81",
           517 => x"39",
           518 => x"39",
           519 => x"80",
           520 => x"81",
           521 => x"55",
           522 => x"2e",
           523 => x"55",
           524 => x"84",
           525 => x"38",
           526 => x"06",
           527 => x"2e",
           528 => x"88",
           529 => x"70",
           530 => x"34",
           531 => x"71",
           532 => x"ec",
           533 => x"3d",
           534 => x"3d",
           535 => x"72",
           536 => x"91",
           537 => x"fc",
           538 => x"51",
           539 => x"81",
           540 => x"85",
           541 => x"83",
           542 => x"72",
           543 => x"0c",
           544 => x"04",
           545 => x"76",
           546 => x"ff",
           547 => x"81",
           548 => x"26",
           549 => x"83",
           550 => x"05",
           551 => x"70",
           552 => x"8a",
           553 => x"33",
           554 => x"70",
           555 => x"fe",
           556 => x"33",
           557 => x"70",
           558 => x"f2",
           559 => x"33",
           560 => x"70",
           561 => x"e6",
           562 => x"22",
           563 => x"74",
           564 => x"80",
           565 => x"13",
           566 => x"52",
           567 => x"26",
           568 => x"81",
           569 => x"98",
           570 => x"22",
           571 => x"bc",
           572 => x"33",
           573 => x"b8",
           574 => x"33",
           575 => x"b4",
           576 => x"33",
           577 => x"b0",
           578 => x"33",
           579 => x"ac",
           580 => x"33",
           581 => x"a8",
           582 => x"c0",
           583 => x"73",
           584 => x"a0",
           585 => x"87",
           586 => x"0c",
           587 => x"81",
           588 => x"86",
           589 => x"f3",
           590 => x"5b",
           591 => x"9c",
           592 => x"0c",
           593 => x"bc",
           594 => x"7b",
           595 => x"98",
           596 => x"79",
           597 => x"87",
           598 => x"08",
           599 => x"1c",
           600 => x"98",
           601 => x"79",
           602 => x"87",
           603 => x"08",
           604 => x"1c",
           605 => x"98",
           606 => x"79",
           607 => x"87",
           608 => x"08",
           609 => x"1c",
           610 => x"98",
           611 => x"79",
           612 => x"80",
           613 => x"83",
           614 => x"59",
           615 => x"ff",
           616 => x"1b",
           617 => x"1b",
           618 => x"1b",
           619 => x"1b",
           620 => x"1b",
           621 => x"83",
           622 => x"52",
           623 => x"51",
           624 => x"8f",
           625 => x"ff",
           626 => x"8f",
           627 => x"30",
           628 => x"51",
           629 => x"0b",
           630 => x"88",
           631 => x"0d",
           632 => x"0d",
           633 => x"81",
           634 => x"70",
           635 => x"57",
           636 => x"c0",
           637 => x"74",
           638 => x"38",
           639 => x"94",
           640 => x"70",
           641 => x"81",
           642 => x"52",
           643 => x"8c",
           644 => x"2a",
           645 => x"51",
           646 => x"38",
           647 => x"70",
           648 => x"51",
           649 => x"8d",
           650 => x"2a",
           651 => x"51",
           652 => x"be",
           653 => x"ff",
           654 => x"c0",
           655 => x"70",
           656 => x"38",
           657 => x"90",
           658 => x"0c",
           659 => x"e0",
           660 => x"0d",
           661 => x"0d",
           662 => x"33",
           663 => x"e9",
           664 => x"81",
           665 => x"55",
           666 => x"94",
           667 => x"80",
           668 => x"87",
           669 => x"51",
           670 => x"96",
           671 => x"06",
           672 => x"70",
           673 => x"38",
           674 => x"70",
           675 => x"51",
           676 => x"72",
           677 => x"81",
           678 => x"70",
           679 => x"38",
           680 => x"70",
           681 => x"51",
           682 => x"38",
           683 => x"06",
           684 => x"94",
           685 => x"80",
           686 => x"87",
           687 => x"52",
           688 => x"87",
           689 => x"f9",
           690 => x"54",
           691 => x"70",
           692 => x"53",
           693 => x"77",
           694 => x"38",
           695 => x"06",
           696 => x"0b",
           697 => x"33",
           698 => x"06",
           699 => x"58",
           700 => x"84",
           701 => x"2e",
           702 => x"c0",
           703 => x"70",
           704 => x"2a",
           705 => x"53",
           706 => x"80",
           707 => x"71",
           708 => x"81",
           709 => x"70",
           710 => x"81",
           711 => x"06",
           712 => x"80",
           713 => x"71",
           714 => x"81",
           715 => x"70",
           716 => x"74",
           717 => x"51",
           718 => x"80",
           719 => x"2e",
           720 => x"c0",
           721 => x"77",
           722 => x"17",
           723 => x"81",
           724 => x"53",
           725 => x"84",
           726 => x"ec",
           727 => x"3d",
           728 => x"3d",
           729 => x"81",
           730 => x"70",
           731 => x"54",
           732 => x"94",
           733 => x"80",
           734 => x"87",
           735 => x"51",
           736 => x"82",
           737 => x"06",
           738 => x"70",
           739 => x"38",
           740 => x"06",
           741 => x"94",
           742 => x"80",
           743 => x"87",
           744 => x"52",
           745 => x"81",
           746 => x"ec",
           747 => x"84",
           748 => x"fe",
           749 => x"0b",
           750 => x"33",
           751 => x"06",
           752 => x"c0",
           753 => x"70",
           754 => x"38",
           755 => x"94",
           756 => x"70",
           757 => x"81",
           758 => x"51",
           759 => x"80",
           760 => x"72",
           761 => x"51",
           762 => x"80",
           763 => x"2e",
           764 => x"c0",
           765 => x"71",
           766 => x"2b",
           767 => x"51",
           768 => x"81",
           769 => x"84",
           770 => x"ff",
           771 => x"c0",
           772 => x"70",
           773 => x"06",
           774 => x"80",
           775 => x"38",
           776 => x"a4",
           777 => x"8c",
           778 => x"9e",
           779 => x"e9",
           780 => x"c0",
           781 => x"81",
           782 => x"87",
           783 => x"08",
           784 => x"0c",
           785 => x"9c",
           786 => x"9c",
           787 => x"9e",
           788 => x"e9",
           789 => x"c0",
           790 => x"81",
           791 => x"87",
           792 => x"08",
           793 => x"0c",
           794 => x"b4",
           795 => x"ac",
           796 => x"9e",
           797 => x"e9",
           798 => x"c0",
           799 => x"81",
           800 => x"87",
           801 => x"08",
           802 => x"0c",
           803 => x"c4",
           804 => x"bc",
           805 => x"9e",
           806 => x"70",
           807 => x"23",
           808 => x"84",
           809 => x"c4",
           810 => x"9e",
           811 => x"e9",
           812 => x"c0",
           813 => x"81",
           814 => x"81",
           815 => x"d0",
           816 => x"87",
           817 => x"08",
           818 => x"0a",
           819 => x"52",
           820 => x"83",
           821 => x"71",
           822 => x"34",
           823 => x"c0",
           824 => x"70",
           825 => x"06",
           826 => x"70",
           827 => x"38",
           828 => x"81",
           829 => x"80",
           830 => x"9e",
           831 => x"90",
           832 => x"51",
           833 => x"80",
           834 => x"81",
           835 => x"e9",
           836 => x"0b",
           837 => x"90",
           838 => x"80",
           839 => x"52",
           840 => x"2e",
           841 => x"52",
           842 => x"d4",
           843 => x"87",
           844 => x"08",
           845 => x"80",
           846 => x"52",
           847 => x"83",
           848 => x"71",
           849 => x"34",
           850 => x"c0",
           851 => x"70",
           852 => x"06",
           853 => x"70",
           854 => x"38",
           855 => x"81",
           856 => x"80",
           857 => x"9e",
           858 => x"84",
           859 => x"51",
           860 => x"80",
           861 => x"81",
           862 => x"e9",
           863 => x"0b",
           864 => x"90",
           865 => x"80",
           866 => x"52",
           867 => x"2e",
           868 => x"52",
           869 => x"d8",
           870 => x"87",
           871 => x"08",
           872 => x"80",
           873 => x"52",
           874 => x"83",
           875 => x"71",
           876 => x"34",
           877 => x"c0",
           878 => x"70",
           879 => x"06",
           880 => x"70",
           881 => x"38",
           882 => x"81",
           883 => x"80",
           884 => x"9e",
           885 => x"a0",
           886 => x"52",
           887 => x"2e",
           888 => x"52",
           889 => x"db",
           890 => x"9e",
           891 => x"98",
           892 => x"8a",
           893 => x"51",
           894 => x"dc",
           895 => x"87",
           896 => x"08",
           897 => x"06",
           898 => x"70",
           899 => x"38",
           900 => x"81",
           901 => x"87",
           902 => x"08",
           903 => x"06",
           904 => x"51",
           905 => x"81",
           906 => x"80",
           907 => x"9e",
           908 => x"88",
           909 => x"52",
           910 => x"83",
           911 => x"71",
           912 => x"34",
           913 => x"90",
           914 => x"06",
           915 => x"81",
           916 => x"83",
           917 => x"fb",
           918 => x"d5",
           919 => x"c7",
           920 => x"d0",
           921 => x"80",
           922 => x"81",
           923 => x"85",
           924 => x"d6",
           925 => x"af",
           926 => x"d2",
           927 => x"80",
           928 => x"81",
           929 => x"81",
           930 => x"11",
           931 => x"d6",
           932 => x"f7",
           933 => x"d7",
           934 => x"80",
           935 => x"81",
           936 => x"81",
           937 => x"11",
           938 => x"d6",
           939 => x"db",
           940 => x"d4",
           941 => x"80",
           942 => x"81",
           943 => x"81",
           944 => x"11",
           945 => x"d6",
           946 => x"bf",
           947 => x"d5",
           948 => x"80",
           949 => x"81",
           950 => x"81",
           951 => x"11",
           952 => x"d7",
           953 => x"a3",
           954 => x"d6",
           955 => x"80",
           956 => x"81",
           957 => x"81",
           958 => x"11",
           959 => x"d7",
           960 => x"87",
           961 => x"db",
           962 => x"80",
           963 => x"81",
           964 => x"52",
           965 => x"51",
           966 => x"81",
           967 => x"54",
           968 => x"8d",
           969 => x"e0",
           970 => x"d7",
           971 => x"db",
           972 => x"dd",
           973 => x"80",
           974 => x"81",
           975 => x"52",
           976 => x"51",
           977 => x"81",
           978 => x"54",
           979 => x"88",
           980 => x"a4",
           981 => x"3f",
           982 => x"33",
           983 => x"2e",
           984 => x"d8",
           985 => x"bf",
           986 => x"d8",
           987 => x"80",
           988 => x"81",
           989 => x"83",
           990 => x"e9",
           991 => x"73",
           992 => x"38",
           993 => x"51",
           994 => x"81",
           995 => x"54",
           996 => x"88",
           997 => x"dc",
           998 => x"3f",
           999 => x"51",
          1000 => x"81",
          1001 => x"52",
          1002 => x"51",
          1003 => x"81",
          1004 => x"52",
          1005 => x"51",
          1006 => x"81",
          1007 => x"52",
          1008 => x"51",
          1009 => x"81",
          1010 => x"82",
          1011 => x"e9",
          1012 => x"81",
          1013 => x"88",
          1014 => x"e9",
          1015 => x"bd",
          1016 => x"75",
          1017 => x"3f",
          1018 => x"08",
          1019 => x"29",
          1020 => x"54",
          1021 => x"e0",
          1022 => x"da",
          1023 => x"8b",
          1024 => x"d7",
          1025 => x"80",
          1026 => x"81",
          1027 => x"56",
          1028 => x"52",
          1029 => x"95",
          1030 => x"e0",
          1031 => x"c0",
          1032 => x"31",
          1033 => x"ec",
          1034 => x"81",
          1035 => x"87",
          1036 => x"e9",
          1037 => x"73",
          1038 => x"38",
          1039 => x"08",
          1040 => x"c0",
          1041 => x"e9",
          1042 => x"ec",
          1043 => x"84",
          1044 => x"71",
          1045 => x"81",
          1046 => x"52",
          1047 => x"51",
          1048 => x"81",
          1049 => x"81",
          1050 => x"3d",
          1051 => x"3d",
          1052 => x"05",
          1053 => x"52",
          1054 => x"ac",
          1055 => x"29",
          1056 => x"d4",
          1057 => x"71",
          1058 => x"db",
          1059 => x"39",
          1060 => x"51",
          1061 => x"db",
          1062 => x"39",
          1063 => x"51",
          1064 => x"db",
          1065 => x"39",
          1066 => x"51",
          1067 => x"84",
          1068 => x"71",
          1069 => x"04",
          1070 => x"c0",
          1071 => x"04",
          1072 => x"08",
          1073 => x"84",
          1074 => x"3d",
          1075 => x"05",
          1076 => x"8a",
          1077 => x"06",
          1078 => x"51",
          1079 => x"ec",
          1080 => x"71",
          1081 => x"38",
          1082 => x"81",
          1083 => x"81",
          1084 => x"f8",
          1085 => x"81",
          1086 => x"52",
          1087 => x"85",
          1088 => x"71",
          1089 => x"0d",
          1090 => x"0d",
          1091 => x"33",
          1092 => x"08",
          1093 => x"f0",
          1094 => x"ff",
          1095 => x"81",
          1096 => x"84",
          1097 => x"fd",
          1098 => x"54",
          1099 => x"81",
          1100 => x"53",
          1101 => x"8e",
          1102 => x"ff",
          1103 => x"14",
          1104 => x"3f",
          1105 => x"3d",
          1106 => x"3d",
          1107 => x"ec",
          1108 => x"81",
          1109 => x"56",
          1110 => x"70",
          1111 => x"53",
          1112 => x"2e",
          1113 => x"81",
          1114 => x"81",
          1115 => x"da",
          1116 => x"74",
          1117 => x"0c",
          1118 => x"04",
          1119 => x"66",
          1120 => x"78",
          1121 => x"5a",
          1122 => x"80",
          1123 => x"38",
          1124 => x"09",
          1125 => x"de",
          1126 => x"7a",
          1127 => x"5c",
          1128 => x"5b",
          1129 => x"09",
          1130 => x"38",
          1131 => x"39",
          1132 => x"09",
          1133 => x"38",
          1134 => x"70",
          1135 => x"33",
          1136 => x"2e",
          1137 => x"92",
          1138 => x"19",
          1139 => x"70",
          1140 => x"33",
          1141 => x"53",
          1142 => x"16",
          1143 => x"26",
          1144 => x"88",
          1145 => x"05",
          1146 => x"05",
          1147 => x"05",
          1148 => x"5b",
          1149 => x"80",
          1150 => x"30",
          1151 => x"80",
          1152 => x"cc",
          1153 => x"70",
          1154 => x"25",
          1155 => x"54",
          1156 => x"53",
          1157 => x"8c",
          1158 => x"07",
          1159 => x"05",
          1160 => x"5a",
          1161 => x"83",
          1162 => x"54",
          1163 => x"27",
          1164 => x"16",
          1165 => x"06",
          1166 => x"80",
          1167 => x"aa",
          1168 => x"cf",
          1169 => x"73",
          1170 => x"81",
          1171 => x"80",
          1172 => x"38",
          1173 => x"2e",
          1174 => x"81",
          1175 => x"80",
          1176 => x"8a",
          1177 => x"39",
          1178 => x"2e",
          1179 => x"73",
          1180 => x"8a",
          1181 => x"d3",
          1182 => x"80",
          1183 => x"80",
          1184 => x"ee",
          1185 => x"39",
          1186 => x"71",
          1187 => x"53",
          1188 => x"54",
          1189 => x"2e",
          1190 => x"15",
          1191 => x"33",
          1192 => x"72",
          1193 => x"81",
          1194 => x"39",
          1195 => x"56",
          1196 => x"27",
          1197 => x"51",
          1198 => x"75",
          1199 => x"72",
          1200 => x"38",
          1201 => x"df",
          1202 => x"16",
          1203 => x"7b",
          1204 => x"38",
          1205 => x"f2",
          1206 => x"77",
          1207 => x"12",
          1208 => x"53",
          1209 => x"5c",
          1210 => x"5c",
          1211 => x"5c",
          1212 => x"5c",
          1213 => x"51",
          1214 => x"fd",
          1215 => x"82",
          1216 => x"06",
          1217 => x"80",
          1218 => x"77",
          1219 => x"53",
          1220 => x"18",
          1221 => x"72",
          1222 => x"c4",
          1223 => x"70",
          1224 => x"25",
          1225 => x"55",
          1226 => x"8d",
          1227 => x"2e",
          1228 => x"30",
          1229 => x"5b",
          1230 => x"8f",
          1231 => x"7b",
          1232 => x"e4",
          1233 => x"ec",
          1234 => x"ff",
          1235 => x"75",
          1236 => x"d9",
          1237 => x"e0",
          1238 => x"74",
          1239 => x"a7",
          1240 => x"80",
          1241 => x"38",
          1242 => x"72",
          1243 => x"54",
          1244 => x"72",
          1245 => x"05",
          1246 => x"17",
          1247 => x"77",
          1248 => x"51",
          1249 => x"9f",
          1250 => x"72",
          1251 => x"79",
          1252 => x"81",
          1253 => x"72",
          1254 => x"38",
          1255 => x"05",
          1256 => x"ad",
          1257 => x"17",
          1258 => x"81",
          1259 => x"b0",
          1260 => x"38",
          1261 => x"81",
          1262 => x"06",
          1263 => x"9f",
          1264 => x"55",
          1265 => x"97",
          1266 => x"f9",
          1267 => x"81",
          1268 => x"8b",
          1269 => x"16",
          1270 => x"73",
          1271 => x"96",
          1272 => x"e0",
          1273 => x"17",
          1274 => x"33",
          1275 => x"f9",
          1276 => x"f2",
          1277 => x"16",
          1278 => x"7b",
          1279 => x"38",
          1280 => x"c6",
          1281 => x"96",
          1282 => x"fd",
          1283 => x"3d",
          1284 => x"05",
          1285 => x"52",
          1286 => x"e0",
          1287 => x"0d",
          1288 => x"0d",
          1289 => x"f8",
          1290 => x"88",
          1291 => x"51",
          1292 => x"81",
          1293 => x"53",
          1294 => x"80",
          1295 => x"f8",
          1296 => x"0d",
          1297 => x"0d",
          1298 => x"08",
          1299 => x"f0",
          1300 => x"88",
          1301 => x"52",
          1302 => x"3f",
          1303 => x"f0",
          1304 => x"0d",
          1305 => x"0d",
          1306 => x"ec",
          1307 => x"56",
          1308 => x"80",
          1309 => x"2e",
          1310 => x"81",
          1311 => x"52",
          1312 => x"ec",
          1313 => x"ff",
          1314 => x"80",
          1315 => x"38",
          1316 => x"b9",
          1317 => x"32",
          1318 => x"80",
          1319 => x"52",
          1320 => x"8b",
          1321 => x"2e",
          1322 => x"14",
          1323 => x"9f",
          1324 => x"38",
          1325 => x"73",
          1326 => x"38",
          1327 => x"72",
          1328 => x"14",
          1329 => x"f8",
          1330 => x"af",
          1331 => x"52",
          1332 => x"8a",
          1333 => x"3f",
          1334 => x"81",
          1335 => x"87",
          1336 => x"fe",
          1337 => x"ec",
          1338 => x"81",
          1339 => x"77",
          1340 => x"53",
          1341 => x"72",
          1342 => x"0c",
          1343 => x"04",
          1344 => x"7a",
          1345 => x"80",
          1346 => x"58",
          1347 => x"33",
          1348 => x"a0",
          1349 => x"06",
          1350 => x"13",
          1351 => x"39",
          1352 => x"09",
          1353 => x"38",
          1354 => x"11",
          1355 => x"08",
          1356 => x"54",
          1357 => x"2e",
          1358 => x"80",
          1359 => x"08",
          1360 => x"0c",
          1361 => x"33",
          1362 => x"80",
          1363 => x"38",
          1364 => x"80",
          1365 => x"38",
          1366 => x"57",
          1367 => x"0c",
          1368 => x"33",
          1369 => x"39",
          1370 => x"74",
          1371 => x"38",
          1372 => x"80",
          1373 => x"89",
          1374 => x"38",
          1375 => x"d0",
          1376 => x"55",
          1377 => x"80",
          1378 => x"39",
          1379 => x"d9",
          1380 => x"80",
          1381 => x"27",
          1382 => x"80",
          1383 => x"89",
          1384 => x"70",
          1385 => x"55",
          1386 => x"70",
          1387 => x"55",
          1388 => x"27",
          1389 => x"14",
          1390 => x"06",
          1391 => x"74",
          1392 => x"73",
          1393 => x"38",
          1394 => x"14",
          1395 => x"05",
          1396 => x"08",
          1397 => x"54",
          1398 => x"39",
          1399 => x"84",
          1400 => x"55",
          1401 => x"81",
          1402 => x"ec",
          1403 => x"3d",
          1404 => x"3d",
          1405 => x"5a",
          1406 => x"7a",
          1407 => x"08",
          1408 => x"53",
          1409 => x"09",
          1410 => x"38",
          1411 => x"0c",
          1412 => x"ad",
          1413 => x"06",
          1414 => x"76",
          1415 => x"0c",
          1416 => x"33",
          1417 => x"73",
          1418 => x"81",
          1419 => x"38",
          1420 => x"05",
          1421 => x"08",
          1422 => x"53",
          1423 => x"2e",
          1424 => x"57",
          1425 => x"2e",
          1426 => x"39",
          1427 => x"13",
          1428 => x"08",
          1429 => x"53",
          1430 => x"55",
          1431 => x"80",
          1432 => x"14",
          1433 => x"88",
          1434 => x"27",
          1435 => x"eb",
          1436 => x"53",
          1437 => x"89",
          1438 => x"38",
          1439 => x"55",
          1440 => x"8a",
          1441 => x"a0",
          1442 => x"c2",
          1443 => x"74",
          1444 => x"e0",
          1445 => x"ff",
          1446 => x"d0",
          1447 => x"ff",
          1448 => x"90",
          1449 => x"38",
          1450 => x"81",
          1451 => x"53",
          1452 => x"ca",
          1453 => x"27",
          1454 => x"77",
          1455 => x"08",
          1456 => x"0c",
          1457 => x"33",
          1458 => x"ff",
          1459 => x"80",
          1460 => x"74",
          1461 => x"79",
          1462 => x"74",
          1463 => x"0c",
          1464 => x"04",
          1465 => x"02",
          1466 => x"51",
          1467 => x"72",
          1468 => x"81",
          1469 => x"33",
          1470 => x"ec",
          1471 => x"3d",
          1472 => x"3d",
          1473 => x"05",
          1474 => x"05",
          1475 => x"56",
          1476 => x"72",
          1477 => x"e0",
          1478 => x"2b",
          1479 => x"8c",
          1480 => x"88",
          1481 => x"2e",
          1482 => x"88",
          1483 => x"0c",
          1484 => x"8c",
          1485 => x"71",
          1486 => x"87",
          1487 => x"0c",
          1488 => x"08",
          1489 => x"51",
          1490 => x"2e",
          1491 => x"c0",
          1492 => x"51",
          1493 => x"71",
          1494 => x"80",
          1495 => x"92",
          1496 => x"98",
          1497 => x"70",
          1498 => x"38",
          1499 => x"e8",
          1500 => x"e9",
          1501 => x"51",
          1502 => x"e0",
          1503 => x"0d",
          1504 => x"0d",
          1505 => x"02",
          1506 => x"05",
          1507 => x"58",
          1508 => x"52",
          1509 => x"3f",
          1510 => x"08",
          1511 => x"54",
          1512 => x"be",
          1513 => x"75",
          1514 => x"c0",
          1515 => x"87",
          1516 => x"12",
          1517 => x"84",
          1518 => x"40",
          1519 => x"85",
          1520 => x"98",
          1521 => x"7d",
          1522 => x"0c",
          1523 => x"85",
          1524 => x"06",
          1525 => x"71",
          1526 => x"38",
          1527 => x"71",
          1528 => x"05",
          1529 => x"19",
          1530 => x"a2",
          1531 => x"71",
          1532 => x"38",
          1533 => x"83",
          1534 => x"38",
          1535 => x"8a",
          1536 => x"98",
          1537 => x"71",
          1538 => x"c0",
          1539 => x"52",
          1540 => x"87",
          1541 => x"80",
          1542 => x"81",
          1543 => x"c0",
          1544 => x"53",
          1545 => x"82",
          1546 => x"71",
          1547 => x"1a",
          1548 => x"84",
          1549 => x"19",
          1550 => x"06",
          1551 => x"79",
          1552 => x"38",
          1553 => x"80",
          1554 => x"87",
          1555 => x"26",
          1556 => x"73",
          1557 => x"06",
          1558 => x"2e",
          1559 => x"52",
          1560 => x"81",
          1561 => x"8f",
          1562 => x"f3",
          1563 => x"62",
          1564 => x"05",
          1565 => x"57",
          1566 => x"83",
          1567 => x"52",
          1568 => x"3f",
          1569 => x"08",
          1570 => x"54",
          1571 => x"2e",
          1572 => x"81",
          1573 => x"74",
          1574 => x"c0",
          1575 => x"87",
          1576 => x"12",
          1577 => x"84",
          1578 => x"5f",
          1579 => x"0b",
          1580 => x"8c",
          1581 => x"0c",
          1582 => x"80",
          1583 => x"70",
          1584 => x"81",
          1585 => x"54",
          1586 => x"8c",
          1587 => x"81",
          1588 => x"7c",
          1589 => x"58",
          1590 => x"70",
          1591 => x"52",
          1592 => x"8a",
          1593 => x"98",
          1594 => x"71",
          1595 => x"c0",
          1596 => x"52",
          1597 => x"87",
          1598 => x"80",
          1599 => x"81",
          1600 => x"c0",
          1601 => x"53",
          1602 => x"82",
          1603 => x"71",
          1604 => x"19",
          1605 => x"81",
          1606 => x"ff",
          1607 => x"19",
          1608 => x"78",
          1609 => x"38",
          1610 => x"80",
          1611 => x"87",
          1612 => x"26",
          1613 => x"73",
          1614 => x"06",
          1615 => x"2e",
          1616 => x"52",
          1617 => x"81",
          1618 => x"8f",
          1619 => x"fa",
          1620 => x"02",
          1621 => x"05",
          1622 => x"05",
          1623 => x"71",
          1624 => x"57",
          1625 => x"81",
          1626 => x"81",
          1627 => x"54",
          1628 => x"38",
          1629 => x"c0",
          1630 => x"81",
          1631 => x"2e",
          1632 => x"71",
          1633 => x"38",
          1634 => x"87",
          1635 => x"11",
          1636 => x"80",
          1637 => x"80",
          1638 => x"83",
          1639 => x"38",
          1640 => x"72",
          1641 => x"2a",
          1642 => x"51",
          1643 => x"80",
          1644 => x"87",
          1645 => x"08",
          1646 => x"38",
          1647 => x"8c",
          1648 => x"96",
          1649 => x"0c",
          1650 => x"8c",
          1651 => x"08",
          1652 => x"51",
          1653 => x"38",
          1654 => x"56",
          1655 => x"80",
          1656 => x"85",
          1657 => x"77",
          1658 => x"83",
          1659 => x"75",
          1660 => x"ec",
          1661 => x"3d",
          1662 => x"3d",
          1663 => x"11",
          1664 => x"71",
          1665 => x"81",
          1666 => x"53",
          1667 => x"0d",
          1668 => x"0d",
          1669 => x"33",
          1670 => x"71",
          1671 => x"88",
          1672 => x"14",
          1673 => x"07",
          1674 => x"33",
          1675 => x"ec",
          1676 => x"53",
          1677 => x"52",
          1678 => x"04",
          1679 => x"73",
          1680 => x"92",
          1681 => x"52",
          1682 => x"81",
          1683 => x"70",
          1684 => x"70",
          1685 => x"3d",
          1686 => x"3d",
          1687 => x"52",
          1688 => x"70",
          1689 => x"34",
          1690 => x"51",
          1691 => x"81",
          1692 => x"70",
          1693 => x"70",
          1694 => x"05",
          1695 => x"88",
          1696 => x"72",
          1697 => x"0d",
          1698 => x"0d",
          1699 => x"54",
          1700 => x"80",
          1701 => x"71",
          1702 => x"53",
          1703 => x"81",
          1704 => x"ff",
          1705 => x"39",
          1706 => x"04",
          1707 => x"75",
          1708 => x"52",
          1709 => x"70",
          1710 => x"34",
          1711 => x"70",
          1712 => x"3d",
          1713 => x"3d",
          1714 => x"79",
          1715 => x"74",
          1716 => x"56",
          1717 => x"81",
          1718 => x"71",
          1719 => x"16",
          1720 => x"52",
          1721 => x"86",
          1722 => x"2e",
          1723 => x"81",
          1724 => x"86",
          1725 => x"fe",
          1726 => x"76",
          1727 => x"39",
          1728 => x"8a",
          1729 => x"51",
          1730 => x"71",
          1731 => x"33",
          1732 => x"0c",
          1733 => x"04",
          1734 => x"ec",
          1735 => x"80",
          1736 => x"e0",
          1737 => x"3d",
          1738 => x"80",
          1739 => x"33",
          1740 => x"7a",
          1741 => x"38",
          1742 => x"16",
          1743 => x"16",
          1744 => x"17",
          1745 => x"fa",
          1746 => x"ec",
          1747 => x"2e",
          1748 => x"b7",
          1749 => x"e0",
          1750 => x"34",
          1751 => x"70",
          1752 => x"31",
          1753 => x"59",
          1754 => x"77",
          1755 => x"82",
          1756 => x"74",
          1757 => x"81",
          1758 => x"81",
          1759 => x"53",
          1760 => x"16",
          1761 => x"e3",
          1762 => x"81",
          1763 => x"ec",
          1764 => x"3d",
          1765 => x"3d",
          1766 => x"56",
          1767 => x"74",
          1768 => x"2e",
          1769 => x"51",
          1770 => x"81",
          1771 => x"57",
          1772 => x"08",
          1773 => x"54",
          1774 => x"16",
          1775 => x"33",
          1776 => x"3f",
          1777 => x"08",
          1778 => x"38",
          1779 => x"57",
          1780 => x"0c",
          1781 => x"e0",
          1782 => x"0d",
          1783 => x"0d",
          1784 => x"57",
          1785 => x"81",
          1786 => x"58",
          1787 => x"08",
          1788 => x"76",
          1789 => x"83",
          1790 => x"06",
          1791 => x"84",
          1792 => x"78",
          1793 => x"81",
          1794 => x"38",
          1795 => x"81",
          1796 => x"52",
          1797 => x"52",
          1798 => x"3f",
          1799 => x"52",
          1800 => x"51",
          1801 => x"84",
          1802 => x"d2",
          1803 => x"fc",
          1804 => x"8a",
          1805 => x"52",
          1806 => x"51",
          1807 => x"90",
          1808 => x"84",
          1809 => x"fc",
          1810 => x"17",
          1811 => x"a0",
          1812 => x"86",
          1813 => x"08",
          1814 => x"b0",
          1815 => x"55",
          1816 => x"81",
          1817 => x"f8",
          1818 => x"84",
          1819 => x"53",
          1820 => x"17",
          1821 => x"d7",
          1822 => x"e0",
          1823 => x"83",
          1824 => x"77",
          1825 => x"0c",
          1826 => x"04",
          1827 => x"77",
          1828 => x"12",
          1829 => x"55",
          1830 => x"56",
          1831 => x"8d",
          1832 => x"22",
          1833 => x"ac",
          1834 => x"57",
          1835 => x"ec",
          1836 => x"3d",
          1837 => x"3d",
          1838 => x"70",
          1839 => x"57",
          1840 => x"81",
          1841 => x"98",
          1842 => x"81",
          1843 => x"74",
          1844 => x"72",
          1845 => x"f5",
          1846 => x"24",
          1847 => x"81",
          1848 => x"81",
          1849 => x"83",
          1850 => x"38",
          1851 => x"76",
          1852 => x"70",
          1853 => x"16",
          1854 => x"74",
          1855 => x"96",
          1856 => x"e0",
          1857 => x"38",
          1858 => x"06",
          1859 => x"33",
          1860 => x"89",
          1861 => x"08",
          1862 => x"54",
          1863 => x"fc",
          1864 => x"ec",
          1865 => x"fe",
          1866 => x"ff",
          1867 => x"11",
          1868 => x"2b",
          1869 => x"81",
          1870 => x"2a",
          1871 => x"51",
          1872 => x"e2",
          1873 => x"ff",
          1874 => x"da",
          1875 => x"2a",
          1876 => x"05",
          1877 => x"fc",
          1878 => x"ec",
          1879 => x"c6",
          1880 => x"83",
          1881 => x"05",
          1882 => x"f9",
          1883 => x"ec",
          1884 => x"ff",
          1885 => x"ae",
          1886 => x"2a",
          1887 => x"05",
          1888 => x"fc",
          1889 => x"ec",
          1890 => x"38",
          1891 => x"83",
          1892 => x"05",
          1893 => x"f8",
          1894 => x"ec",
          1895 => x"0a",
          1896 => x"39",
          1897 => x"81",
          1898 => x"89",
          1899 => x"f8",
          1900 => x"7c",
          1901 => x"56",
          1902 => x"77",
          1903 => x"38",
          1904 => x"08",
          1905 => x"38",
          1906 => x"72",
          1907 => x"9d",
          1908 => x"24",
          1909 => x"81",
          1910 => x"82",
          1911 => x"83",
          1912 => x"38",
          1913 => x"76",
          1914 => x"70",
          1915 => x"18",
          1916 => x"76",
          1917 => x"9e",
          1918 => x"e0",
          1919 => x"ec",
          1920 => x"d9",
          1921 => x"ff",
          1922 => x"05",
          1923 => x"81",
          1924 => x"54",
          1925 => x"80",
          1926 => x"77",
          1927 => x"f0",
          1928 => x"8f",
          1929 => x"51",
          1930 => x"34",
          1931 => x"17",
          1932 => x"2a",
          1933 => x"05",
          1934 => x"fa",
          1935 => x"ec",
          1936 => x"81",
          1937 => x"81",
          1938 => x"83",
          1939 => x"b4",
          1940 => x"2a",
          1941 => x"8f",
          1942 => x"2a",
          1943 => x"f0",
          1944 => x"06",
          1945 => x"72",
          1946 => x"ec",
          1947 => x"2a",
          1948 => x"05",
          1949 => x"fa",
          1950 => x"ec",
          1951 => x"81",
          1952 => x"80",
          1953 => x"83",
          1954 => x"52",
          1955 => x"fe",
          1956 => x"b4",
          1957 => x"a4",
          1958 => x"76",
          1959 => x"17",
          1960 => x"75",
          1961 => x"3f",
          1962 => x"08",
          1963 => x"e0",
          1964 => x"77",
          1965 => x"77",
          1966 => x"fc",
          1967 => x"b4",
          1968 => x"51",
          1969 => x"c9",
          1970 => x"e0",
          1971 => x"06",
          1972 => x"72",
          1973 => x"3f",
          1974 => x"17",
          1975 => x"ec",
          1976 => x"3d",
          1977 => x"3d",
          1978 => x"7e",
          1979 => x"56",
          1980 => x"75",
          1981 => x"74",
          1982 => x"27",
          1983 => x"80",
          1984 => x"ff",
          1985 => x"75",
          1986 => x"3f",
          1987 => x"08",
          1988 => x"e0",
          1989 => x"38",
          1990 => x"54",
          1991 => x"81",
          1992 => x"39",
          1993 => x"08",
          1994 => x"39",
          1995 => x"51",
          1996 => x"81",
          1997 => x"58",
          1998 => x"08",
          1999 => x"c7",
          2000 => x"e0",
          2001 => x"d2",
          2002 => x"e0",
          2003 => x"cf",
          2004 => x"74",
          2005 => x"fc",
          2006 => x"ec",
          2007 => x"38",
          2008 => x"fe",
          2009 => x"08",
          2010 => x"74",
          2011 => x"38",
          2012 => x"17",
          2013 => x"33",
          2014 => x"73",
          2015 => x"77",
          2016 => x"26",
          2017 => x"80",
          2018 => x"ec",
          2019 => x"3d",
          2020 => x"3d",
          2021 => x"71",
          2022 => x"5b",
          2023 => x"8c",
          2024 => x"77",
          2025 => x"38",
          2026 => x"78",
          2027 => x"81",
          2028 => x"79",
          2029 => x"f9",
          2030 => x"55",
          2031 => x"e0",
          2032 => x"e0",
          2033 => x"e0",
          2034 => x"ec",
          2035 => x"2e",
          2036 => x"98",
          2037 => x"ec",
          2038 => x"82",
          2039 => x"58",
          2040 => x"70",
          2041 => x"80",
          2042 => x"38",
          2043 => x"09",
          2044 => x"e2",
          2045 => x"56",
          2046 => x"76",
          2047 => x"82",
          2048 => x"7a",
          2049 => x"3f",
          2050 => x"ec",
          2051 => x"2e",
          2052 => x"86",
          2053 => x"e0",
          2054 => x"ec",
          2055 => x"70",
          2056 => x"07",
          2057 => x"7c",
          2058 => x"e0",
          2059 => x"51",
          2060 => x"81",
          2061 => x"ec",
          2062 => x"2e",
          2063 => x"17",
          2064 => x"74",
          2065 => x"73",
          2066 => x"27",
          2067 => x"58",
          2068 => x"80",
          2069 => x"56",
          2070 => x"98",
          2071 => x"26",
          2072 => x"56",
          2073 => x"81",
          2074 => x"52",
          2075 => x"c6",
          2076 => x"e0",
          2077 => x"b8",
          2078 => x"81",
          2079 => x"81",
          2080 => x"06",
          2081 => x"ec",
          2082 => x"81",
          2083 => x"09",
          2084 => x"72",
          2085 => x"70",
          2086 => x"51",
          2087 => x"80",
          2088 => x"78",
          2089 => x"06",
          2090 => x"73",
          2091 => x"39",
          2092 => x"52",
          2093 => x"f7",
          2094 => x"e0",
          2095 => x"e0",
          2096 => x"81",
          2097 => x"07",
          2098 => x"55",
          2099 => x"2e",
          2100 => x"80",
          2101 => x"75",
          2102 => x"76",
          2103 => x"3f",
          2104 => x"08",
          2105 => x"38",
          2106 => x"0c",
          2107 => x"fe",
          2108 => x"08",
          2109 => x"74",
          2110 => x"ff",
          2111 => x"0c",
          2112 => x"81",
          2113 => x"84",
          2114 => x"39",
          2115 => x"81",
          2116 => x"8c",
          2117 => x"8c",
          2118 => x"e0",
          2119 => x"39",
          2120 => x"55",
          2121 => x"e0",
          2122 => x"0d",
          2123 => x"0d",
          2124 => x"55",
          2125 => x"81",
          2126 => x"58",
          2127 => x"ec",
          2128 => x"d8",
          2129 => x"74",
          2130 => x"3f",
          2131 => x"08",
          2132 => x"08",
          2133 => x"59",
          2134 => x"77",
          2135 => x"70",
          2136 => x"c8",
          2137 => x"84",
          2138 => x"56",
          2139 => x"58",
          2140 => x"97",
          2141 => x"75",
          2142 => x"52",
          2143 => x"51",
          2144 => x"81",
          2145 => x"80",
          2146 => x"8a",
          2147 => x"32",
          2148 => x"72",
          2149 => x"2a",
          2150 => x"56",
          2151 => x"e0",
          2152 => x"0d",
          2153 => x"0d",
          2154 => x"08",
          2155 => x"74",
          2156 => x"26",
          2157 => x"74",
          2158 => x"72",
          2159 => x"74",
          2160 => x"88",
          2161 => x"73",
          2162 => x"33",
          2163 => x"27",
          2164 => x"16",
          2165 => x"9b",
          2166 => x"2a",
          2167 => x"88",
          2168 => x"58",
          2169 => x"80",
          2170 => x"16",
          2171 => x"0c",
          2172 => x"8a",
          2173 => x"89",
          2174 => x"72",
          2175 => x"38",
          2176 => x"51",
          2177 => x"81",
          2178 => x"54",
          2179 => x"08",
          2180 => x"38",
          2181 => x"ec",
          2182 => x"8b",
          2183 => x"08",
          2184 => x"08",
          2185 => x"82",
          2186 => x"74",
          2187 => x"cb",
          2188 => x"75",
          2189 => x"3f",
          2190 => x"08",
          2191 => x"73",
          2192 => x"98",
          2193 => x"82",
          2194 => x"2e",
          2195 => x"39",
          2196 => x"39",
          2197 => x"13",
          2198 => x"74",
          2199 => x"16",
          2200 => x"18",
          2201 => x"77",
          2202 => x"0c",
          2203 => x"04",
          2204 => x"7a",
          2205 => x"12",
          2206 => x"59",
          2207 => x"80",
          2208 => x"86",
          2209 => x"98",
          2210 => x"14",
          2211 => x"55",
          2212 => x"81",
          2213 => x"83",
          2214 => x"77",
          2215 => x"81",
          2216 => x"0c",
          2217 => x"55",
          2218 => x"76",
          2219 => x"17",
          2220 => x"74",
          2221 => x"9b",
          2222 => x"39",
          2223 => x"ff",
          2224 => x"2a",
          2225 => x"81",
          2226 => x"52",
          2227 => x"e6",
          2228 => x"e0",
          2229 => x"55",
          2230 => x"ec",
          2231 => x"80",
          2232 => x"55",
          2233 => x"08",
          2234 => x"f4",
          2235 => x"08",
          2236 => x"08",
          2237 => x"38",
          2238 => x"77",
          2239 => x"84",
          2240 => x"39",
          2241 => x"52",
          2242 => x"86",
          2243 => x"e0",
          2244 => x"55",
          2245 => x"08",
          2246 => x"c4",
          2247 => x"81",
          2248 => x"81",
          2249 => x"81",
          2250 => x"e0",
          2251 => x"b0",
          2252 => x"e0",
          2253 => x"51",
          2254 => x"81",
          2255 => x"a0",
          2256 => x"15",
          2257 => x"75",
          2258 => x"3f",
          2259 => x"08",
          2260 => x"76",
          2261 => x"77",
          2262 => x"9c",
          2263 => x"55",
          2264 => x"e0",
          2265 => x"0d",
          2266 => x"0d",
          2267 => x"08",
          2268 => x"80",
          2269 => x"fc",
          2270 => x"ec",
          2271 => x"81",
          2272 => x"80",
          2273 => x"ec",
          2274 => x"98",
          2275 => x"78",
          2276 => x"3f",
          2277 => x"08",
          2278 => x"e0",
          2279 => x"38",
          2280 => x"08",
          2281 => x"70",
          2282 => x"58",
          2283 => x"2e",
          2284 => x"83",
          2285 => x"81",
          2286 => x"55",
          2287 => x"81",
          2288 => x"07",
          2289 => x"2e",
          2290 => x"16",
          2291 => x"2e",
          2292 => x"88",
          2293 => x"81",
          2294 => x"56",
          2295 => x"51",
          2296 => x"81",
          2297 => x"54",
          2298 => x"08",
          2299 => x"9b",
          2300 => x"2e",
          2301 => x"83",
          2302 => x"73",
          2303 => x"0c",
          2304 => x"04",
          2305 => x"76",
          2306 => x"54",
          2307 => x"81",
          2308 => x"83",
          2309 => x"76",
          2310 => x"53",
          2311 => x"2e",
          2312 => x"90",
          2313 => x"51",
          2314 => x"81",
          2315 => x"90",
          2316 => x"53",
          2317 => x"e0",
          2318 => x"0d",
          2319 => x"0d",
          2320 => x"83",
          2321 => x"54",
          2322 => x"55",
          2323 => x"3f",
          2324 => x"51",
          2325 => x"2e",
          2326 => x"8b",
          2327 => x"2a",
          2328 => x"51",
          2329 => x"86",
          2330 => x"f7",
          2331 => x"7d",
          2332 => x"75",
          2333 => x"98",
          2334 => x"2e",
          2335 => x"98",
          2336 => x"78",
          2337 => x"3f",
          2338 => x"08",
          2339 => x"e0",
          2340 => x"38",
          2341 => x"70",
          2342 => x"73",
          2343 => x"58",
          2344 => x"8b",
          2345 => x"bf",
          2346 => x"ff",
          2347 => x"53",
          2348 => x"34",
          2349 => x"08",
          2350 => x"e5",
          2351 => x"81",
          2352 => x"2e",
          2353 => x"70",
          2354 => x"57",
          2355 => x"9e",
          2356 => x"2e",
          2357 => x"ec",
          2358 => x"df",
          2359 => x"72",
          2360 => x"81",
          2361 => x"76",
          2362 => x"2e",
          2363 => x"52",
          2364 => x"fc",
          2365 => x"e0",
          2366 => x"ec",
          2367 => x"38",
          2368 => x"fe",
          2369 => x"39",
          2370 => x"16",
          2371 => x"ec",
          2372 => x"3d",
          2373 => x"3d",
          2374 => x"08",
          2375 => x"52",
          2376 => x"c5",
          2377 => x"e0",
          2378 => x"ec",
          2379 => x"38",
          2380 => x"52",
          2381 => x"de",
          2382 => x"e0",
          2383 => x"ec",
          2384 => x"38",
          2385 => x"ec",
          2386 => x"9c",
          2387 => x"ea",
          2388 => x"53",
          2389 => x"9c",
          2390 => x"ea",
          2391 => x"0b",
          2392 => x"74",
          2393 => x"0c",
          2394 => x"04",
          2395 => x"75",
          2396 => x"12",
          2397 => x"53",
          2398 => x"9a",
          2399 => x"e0",
          2400 => x"9c",
          2401 => x"e5",
          2402 => x"0b",
          2403 => x"85",
          2404 => x"fa",
          2405 => x"7a",
          2406 => x"0b",
          2407 => x"98",
          2408 => x"2e",
          2409 => x"80",
          2410 => x"55",
          2411 => x"17",
          2412 => x"33",
          2413 => x"51",
          2414 => x"2e",
          2415 => x"85",
          2416 => x"06",
          2417 => x"e5",
          2418 => x"2e",
          2419 => x"8b",
          2420 => x"70",
          2421 => x"34",
          2422 => x"71",
          2423 => x"05",
          2424 => x"15",
          2425 => x"27",
          2426 => x"15",
          2427 => x"80",
          2428 => x"34",
          2429 => x"52",
          2430 => x"88",
          2431 => x"17",
          2432 => x"52",
          2433 => x"3f",
          2434 => x"08",
          2435 => x"12",
          2436 => x"3f",
          2437 => x"08",
          2438 => x"98",
          2439 => x"da",
          2440 => x"e0",
          2441 => x"23",
          2442 => x"04",
          2443 => x"7f",
          2444 => x"5b",
          2445 => x"33",
          2446 => x"73",
          2447 => x"38",
          2448 => x"80",
          2449 => x"38",
          2450 => x"8c",
          2451 => x"08",
          2452 => x"aa",
          2453 => x"41",
          2454 => x"33",
          2455 => x"73",
          2456 => x"81",
          2457 => x"81",
          2458 => x"dc",
          2459 => x"70",
          2460 => x"07",
          2461 => x"73",
          2462 => x"88",
          2463 => x"70",
          2464 => x"73",
          2465 => x"38",
          2466 => x"ab",
          2467 => x"52",
          2468 => x"91",
          2469 => x"e0",
          2470 => x"98",
          2471 => x"61",
          2472 => x"5a",
          2473 => x"a0",
          2474 => x"e7",
          2475 => x"70",
          2476 => x"79",
          2477 => x"73",
          2478 => x"81",
          2479 => x"38",
          2480 => x"33",
          2481 => x"ae",
          2482 => x"70",
          2483 => x"82",
          2484 => x"51",
          2485 => x"54",
          2486 => x"79",
          2487 => x"74",
          2488 => x"57",
          2489 => x"af",
          2490 => x"70",
          2491 => x"51",
          2492 => x"dc",
          2493 => x"73",
          2494 => x"38",
          2495 => x"82",
          2496 => x"19",
          2497 => x"54",
          2498 => x"82",
          2499 => x"54",
          2500 => x"78",
          2501 => x"81",
          2502 => x"54",
          2503 => x"81",
          2504 => x"af",
          2505 => x"77",
          2506 => x"70",
          2507 => x"25",
          2508 => x"07",
          2509 => x"51",
          2510 => x"2e",
          2511 => x"39",
          2512 => x"80",
          2513 => x"33",
          2514 => x"73",
          2515 => x"81",
          2516 => x"81",
          2517 => x"dc",
          2518 => x"70",
          2519 => x"07",
          2520 => x"73",
          2521 => x"b5",
          2522 => x"2e",
          2523 => x"83",
          2524 => x"76",
          2525 => x"07",
          2526 => x"2e",
          2527 => x"8b",
          2528 => x"77",
          2529 => x"30",
          2530 => x"71",
          2531 => x"53",
          2532 => x"55",
          2533 => x"38",
          2534 => x"5c",
          2535 => x"75",
          2536 => x"73",
          2537 => x"38",
          2538 => x"06",
          2539 => x"11",
          2540 => x"75",
          2541 => x"3f",
          2542 => x"08",
          2543 => x"38",
          2544 => x"33",
          2545 => x"54",
          2546 => x"e6",
          2547 => x"ec",
          2548 => x"2e",
          2549 => x"ff",
          2550 => x"74",
          2551 => x"38",
          2552 => x"75",
          2553 => x"17",
          2554 => x"57",
          2555 => x"a7",
          2556 => x"81",
          2557 => x"e5",
          2558 => x"ec",
          2559 => x"38",
          2560 => x"54",
          2561 => x"89",
          2562 => x"70",
          2563 => x"57",
          2564 => x"54",
          2565 => x"81",
          2566 => x"f7",
          2567 => x"7e",
          2568 => x"2e",
          2569 => x"33",
          2570 => x"e5",
          2571 => x"06",
          2572 => x"7a",
          2573 => x"a0",
          2574 => x"38",
          2575 => x"55",
          2576 => x"84",
          2577 => x"39",
          2578 => x"8b",
          2579 => x"7b",
          2580 => x"7a",
          2581 => x"3f",
          2582 => x"08",
          2583 => x"e0",
          2584 => x"38",
          2585 => x"52",
          2586 => x"aa",
          2587 => x"e0",
          2588 => x"ec",
          2589 => x"c2",
          2590 => x"08",
          2591 => x"55",
          2592 => x"ff",
          2593 => x"15",
          2594 => x"54",
          2595 => x"34",
          2596 => x"70",
          2597 => x"81",
          2598 => x"58",
          2599 => x"8b",
          2600 => x"74",
          2601 => x"3f",
          2602 => x"08",
          2603 => x"38",
          2604 => x"51",
          2605 => x"ff",
          2606 => x"ab",
          2607 => x"55",
          2608 => x"bb",
          2609 => x"2e",
          2610 => x"80",
          2611 => x"85",
          2612 => x"06",
          2613 => x"58",
          2614 => x"80",
          2615 => x"75",
          2616 => x"73",
          2617 => x"b5",
          2618 => x"0b",
          2619 => x"80",
          2620 => x"39",
          2621 => x"54",
          2622 => x"85",
          2623 => x"75",
          2624 => x"81",
          2625 => x"73",
          2626 => x"1b",
          2627 => x"2a",
          2628 => x"51",
          2629 => x"80",
          2630 => x"90",
          2631 => x"ff",
          2632 => x"05",
          2633 => x"f5",
          2634 => x"ec",
          2635 => x"1c",
          2636 => x"39",
          2637 => x"e0",
          2638 => x"0d",
          2639 => x"0d",
          2640 => x"7b",
          2641 => x"73",
          2642 => x"55",
          2643 => x"2e",
          2644 => x"75",
          2645 => x"57",
          2646 => x"26",
          2647 => x"ba",
          2648 => x"70",
          2649 => x"ba",
          2650 => x"06",
          2651 => x"73",
          2652 => x"70",
          2653 => x"51",
          2654 => x"89",
          2655 => x"82",
          2656 => x"ff",
          2657 => x"56",
          2658 => x"2e",
          2659 => x"80",
          2660 => x"a0",
          2661 => x"08",
          2662 => x"76",
          2663 => x"58",
          2664 => x"81",
          2665 => x"ff",
          2666 => x"53",
          2667 => x"26",
          2668 => x"13",
          2669 => x"06",
          2670 => x"9f",
          2671 => x"99",
          2672 => x"e0",
          2673 => x"ff",
          2674 => x"72",
          2675 => x"2a",
          2676 => x"72",
          2677 => x"06",
          2678 => x"ff",
          2679 => x"30",
          2680 => x"70",
          2681 => x"07",
          2682 => x"9f",
          2683 => x"54",
          2684 => x"80",
          2685 => x"81",
          2686 => x"59",
          2687 => x"25",
          2688 => x"8b",
          2689 => x"24",
          2690 => x"76",
          2691 => x"78",
          2692 => x"81",
          2693 => x"51",
          2694 => x"e0",
          2695 => x"0d",
          2696 => x"0d",
          2697 => x"0b",
          2698 => x"ff",
          2699 => x"0c",
          2700 => x"51",
          2701 => x"84",
          2702 => x"e0",
          2703 => x"38",
          2704 => x"51",
          2705 => x"81",
          2706 => x"83",
          2707 => x"54",
          2708 => x"82",
          2709 => x"09",
          2710 => x"e3",
          2711 => x"b4",
          2712 => x"57",
          2713 => x"2e",
          2714 => x"83",
          2715 => x"74",
          2716 => x"70",
          2717 => x"25",
          2718 => x"51",
          2719 => x"38",
          2720 => x"2e",
          2721 => x"b5",
          2722 => x"81",
          2723 => x"80",
          2724 => x"e0",
          2725 => x"ec",
          2726 => x"81",
          2727 => x"80",
          2728 => x"85",
          2729 => x"e4",
          2730 => x"16",
          2731 => x"3f",
          2732 => x"08",
          2733 => x"e0",
          2734 => x"83",
          2735 => x"74",
          2736 => x"0c",
          2737 => x"04",
          2738 => x"61",
          2739 => x"80",
          2740 => x"58",
          2741 => x"0c",
          2742 => x"e1",
          2743 => x"e0",
          2744 => x"56",
          2745 => x"ec",
          2746 => x"86",
          2747 => x"ec",
          2748 => x"29",
          2749 => x"05",
          2750 => x"53",
          2751 => x"80",
          2752 => x"38",
          2753 => x"76",
          2754 => x"74",
          2755 => x"72",
          2756 => x"38",
          2757 => x"51",
          2758 => x"81",
          2759 => x"81",
          2760 => x"81",
          2761 => x"72",
          2762 => x"80",
          2763 => x"38",
          2764 => x"70",
          2765 => x"53",
          2766 => x"86",
          2767 => x"a7",
          2768 => x"34",
          2769 => x"34",
          2770 => x"14",
          2771 => x"b2",
          2772 => x"e0",
          2773 => x"06",
          2774 => x"54",
          2775 => x"72",
          2776 => x"76",
          2777 => x"38",
          2778 => x"70",
          2779 => x"53",
          2780 => x"85",
          2781 => x"70",
          2782 => x"5b",
          2783 => x"81",
          2784 => x"81",
          2785 => x"76",
          2786 => x"81",
          2787 => x"38",
          2788 => x"56",
          2789 => x"83",
          2790 => x"70",
          2791 => x"80",
          2792 => x"83",
          2793 => x"dc",
          2794 => x"ec",
          2795 => x"76",
          2796 => x"05",
          2797 => x"16",
          2798 => x"56",
          2799 => x"d7",
          2800 => x"8d",
          2801 => x"72",
          2802 => x"54",
          2803 => x"57",
          2804 => x"95",
          2805 => x"73",
          2806 => x"3f",
          2807 => x"08",
          2808 => x"57",
          2809 => x"89",
          2810 => x"56",
          2811 => x"d7",
          2812 => x"76",
          2813 => x"f1",
          2814 => x"76",
          2815 => x"e9",
          2816 => x"51",
          2817 => x"81",
          2818 => x"83",
          2819 => x"53",
          2820 => x"2e",
          2821 => x"84",
          2822 => x"ca",
          2823 => x"da",
          2824 => x"e0",
          2825 => x"ff",
          2826 => x"8d",
          2827 => x"14",
          2828 => x"3f",
          2829 => x"08",
          2830 => x"15",
          2831 => x"14",
          2832 => x"34",
          2833 => x"33",
          2834 => x"81",
          2835 => x"54",
          2836 => x"72",
          2837 => x"91",
          2838 => x"ff",
          2839 => x"29",
          2840 => x"33",
          2841 => x"72",
          2842 => x"72",
          2843 => x"38",
          2844 => x"06",
          2845 => x"2e",
          2846 => x"56",
          2847 => x"80",
          2848 => x"da",
          2849 => x"ec",
          2850 => x"81",
          2851 => x"88",
          2852 => x"8f",
          2853 => x"56",
          2854 => x"38",
          2855 => x"51",
          2856 => x"81",
          2857 => x"83",
          2858 => x"55",
          2859 => x"80",
          2860 => x"da",
          2861 => x"ec",
          2862 => x"80",
          2863 => x"da",
          2864 => x"ec",
          2865 => x"ff",
          2866 => x"8d",
          2867 => x"2e",
          2868 => x"88",
          2869 => x"14",
          2870 => x"05",
          2871 => x"75",
          2872 => x"38",
          2873 => x"52",
          2874 => x"51",
          2875 => x"3f",
          2876 => x"08",
          2877 => x"e0",
          2878 => x"82",
          2879 => x"ec",
          2880 => x"ff",
          2881 => x"26",
          2882 => x"57",
          2883 => x"f5",
          2884 => x"82",
          2885 => x"f5",
          2886 => x"81",
          2887 => x"8d",
          2888 => x"2e",
          2889 => x"82",
          2890 => x"16",
          2891 => x"16",
          2892 => x"70",
          2893 => x"7a",
          2894 => x"0c",
          2895 => x"83",
          2896 => x"06",
          2897 => x"de",
          2898 => x"ae",
          2899 => x"e0",
          2900 => x"ff",
          2901 => x"56",
          2902 => x"38",
          2903 => x"38",
          2904 => x"51",
          2905 => x"81",
          2906 => x"a8",
          2907 => x"82",
          2908 => x"39",
          2909 => x"80",
          2910 => x"38",
          2911 => x"15",
          2912 => x"53",
          2913 => x"8d",
          2914 => x"15",
          2915 => x"76",
          2916 => x"51",
          2917 => x"13",
          2918 => x"8d",
          2919 => x"15",
          2920 => x"c5",
          2921 => x"90",
          2922 => x"0b",
          2923 => x"ff",
          2924 => x"15",
          2925 => x"2e",
          2926 => x"81",
          2927 => x"e4",
          2928 => x"b6",
          2929 => x"e0",
          2930 => x"ff",
          2931 => x"81",
          2932 => x"06",
          2933 => x"81",
          2934 => x"51",
          2935 => x"81",
          2936 => x"80",
          2937 => x"ec",
          2938 => x"15",
          2939 => x"14",
          2940 => x"3f",
          2941 => x"08",
          2942 => x"06",
          2943 => x"d4",
          2944 => x"81",
          2945 => x"38",
          2946 => x"d8",
          2947 => x"ec",
          2948 => x"8b",
          2949 => x"2e",
          2950 => x"b3",
          2951 => x"14",
          2952 => x"3f",
          2953 => x"08",
          2954 => x"e4",
          2955 => x"81",
          2956 => x"84",
          2957 => x"d7",
          2958 => x"ec",
          2959 => x"15",
          2960 => x"14",
          2961 => x"3f",
          2962 => x"08",
          2963 => x"76",
          2964 => x"ed",
          2965 => x"05",
          2966 => x"ed",
          2967 => x"86",
          2968 => x"0b",
          2969 => x"80",
          2970 => x"ec",
          2971 => x"3d",
          2972 => x"3d",
          2973 => x"89",
          2974 => x"2e",
          2975 => x"08",
          2976 => x"2e",
          2977 => x"33",
          2978 => x"2e",
          2979 => x"13",
          2980 => x"22",
          2981 => x"76",
          2982 => x"06",
          2983 => x"13",
          2984 => x"c0",
          2985 => x"e0",
          2986 => x"52",
          2987 => x"71",
          2988 => x"55",
          2989 => x"53",
          2990 => x"0c",
          2991 => x"ec",
          2992 => x"3d",
          2993 => x"3d",
          2994 => x"05",
          2995 => x"89",
          2996 => x"52",
          2997 => x"3f",
          2998 => x"0b",
          2999 => x"08",
          3000 => x"81",
          3001 => x"84",
          3002 => x"fc",
          3003 => x"55",
          3004 => x"2e",
          3005 => x"74",
          3006 => x"73",
          3007 => x"38",
          3008 => x"78",
          3009 => x"54",
          3010 => x"92",
          3011 => x"89",
          3012 => x"84",
          3013 => x"b0",
          3014 => x"e0",
          3015 => x"81",
          3016 => x"88",
          3017 => x"eb",
          3018 => x"02",
          3019 => x"e7",
          3020 => x"59",
          3021 => x"80",
          3022 => x"38",
          3023 => x"70",
          3024 => x"d0",
          3025 => x"3d",
          3026 => x"58",
          3027 => x"81",
          3028 => x"55",
          3029 => x"08",
          3030 => x"7a",
          3031 => x"8c",
          3032 => x"56",
          3033 => x"81",
          3034 => x"55",
          3035 => x"08",
          3036 => x"80",
          3037 => x"70",
          3038 => x"57",
          3039 => x"83",
          3040 => x"77",
          3041 => x"73",
          3042 => x"ab",
          3043 => x"2e",
          3044 => x"84",
          3045 => x"06",
          3046 => x"51",
          3047 => x"81",
          3048 => x"55",
          3049 => x"b2",
          3050 => x"06",
          3051 => x"b8",
          3052 => x"2a",
          3053 => x"51",
          3054 => x"2e",
          3055 => x"55",
          3056 => x"77",
          3057 => x"74",
          3058 => x"77",
          3059 => x"81",
          3060 => x"73",
          3061 => x"af",
          3062 => x"7a",
          3063 => x"3f",
          3064 => x"08",
          3065 => x"b2",
          3066 => x"8e",
          3067 => x"ea",
          3068 => x"a0",
          3069 => x"34",
          3070 => x"52",
          3071 => x"bd",
          3072 => x"62",
          3073 => x"d4",
          3074 => x"54",
          3075 => x"15",
          3076 => x"2e",
          3077 => x"7a",
          3078 => x"51",
          3079 => x"75",
          3080 => x"d4",
          3081 => x"be",
          3082 => x"e0",
          3083 => x"ec",
          3084 => x"ca",
          3085 => x"74",
          3086 => x"02",
          3087 => x"70",
          3088 => x"81",
          3089 => x"56",
          3090 => x"86",
          3091 => x"82",
          3092 => x"81",
          3093 => x"06",
          3094 => x"80",
          3095 => x"75",
          3096 => x"73",
          3097 => x"38",
          3098 => x"92",
          3099 => x"7a",
          3100 => x"3f",
          3101 => x"08",
          3102 => x"8c",
          3103 => x"55",
          3104 => x"08",
          3105 => x"77",
          3106 => x"81",
          3107 => x"73",
          3108 => x"38",
          3109 => x"07",
          3110 => x"11",
          3111 => x"0c",
          3112 => x"0c",
          3113 => x"52",
          3114 => x"3f",
          3115 => x"08",
          3116 => x"08",
          3117 => x"63",
          3118 => x"5a",
          3119 => x"81",
          3120 => x"81",
          3121 => x"8c",
          3122 => x"7a",
          3123 => x"17",
          3124 => x"23",
          3125 => x"34",
          3126 => x"1a",
          3127 => x"9c",
          3128 => x"0b",
          3129 => x"77",
          3130 => x"81",
          3131 => x"73",
          3132 => x"8d",
          3133 => x"e0",
          3134 => x"81",
          3135 => x"ec",
          3136 => x"1a",
          3137 => x"22",
          3138 => x"7b",
          3139 => x"a8",
          3140 => x"78",
          3141 => x"3f",
          3142 => x"08",
          3143 => x"e0",
          3144 => x"83",
          3145 => x"81",
          3146 => x"ff",
          3147 => x"06",
          3148 => x"55",
          3149 => x"56",
          3150 => x"76",
          3151 => x"51",
          3152 => x"27",
          3153 => x"70",
          3154 => x"5a",
          3155 => x"76",
          3156 => x"74",
          3157 => x"83",
          3158 => x"73",
          3159 => x"38",
          3160 => x"51",
          3161 => x"81",
          3162 => x"85",
          3163 => x"8e",
          3164 => x"2a",
          3165 => x"08",
          3166 => x"0c",
          3167 => x"79",
          3168 => x"73",
          3169 => x"0c",
          3170 => x"04",
          3171 => x"60",
          3172 => x"40",
          3173 => x"80",
          3174 => x"3d",
          3175 => x"78",
          3176 => x"3f",
          3177 => x"08",
          3178 => x"e0",
          3179 => x"91",
          3180 => x"74",
          3181 => x"38",
          3182 => x"c4",
          3183 => x"33",
          3184 => x"87",
          3185 => x"2e",
          3186 => x"95",
          3187 => x"91",
          3188 => x"56",
          3189 => x"81",
          3190 => x"34",
          3191 => x"a0",
          3192 => x"08",
          3193 => x"31",
          3194 => x"27",
          3195 => x"5c",
          3196 => x"82",
          3197 => x"19",
          3198 => x"ff",
          3199 => x"74",
          3200 => x"7e",
          3201 => x"ff",
          3202 => x"2a",
          3203 => x"79",
          3204 => x"87",
          3205 => x"08",
          3206 => x"98",
          3207 => x"78",
          3208 => x"3f",
          3209 => x"08",
          3210 => x"27",
          3211 => x"74",
          3212 => x"a3",
          3213 => x"1a",
          3214 => x"08",
          3215 => x"d4",
          3216 => x"ec",
          3217 => x"2e",
          3218 => x"81",
          3219 => x"1a",
          3220 => x"59",
          3221 => x"2e",
          3222 => x"77",
          3223 => x"11",
          3224 => x"55",
          3225 => x"85",
          3226 => x"31",
          3227 => x"76",
          3228 => x"81",
          3229 => x"ca",
          3230 => x"ec",
          3231 => x"d7",
          3232 => x"11",
          3233 => x"74",
          3234 => x"38",
          3235 => x"77",
          3236 => x"78",
          3237 => x"84",
          3238 => x"16",
          3239 => x"08",
          3240 => x"2b",
          3241 => x"cf",
          3242 => x"89",
          3243 => x"39",
          3244 => x"0c",
          3245 => x"83",
          3246 => x"80",
          3247 => x"55",
          3248 => x"83",
          3249 => x"9c",
          3250 => x"7e",
          3251 => x"3f",
          3252 => x"08",
          3253 => x"75",
          3254 => x"08",
          3255 => x"1f",
          3256 => x"7c",
          3257 => x"3f",
          3258 => x"7e",
          3259 => x"0c",
          3260 => x"1b",
          3261 => x"1c",
          3262 => x"fd",
          3263 => x"56",
          3264 => x"e0",
          3265 => x"0d",
          3266 => x"0d",
          3267 => x"64",
          3268 => x"58",
          3269 => x"90",
          3270 => x"52",
          3271 => x"d2",
          3272 => x"e0",
          3273 => x"ec",
          3274 => x"38",
          3275 => x"55",
          3276 => x"86",
          3277 => x"83",
          3278 => x"18",
          3279 => x"2a",
          3280 => x"51",
          3281 => x"56",
          3282 => x"83",
          3283 => x"39",
          3284 => x"19",
          3285 => x"83",
          3286 => x"0b",
          3287 => x"81",
          3288 => x"39",
          3289 => x"7c",
          3290 => x"74",
          3291 => x"38",
          3292 => x"7b",
          3293 => x"ec",
          3294 => x"08",
          3295 => x"06",
          3296 => x"81",
          3297 => x"8a",
          3298 => x"05",
          3299 => x"06",
          3300 => x"bf",
          3301 => x"38",
          3302 => x"55",
          3303 => x"7a",
          3304 => x"98",
          3305 => x"77",
          3306 => x"3f",
          3307 => x"08",
          3308 => x"e0",
          3309 => x"82",
          3310 => x"81",
          3311 => x"38",
          3312 => x"ff",
          3313 => x"98",
          3314 => x"18",
          3315 => x"74",
          3316 => x"7e",
          3317 => x"08",
          3318 => x"2e",
          3319 => x"8d",
          3320 => x"ce",
          3321 => x"ec",
          3322 => x"ee",
          3323 => x"08",
          3324 => x"d1",
          3325 => x"ec",
          3326 => x"2e",
          3327 => x"81",
          3328 => x"1b",
          3329 => x"5a",
          3330 => x"2e",
          3331 => x"78",
          3332 => x"11",
          3333 => x"55",
          3334 => x"85",
          3335 => x"31",
          3336 => x"76",
          3337 => x"81",
          3338 => x"c8",
          3339 => x"ec",
          3340 => x"a6",
          3341 => x"11",
          3342 => x"56",
          3343 => x"27",
          3344 => x"80",
          3345 => x"08",
          3346 => x"2b",
          3347 => x"b4",
          3348 => x"b5",
          3349 => x"80",
          3350 => x"34",
          3351 => x"56",
          3352 => x"8c",
          3353 => x"19",
          3354 => x"38",
          3355 => x"b6",
          3356 => x"e0",
          3357 => x"38",
          3358 => x"12",
          3359 => x"9c",
          3360 => x"18",
          3361 => x"06",
          3362 => x"31",
          3363 => x"76",
          3364 => x"7b",
          3365 => x"08",
          3366 => x"cd",
          3367 => x"ec",
          3368 => x"b6",
          3369 => x"7c",
          3370 => x"08",
          3371 => x"1f",
          3372 => x"cb",
          3373 => x"55",
          3374 => x"16",
          3375 => x"31",
          3376 => x"7f",
          3377 => x"94",
          3378 => x"70",
          3379 => x"8c",
          3380 => x"58",
          3381 => x"76",
          3382 => x"75",
          3383 => x"19",
          3384 => x"39",
          3385 => x"80",
          3386 => x"74",
          3387 => x"80",
          3388 => x"ec",
          3389 => x"3d",
          3390 => x"3d",
          3391 => x"3d",
          3392 => x"70",
          3393 => x"ea",
          3394 => x"e0",
          3395 => x"ec",
          3396 => x"fb",
          3397 => x"33",
          3398 => x"70",
          3399 => x"55",
          3400 => x"2e",
          3401 => x"a0",
          3402 => x"78",
          3403 => x"3f",
          3404 => x"08",
          3405 => x"e0",
          3406 => x"38",
          3407 => x"8b",
          3408 => x"07",
          3409 => x"8b",
          3410 => x"16",
          3411 => x"52",
          3412 => x"dd",
          3413 => x"16",
          3414 => x"15",
          3415 => x"3f",
          3416 => x"0a",
          3417 => x"51",
          3418 => x"76",
          3419 => x"51",
          3420 => x"78",
          3421 => x"83",
          3422 => x"51",
          3423 => x"81",
          3424 => x"90",
          3425 => x"bf",
          3426 => x"73",
          3427 => x"76",
          3428 => x"0c",
          3429 => x"04",
          3430 => x"76",
          3431 => x"fe",
          3432 => x"ec",
          3433 => x"81",
          3434 => x"9c",
          3435 => x"fc",
          3436 => x"51",
          3437 => x"81",
          3438 => x"53",
          3439 => x"08",
          3440 => x"ec",
          3441 => x"0c",
          3442 => x"e0",
          3443 => x"0d",
          3444 => x"0d",
          3445 => x"e6",
          3446 => x"52",
          3447 => x"ec",
          3448 => x"8b",
          3449 => x"e0",
          3450 => x"90",
          3451 => x"71",
          3452 => x"0c",
          3453 => x"04",
          3454 => x"80",
          3455 => x"d0",
          3456 => x"3d",
          3457 => x"3f",
          3458 => x"08",
          3459 => x"e0",
          3460 => x"38",
          3461 => x"52",
          3462 => x"05",
          3463 => x"3f",
          3464 => x"08",
          3465 => x"e0",
          3466 => x"02",
          3467 => x"33",
          3468 => x"55",
          3469 => x"25",
          3470 => x"7a",
          3471 => x"54",
          3472 => x"a2",
          3473 => x"84",
          3474 => x"06",
          3475 => x"73",
          3476 => x"38",
          3477 => x"70",
          3478 => x"a8",
          3479 => x"e0",
          3480 => x"0c",
          3481 => x"ec",
          3482 => x"2e",
          3483 => x"83",
          3484 => x"74",
          3485 => x"0c",
          3486 => x"04",
          3487 => x"6f",
          3488 => x"80",
          3489 => x"53",
          3490 => x"b8",
          3491 => x"3d",
          3492 => x"3f",
          3493 => x"08",
          3494 => x"e0",
          3495 => x"38",
          3496 => x"7c",
          3497 => x"47",
          3498 => x"54",
          3499 => x"81",
          3500 => x"52",
          3501 => x"52",
          3502 => x"3f",
          3503 => x"08",
          3504 => x"e0",
          3505 => x"38",
          3506 => x"51",
          3507 => x"81",
          3508 => x"57",
          3509 => x"08",
          3510 => x"69",
          3511 => x"da",
          3512 => x"ec",
          3513 => x"76",
          3514 => x"d5",
          3515 => x"ec",
          3516 => x"81",
          3517 => x"82",
          3518 => x"52",
          3519 => x"eb",
          3520 => x"e0",
          3521 => x"ec",
          3522 => x"38",
          3523 => x"51",
          3524 => x"73",
          3525 => x"08",
          3526 => x"76",
          3527 => x"d6",
          3528 => x"ec",
          3529 => x"81",
          3530 => x"80",
          3531 => x"76",
          3532 => x"81",
          3533 => x"82",
          3534 => x"39",
          3535 => x"38",
          3536 => x"bc",
          3537 => x"51",
          3538 => x"76",
          3539 => x"11",
          3540 => x"51",
          3541 => x"73",
          3542 => x"38",
          3543 => x"55",
          3544 => x"16",
          3545 => x"56",
          3546 => x"38",
          3547 => x"73",
          3548 => x"90",
          3549 => x"2e",
          3550 => x"16",
          3551 => x"ff",
          3552 => x"ff",
          3553 => x"58",
          3554 => x"74",
          3555 => x"75",
          3556 => x"18",
          3557 => x"58",
          3558 => x"fe",
          3559 => x"7b",
          3560 => x"06",
          3561 => x"18",
          3562 => x"58",
          3563 => x"80",
          3564 => x"90",
          3565 => x"29",
          3566 => x"05",
          3567 => x"33",
          3568 => x"56",
          3569 => x"2e",
          3570 => x"16",
          3571 => x"33",
          3572 => x"73",
          3573 => x"16",
          3574 => x"26",
          3575 => x"55",
          3576 => x"91",
          3577 => x"54",
          3578 => x"70",
          3579 => x"34",
          3580 => x"ec",
          3581 => x"70",
          3582 => x"34",
          3583 => x"09",
          3584 => x"38",
          3585 => x"39",
          3586 => x"19",
          3587 => x"33",
          3588 => x"05",
          3589 => x"78",
          3590 => x"80",
          3591 => x"81",
          3592 => x"9e",
          3593 => x"f7",
          3594 => x"7d",
          3595 => x"05",
          3596 => x"57",
          3597 => x"3f",
          3598 => x"08",
          3599 => x"e0",
          3600 => x"38",
          3601 => x"53",
          3602 => x"38",
          3603 => x"54",
          3604 => x"92",
          3605 => x"33",
          3606 => x"70",
          3607 => x"54",
          3608 => x"38",
          3609 => x"15",
          3610 => x"70",
          3611 => x"58",
          3612 => x"82",
          3613 => x"8a",
          3614 => x"89",
          3615 => x"53",
          3616 => x"b7",
          3617 => x"ff",
          3618 => x"99",
          3619 => x"ec",
          3620 => x"15",
          3621 => x"53",
          3622 => x"99",
          3623 => x"ec",
          3624 => x"26",
          3625 => x"30",
          3626 => x"70",
          3627 => x"77",
          3628 => x"18",
          3629 => x"51",
          3630 => x"88",
          3631 => x"73",
          3632 => x"52",
          3633 => x"ca",
          3634 => x"e0",
          3635 => x"ec",
          3636 => x"2e",
          3637 => x"81",
          3638 => x"ff",
          3639 => x"38",
          3640 => x"08",
          3641 => x"73",
          3642 => x"73",
          3643 => x"9c",
          3644 => x"27",
          3645 => x"75",
          3646 => x"16",
          3647 => x"17",
          3648 => x"33",
          3649 => x"70",
          3650 => x"55",
          3651 => x"80",
          3652 => x"73",
          3653 => x"cc",
          3654 => x"ec",
          3655 => x"81",
          3656 => x"94",
          3657 => x"e0",
          3658 => x"39",
          3659 => x"51",
          3660 => x"81",
          3661 => x"54",
          3662 => x"be",
          3663 => x"27",
          3664 => x"53",
          3665 => x"08",
          3666 => x"73",
          3667 => x"ff",
          3668 => x"15",
          3669 => x"16",
          3670 => x"ff",
          3671 => x"80",
          3672 => x"73",
          3673 => x"c6",
          3674 => x"ec",
          3675 => x"38",
          3676 => x"16",
          3677 => x"80",
          3678 => x"0b",
          3679 => x"81",
          3680 => x"75",
          3681 => x"ec",
          3682 => x"58",
          3683 => x"54",
          3684 => x"74",
          3685 => x"73",
          3686 => x"90",
          3687 => x"c0",
          3688 => x"90",
          3689 => x"83",
          3690 => x"72",
          3691 => x"38",
          3692 => x"08",
          3693 => x"77",
          3694 => x"80",
          3695 => x"ec",
          3696 => x"3d",
          3697 => x"3d",
          3698 => x"89",
          3699 => x"2e",
          3700 => x"80",
          3701 => x"fc",
          3702 => x"3d",
          3703 => x"e1",
          3704 => x"ec",
          3705 => x"81",
          3706 => x"80",
          3707 => x"76",
          3708 => x"75",
          3709 => x"3f",
          3710 => x"08",
          3711 => x"e0",
          3712 => x"38",
          3713 => x"70",
          3714 => x"57",
          3715 => x"a2",
          3716 => x"33",
          3717 => x"70",
          3718 => x"55",
          3719 => x"2e",
          3720 => x"16",
          3721 => x"51",
          3722 => x"81",
          3723 => x"88",
          3724 => x"54",
          3725 => x"84",
          3726 => x"52",
          3727 => x"e5",
          3728 => x"e0",
          3729 => x"84",
          3730 => x"06",
          3731 => x"55",
          3732 => x"80",
          3733 => x"80",
          3734 => x"54",
          3735 => x"e0",
          3736 => x"0d",
          3737 => x"0d",
          3738 => x"fc",
          3739 => x"52",
          3740 => x"3f",
          3741 => x"08",
          3742 => x"ec",
          3743 => x"0c",
          3744 => x"04",
          3745 => x"77",
          3746 => x"fc",
          3747 => x"53",
          3748 => x"de",
          3749 => x"e0",
          3750 => x"ec",
          3751 => x"df",
          3752 => x"38",
          3753 => x"08",
          3754 => x"cd",
          3755 => x"ec",
          3756 => x"80",
          3757 => x"ec",
          3758 => x"73",
          3759 => x"3f",
          3760 => x"08",
          3761 => x"e0",
          3762 => x"09",
          3763 => x"38",
          3764 => x"39",
          3765 => x"08",
          3766 => x"52",
          3767 => x"b3",
          3768 => x"73",
          3769 => x"3f",
          3770 => x"08",
          3771 => x"30",
          3772 => x"9f",
          3773 => x"ec",
          3774 => x"51",
          3775 => x"72",
          3776 => x"0c",
          3777 => x"04",
          3778 => x"65",
          3779 => x"89",
          3780 => x"96",
          3781 => x"df",
          3782 => x"ec",
          3783 => x"81",
          3784 => x"b2",
          3785 => x"75",
          3786 => x"3f",
          3787 => x"08",
          3788 => x"e0",
          3789 => x"02",
          3790 => x"33",
          3791 => x"55",
          3792 => x"25",
          3793 => x"55",
          3794 => x"80",
          3795 => x"76",
          3796 => x"d4",
          3797 => x"81",
          3798 => x"94",
          3799 => x"f0",
          3800 => x"65",
          3801 => x"53",
          3802 => x"05",
          3803 => x"51",
          3804 => x"81",
          3805 => x"5b",
          3806 => x"08",
          3807 => x"7c",
          3808 => x"08",
          3809 => x"fe",
          3810 => x"08",
          3811 => x"55",
          3812 => x"91",
          3813 => x"0c",
          3814 => x"81",
          3815 => x"39",
          3816 => x"c7",
          3817 => x"e0",
          3818 => x"55",
          3819 => x"2e",
          3820 => x"bf",
          3821 => x"5f",
          3822 => x"92",
          3823 => x"51",
          3824 => x"81",
          3825 => x"ff",
          3826 => x"81",
          3827 => x"81",
          3828 => x"81",
          3829 => x"30",
          3830 => x"e0",
          3831 => x"25",
          3832 => x"19",
          3833 => x"5a",
          3834 => x"08",
          3835 => x"38",
          3836 => x"a4",
          3837 => x"ec",
          3838 => x"58",
          3839 => x"77",
          3840 => x"7d",
          3841 => x"bf",
          3842 => x"ec",
          3843 => x"81",
          3844 => x"80",
          3845 => x"70",
          3846 => x"ff",
          3847 => x"56",
          3848 => x"2e",
          3849 => x"9e",
          3850 => x"51",
          3851 => x"3f",
          3852 => x"08",
          3853 => x"06",
          3854 => x"80",
          3855 => x"19",
          3856 => x"54",
          3857 => x"14",
          3858 => x"c5",
          3859 => x"e0",
          3860 => x"06",
          3861 => x"80",
          3862 => x"19",
          3863 => x"54",
          3864 => x"06",
          3865 => x"79",
          3866 => x"78",
          3867 => x"79",
          3868 => x"84",
          3869 => x"07",
          3870 => x"84",
          3871 => x"81",
          3872 => x"92",
          3873 => x"f9",
          3874 => x"8a",
          3875 => x"53",
          3876 => x"e3",
          3877 => x"ec",
          3878 => x"81",
          3879 => x"81",
          3880 => x"17",
          3881 => x"81",
          3882 => x"17",
          3883 => x"2a",
          3884 => x"51",
          3885 => x"55",
          3886 => x"81",
          3887 => x"17",
          3888 => x"8c",
          3889 => x"81",
          3890 => x"9b",
          3891 => x"e0",
          3892 => x"17",
          3893 => x"51",
          3894 => x"81",
          3895 => x"74",
          3896 => x"56",
          3897 => x"98",
          3898 => x"76",
          3899 => x"c6",
          3900 => x"e0",
          3901 => x"09",
          3902 => x"38",
          3903 => x"ec",
          3904 => x"2e",
          3905 => x"85",
          3906 => x"a3",
          3907 => x"38",
          3908 => x"ec",
          3909 => x"15",
          3910 => x"38",
          3911 => x"53",
          3912 => x"08",
          3913 => x"c3",
          3914 => x"ec",
          3915 => x"94",
          3916 => x"18",
          3917 => x"33",
          3918 => x"54",
          3919 => x"34",
          3920 => x"85",
          3921 => x"18",
          3922 => x"74",
          3923 => x"0c",
          3924 => x"04",
          3925 => x"82",
          3926 => x"ff",
          3927 => x"a1",
          3928 => x"e4",
          3929 => x"e0",
          3930 => x"ec",
          3931 => x"f5",
          3932 => x"a1",
          3933 => x"95",
          3934 => x"58",
          3935 => x"81",
          3936 => x"55",
          3937 => x"08",
          3938 => x"02",
          3939 => x"33",
          3940 => x"70",
          3941 => x"55",
          3942 => x"73",
          3943 => x"75",
          3944 => x"80",
          3945 => x"bd",
          3946 => x"d6",
          3947 => x"81",
          3948 => x"87",
          3949 => x"ad",
          3950 => x"78",
          3951 => x"3f",
          3952 => x"08",
          3953 => x"70",
          3954 => x"55",
          3955 => x"2e",
          3956 => x"78",
          3957 => x"e0",
          3958 => x"08",
          3959 => x"38",
          3960 => x"ec",
          3961 => x"76",
          3962 => x"70",
          3963 => x"b5",
          3964 => x"e0",
          3965 => x"ec",
          3966 => x"e9",
          3967 => x"e0",
          3968 => x"51",
          3969 => x"81",
          3970 => x"55",
          3971 => x"08",
          3972 => x"55",
          3973 => x"81",
          3974 => x"84",
          3975 => x"81",
          3976 => x"80",
          3977 => x"51",
          3978 => x"81",
          3979 => x"81",
          3980 => x"30",
          3981 => x"e0",
          3982 => x"25",
          3983 => x"75",
          3984 => x"38",
          3985 => x"8f",
          3986 => x"75",
          3987 => x"c1",
          3988 => x"ec",
          3989 => x"74",
          3990 => x"51",
          3991 => x"3f",
          3992 => x"08",
          3993 => x"ec",
          3994 => x"3d",
          3995 => x"3d",
          3996 => x"99",
          3997 => x"52",
          3998 => x"d8",
          3999 => x"ec",
          4000 => x"81",
          4001 => x"82",
          4002 => x"5e",
          4003 => x"3d",
          4004 => x"cf",
          4005 => x"ec",
          4006 => x"81",
          4007 => x"86",
          4008 => x"82",
          4009 => x"ec",
          4010 => x"2e",
          4011 => x"82",
          4012 => x"80",
          4013 => x"70",
          4014 => x"06",
          4015 => x"54",
          4016 => x"38",
          4017 => x"52",
          4018 => x"52",
          4019 => x"3f",
          4020 => x"08",
          4021 => x"81",
          4022 => x"83",
          4023 => x"81",
          4024 => x"81",
          4025 => x"06",
          4026 => x"54",
          4027 => x"08",
          4028 => x"81",
          4029 => x"81",
          4030 => x"39",
          4031 => x"38",
          4032 => x"08",
          4033 => x"c4",
          4034 => x"ec",
          4035 => x"81",
          4036 => x"81",
          4037 => x"53",
          4038 => x"19",
          4039 => x"8c",
          4040 => x"ae",
          4041 => x"34",
          4042 => x"0b",
          4043 => x"82",
          4044 => x"52",
          4045 => x"51",
          4046 => x"3f",
          4047 => x"b4",
          4048 => x"c9",
          4049 => x"53",
          4050 => x"53",
          4051 => x"51",
          4052 => x"3f",
          4053 => x"0b",
          4054 => x"34",
          4055 => x"80",
          4056 => x"51",
          4057 => x"78",
          4058 => x"83",
          4059 => x"51",
          4060 => x"81",
          4061 => x"54",
          4062 => x"08",
          4063 => x"88",
          4064 => x"64",
          4065 => x"ff",
          4066 => x"75",
          4067 => x"78",
          4068 => x"3f",
          4069 => x"0b",
          4070 => x"78",
          4071 => x"83",
          4072 => x"51",
          4073 => x"3f",
          4074 => x"08",
          4075 => x"80",
          4076 => x"76",
          4077 => x"ae",
          4078 => x"ec",
          4079 => x"3d",
          4080 => x"3d",
          4081 => x"84",
          4082 => x"f1",
          4083 => x"a8",
          4084 => x"05",
          4085 => x"51",
          4086 => x"81",
          4087 => x"55",
          4088 => x"08",
          4089 => x"78",
          4090 => x"08",
          4091 => x"70",
          4092 => x"b8",
          4093 => x"e0",
          4094 => x"ec",
          4095 => x"b9",
          4096 => x"9b",
          4097 => x"a0",
          4098 => x"55",
          4099 => x"38",
          4100 => x"3d",
          4101 => x"3d",
          4102 => x"51",
          4103 => x"3f",
          4104 => x"52",
          4105 => x"52",
          4106 => x"dd",
          4107 => x"08",
          4108 => x"cb",
          4109 => x"ec",
          4110 => x"81",
          4111 => x"95",
          4112 => x"2e",
          4113 => x"88",
          4114 => x"3d",
          4115 => x"38",
          4116 => x"e5",
          4117 => x"e0",
          4118 => x"09",
          4119 => x"b8",
          4120 => x"c9",
          4121 => x"ec",
          4122 => x"81",
          4123 => x"81",
          4124 => x"56",
          4125 => x"3d",
          4126 => x"52",
          4127 => x"ff",
          4128 => x"02",
          4129 => x"8b",
          4130 => x"16",
          4131 => x"2a",
          4132 => x"51",
          4133 => x"89",
          4134 => x"07",
          4135 => x"17",
          4136 => x"81",
          4137 => x"34",
          4138 => x"70",
          4139 => x"81",
          4140 => x"55",
          4141 => x"80",
          4142 => x"64",
          4143 => x"38",
          4144 => x"51",
          4145 => x"81",
          4146 => x"52",
          4147 => x"b7",
          4148 => x"55",
          4149 => x"08",
          4150 => x"dd",
          4151 => x"e0",
          4152 => x"51",
          4153 => x"3f",
          4154 => x"08",
          4155 => x"11",
          4156 => x"81",
          4157 => x"80",
          4158 => x"16",
          4159 => x"ae",
          4160 => x"06",
          4161 => x"53",
          4162 => x"51",
          4163 => x"78",
          4164 => x"83",
          4165 => x"39",
          4166 => x"08",
          4167 => x"51",
          4168 => x"81",
          4169 => x"55",
          4170 => x"08",
          4171 => x"51",
          4172 => x"3f",
          4173 => x"08",
          4174 => x"ec",
          4175 => x"3d",
          4176 => x"3d",
          4177 => x"db",
          4178 => x"84",
          4179 => x"05",
          4180 => x"82",
          4181 => x"d0",
          4182 => x"3d",
          4183 => x"3f",
          4184 => x"08",
          4185 => x"e0",
          4186 => x"38",
          4187 => x"52",
          4188 => x"05",
          4189 => x"3f",
          4190 => x"08",
          4191 => x"e0",
          4192 => x"02",
          4193 => x"33",
          4194 => x"54",
          4195 => x"aa",
          4196 => x"06",
          4197 => x"8b",
          4198 => x"06",
          4199 => x"07",
          4200 => x"56",
          4201 => x"34",
          4202 => x"0b",
          4203 => x"78",
          4204 => x"a9",
          4205 => x"e0",
          4206 => x"81",
          4207 => x"95",
          4208 => x"ef",
          4209 => x"56",
          4210 => x"3d",
          4211 => x"94",
          4212 => x"f4",
          4213 => x"e0",
          4214 => x"ec",
          4215 => x"cb",
          4216 => x"63",
          4217 => x"d4",
          4218 => x"c0",
          4219 => x"e0",
          4220 => x"ec",
          4221 => x"38",
          4222 => x"05",
          4223 => x"06",
          4224 => x"73",
          4225 => x"16",
          4226 => x"22",
          4227 => x"07",
          4228 => x"1f",
          4229 => x"c2",
          4230 => x"81",
          4231 => x"34",
          4232 => x"b3",
          4233 => x"ec",
          4234 => x"74",
          4235 => x"0c",
          4236 => x"04",
          4237 => x"69",
          4238 => x"80",
          4239 => x"d0",
          4240 => x"3d",
          4241 => x"3f",
          4242 => x"08",
          4243 => x"08",
          4244 => x"ec",
          4245 => x"80",
          4246 => x"57",
          4247 => x"81",
          4248 => x"70",
          4249 => x"55",
          4250 => x"80",
          4251 => x"5d",
          4252 => x"52",
          4253 => x"52",
          4254 => x"a9",
          4255 => x"e0",
          4256 => x"ec",
          4257 => x"d1",
          4258 => x"73",
          4259 => x"3f",
          4260 => x"08",
          4261 => x"e0",
          4262 => x"81",
          4263 => x"81",
          4264 => x"65",
          4265 => x"78",
          4266 => x"7b",
          4267 => x"55",
          4268 => x"34",
          4269 => x"8a",
          4270 => x"38",
          4271 => x"1a",
          4272 => x"34",
          4273 => x"9e",
          4274 => x"70",
          4275 => x"51",
          4276 => x"a0",
          4277 => x"8e",
          4278 => x"2e",
          4279 => x"86",
          4280 => x"34",
          4281 => x"30",
          4282 => x"80",
          4283 => x"7a",
          4284 => x"c1",
          4285 => x"2e",
          4286 => x"a0",
          4287 => x"51",
          4288 => x"3f",
          4289 => x"08",
          4290 => x"e0",
          4291 => x"7b",
          4292 => x"55",
          4293 => x"73",
          4294 => x"38",
          4295 => x"73",
          4296 => x"38",
          4297 => x"15",
          4298 => x"ff",
          4299 => x"81",
          4300 => x"7b",
          4301 => x"ec",
          4302 => x"3d",
          4303 => x"3d",
          4304 => x"9c",
          4305 => x"05",
          4306 => x"51",
          4307 => x"81",
          4308 => x"81",
          4309 => x"56",
          4310 => x"e0",
          4311 => x"38",
          4312 => x"52",
          4313 => x"52",
          4314 => x"c0",
          4315 => x"70",
          4316 => x"ff",
          4317 => x"55",
          4318 => x"27",
          4319 => x"78",
          4320 => x"ff",
          4321 => x"05",
          4322 => x"55",
          4323 => x"3f",
          4324 => x"08",
          4325 => x"38",
          4326 => x"70",
          4327 => x"ff",
          4328 => x"81",
          4329 => x"80",
          4330 => x"74",
          4331 => x"07",
          4332 => x"4e",
          4333 => x"81",
          4334 => x"55",
          4335 => x"70",
          4336 => x"06",
          4337 => x"99",
          4338 => x"e0",
          4339 => x"ff",
          4340 => x"54",
          4341 => x"27",
          4342 => x"db",
          4343 => x"55",
          4344 => x"a3",
          4345 => x"81",
          4346 => x"ff",
          4347 => x"81",
          4348 => x"93",
          4349 => x"75",
          4350 => x"76",
          4351 => x"38",
          4352 => x"77",
          4353 => x"86",
          4354 => x"39",
          4355 => x"27",
          4356 => x"88",
          4357 => x"78",
          4358 => x"5a",
          4359 => x"57",
          4360 => x"81",
          4361 => x"81",
          4362 => x"33",
          4363 => x"06",
          4364 => x"57",
          4365 => x"fe",
          4366 => x"3d",
          4367 => x"55",
          4368 => x"2e",
          4369 => x"76",
          4370 => x"38",
          4371 => x"55",
          4372 => x"33",
          4373 => x"a0",
          4374 => x"06",
          4375 => x"17",
          4376 => x"38",
          4377 => x"43",
          4378 => x"3d",
          4379 => x"ff",
          4380 => x"81",
          4381 => x"54",
          4382 => x"08",
          4383 => x"81",
          4384 => x"ff",
          4385 => x"81",
          4386 => x"54",
          4387 => x"08",
          4388 => x"80",
          4389 => x"54",
          4390 => x"80",
          4391 => x"ec",
          4392 => x"2e",
          4393 => x"80",
          4394 => x"54",
          4395 => x"80",
          4396 => x"52",
          4397 => x"bd",
          4398 => x"ec",
          4399 => x"81",
          4400 => x"b1",
          4401 => x"81",
          4402 => x"52",
          4403 => x"ab",
          4404 => x"54",
          4405 => x"15",
          4406 => x"78",
          4407 => x"ff",
          4408 => x"79",
          4409 => x"83",
          4410 => x"51",
          4411 => x"3f",
          4412 => x"08",
          4413 => x"74",
          4414 => x"0c",
          4415 => x"04",
          4416 => x"60",
          4417 => x"05",
          4418 => x"33",
          4419 => x"05",
          4420 => x"40",
          4421 => x"da",
          4422 => x"e0",
          4423 => x"ec",
          4424 => x"bd",
          4425 => x"33",
          4426 => x"b5",
          4427 => x"2e",
          4428 => x"1a",
          4429 => x"90",
          4430 => x"33",
          4431 => x"70",
          4432 => x"55",
          4433 => x"38",
          4434 => x"97",
          4435 => x"82",
          4436 => x"58",
          4437 => x"7e",
          4438 => x"70",
          4439 => x"55",
          4440 => x"56",
          4441 => x"c5",
          4442 => x"7d",
          4443 => x"70",
          4444 => x"2a",
          4445 => x"08",
          4446 => x"08",
          4447 => x"5d",
          4448 => x"77",
          4449 => x"98",
          4450 => x"26",
          4451 => x"57",
          4452 => x"59",
          4453 => x"52",
          4454 => x"ae",
          4455 => x"15",
          4456 => x"98",
          4457 => x"26",
          4458 => x"55",
          4459 => x"08",
          4460 => x"99",
          4461 => x"e0",
          4462 => x"ff",
          4463 => x"ec",
          4464 => x"38",
          4465 => x"75",
          4466 => x"81",
          4467 => x"93",
          4468 => x"80",
          4469 => x"2e",
          4470 => x"ff",
          4471 => x"58",
          4472 => x"7d",
          4473 => x"38",
          4474 => x"55",
          4475 => x"b4",
          4476 => x"56",
          4477 => x"09",
          4478 => x"38",
          4479 => x"53",
          4480 => x"51",
          4481 => x"3f",
          4482 => x"08",
          4483 => x"e0",
          4484 => x"38",
          4485 => x"ff",
          4486 => x"5c",
          4487 => x"84",
          4488 => x"5c",
          4489 => x"12",
          4490 => x"80",
          4491 => x"78",
          4492 => x"7c",
          4493 => x"90",
          4494 => x"c0",
          4495 => x"90",
          4496 => x"15",
          4497 => x"90",
          4498 => x"54",
          4499 => x"91",
          4500 => x"31",
          4501 => x"84",
          4502 => x"07",
          4503 => x"16",
          4504 => x"73",
          4505 => x"0c",
          4506 => x"04",
          4507 => x"6b",
          4508 => x"05",
          4509 => x"33",
          4510 => x"5a",
          4511 => x"bd",
          4512 => x"80",
          4513 => x"e0",
          4514 => x"f8",
          4515 => x"e0",
          4516 => x"81",
          4517 => x"70",
          4518 => x"74",
          4519 => x"38",
          4520 => x"81",
          4521 => x"81",
          4522 => x"81",
          4523 => x"ff",
          4524 => x"81",
          4525 => x"81",
          4526 => x"81",
          4527 => x"83",
          4528 => x"c0",
          4529 => x"2a",
          4530 => x"51",
          4531 => x"74",
          4532 => x"99",
          4533 => x"53",
          4534 => x"51",
          4535 => x"3f",
          4536 => x"08",
          4537 => x"55",
          4538 => x"92",
          4539 => x"80",
          4540 => x"38",
          4541 => x"06",
          4542 => x"2e",
          4543 => x"48",
          4544 => x"87",
          4545 => x"79",
          4546 => x"78",
          4547 => x"26",
          4548 => x"19",
          4549 => x"74",
          4550 => x"38",
          4551 => x"e4",
          4552 => x"2a",
          4553 => x"70",
          4554 => x"59",
          4555 => x"7a",
          4556 => x"56",
          4557 => x"80",
          4558 => x"51",
          4559 => x"74",
          4560 => x"99",
          4561 => x"53",
          4562 => x"51",
          4563 => x"3f",
          4564 => x"ec",
          4565 => x"ac",
          4566 => x"2a",
          4567 => x"81",
          4568 => x"43",
          4569 => x"83",
          4570 => x"66",
          4571 => x"60",
          4572 => x"90",
          4573 => x"31",
          4574 => x"80",
          4575 => x"8a",
          4576 => x"56",
          4577 => x"26",
          4578 => x"77",
          4579 => x"81",
          4580 => x"74",
          4581 => x"38",
          4582 => x"55",
          4583 => x"83",
          4584 => x"81",
          4585 => x"80",
          4586 => x"38",
          4587 => x"55",
          4588 => x"5e",
          4589 => x"89",
          4590 => x"5a",
          4591 => x"09",
          4592 => x"e1",
          4593 => x"38",
          4594 => x"57",
          4595 => x"dd",
          4596 => x"5a",
          4597 => x"9d",
          4598 => x"26",
          4599 => x"dd",
          4600 => x"10",
          4601 => x"22",
          4602 => x"74",
          4603 => x"38",
          4604 => x"ee",
          4605 => x"66",
          4606 => x"b1",
          4607 => x"e0",
          4608 => x"84",
          4609 => x"89",
          4610 => x"a0",
          4611 => x"81",
          4612 => x"fc",
          4613 => x"56",
          4614 => x"f0",
          4615 => x"80",
          4616 => x"d3",
          4617 => x"38",
          4618 => x"57",
          4619 => x"dd",
          4620 => x"5a",
          4621 => x"9d",
          4622 => x"26",
          4623 => x"dd",
          4624 => x"10",
          4625 => x"22",
          4626 => x"74",
          4627 => x"38",
          4628 => x"ee",
          4629 => x"66",
          4630 => x"d1",
          4631 => x"e0",
          4632 => x"05",
          4633 => x"e0",
          4634 => x"26",
          4635 => x"0b",
          4636 => x"08",
          4637 => x"e0",
          4638 => x"11",
          4639 => x"05",
          4640 => x"83",
          4641 => x"2a",
          4642 => x"a0",
          4643 => x"7d",
          4644 => x"69",
          4645 => x"05",
          4646 => x"72",
          4647 => x"5c",
          4648 => x"59",
          4649 => x"2e",
          4650 => x"89",
          4651 => x"60",
          4652 => x"84",
          4653 => x"5d",
          4654 => x"18",
          4655 => x"68",
          4656 => x"74",
          4657 => x"af",
          4658 => x"31",
          4659 => x"53",
          4660 => x"52",
          4661 => x"d5",
          4662 => x"e0",
          4663 => x"83",
          4664 => x"06",
          4665 => x"ec",
          4666 => x"ff",
          4667 => x"dd",
          4668 => x"83",
          4669 => x"2a",
          4670 => x"be",
          4671 => x"39",
          4672 => x"09",
          4673 => x"c5",
          4674 => x"f5",
          4675 => x"e0",
          4676 => x"38",
          4677 => x"79",
          4678 => x"80",
          4679 => x"38",
          4680 => x"96",
          4681 => x"06",
          4682 => x"2e",
          4683 => x"5e",
          4684 => x"81",
          4685 => x"9f",
          4686 => x"38",
          4687 => x"38",
          4688 => x"81",
          4689 => x"fc",
          4690 => x"ab",
          4691 => x"7d",
          4692 => x"81",
          4693 => x"7d",
          4694 => x"78",
          4695 => x"74",
          4696 => x"8e",
          4697 => x"9c",
          4698 => x"53",
          4699 => x"51",
          4700 => x"3f",
          4701 => x"db",
          4702 => x"51",
          4703 => x"3f",
          4704 => x"8b",
          4705 => x"a1",
          4706 => x"8d",
          4707 => x"83",
          4708 => x"52",
          4709 => x"ff",
          4710 => x"81",
          4711 => x"34",
          4712 => x"70",
          4713 => x"2a",
          4714 => x"54",
          4715 => x"1b",
          4716 => x"88",
          4717 => x"74",
          4718 => x"26",
          4719 => x"83",
          4720 => x"52",
          4721 => x"ff",
          4722 => x"8a",
          4723 => x"a0",
          4724 => x"a1",
          4725 => x"0b",
          4726 => x"bf",
          4727 => x"51",
          4728 => x"3f",
          4729 => x"9a",
          4730 => x"a0",
          4731 => x"52",
          4732 => x"ff",
          4733 => x"7d",
          4734 => x"81",
          4735 => x"38",
          4736 => x"0a",
          4737 => x"1b",
          4738 => x"ce",
          4739 => x"a4",
          4740 => x"a0",
          4741 => x"52",
          4742 => x"ff",
          4743 => x"81",
          4744 => x"51",
          4745 => x"3f",
          4746 => x"1b",
          4747 => x"8c",
          4748 => x"0b",
          4749 => x"34",
          4750 => x"c2",
          4751 => x"53",
          4752 => x"52",
          4753 => x"51",
          4754 => x"88",
          4755 => x"a7",
          4756 => x"a0",
          4757 => x"83",
          4758 => x"52",
          4759 => x"ff",
          4760 => x"ff",
          4761 => x"1c",
          4762 => x"a6",
          4763 => x"53",
          4764 => x"52",
          4765 => x"ff",
          4766 => x"82",
          4767 => x"83",
          4768 => x"52",
          4769 => x"b4",
          4770 => x"60",
          4771 => x"7e",
          4772 => x"d7",
          4773 => x"81",
          4774 => x"83",
          4775 => x"83",
          4776 => x"06",
          4777 => x"75",
          4778 => x"05",
          4779 => x"7e",
          4780 => x"b7",
          4781 => x"53",
          4782 => x"51",
          4783 => x"3f",
          4784 => x"a4",
          4785 => x"51",
          4786 => x"3f",
          4787 => x"e4",
          4788 => x"e4",
          4789 => x"9f",
          4790 => x"18",
          4791 => x"1b",
          4792 => x"f6",
          4793 => x"83",
          4794 => x"ff",
          4795 => x"82",
          4796 => x"78",
          4797 => x"c4",
          4798 => x"60",
          4799 => x"7a",
          4800 => x"ff",
          4801 => x"75",
          4802 => x"53",
          4803 => x"51",
          4804 => x"3f",
          4805 => x"52",
          4806 => x"9f",
          4807 => x"56",
          4808 => x"83",
          4809 => x"06",
          4810 => x"52",
          4811 => x"9e",
          4812 => x"52",
          4813 => x"ff",
          4814 => x"f0",
          4815 => x"1b",
          4816 => x"87",
          4817 => x"55",
          4818 => x"83",
          4819 => x"74",
          4820 => x"ff",
          4821 => x"7c",
          4822 => x"74",
          4823 => x"38",
          4824 => x"54",
          4825 => x"52",
          4826 => x"99",
          4827 => x"ec",
          4828 => x"87",
          4829 => x"53",
          4830 => x"08",
          4831 => x"ff",
          4832 => x"76",
          4833 => x"31",
          4834 => x"cd",
          4835 => x"58",
          4836 => x"ff",
          4837 => x"55",
          4838 => x"83",
          4839 => x"61",
          4840 => x"26",
          4841 => x"57",
          4842 => x"53",
          4843 => x"51",
          4844 => x"3f",
          4845 => x"08",
          4846 => x"76",
          4847 => x"31",
          4848 => x"db",
          4849 => x"7d",
          4850 => x"38",
          4851 => x"83",
          4852 => x"8a",
          4853 => x"7d",
          4854 => x"38",
          4855 => x"81",
          4856 => x"80",
          4857 => x"80",
          4858 => x"7a",
          4859 => x"bc",
          4860 => x"d5",
          4861 => x"ff",
          4862 => x"83",
          4863 => x"77",
          4864 => x"0b",
          4865 => x"81",
          4866 => x"34",
          4867 => x"34",
          4868 => x"34",
          4869 => x"56",
          4870 => x"52",
          4871 => x"f2",
          4872 => x"0b",
          4873 => x"81",
          4874 => x"82",
          4875 => x"56",
          4876 => x"34",
          4877 => x"08",
          4878 => x"60",
          4879 => x"1b",
          4880 => x"96",
          4881 => x"83",
          4882 => x"ff",
          4883 => x"81",
          4884 => x"7a",
          4885 => x"ff",
          4886 => x"81",
          4887 => x"e0",
          4888 => x"80",
          4889 => x"7e",
          4890 => x"e3",
          4891 => x"81",
          4892 => x"90",
          4893 => x"8e",
          4894 => x"81",
          4895 => x"81",
          4896 => x"56",
          4897 => x"e0",
          4898 => x"0d",
          4899 => x"0d",
          4900 => x"59",
          4901 => x"ff",
          4902 => x"57",
          4903 => x"b4",
          4904 => x"f8",
          4905 => x"81",
          4906 => x"52",
          4907 => x"dc",
          4908 => x"2e",
          4909 => x"9c",
          4910 => x"33",
          4911 => x"2e",
          4912 => x"76",
          4913 => x"58",
          4914 => x"57",
          4915 => x"09",
          4916 => x"38",
          4917 => x"78",
          4918 => x"38",
          4919 => x"81",
          4920 => x"8d",
          4921 => x"fa",
          4922 => x"70",
          4923 => x"56",
          4924 => x"2e",
          4925 => x"8e",
          4926 => x"0c",
          4927 => x"53",
          4928 => x"81",
          4929 => x"75",
          4930 => x"73",
          4931 => x"38",
          4932 => x"30",
          4933 => x"77",
          4934 => x"72",
          4935 => x"a0",
          4936 => x"06",
          4937 => x"75",
          4938 => x"57",
          4939 => x"75",
          4940 => x"e9",
          4941 => x"08",
          4942 => x"52",
          4943 => x"f6",
          4944 => x"e0",
          4945 => x"84",
          4946 => x"72",
          4947 => x"a9",
          4948 => x"70",
          4949 => x"57",
          4950 => x"27",
          4951 => x"53",
          4952 => x"e0",
          4953 => x"0d",
          4954 => x"0d",
          4955 => x"93",
          4956 => x"38",
          4957 => x"81",
          4958 => x"52",
          4959 => x"81",
          4960 => x"81",
          4961 => x"df",
          4962 => x"f9",
          4963 => x"9c",
          4964 => x"39",
          4965 => x"51",
          4966 => x"81",
          4967 => x"80",
          4968 => x"df",
          4969 => x"dd",
          4970 => x"e4",
          4971 => x"39",
          4972 => x"51",
          4973 => x"81",
          4974 => x"80",
          4975 => x"e0",
          4976 => x"c1",
          4977 => x"bc",
          4978 => x"81",
          4979 => x"b5",
          4980 => x"ec",
          4981 => x"81",
          4982 => x"a9",
          4983 => x"ac",
          4984 => x"81",
          4985 => x"9d",
          4986 => x"e0",
          4987 => x"81",
          4988 => x"91",
          4989 => x"90",
          4990 => x"81",
          4991 => x"85",
          4992 => x"b4",
          4993 => x"9f",
          4994 => x"0d",
          4995 => x"0d",
          4996 => x"56",
          4997 => x"26",
          4998 => x"52",
          4999 => x"29",
          5000 => x"87",
          5001 => x"51",
          5002 => x"3f",
          5003 => x"08",
          5004 => x"fe",
          5005 => x"81",
          5006 => x"54",
          5007 => x"52",
          5008 => x"51",
          5009 => x"3f",
          5010 => x"04",
          5011 => x"66",
          5012 => x"80",
          5013 => x"5b",
          5014 => x"78",
          5015 => x"07",
          5016 => x"57",
          5017 => x"56",
          5018 => x"26",
          5019 => x"56",
          5020 => x"70",
          5021 => x"51",
          5022 => x"74",
          5023 => x"81",
          5024 => x"8c",
          5025 => x"56",
          5026 => x"81",
          5027 => x"57",
          5028 => x"08",
          5029 => x"ec",
          5030 => x"c0",
          5031 => x"81",
          5032 => x"59",
          5033 => x"05",
          5034 => x"53",
          5035 => x"51",
          5036 => x"81",
          5037 => x"57",
          5038 => x"08",
          5039 => x"55",
          5040 => x"89",
          5041 => x"75",
          5042 => x"d8",
          5043 => x"d8",
          5044 => x"c4",
          5045 => x"70",
          5046 => x"25",
          5047 => x"9f",
          5048 => x"51",
          5049 => x"74",
          5050 => x"38",
          5051 => x"53",
          5052 => x"88",
          5053 => x"51",
          5054 => x"76",
          5055 => x"ec",
          5056 => x"3d",
          5057 => x"3d",
          5058 => x"84",
          5059 => x"33",
          5060 => x"57",
          5061 => x"52",
          5062 => x"b0",
          5063 => x"e0",
          5064 => x"75",
          5065 => x"38",
          5066 => x"98",
          5067 => x"60",
          5068 => x"81",
          5069 => x"7e",
          5070 => x"77",
          5071 => x"e0",
          5072 => x"39",
          5073 => x"81",
          5074 => x"89",
          5075 => x"f3",
          5076 => x"61",
          5077 => x"05",
          5078 => x"33",
          5079 => x"68",
          5080 => x"5c",
          5081 => x"7a",
          5082 => x"f0",
          5083 => x"9b",
          5084 => x"f8",
          5085 => x"af",
          5086 => x"74",
          5087 => x"fc",
          5088 => x"2e",
          5089 => x"a0",
          5090 => x"80",
          5091 => x"18",
          5092 => x"27",
          5093 => x"22",
          5094 => x"fc",
          5095 => x"eb",
          5096 => x"81",
          5097 => x"ff",
          5098 => x"82",
          5099 => x"c3",
          5100 => x"53",
          5101 => x"8e",
          5102 => x"52",
          5103 => x"51",
          5104 => x"3f",
          5105 => x"e3",
          5106 => x"82",
          5107 => x"15",
          5108 => x"74",
          5109 => x"7a",
          5110 => x"72",
          5111 => x"e3",
          5112 => x"88",
          5113 => x"39",
          5114 => x"51",
          5115 => x"3f",
          5116 => x"a0",
          5117 => x"d2",
          5118 => x"39",
          5119 => x"51",
          5120 => x"3f",
          5121 => x"79",
          5122 => x"74",
          5123 => x"55",
          5124 => x"72",
          5125 => x"38",
          5126 => x"53",
          5127 => x"83",
          5128 => x"75",
          5129 => x"81",
          5130 => x"53",
          5131 => x"8b",
          5132 => x"fe",
          5133 => x"73",
          5134 => x"a0",
          5135 => x"8a",
          5136 => x"55",
          5137 => x"e3",
          5138 => x"81",
          5139 => x"18",
          5140 => x"58",
          5141 => x"3f",
          5142 => x"08",
          5143 => x"98",
          5144 => x"76",
          5145 => x"81",
          5146 => x"fe",
          5147 => x"81",
          5148 => x"98",
          5149 => x"2c",
          5150 => x"70",
          5151 => x"32",
          5152 => x"72",
          5153 => x"07",
          5154 => x"58",
          5155 => x"57",
          5156 => x"d7",
          5157 => x"2e",
          5158 => x"85",
          5159 => x"8c",
          5160 => x"53",
          5161 => x"fd",
          5162 => x"53",
          5163 => x"e0",
          5164 => x"0d",
          5165 => x"0d",
          5166 => x"33",
          5167 => x"53",
          5168 => x"52",
          5169 => x"c3",
          5170 => x"c0",
          5171 => x"ff",
          5172 => x"e3",
          5173 => x"e3",
          5174 => x"e9",
          5175 => x"81",
          5176 => x"ff",
          5177 => x"74",
          5178 => x"38",
          5179 => x"3f",
          5180 => x"04",
          5181 => x"87",
          5182 => x"08",
          5183 => x"b8",
          5184 => x"fe",
          5185 => x"81",
          5186 => x"fe",
          5187 => x"80",
          5188 => x"b3",
          5189 => x"2a",
          5190 => x"51",
          5191 => x"2e",
          5192 => x"51",
          5193 => x"3f",
          5194 => x"51",
          5195 => x"3f",
          5196 => x"f1",
          5197 => x"82",
          5198 => x"06",
          5199 => x"80",
          5200 => x"81",
          5201 => x"ff",
          5202 => x"90",
          5203 => x"f7",
          5204 => x"fe",
          5205 => x"72",
          5206 => x"81",
          5207 => x"71",
          5208 => x"38",
          5209 => x"f0",
          5210 => x"e4",
          5211 => x"f2",
          5212 => x"51",
          5213 => x"3f",
          5214 => x"70",
          5215 => x"52",
          5216 => x"95",
          5217 => x"fe",
          5218 => x"81",
          5219 => x"fe",
          5220 => x"80",
          5221 => x"af",
          5222 => x"2a",
          5223 => x"51",
          5224 => x"2e",
          5225 => x"51",
          5226 => x"3f",
          5227 => x"51",
          5228 => x"3f",
          5229 => x"f0",
          5230 => x"86",
          5231 => x"06",
          5232 => x"80",
          5233 => x"81",
          5234 => x"fb",
          5235 => x"dc",
          5236 => x"f3",
          5237 => x"fe",
          5238 => x"72",
          5239 => x"81",
          5240 => x"71",
          5241 => x"38",
          5242 => x"ef",
          5243 => x"e4",
          5244 => x"f1",
          5245 => x"51",
          5246 => x"3f",
          5247 => x"70",
          5248 => x"52",
          5249 => x"95",
          5250 => x"fe",
          5251 => x"81",
          5252 => x"fe",
          5253 => x"80",
          5254 => x"ab",
          5255 => x"a0",
          5256 => x"0d",
          5257 => x"0d",
          5258 => x"55",
          5259 => x"52",
          5260 => x"e8",
          5261 => x"e9",
          5262 => x"73",
          5263 => x"53",
          5264 => x"52",
          5265 => x"51",
          5266 => x"3f",
          5267 => x"08",
          5268 => x"ec",
          5269 => x"80",
          5270 => x"31",
          5271 => x"73",
          5272 => x"34",
          5273 => x"33",
          5274 => x"2e",
          5275 => x"ac",
          5276 => x"e4",
          5277 => x"75",
          5278 => x"3f",
          5279 => x"08",
          5280 => x"38",
          5281 => x"08",
          5282 => x"9b",
          5283 => x"82",
          5284 => x"c6",
          5285 => x"0b",
          5286 => x"34",
          5287 => x"33",
          5288 => x"2e",
          5289 => x"89",
          5290 => x"75",
          5291 => x"b5",
          5292 => x"81",
          5293 => x"87",
          5294 => x"ce",
          5295 => x"70",
          5296 => x"e0",
          5297 => x"81",
          5298 => x"ff",
          5299 => x"81",
          5300 => x"81",
          5301 => x"78",
          5302 => x"81",
          5303 => x"81",
          5304 => x"96",
          5305 => x"59",
          5306 => x"3f",
          5307 => x"52",
          5308 => x"51",
          5309 => x"3f",
          5310 => x"08",
          5311 => x"38",
          5312 => x"51",
          5313 => x"81",
          5314 => x"81",
          5315 => x"fe",
          5316 => x"96",
          5317 => x"5a",
          5318 => x"79",
          5319 => x"3f",
          5320 => x"84",
          5321 => x"bf",
          5322 => x"e0",
          5323 => x"70",
          5324 => x"59",
          5325 => x"2e",
          5326 => x"78",
          5327 => x"b2",
          5328 => x"2e",
          5329 => x"78",
          5330 => x"38",
          5331 => x"ff",
          5332 => x"bc",
          5333 => x"38",
          5334 => x"78",
          5335 => x"83",
          5336 => x"80",
          5337 => x"dd",
          5338 => x"2e",
          5339 => x"8a",
          5340 => x"80",
          5341 => x"ea",
          5342 => x"f9",
          5343 => x"78",
          5344 => x"88",
          5345 => x"80",
          5346 => x"b1",
          5347 => x"39",
          5348 => x"2e",
          5349 => x"78",
          5350 => x"8b",
          5351 => x"82",
          5352 => x"38",
          5353 => x"78",
          5354 => x"8a",
          5355 => x"93",
          5356 => x"ff",
          5357 => x"ff",
          5358 => x"ff",
          5359 => x"81",
          5360 => x"80",
          5361 => x"38",
          5362 => x"fc",
          5363 => x"84",
          5364 => x"82",
          5365 => x"ec",
          5366 => x"2e",
          5367 => x"b4",
          5368 => x"11",
          5369 => x"05",
          5370 => x"94",
          5371 => x"e0",
          5372 => x"81",
          5373 => x"42",
          5374 => x"51",
          5375 => x"3f",
          5376 => x"5a",
          5377 => x"81",
          5378 => x"59",
          5379 => x"84",
          5380 => x"7a",
          5381 => x"38",
          5382 => x"b4",
          5383 => x"11",
          5384 => x"05",
          5385 => x"d8",
          5386 => x"e0",
          5387 => x"fd",
          5388 => x"3d",
          5389 => x"53",
          5390 => x"51",
          5391 => x"3f",
          5392 => x"08",
          5393 => x"c3",
          5394 => x"fe",
          5395 => x"ff",
          5396 => x"ff",
          5397 => x"81",
          5398 => x"80",
          5399 => x"38",
          5400 => x"51",
          5401 => x"3f",
          5402 => x"63",
          5403 => x"38",
          5404 => x"70",
          5405 => x"33",
          5406 => x"81",
          5407 => x"39",
          5408 => x"80",
          5409 => x"84",
          5410 => x"80",
          5411 => x"ec",
          5412 => x"2e",
          5413 => x"b4",
          5414 => x"11",
          5415 => x"05",
          5416 => x"dc",
          5417 => x"e0",
          5418 => x"fc",
          5419 => x"3d",
          5420 => x"53",
          5421 => x"51",
          5422 => x"3f",
          5423 => x"08",
          5424 => x"c7",
          5425 => x"b0",
          5426 => x"db",
          5427 => x"79",
          5428 => x"38",
          5429 => x"7b",
          5430 => x"5b",
          5431 => x"92",
          5432 => x"7a",
          5433 => x"53",
          5434 => x"e6",
          5435 => x"fe",
          5436 => x"1a",
          5437 => x"43",
          5438 => x"81",
          5439 => x"82",
          5440 => x"3d",
          5441 => x"53",
          5442 => x"51",
          5443 => x"3f",
          5444 => x"08",
          5445 => x"81",
          5446 => x"59",
          5447 => x"89",
          5448 => x"8c",
          5449 => x"cd",
          5450 => x"d5",
          5451 => x"80",
          5452 => x"81",
          5453 => x"44",
          5454 => x"e9",
          5455 => x"78",
          5456 => x"38",
          5457 => x"08",
          5458 => x"81",
          5459 => x"59",
          5460 => x"88",
          5461 => x"a4",
          5462 => x"39",
          5463 => x"33",
          5464 => x"2e",
          5465 => x"e9",
          5466 => x"89",
          5467 => x"bc",
          5468 => x"05",
          5469 => x"fe",
          5470 => x"ff",
          5471 => x"fe",
          5472 => x"81",
          5473 => x"80",
          5474 => x"e9",
          5475 => x"78",
          5476 => x"38",
          5477 => x"08",
          5478 => x"39",
          5479 => x"33",
          5480 => x"2e",
          5481 => x"e9",
          5482 => x"bb",
          5483 => x"d6",
          5484 => x"80",
          5485 => x"81",
          5486 => x"43",
          5487 => x"e9",
          5488 => x"78",
          5489 => x"38",
          5490 => x"08",
          5491 => x"81",
          5492 => x"59",
          5493 => x"88",
          5494 => x"b0",
          5495 => x"39",
          5496 => x"08",
          5497 => x"b4",
          5498 => x"11",
          5499 => x"05",
          5500 => x"8c",
          5501 => x"e0",
          5502 => x"a7",
          5503 => x"5c",
          5504 => x"2e",
          5505 => x"5c",
          5506 => x"70",
          5507 => x"07",
          5508 => x"7f",
          5509 => x"5a",
          5510 => x"2e",
          5511 => x"a0",
          5512 => x"88",
          5513 => x"dc",
          5514 => x"fb",
          5515 => x"63",
          5516 => x"62",
          5517 => x"f2",
          5518 => x"e6",
          5519 => x"f5",
          5520 => x"c7",
          5521 => x"ff",
          5522 => x"ff",
          5523 => x"fe",
          5524 => x"81",
          5525 => x"80",
          5526 => x"38",
          5527 => x"fc",
          5528 => x"84",
          5529 => x"fd",
          5530 => x"ec",
          5531 => x"2e",
          5532 => x"59",
          5533 => x"05",
          5534 => x"63",
          5535 => x"b4",
          5536 => x"11",
          5537 => x"05",
          5538 => x"f4",
          5539 => x"e0",
          5540 => x"f8",
          5541 => x"70",
          5542 => x"81",
          5543 => x"fe",
          5544 => x"80",
          5545 => x"51",
          5546 => x"3f",
          5547 => x"33",
          5548 => x"2e",
          5549 => x"9f",
          5550 => x"38",
          5551 => x"fc",
          5552 => x"84",
          5553 => x"fc",
          5554 => x"ec",
          5555 => x"2e",
          5556 => x"59",
          5557 => x"05",
          5558 => x"63",
          5559 => x"ff",
          5560 => x"e7",
          5561 => x"f4",
          5562 => x"aa",
          5563 => x"fe",
          5564 => x"ff",
          5565 => x"fe",
          5566 => x"81",
          5567 => x"80",
          5568 => x"38",
          5569 => x"f0",
          5570 => x"84",
          5571 => x"fd",
          5572 => x"ec",
          5573 => x"2e",
          5574 => x"59",
          5575 => x"22",
          5576 => x"05",
          5577 => x"41",
          5578 => x"f0",
          5579 => x"84",
          5580 => x"fd",
          5581 => x"ec",
          5582 => x"38",
          5583 => x"60",
          5584 => x"52",
          5585 => x"51",
          5586 => x"3f",
          5587 => x"79",
          5588 => x"91",
          5589 => x"79",
          5590 => x"ae",
          5591 => x"38",
          5592 => x"87",
          5593 => x"05",
          5594 => x"b4",
          5595 => x"11",
          5596 => x"05",
          5597 => x"fa",
          5598 => x"e0",
          5599 => x"92",
          5600 => x"02",
          5601 => x"79",
          5602 => x"5b",
          5603 => x"ff",
          5604 => x"e7",
          5605 => x"f3",
          5606 => x"a3",
          5607 => x"fe",
          5608 => x"ff",
          5609 => x"fe",
          5610 => x"81",
          5611 => x"80",
          5612 => x"38",
          5613 => x"f0",
          5614 => x"84",
          5615 => x"fc",
          5616 => x"ec",
          5617 => x"2e",
          5618 => x"60",
          5619 => x"60",
          5620 => x"b4",
          5621 => x"11",
          5622 => x"05",
          5623 => x"92",
          5624 => x"e0",
          5625 => x"f6",
          5626 => x"70",
          5627 => x"81",
          5628 => x"fe",
          5629 => x"80",
          5630 => x"51",
          5631 => x"3f",
          5632 => x"33",
          5633 => x"2e",
          5634 => x"9f",
          5635 => x"38",
          5636 => x"f0",
          5637 => x"84",
          5638 => x"fb",
          5639 => x"ec",
          5640 => x"2e",
          5641 => x"60",
          5642 => x"60",
          5643 => x"ff",
          5644 => x"e7",
          5645 => x"f1",
          5646 => x"ae",
          5647 => x"ff",
          5648 => x"ff",
          5649 => x"fe",
          5650 => x"81",
          5651 => x"80",
          5652 => x"38",
          5653 => x"e7",
          5654 => x"f7",
          5655 => x"59",
          5656 => x"3d",
          5657 => x"53",
          5658 => x"51",
          5659 => x"3f",
          5660 => x"08",
          5661 => x"93",
          5662 => x"81",
          5663 => x"fe",
          5664 => x"63",
          5665 => x"81",
          5666 => x"80",
          5667 => x"38",
          5668 => x"08",
          5669 => x"dc",
          5670 => x"ef",
          5671 => x"39",
          5672 => x"51",
          5673 => x"3f",
          5674 => x"3f",
          5675 => x"81",
          5676 => x"fe",
          5677 => x"80",
          5678 => x"39",
          5679 => x"3f",
          5680 => x"64",
          5681 => x"59",
          5682 => x"f4",
          5683 => x"7d",
          5684 => x"80",
          5685 => x"38",
          5686 => x"84",
          5687 => x"de",
          5688 => x"ec",
          5689 => x"81",
          5690 => x"2e",
          5691 => x"82",
          5692 => x"7a",
          5693 => x"38",
          5694 => x"7a",
          5695 => x"38",
          5696 => x"81",
          5697 => x"7b",
          5698 => x"ac",
          5699 => x"81",
          5700 => x"b4",
          5701 => x"05",
          5702 => x"85",
          5703 => x"81",
          5704 => x"b4",
          5705 => x"05",
          5706 => x"f5",
          5707 => x"7b",
          5708 => x"ac",
          5709 => x"81",
          5710 => x"b4",
          5711 => x"05",
          5712 => x"dd",
          5713 => x"7b",
          5714 => x"81",
          5715 => x"b4",
          5716 => x"05",
          5717 => x"c9",
          5718 => x"8c",
          5719 => x"94",
          5720 => x"64",
          5721 => x"81",
          5722 => x"54",
          5723 => x"53",
          5724 => x"52",
          5725 => x"b0",
          5726 => x"8a",
          5727 => x"e0",
          5728 => x"e0",
          5729 => x"30",
          5730 => x"80",
          5731 => x"5b",
          5732 => x"7a",
          5733 => x"38",
          5734 => x"7a",
          5735 => x"80",
          5736 => x"81",
          5737 => x"ff",
          5738 => x"7a",
          5739 => x"7d",
          5740 => x"81",
          5741 => x"78",
          5742 => x"ff",
          5743 => x"06",
          5744 => x"81",
          5745 => x"fe",
          5746 => x"f2",
          5747 => x"3d",
          5748 => x"81",
          5749 => x"87",
          5750 => x"70",
          5751 => x"87",
          5752 => x"72",
          5753 => x"c5",
          5754 => x"e0",
          5755 => x"75",
          5756 => x"87",
          5757 => x"73",
          5758 => x"b1",
          5759 => x"ec",
          5760 => x"75",
          5761 => x"94",
          5762 => x"54",
          5763 => x"80",
          5764 => x"fe",
          5765 => x"81",
          5766 => x"90",
          5767 => x"55",
          5768 => x"80",
          5769 => x"fe",
          5770 => x"72",
          5771 => x"08",
          5772 => x"8c",
          5773 => x"87",
          5774 => x"0c",
          5775 => x"0b",
          5776 => x"94",
          5777 => x"0b",
          5778 => x"0c",
          5779 => x"81",
          5780 => x"fe",
          5781 => x"fe",
          5782 => x"81",
          5783 => x"fe",
          5784 => x"81",
          5785 => x"fe",
          5786 => x"81",
          5787 => x"fe",
          5788 => x"81",
          5789 => x"3f",
          5790 => x"80",
          5791 => x"00",
          5792 => x"00",
          5793 => x"00",
          5794 => x"00",
          5795 => x"00",
          5796 => x"00",
          5797 => x"00",
          5798 => x"00",
          5799 => x"00",
          5800 => x"00",
          5801 => x"00",
          5802 => x"00",
          5803 => x"00",
          5804 => x"00",
          5805 => x"00",
          5806 => x"00",
          5807 => x"00",
          5808 => x"00",
          5809 => x"00",
          5810 => x"00",
          5811 => x"00",
          5812 => x"00",
          5813 => x"00",
          5814 => x"00",
          5815 => x"00",
          5816 => x"64",
          5817 => x"2f",
          5818 => x"25",
          5819 => x"64",
          5820 => x"2e",
          5821 => x"64",
          5822 => x"6f",
          5823 => x"6f",
          5824 => x"67",
          5825 => x"74",
          5826 => x"00",
          5827 => x"28",
          5828 => x"6d",
          5829 => x"43",
          5830 => x"6e",
          5831 => x"29",
          5832 => x"0a",
          5833 => x"69",
          5834 => x"20",
          5835 => x"6c",
          5836 => x"6e",
          5837 => x"3a",
          5838 => x"20",
          5839 => x"42",
          5840 => x"52",
          5841 => x"20",
          5842 => x"38",
          5843 => x"30",
          5844 => x"2e",
          5845 => x"20",
          5846 => x"44",
          5847 => x"20",
          5848 => x"20",
          5849 => x"38",
          5850 => x"30",
          5851 => x"2e",
          5852 => x"20",
          5853 => x"4e",
          5854 => x"42",
          5855 => x"20",
          5856 => x"38",
          5857 => x"30",
          5858 => x"2e",
          5859 => x"20",
          5860 => x"52",
          5861 => x"20",
          5862 => x"20",
          5863 => x"38",
          5864 => x"30",
          5865 => x"2e",
          5866 => x"20",
          5867 => x"41",
          5868 => x"20",
          5869 => x"20",
          5870 => x"38",
          5871 => x"30",
          5872 => x"2e",
          5873 => x"20",
          5874 => x"44",
          5875 => x"52",
          5876 => x"20",
          5877 => x"76",
          5878 => x"73",
          5879 => x"30",
          5880 => x"2e",
          5881 => x"20",
          5882 => x"49",
          5883 => x"31",
          5884 => x"20",
          5885 => x"6d",
          5886 => x"20",
          5887 => x"30",
          5888 => x"2e",
          5889 => x"20",
          5890 => x"4e",
          5891 => x"43",
          5892 => x"20",
          5893 => x"61",
          5894 => x"6c",
          5895 => x"30",
          5896 => x"2e",
          5897 => x"20",
          5898 => x"49",
          5899 => x"4f",
          5900 => x"42",
          5901 => x"00",
          5902 => x"20",
          5903 => x"42",
          5904 => x"43",
          5905 => x"20",
          5906 => x"4f",
          5907 => x"0a",
          5908 => x"20",
          5909 => x"53",
          5910 => x"00",
          5911 => x"20",
          5912 => x"50",
          5913 => x"00",
          5914 => x"64",
          5915 => x"73",
          5916 => x"3a",
          5917 => x"20",
          5918 => x"50",
          5919 => x"65",
          5920 => x"20",
          5921 => x"74",
          5922 => x"41",
          5923 => x"65",
          5924 => x"3d",
          5925 => x"38",
          5926 => x"00",
          5927 => x"20",
          5928 => x"50",
          5929 => x"65",
          5930 => x"79",
          5931 => x"61",
          5932 => x"41",
          5933 => x"65",
          5934 => x"3d",
          5935 => x"38",
          5936 => x"00",
          5937 => x"20",
          5938 => x"74",
          5939 => x"20",
          5940 => x"72",
          5941 => x"64",
          5942 => x"73",
          5943 => x"20",
          5944 => x"3d",
          5945 => x"38",
          5946 => x"00",
          5947 => x"69",
          5948 => x"0a",
          5949 => x"20",
          5950 => x"50",
          5951 => x"64",
          5952 => x"20",
          5953 => x"20",
          5954 => x"20",
          5955 => x"20",
          5956 => x"3d",
          5957 => x"34",
          5958 => x"00",
          5959 => x"20",
          5960 => x"79",
          5961 => x"6d",
          5962 => x"6f",
          5963 => x"46",
          5964 => x"20",
          5965 => x"20",
          5966 => x"3d",
          5967 => x"2e",
          5968 => x"64",
          5969 => x"0a",
          5970 => x"20",
          5971 => x"44",
          5972 => x"20",
          5973 => x"63",
          5974 => x"72",
          5975 => x"20",
          5976 => x"20",
          5977 => x"3d",
          5978 => x"2e",
          5979 => x"64",
          5980 => x"0a",
          5981 => x"20",
          5982 => x"69",
          5983 => x"6f",
          5984 => x"53",
          5985 => x"4d",
          5986 => x"6f",
          5987 => x"46",
          5988 => x"3d",
          5989 => x"2e",
          5990 => x"64",
          5991 => x"0a",
          5992 => x"6d",
          5993 => x"00",
          5994 => x"65",
          5995 => x"6d",
          5996 => x"6c",
          5997 => x"00",
          5998 => x"56",
          5999 => x"56",
          6000 => x"6e",
          6001 => x"6e",
          6002 => x"77",
          6003 => x"44",
          6004 => x"2a",
          6005 => x"3b",
          6006 => x"3f",
          6007 => x"7f",
          6008 => x"41",
          6009 => x"41",
          6010 => x"00",
          6011 => x"fe",
          6012 => x"44",
          6013 => x"2e",
          6014 => x"4f",
          6015 => x"4d",
          6016 => x"20",
          6017 => x"54",
          6018 => x"20",
          6019 => x"4f",
          6020 => x"4d",
          6021 => x"20",
          6022 => x"54",
          6023 => x"20",
          6024 => x"00",
          6025 => x"00",
          6026 => x"00",
          6027 => x"00",
          6028 => x"9a",
          6029 => x"41",
          6030 => x"45",
          6031 => x"49",
          6032 => x"92",
          6033 => x"4f",
          6034 => x"99",
          6035 => x"9d",
          6036 => x"49",
          6037 => x"a5",
          6038 => x"a9",
          6039 => x"ad",
          6040 => x"b1",
          6041 => x"b5",
          6042 => x"b9",
          6043 => x"bd",
          6044 => x"c1",
          6045 => x"c5",
          6046 => x"c9",
          6047 => x"cd",
          6048 => x"d1",
          6049 => x"d5",
          6050 => x"d9",
          6051 => x"dd",
          6052 => x"e1",
          6053 => x"e5",
          6054 => x"e9",
          6055 => x"ed",
          6056 => x"f1",
          6057 => x"f5",
          6058 => x"f9",
          6059 => x"fd",
          6060 => x"2e",
          6061 => x"5b",
          6062 => x"22",
          6063 => x"3e",
          6064 => x"00",
          6065 => x"01",
          6066 => x"10",
          6067 => x"00",
          6068 => x"00",
          6069 => x"01",
          6070 => x"04",
          6071 => x"10",
          6072 => x"00",
          6073 => x"69",
          6074 => x"00",
          6075 => x"69",
          6076 => x"6c",
          6077 => x"69",
          6078 => x"00",
          6079 => x"6c",
          6080 => x"00",
          6081 => x"65",
          6082 => x"00",
          6083 => x"63",
          6084 => x"72",
          6085 => x"63",
          6086 => x"00",
          6087 => x"64",
          6088 => x"00",
          6089 => x"64",
          6090 => x"00",
          6091 => x"65",
          6092 => x"65",
          6093 => x"65",
          6094 => x"69",
          6095 => x"69",
          6096 => x"66",
          6097 => x"66",
          6098 => x"61",
          6099 => x"00",
          6100 => x"6d",
          6101 => x"65",
          6102 => x"72",
          6103 => x"65",
          6104 => x"00",
          6105 => x"6e",
          6106 => x"00",
          6107 => x"65",
          6108 => x"00",
          6109 => x"62",
          6110 => x"63",
          6111 => x"69",
          6112 => x"45",
          6113 => x"72",
          6114 => x"6e",
          6115 => x"6e",
          6116 => x"65",
          6117 => x"72",
          6118 => x"00",
          6119 => x"69",
          6120 => x"6e",
          6121 => x"72",
          6122 => x"79",
          6123 => x"00",
          6124 => x"6f",
          6125 => x"6c",
          6126 => x"6f",
          6127 => x"2e",
          6128 => x"6f",
          6129 => x"74",
          6130 => x"6f",
          6131 => x"2e",
          6132 => x"6e",
          6133 => x"69",
          6134 => x"69",
          6135 => x"61",
          6136 => x"0a",
          6137 => x"63",
          6138 => x"73",
          6139 => x"6e",
          6140 => x"2e",
          6141 => x"69",
          6142 => x"61",
          6143 => x"61",
          6144 => x"65",
          6145 => x"74",
          6146 => x"00",
          6147 => x"69",
          6148 => x"68",
          6149 => x"6c",
          6150 => x"6e",
          6151 => x"69",
          6152 => x"00",
          6153 => x"44",
          6154 => x"20",
          6155 => x"74",
          6156 => x"72",
          6157 => x"63",
          6158 => x"2e",
          6159 => x"72",
          6160 => x"20",
          6161 => x"62",
          6162 => x"69",
          6163 => x"6e",
          6164 => x"69",
          6165 => x"00",
          6166 => x"69",
          6167 => x"6e",
          6168 => x"65",
          6169 => x"6c",
          6170 => x"0a",
          6171 => x"6f",
          6172 => x"6d",
          6173 => x"69",
          6174 => x"20",
          6175 => x"65",
          6176 => x"74",
          6177 => x"66",
          6178 => x"64",
          6179 => x"20",
          6180 => x"6b",
          6181 => x"00",
          6182 => x"6f",
          6183 => x"74",
          6184 => x"6f",
          6185 => x"64",
          6186 => x"00",
          6187 => x"69",
          6188 => x"75",
          6189 => x"6f",
          6190 => x"61",
          6191 => x"6e",
          6192 => x"6e",
          6193 => x"6c",
          6194 => x"0a",
          6195 => x"69",
          6196 => x"69",
          6197 => x"6f",
          6198 => x"64",
          6199 => x"00",
          6200 => x"6e",
          6201 => x"66",
          6202 => x"65",
          6203 => x"6d",
          6204 => x"72",
          6205 => x"00",
          6206 => x"6f",
          6207 => x"61",
          6208 => x"6f",
          6209 => x"20",
          6210 => x"65",
          6211 => x"00",
          6212 => x"61",
          6213 => x"65",
          6214 => x"73",
          6215 => x"63",
          6216 => x"65",
          6217 => x"0a",
          6218 => x"75",
          6219 => x"73",
          6220 => x"00",
          6221 => x"6e",
          6222 => x"77",
          6223 => x"72",
          6224 => x"2e",
          6225 => x"25",
          6226 => x"62",
          6227 => x"73",
          6228 => x"20",
          6229 => x"25",
          6230 => x"62",
          6231 => x"73",
          6232 => x"63",
          6233 => x"00",
          6234 => x"65",
          6235 => x"00",
          6236 => x"30",
          6237 => x"00",
          6238 => x"20",
          6239 => x"30",
          6240 => x"00",
          6241 => x"20",
          6242 => x"20",
          6243 => x"00",
          6244 => x"30",
          6245 => x"00",
          6246 => x"20",
          6247 => x"7c",
          6248 => x"0d",
          6249 => x"4f",
          6250 => x"2a",
          6251 => x"73",
          6252 => x"00",
          6253 => x"30",
          6254 => x"2f",
          6255 => x"30",
          6256 => x"31",
          6257 => x"00",
          6258 => x"5a",
          6259 => x"20",
          6260 => x"20",
          6261 => x"78",
          6262 => x"73",
          6263 => x"20",
          6264 => x"0a",
          6265 => x"50",
          6266 => x"6e",
          6267 => x"72",
          6268 => x"20",
          6269 => x"64",
          6270 => x"0a",
          6271 => x"69",
          6272 => x"20",
          6273 => x"65",
          6274 => x"70",
          6275 => x"00",
          6276 => x"53",
          6277 => x"6e",
          6278 => x"72",
          6279 => x"0a",
          6280 => x"4f",
          6281 => x"20",
          6282 => x"69",
          6283 => x"72",
          6284 => x"74",
          6285 => x"4f",
          6286 => x"20",
          6287 => x"69",
          6288 => x"72",
          6289 => x"74",
          6290 => x"41",
          6291 => x"20",
          6292 => x"69",
          6293 => x"72",
          6294 => x"74",
          6295 => x"41",
          6296 => x"20",
          6297 => x"69",
          6298 => x"72",
          6299 => x"74",
          6300 => x"41",
          6301 => x"20",
          6302 => x"69",
          6303 => x"72",
          6304 => x"74",
          6305 => x"41",
          6306 => x"20",
          6307 => x"69",
          6308 => x"72",
          6309 => x"74",
          6310 => x"65",
          6311 => x"6e",
          6312 => x"70",
          6313 => x"6d",
          6314 => x"2e",
          6315 => x"00",
          6316 => x"6e",
          6317 => x"69",
          6318 => x"74",
          6319 => x"72",
          6320 => x"0a",
          6321 => x"75",
          6322 => x"78",
          6323 => x"62",
          6324 => x"00",
          6325 => x"3a",
          6326 => x"61",
          6327 => x"64",
          6328 => x"20",
          6329 => x"74",
          6330 => x"69",
          6331 => x"73",
          6332 => x"61",
          6333 => x"30",
          6334 => x"6c",
          6335 => x"65",
          6336 => x"69",
          6337 => x"61",
          6338 => x"6c",
          6339 => x"0a",
          6340 => x"20",
          6341 => x"6c",
          6342 => x"69",
          6343 => x"2e",
          6344 => x"00",
          6345 => x"6f",
          6346 => x"6e",
          6347 => x"2e",
          6348 => x"6f",
          6349 => x"72",
          6350 => x"2e",
          6351 => x"00",
          6352 => x"30",
          6353 => x"28",
          6354 => x"78",
          6355 => x"25",
          6356 => x"78",
          6357 => x"38",
          6358 => x"00",
          6359 => x"75",
          6360 => x"4d",
          6361 => x"72",
          6362 => x"00",
          6363 => x"43",
          6364 => x"6c",
          6365 => x"2e",
          6366 => x"30",
          6367 => x"25",
          6368 => x"2d",
          6369 => x"3f",
          6370 => x"00",
          6371 => x"30",
          6372 => x"25",
          6373 => x"2d",
          6374 => x"30",
          6375 => x"25",
          6376 => x"2d",
          6377 => x"78",
          6378 => x"74",
          6379 => x"20",
          6380 => x"65",
          6381 => x"25",
          6382 => x"20",
          6383 => x"0a",
          6384 => x"61",
          6385 => x"6e",
          6386 => x"6f",
          6387 => x"40",
          6388 => x"38",
          6389 => x"2e",
          6390 => x"00",
          6391 => x"61",
          6392 => x"72",
          6393 => x"72",
          6394 => x"20",
          6395 => x"65",
          6396 => x"64",
          6397 => x"00",
          6398 => x"65",
          6399 => x"72",
          6400 => x"67",
          6401 => x"70",
          6402 => x"61",
          6403 => x"6e",
          6404 => x"0a",
          6405 => x"6f",
          6406 => x"72",
          6407 => x"6f",
          6408 => x"67",
          6409 => x"0a",
          6410 => x"50",
          6411 => x"69",
          6412 => x"64",
          6413 => x"73",
          6414 => x"2e",
          6415 => x"00",
          6416 => x"64",
          6417 => x"73",
          6418 => x"00",
          6419 => x"64",
          6420 => x"73",
          6421 => x"61",
          6422 => x"6f",
          6423 => x"6e",
          6424 => x"00",
          6425 => x"75",
          6426 => x"6e",
          6427 => x"2e",
          6428 => x"6e",
          6429 => x"69",
          6430 => x"69",
          6431 => x"72",
          6432 => x"74",
          6433 => x"2e",
          6434 => x"00",
          6435 => x"00",
          6436 => x"00",
          6437 => x"00",
          6438 => x"00",
          6439 => x"01",
          6440 => x"00",
          6441 => x"01",
          6442 => x"81",
          6443 => x"00",
          6444 => x"7f",
          6445 => x"00",
          6446 => x"00",
          6447 => x"00",
          6448 => x"00",
          6449 => x"f5",
          6450 => x"f5",
          6451 => x"f5",
          6452 => x"00",
          6453 => x"01",
          6454 => x"01",
          6455 => x"01",
          6456 => x"00",
          6457 => x"00",
          6458 => x"00",
          6459 => x"00",
          6460 => x"00",
          6461 => x"02",
          6462 => x"00",
          6463 => x"00",
          6464 => x"00",
          6465 => x"04",
          6466 => x"00",
          6467 => x"00",
          6468 => x"00",
          6469 => x"14",
          6470 => x"00",
          6471 => x"00",
          6472 => x"00",
          6473 => x"2b",
          6474 => x"00",
          6475 => x"00",
          6476 => x"00",
          6477 => x"30",
          6478 => x"00",
          6479 => x"00",
          6480 => x"00",
          6481 => x"3c",
          6482 => x"00",
          6483 => x"00",
          6484 => x"00",
          6485 => x"3d",
          6486 => x"00",
          6487 => x"00",
          6488 => x"00",
          6489 => x"3f",
          6490 => x"00",
          6491 => x"00",
          6492 => x"00",
          6493 => x"40",
          6494 => x"00",
          6495 => x"00",
          6496 => x"00",
          6497 => x"41",
          6498 => x"00",
          6499 => x"00",
          6500 => x"00",
          6501 => x"42",
          6502 => x"00",
          6503 => x"00",
          6504 => x"00",
          6505 => x"43",
          6506 => x"00",
          6507 => x"00",
          6508 => x"00",
          6509 => x"50",
          6510 => x"00",
          6511 => x"00",
          6512 => x"00",
          6513 => x"51",
          6514 => x"00",
          6515 => x"00",
          6516 => x"00",
          6517 => x"54",
          6518 => x"00",
          6519 => x"00",
          6520 => x"00",
          6521 => x"55",
          6522 => x"00",
          6523 => x"00",
          6524 => x"00",
          6525 => x"79",
          6526 => x"00",
          6527 => x"00",
          6528 => x"00",
          6529 => x"78",
          6530 => x"00",
          6531 => x"00",
          6532 => x"00",
          6533 => x"82",
          6534 => x"00",
          6535 => x"00",
          6536 => x"00",
          6537 => x"83",
          6538 => x"00",
          6539 => x"00",
          6540 => x"00",
          6541 => x"85",
          6542 => x"00",
          6543 => x"00",
          6544 => x"00",
          6545 => x"87",
          6546 => x"00",
          6547 => x"00",
          6548 => x"00",
          6549 => x"8c",
          6550 => x"00",
          6551 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"80",
             2 => x"0b",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"80",
            10 => x"0b",
            11 => x"0b",
            12 => x"93",
            13 => x"0b",
            14 => x"0b",
            15 => x"b3",
            16 => x"0b",
            17 => x"0b",
            18 => x"d3",
            19 => x"0b",
            20 => x"0b",
            21 => x"f3",
            22 => x"0b",
            23 => x"0b",
            24 => x"93",
            25 => x"0b",
            26 => x"0b",
            27 => x"b3",
            28 => x"0b",
            29 => x"0b",
            30 => x"d2",
            31 => x"0b",
            32 => x"0b",
            33 => x"f0",
            34 => x"0b",
            35 => x"0b",
            36 => x"8e",
            37 => x"0b",
            38 => x"0b",
            39 => x"ae",
            40 => x"0b",
            41 => x"0b",
            42 => x"ce",
            43 => x"0b",
            44 => x"0b",
            45 => x"ee",
            46 => x"0b",
            47 => x"0b",
            48 => x"8e",
            49 => x"0b",
            50 => x"0b",
            51 => x"ae",
            52 => x"0b",
            53 => x"0b",
            54 => x"ce",
            55 => x"0b",
            56 => x"0b",
            57 => x"ee",
            58 => x"0b",
            59 => x"0b",
            60 => x"8e",
            61 => x"0b",
            62 => x"0b",
            63 => x"ae",
            64 => x"0b",
            65 => x"0b",
            66 => x"ce",
            67 => x"0b",
            68 => x"0b",
            69 => x"ee",
            70 => x"0b",
            71 => x"0b",
            72 => x"8e",
            73 => x"0b",
            74 => x"0b",
            75 => x"ae",
            76 => x"0b",
            77 => x"0b",
            78 => x"ce",
            79 => x"0b",
            80 => x"0b",
            81 => x"ec",
            82 => x"0b",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"00",
           129 => x"81",
           130 => x"b4",
           131 => x"ec",
           132 => x"80",
           133 => x"ec",
           134 => x"c1",
           135 => x"ec",
           136 => x"80",
           137 => x"ec",
           138 => x"c2",
           139 => x"ec",
           140 => x"80",
           141 => x"ec",
           142 => x"c2",
           143 => x"ec",
           144 => x"80",
           145 => x"ec",
           146 => x"c8",
           147 => x"ec",
           148 => x"80",
           149 => x"ec",
           150 => x"c9",
           151 => x"ec",
           152 => x"80",
           153 => x"ec",
           154 => x"c2",
           155 => x"ec",
           156 => x"80",
           157 => x"ec",
           158 => x"c9",
           159 => x"ec",
           160 => x"80",
           161 => x"ec",
           162 => x"cb",
           163 => x"ec",
           164 => x"80",
           165 => x"ec",
           166 => x"c8",
           167 => x"ec",
           168 => x"80",
           169 => x"ec",
           170 => x"c8",
           171 => x"ec",
           172 => x"80",
           173 => x"ec",
           174 => x"c8",
           175 => x"ec",
           176 => x"80",
           177 => x"ec",
           178 => x"e0",
           179 => x"ec",
           180 => x"90",
           181 => x"ec",
           182 => x"2d",
           183 => x"08",
           184 => x"04",
           185 => x"0c",
           186 => x"81",
           187 => x"83",
           188 => x"81",
           189 => x"b1",
           190 => x"ec",
           191 => x"80",
           192 => x"ec",
           193 => x"b5",
           194 => x"ec",
           195 => x"90",
           196 => x"ec",
           197 => x"a5",
           198 => x"ec",
           199 => x"90",
           200 => x"ec",
           201 => x"96",
           202 => x"ec",
           203 => x"90",
           204 => x"ec",
           205 => x"8a",
           206 => x"ec",
           207 => x"90",
           208 => x"ec",
           209 => x"87",
           210 => x"ec",
           211 => x"90",
           212 => x"ec",
           213 => x"a5",
           214 => x"ec",
           215 => x"90",
           216 => x"ec",
           217 => x"85",
           218 => x"ec",
           219 => x"90",
           220 => x"ec",
           221 => x"f8",
           222 => x"ec",
           223 => x"90",
           224 => x"ec",
           225 => x"c4",
           226 => x"ec",
           227 => x"90",
           228 => x"ec",
           229 => x"e3",
           230 => x"ec",
           231 => x"90",
           232 => x"ec",
           233 => x"82",
           234 => x"ec",
           235 => x"90",
           236 => x"ec",
           237 => x"ec",
           238 => x"ec",
           239 => x"90",
           240 => x"ec",
           241 => x"d2",
           242 => x"ec",
           243 => x"90",
           244 => x"ec",
           245 => x"c0",
           246 => x"ec",
           247 => x"90",
           248 => x"ec",
           249 => x"86",
           250 => x"ec",
           251 => x"90",
           252 => x"ec",
           253 => x"c0",
           254 => x"ec",
           255 => x"90",
           256 => x"ec",
           257 => x"c1",
           258 => x"ec",
           259 => x"90",
           260 => x"ec",
           261 => x"f6",
           262 => x"ec",
           263 => x"90",
           264 => x"ec",
           265 => x"cf",
           266 => x"ec",
           267 => x"90",
           268 => x"ec",
           269 => x"fa",
           270 => x"ec",
           271 => x"90",
           272 => x"ec",
           273 => x"dd",
           274 => x"ec",
           275 => x"90",
           276 => x"ec",
           277 => x"b2",
           278 => x"ec",
           279 => x"90",
           280 => x"ec",
           281 => x"bc",
           282 => x"ec",
           283 => x"90",
           284 => x"ec",
           285 => x"fe",
           286 => x"ec",
           287 => x"90",
           288 => x"ec",
           289 => x"c4",
           290 => x"ec",
           291 => x"90",
           292 => x"ec",
           293 => x"ea",
           294 => x"ec",
           295 => x"90",
           296 => x"ec",
           297 => x"ff",
           298 => x"ec",
           299 => x"90",
           300 => x"ec",
           301 => x"e9",
           302 => x"ec",
           303 => x"90",
           304 => x"ec",
           305 => x"cd",
           306 => x"ec",
           307 => x"90",
           308 => x"ec",
           309 => x"2d",
           310 => x"08",
           311 => x"04",
           312 => x"0c",
           313 => x"81",
           314 => x"83",
           315 => x"81",
           316 => x"b3",
           317 => x"ec",
           318 => x"80",
           319 => x"ec",
           320 => x"ba",
           321 => x"ec",
           322 => x"80",
           323 => x"ec",
           324 => x"84",
           325 => x"38",
           326 => x"84",
           327 => x"0b",
           328 => x"8e",
           329 => x"51",
           330 => x"04",
           331 => x"ec",
           332 => x"81",
           333 => x"fd",
           334 => x"53",
           335 => x"08",
           336 => x"52",
           337 => x"08",
           338 => x"51",
           339 => x"81",
           340 => x"70",
           341 => x"0c",
           342 => x"0d",
           343 => x"0c",
           344 => x"ec",
           345 => x"ec",
           346 => x"3d",
           347 => x"81",
           348 => x"8c",
           349 => x"81",
           350 => x"88",
           351 => x"93",
           352 => x"e0",
           353 => x"ec",
           354 => x"85",
           355 => x"ec",
           356 => x"81",
           357 => x"02",
           358 => x"0c",
           359 => x"81",
           360 => x"ec",
           361 => x"0c",
           362 => x"ec",
           363 => x"05",
           364 => x"ec",
           365 => x"08",
           366 => x"08",
           367 => x"27",
           368 => x"ec",
           369 => x"05",
           370 => x"ae",
           371 => x"81",
           372 => x"8c",
           373 => x"a2",
           374 => x"ec",
           375 => x"08",
           376 => x"ec",
           377 => x"0c",
           378 => x"08",
           379 => x"10",
           380 => x"08",
           381 => x"ff",
           382 => x"ec",
           383 => x"05",
           384 => x"80",
           385 => x"ec",
           386 => x"05",
           387 => x"ec",
           388 => x"08",
           389 => x"81",
           390 => x"88",
           391 => x"ec",
           392 => x"05",
           393 => x"ec",
           394 => x"05",
           395 => x"ec",
           396 => x"08",
           397 => x"08",
           398 => x"07",
           399 => x"08",
           400 => x"81",
           401 => x"fc",
           402 => x"2a",
           403 => x"08",
           404 => x"81",
           405 => x"8c",
           406 => x"2a",
           407 => x"08",
           408 => x"ff",
           409 => x"ec",
           410 => x"05",
           411 => x"93",
           412 => x"ec",
           413 => x"08",
           414 => x"ec",
           415 => x"0c",
           416 => x"81",
           417 => x"f8",
           418 => x"81",
           419 => x"f4",
           420 => x"81",
           421 => x"f4",
           422 => x"ec",
           423 => x"3d",
           424 => x"ec",
           425 => x"3d",
           426 => x"71",
           427 => x"9f",
           428 => x"55",
           429 => x"72",
           430 => x"74",
           431 => x"70",
           432 => x"38",
           433 => x"71",
           434 => x"38",
           435 => x"81",
           436 => x"ff",
           437 => x"ff",
           438 => x"06",
           439 => x"81",
           440 => x"86",
           441 => x"74",
           442 => x"75",
           443 => x"90",
           444 => x"54",
           445 => x"27",
           446 => x"71",
           447 => x"53",
           448 => x"70",
           449 => x"0c",
           450 => x"84",
           451 => x"72",
           452 => x"05",
           453 => x"12",
           454 => x"26",
           455 => x"72",
           456 => x"72",
           457 => x"05",
           458 => x"12",
           459 => x"26",
           460 => x"53",
           461 => x"fb",
           462 => x"79",
           463 => x"83",
           464 => x"52",
           465 => x"71",
           466 => x"54",
           467 => x"73",
           468 => x"c6",
           469 => x"54",
           470 => x"70",
           471 => x"52",
           472 => x"2e",
           473 => x"33",
           474 => x"2e",
           475 => x"95",
           476 => x"81",
           477 => x"70",
           478 => x"54",
           479 => x"70",
           480 => x"33",
           481 => x"ff",
           482 => x"ff",
           483 => x"31",
           484 => x"0c",
           485 => x"3d",
           486 => x"09",
           487 => x"fd",
           488 => x"70",
           489 => x"81",
           490 => x"51",
           491 => x"38",
           492 => x"16",
           493 => x"56",
           494 => x"08",
           495 => x"73",
           496 => x"ff",
           497 => x"0b",
           498 => x"0c",
           499 => x"04",
           500 => x"80",
           501 => x"71",
           502 => x"87",
           503 => x"ec",
           504 => x"ff",
           505 => x"ff",
           506 => x"72",
           507 => x"38",
           508 => x"e0",
           509 => x"0d",
           510 => x"0d",
           511 => x"70",
           512 => x"71",
           513 => x"ca",
           514 => x"51",
           515 => x"09",
           516 => x"38",
           517 => x"f1",
           518 => x"84",
           519 => x"53",
           520 => x"70",
           521 => x"53",
           522 => x"a0",
           523 => x"81",
           524 => x"2e",
           525 => x"e5",
           526 => x"ff",
           527 => x"a0",
           528 => x"06",
           529 => x"73",
           530 => x"55",
           531 => x"0c",
           532 => x"81",
           533 => x"87",
           534 => x"fc",
           535 => x"53",
           536 => x"2e",
           537 => x"3d",
           538 => x"72",
           539 => x"3f",
           540 => x"08",
           541 => x"53",
           542 => x"53",
           543 => x"e0",
           544 => x"0d",
           545 => x"0d",
           546 => x"33",
           547 => x"53",
           548 => x"8b",
           549 => x"38",
           550 => x"ff",
           551 => x"52",
           552 => x"81",
           553 => x"13",
           554 => x"52",
           555 => x"80",
           556 => x"13",
           557 => x"52",
           558 => x"80",
           559 => x"13",
           560 => x"52",
           561 => x"80",
           562 => x"13",
           563 => x"52",
           564 => x"26",
           565 => x"8a",
           566 => x"87",
           567 => x"e7",
           568 => x"38",
           569 => x"c0",
           570 => x"72",
           571 => x"98",
           572 => x"13",
           573 => x"98",
           574 => x"13",
           575 => x"98",
           576 => x"13",
           577 => x"98",
           578 => x"13",
           579 => x"98",
           580 => x"13",
           581 => x"98",
           582 => x"87",
           583 => x"0c",
           584 => x"98",
           585 => x"0b",
           586 => x"9c",
           587 => x"71",
           588 => x"0c",
           589 => x"04",
           590 => x"7f",
           591 => x"98",
           592 => x"7d",
           593 => x"98",
           594 => x"7d",
           595 => x"c0",
           596 => x"5a",
           597 => x"34",
           598 => x"b4",
           599 => x"83",
           600 => x"c0",
           601 => x"5a",
           602 => x"34",
           603 => x"ac",
           604 => x"85",
           605 => x"c0",
           606 => x"5a",
           607 => x"34",
           608 => x"a4",
           609 => x"88",
           610 => x"c0",
           611 => x"5a",
           612 => x"23",
           613 => x"79",
           614 => x"06",
           615 => x"ff",
           616 => x"86",
           617 => x"85",
           618 => x"84",
           619 => x"83",
           620 => x"82",
           621 => x"7d",
           622 => x"06",
           623 => x"e0",
           624 => x"3f",
           625 => x"04",
           626 => x"02",
           627 => x"70",
           628 => x"2a",
           629 => x"70",
           630 => x"e9",
           631 => x"3d",
           632 => x"3d",
           633 => x"0b",
           634 => x"33",
           635 => x"06",
           636 => x"87",
           637 => x"51",
           638 => x"86",
           639 => x"94",
           640 => x"08",
           641 => x"70",
           642 => x"54",
           643 => x"2e",
           644 => x"91",
           645 => x"06",
           646 => x"d7",
           647 => x"32",
           648 => x"51",
           649 => x"2e",
           650 => x"93",
           651 => x"06",
           652 => x"ff",
           653 => x"81",
           654 => x"87",
           655 => x"52",
           656 => x"86",
           657 => x"94",
           658 => x"72",
           659 => x"ec",
           660 => x"3d",
           661 => x"3d",
           662 => x"05",
           663 => x"81",
           664 => x"70",
           665 => x"57",
           666 => x"c0",
           667 => x"74",
           668 => x"38",
           669 => x"94",
           670 => x"70",
           671 => x"81",
           672 => x"52",
           673 => x"8c",
           674 => x"2a",
           675 => x"51",
           676 => x"38",
           677 => x"70",
           678 => x"51",
           679 => x"8d",
           680 => x"2a",
           681 => x"51",
           682 => x"be",
           683 => x"ff",
           684 => x"c0",
           685 => x"70",
           686 => x"38",
           687 => x"90",
           688 => x"0c",
           689 => x"04",
           690 => x"79",
           691 => x"33",
           692 => x"06",
           693 => x"70",
           694 => x"fe",
           695 => x"ff",
           696 => x"0b",
           697 => x"88",
           698 => x"ff",
           699 => x"55",
           700 => x"94",
           701 => x"80",
           702 => x"87",
           703 => x"51",
           704 => x"96",
           705 => x"06",
           706 => x"70",
           707 => x"38",
           708 => x"70",
           709 => x"51",
           710 => x"72",
           711 => x"81",
           712 => x"70",
           713 => x"38",
           714 => x"70",
           715 => x"51",
           716 => x"38",
           717 => x"06",
           718 => x"94",
           719 => x"80",
           720 => x"87",
           721 => x"52",
           722 => x"81",
           723 => x"70",
           724 => x"53",
           725 => x"ff",
           726 => x"81",
           727 => x"89",
           728 => x"fe",
           729 => x"0b",
           730 => x"33",
           731 => x"06",
           732 => x"c0",
           733 => x"72",
           734 => x"38",
           735 => x"94",
           736 => x"70",
           737 => x"81",
           738 => x"51",
           739 => x"e2",
           740 => x"ff",
           741 => x"c0",
           742 => x"70",
           743 => x"38",
           744 => x"90",
           745 => x"70",
           746 => x"81",
           747 => x"51",
           748 => x"04",
           749 => x"0b",
           750 => x"88",
           751 => x"ff",
           752 => x"87",
           753 => x"52",
           754 => x"86",
           755 => x"94",
           756 => x"08",
           757 => x"70",
           758 => x"51",
           759 => x"70",
           760 => x"38",
           761 => x"06",
           762 => x"94",
           763 => x"80",
           764 => x"87",
           765 => x"52",
           766 => x"98",
           767 => x"2c",
           768 => x"71",
           769 => x"0c",
           770 => x"04",
           771 => x"87",
           772 => x"08",
           773 => x"8a",
           774 => x"70",
           775 => x"b4",
           776 => x"9e",
           777 => x"e9",
           778 => x"c0",
           779 => x"81",
           780 => x"87",
           781 => x"08",
           782 => x"0c",
           783 => x"98",
           784 => x"98",
           785 => x"9e",
           786 => x"e9",
           787 => x"c0",
           788 => x"81",
           789 => x"87",
           790 => x"08",
           791 => x"0c",
           792 => x"b0",
           793 => x"a8",
           794 => x"9e",
           795 => x"e9",
           796 => x"c0",
           797 => x"81",
           798 => x"87",
           799 => x"08",
           800 => x"0c",
           801 => x"c0",
           802 => x"b8",
           803 => x"9e",
           804 => x"e9",
           805 => x"c0",
           806 => x"51",
           807 => x"c0",
           808 => x"9e",
           809 => x"e9",
           810 => x"c0",
           811 => x"81",
           812 => x"87",
           813 => x"08",
           814 => x"0c",
           815 => x"e9",
           816 => x"0b",
           817 => x"90",
           818 => x"80",
           819 => x"52",
           820 => x"2e",
           821 => x"52",
           822 => x"d1",
           823 => x"87",
           824 => x"08",
           825 => x"0a",
           826 => x"52",
           827 => x"83",
           828 => x"71",
           829 => x"34",
           830 => x"c0",
           831 => x"70",
           832 => x"06",
           833 => x"70",
           834 => x"38",
           835 => x"81",
           836 => x"80",
           837 => x"9e",
           838 => x"88",
           839 => x"51",
           840 => x"80",
           841 => x"81",
           842 => x"e9",
           843 => x"0b",
           844 => x"90",
           845 => x"80",
           846 => x"52",
           847 => x"2e",
           848 => x"52",
           849 => x"d5",
           850 => x"87",
           851 => x"08",
           852 => x"80",
           853 => x"52",
           854 => x"83",
           855 => x"71",
           856 => x"34",
           857 => x"c0",
           858 => x"70",
           859 => x"06",
           860 => x"70",
           861 => x"38",
           862 => x"81",
           863 => x"80",
           864 => x"9e",
           865 => x"82",
           866 => x"51",
           867 => x"80",
           868 => x"81",
           869 => x"e9",
           870 => x"0b",
           871 => x"90",
           872 => x"80",
           873 => x"52",
           874 => x"2e",
           875 => x"52",
           876 => x"d9",
           877 => x"87",
           878 => x"08",
           879 => x"80",
           880 => x"52",
           881 => x"83",
           882 => x"71",
           883 => x"34",
           884 => x"c0",
           885 => x"70",
           886 => x"51",
           887 => x"80",
           888 => x"81",
           889 => x"e9",
           890 => x"c0",
           891 => x"70",
           892 => x"70",
           893 => x"51",
           894 => x"e9",
           895 => x"0b",
           896 => x"90",
           897 => x"80",
           898 => x"52",
           899 => x"83",
           900 => x"71",
           901 => x"34",
           902 => x"90",
           903 => x"f0",
           904 => x"2a",
           905 => x"70",
           906 => x"34",
           907 => x"c0",
           908 => x"70",
           909 => x"52",
           910 => x"2e",
           911 => x"52",
           912 => x"df",
           913 => x"9e",
           914 => x"87",
           915 => x"70",
           916 => x"34",
           917 => x"04",
           918 => x"81",
           919 => x"85",
           920 => x"e9",
           921 => x"73",
           922 => x"38",
           923 => x"51",
           924 => x"81",
           925 => x"85",
           926 => x"e9",
           927 => x"73",
           928 => x"38",
           929 => x"08",
           930 => x"08",
           931 => x"81",
           932 => x"8a",
           933 => x"e9",
           934 => x"73",
           935 => x"38",
           936 => x"08",
           937 => x"08",
           938 => x"81",
           939 => x"8a",
           940 => x"e9",
           941 => x"73",
           942 => x"38",
           943 => x"08",
           944 => x"08",
           945 => x"81",
           946 => x"8a",
           947 => x"e9",
           948 => x"73",
           949 => x"38",
           950 => x"08",
           951 => x"08",
           952 => x"81",
           953 => x"8a",
           954 => x"e9",
           955 => x"73",
           956 => x"38",
           957 => x"08",
           958 => x"08",
           959 => x"81",
           960 => x"8a",
           961 => x"e9",
           962 => x"73",
           963 => x"38",
           964 => x"33",
           965 => x"c4",
           966 => x"3f",
           967 => x"33",
           968 => x"2e",
           969 => x"e9",
           970 => x"81",
           971 => x"89",
           972 => x"e9",
           973 => x"73",
           974 => x"38",
           975 => x"33",
           976 => x"84",
           977 => x"3f",
           978 => x"33",
           979 => x"2e",
           980 => x"d8",
           981 => x"d0",
           982 => x"d3",
           983 => x"80",
           984 => x"81",
           985 => x"83",
           986 => x"e9",
           987 => x"73",
           988 => x"38",
           989 => x"51",
           990 => x"81",
           991 => x"54",
           992 => x"88",
           993 => x"d0",
           994 => x"3f",
           995 => x"33",
           996 => x"2e",
           997 => x"d8",
           998 => x"8c",
           999 => x"e8",
          1000 => x"3f",
          1001 => x"08",
          1002 => x"f4",
          1003 => x"3f",
          1004 => x"08",
          1005 => x"9c",
          1006 => x"3f",
          1007 => x"08",
          1008 => x"c4",
          1009 => x"3f",
          1010 => x"51",
          1011 => x"81",
          1012 => x"52",
          1013 => x"51",
          1014 => x"81",
          1015 => x"56",
          1016 => x"52",
          1017 => x"c6",
          1018 => x"e0",
          1019 => x"c0",
          1020 => x"31",
          1021 => x"ec",
          1022 => x"81",
          1023 => x"88",
          1024 => x"e9",
          1025 => x"73",
          1026 => x"38",
          1027 => x"08",
          1028 => x"c0",
          1029 => x"ea",
          1030 => x"ec",
          1031 => x"84",
          1032 => x"71",
          1033 => x"81",
          1034 => x"52",
          1035 => x"51",
          1036 => x"81",
          1037 => x"54",
          1038 => x"a8",
          1039 => x"cc",
          1040 => x"84",
          1041 => x"51",
          1042 => x"81",
          1043 => x"bd",
          1044 => x"76",
          1045 => x"54",
          1046 => x"08",
          1047 => x"f4",
          1048 => x"3f",
          1049 => x"51",
          1050 => x"87",
          1051 => x"fe",
          1052 => x"92",
          1053 => x"05",
          1054 => x"26",
          1055 => x"84",
          1056 => x"81",
          1057 => x"52",
          1058 => x"81",
          1059 => x"9d",
          1060 => x"a8",
          1061 => x"81",
          1062 => x"91",
          1063 => x"b8",
          1064 => x"81",
          1065 => x"85",
          1066 => x"c4",
          1067 => x"3f",
          1068 => x"04",
          1069 => x"0c",
          1070 => x"87",
          1071 => x"0c",
          1072 => x"e4",
          1073 => x"96",
          1074 => x"fe",
          1075 => x"93",
          1076 => x"72",
          1077 => x"81",
          1078 => x"8d",
          1079 => x"81",
          1080 => x"52",
          1081 => x"90",
          1082 => x"34",
          1083 => x"08",
          1084 => x"ec",
          1085 => x"39",
          1086 => x"08",
          1087 => x"2e",
          1088 => x"51",
          1089 => x"3d",
          1090 => x"3d",
          1091 => x"05",
          1092 => x"f0",
          1093 => x"ec",
          1094 => x"51",
          1095 => x"72",
          1096 => x"0c",
          1097 => x"04",
          1098 => x"75",
          1099 => x"70",
          1100 => x"53",
          1101 => x"2e",
          1102 => x"81",
          1103 => x"81",
          1104 => x"87",
          1105 => x"85",
          1106 => x"fc",
          1107 => x"81",
          1108 => x"78",
          1109 => x"0c",
          1110 => x"33",
          1111 => x"06",
          1112 => x"80",
          1113 => x"72",
          1114 => x"51",
          1115 => x"fe",
          1116 => x"39",
          1117 => x"f0",
          1118 => x"0d",
          1119 => x"0d",
          1120 => x"59",
          1121 => x"05",
          1122 => x"75",
          1123 => x"f8",
          1124 => x"2e",
          1125 => x"82",
          1126 => x"70",
          1127 => x"05",
          1128 => x"5b",
          1129 => x"2e",
          1130 => x"85",
          1131 => x"8b",
          1132 => x"2e",
          1133 => x"8a",
          1134 => x"78",
          1135 => x"5a",
          1136 => x"aa",
          1137 => x"06",
          1138 => x"84",
          1139 => x"7b",
          1140 => x"5d",
          1141 => x"59",
          1142 => x"d0",
          1143 => x"89",
          1144 => x"7a",
          1145 => x"10",
          1146 => x"d0",
          1147 => x"81",
          1148 => x"57",
          1149 => x"75",
          1150 => x"70",
          1151 => x"07",
          1152 => x"80",
          1153 => x"30",
          1154 => x"80",
          1155 => x"53",
          1156 => x"55",
          1157 => x"2e",
          1158 => x"84",
          1159 => x"81",
          1160 => x"57",
          1161 => x"2e",
          1162 => x"75",
          1163 => x"76",
          1164 => x"e0",
          1165 => x"ff",
          1166 => x"73",
          1167 => x"81",
          1168 => x"80",
          1169 => x"38",
          1170 => x"2e",
          1171 => x"73",
          1172 => x"8b",
          1173 => x"c2",
          1174 => x"38",
          1175 => x"73",
          1176 => x"81",
          1177 => x"8f",
          1178 => x"d5",
          1179 => x"38",
          1180 => x"24",
          1181 => x"80",
          1182 => x"38",
          1183 => x"73",
          1184 => x"80",
          1185 => x"ef",
          1186 => x"19",
          1187 => x"59",
          1188 => x"33",
          1189 => x"75",
          1190 => x"81",
          1191 => x"70",
          1192 => x"55",
          1193 => x"79",
          1194 => x"90",
          1195 => x"16",
          1196 => x"7b",
          1197 => x"a0",
          1198 => x"3f",
          1199 => x"53",
          1200 => x"e9",
          1201 => x"fc",
          1202 => x"81",
          1203 => x"72",
          1204 => x"b0",
          1205 => x"fb",
          1206 => x"39",
          1207 => x"83",
          1208 => x"59",
          1209 => x"82",
          1210 => x"88",
          1211 => x"8a",
          1212 => x"90",
          1213 => x"75",
          1214 => x"3f",
          1215 => x"79",
          1216 => x"81",
          1217 => x"72",
          1218 => x"38",
          1219 => x"59",
          1220 => x"84",
          1221 => x"58",
          1222 => x"80",
          1223 => x"30",
          1224 => x"80",
          1225 => x"55",
          1226 => x"25",
          1227 => x"80",
          1228 => x"74",
          1229 => x"07",
          1230 => x"0b",
          1231 => x"57",
          1232 => x"51",
          1233 => x"81",
          1234 => x"81",
          1235 => x"53",
          1236 => x"e3",
          1237 => x"ec",
          1238 => x"89",
          1239 => x"38",
          1240 => x"75",
          1241 => x"84",
          1242 => x"53",
          1243 => x"06",
          1244 => x"53",
          1245 => x"81",
          1246 => x"81",
          1247 => x"70",
          1248 => x"2a",
          1249 => x"76",
          1250 => x"38",
          1251 => x"38",
          1252 => x"70",
          1253 => x"53",
          1254 => x"8e",
          1255 => x"77",
          1256 => x"53",
          1257 => x"81",
          1258 => x"7a",
          1259 => x"55",
          1260 => x"83",
          1261 => x"79",
          1262 => x"81",
          1263 => x"72",
          1264 => x"17",
          1265 => x"27",
          1266 => x"51",
          1267 => x"75",
          1268 => x"72",
          1269 => x"81",
          1270 => x"7a",
          1271 => x"38",
          1272 => x"05",
          1273 => x"ff",
          1274 => x"70",
          1275 => x"57",
          1276 => x"76",
          1277 => x"81",
          1278 => x"72",
          1279 => x"84",
          1280 => x"f9",
          1281 => x"39",
          1282 => x"04",
          1283 => x"86",
          1284 => x"84",
          1285 => x"55",
          1286 => x"fa",
          1287 => x"3d",
          1288 => x"3d",
          1289 => x"ec",
          1290 => x"3d",
          1291 => x"75",
          1292 => x"3f",
          1293 => x"08",
          1294 => x"34",
          1295 => x"ec",
          1296 => x"3d",
          1297 => x"3d",
          1298 => x"f0",
          1299 => x"ec",
          1300 => x"3d",
          1301 => x"77",
          1302 => x"a1",
          1303 => x"ec",
          1304 => x"3d",
          1305 => x"3d",
          1306 => x"81",
          1307 => x"70",
          1308 => x"55",
          1309 => x"80",
          1310 => x"38",
          1311 => x"08",
          1312 => x"81",
          1313 => x"81",
          1314 => x"72",
          1315 => x"cb",
          1316 => x"2e",
          1317 => x"88",
          1318 => x"70",
          1319 => x"51",
          1320 => x"2e",
          1321 => x"80",
          1322 => x"ff",
          1323 => x"39",
          1324 => x"c8",
          1325 => x"52",
          1326 => x"c0",
          1327 => x"52",
          1328 => x"81",
          1329 => x"51",
          1330 => x"ff",
          1331 => x"15",
          1332 => x"34",
          1333 => x"f3",
          1334 => x"72",
          1335 => x"0c",
          1336 => x"04",
          1337 => x"81",
          1338 => x"75",
          1339 => x"0c",
          1340 => x"52",
          1341 => x"3f",
          1342 => x"f4",
          1343 => x"0d",
          1344 => x"0d",
          1345 => x"56",
          1346 => x"0c",
          1347 => x"70",
          1348 => x"73",
          1349 => x"81",
          1350 => x"81",
          1351 => x"ed",
          1352 => x"2e",
          1353 => x"8e",
          1354 => x"08",
          1355 => x"76",
          1356 => x"56",
          1357 => x"b0",
          1358 => x"06",
          1359 => x"75",
          1360 => x"76",
          1361 => x"70",
          1362 => x"73",
          1363 => x"8b",
          1364 => x"73",
          1365 => x"85",
          1366 => x"82",
          1367 => x"76",
          1368 => x"70",
          1369 => x"ac",
          1370 => x"a0",
          1371 => x"fa",
          1372 => x"53",
          1373 => x"57",
          1374 => x"98",
          1375 => x"39",
          1376 => x"80",
          1377 => x"26",
          1378 => x"86",
          1379 => x"80",
          1380 => x"57",
          1381 => x"74",
          1382 => x"38",
          1383 => x"27",
          1384 => x"14",
          1385 => x"06",
          1386 => x"14",
          1387 => x"06",
          1388 => x"74",
          1389 => x"f9",
          1390 => x"ff",
          1391 => x"89",
          1392 => x"38",
          1393 => x"c5",
          1394 => x"29",
          1395 => x"81",
          1396 => x"76",
          1397 => x"56",
          1398 => x"ba",
          1399 => x"2e",
          1400 => x"30",
          1401 => x"0c",
          1402 => x"81",
          1403 => x"8a",
          1404 => x"f8",
          1405 => x"7c",
          1406 => x"70",
          1407 => x"75",
          1408 => x"55",
          1409 => x"2e",
          1410 => x"87",
          1411 => x"76",
          1412 => x"73",
          1413 => x"81",
          1414 => x"81",
          1415 => x"77",
          1416 => x"70",
          1417 => x"58",
          1418 => x"09",
          1419 => x"c2",
          1420 => x"81",
          1421 => x"75",
          1422 => x"55",
          1423 => x"e2",
          1424 => x"90",
          1425 => x"f8",
          1426 => x"8f",
          1427 => x"81",
          1428 => x"75",
          1429 => x"55",
          1430 => x"81",
          1431 => x"27",
          1432 => x"d0",
          1433 => x"55",
          1434 => x"73",
          1435 => x"80",
          1436 => x"14",
          1437 => x"72",
          1438 => x"e0",
          1439 => x"80",
          1440 => x"39",
          1441 => x"55",
          1442 => x"80",
          1443 => x"e0",
          1444 => x"38",
          1445 => x"81",
          1446 => x"53",
          1447 => x"81",
          1448 => x"53",
          1449 => x"8e",
          1450 => x"70",
          1451 => x"55",
          1452 => x"27",
          1453 => x"77",
          1454 => x"74",
          1455 => x"76",
          1456 => x"77",
          1457 => x"70",
          1458 => x"55",
          1459 => x"77",
          1460 => x"38",
          1461 => x"74",
          1462 => x"55",
          1463 => x"e0",
          1464 => x"0d",
          1465 => x"0d",
          1466 => x"33",
          1467 => x"70",
          1468 => x"38",
          1469 => x"11",
          1470 => x"81",
          1471 => x"83",
          1472 => x"fc",
          1473 => x"9b",
          1474 => x"84",
          1475 => x"33",
          1476 => x"51",
          1477 => x"80",
          1478 => x"84",
          1479 => x"92",
          1480 => x"51",
          1481 => x"80",
          1482 => x"81",
          1483 => x"72",
          1484 => x"92",
          1485 => x"81",
          1486 => x"0b",
          1487 => x"8c",
          1488 => x"71",
          1489 => x"06",
          1490 => x"80",
          1491 => x"87",
          1492 => x"08",
          1493 => x"38",
          1494 => x"80",
          1495 => x"71",
          1496 => x"c0",
          1497 => x"51",
          1498 => x"87",
          1499 => x"e9",
          1500 => x"81",
          1501 => x"33",
          1502 => x"ec",
          1503 => x"3d",
          1504 => x"3d",
          1505 => x"64",
          1506 => x"bf",
          1507 => x"40",
          1508 => x"74",
          1509 => x"cd",
          1510 => x"e0",
          1511 => x"7a",
          1512 => x"81",
          1513 => x"72",
          1514 => x"87",
          1515 => x"11",
          1516 => x"8c",
          1517 => x"92",
          1518 => x"5a",
          1519 => x"58",
          1520 => x"c0",
          1521 => x"76",
          1522 => x"76",
          1523 => x"70",
          1524 => x"81",
          1525 => x"54",
          1526 => x"8e",
          1527 => x"52",
          1528 => x"81",
          1529 => x"81",
          1530 => x"74",
          1531 => x"53",
          1532 => x"83",
          1533 => x"78",
          1534 => x"8f",
          1535 => x"2e",
          1536 => x"c0",
          1537 => x"52",
          1538 => x"87",
          1539 => x"08",
          1540 => x"2e",
          1541 => x"84",
          1542 => x"38",
          1543 => x"87",
          1544 => x"15",
          1545 => x"70",
          1546 => x"52",
          1547 => x"ff",
          1548 => x"39",
          1549 => x"81",
          1550 => x"ff",
          1551 => x"57",
          1552 => x"90",
          1553 => x"80",
          1554 => x"71",
          1555 => x"78",
          1556 => x"38",
          1557 => x"80",
          1558 => x"80",
          1559 => x"81",
          1560 => x"72",
          1561 => x"0c",
          1562 => x"04",
          1563 => x"60",
          1564 => x"8c",
          1565 => x"33",
          1566 => x"5b",
          1567 => x"74",
          1568 => x"e1",
          1569 => x"e0",
          1570 => x"79",
          1571 => x"78",
          1572 => x"06",
          1573 => x"77",
          1574 => x"87",
          1575 => x"11",
          1576 => x"8c",
          1577 => x"92",
          1578 => x"59",
          1579 => x"85",
          1580 => x"98",
          1581 => x"7d",
          1582 => x"0c",
          1583 => x"08",
          1584 => x"70",
          1585 => x"53",
          1586 => x"2e",
          1587 => x"70",
          1588 => x"33",
          1589 => x"18",
          1590 => x"2a",
          1591 => x"51",
          1592 => x"2e",
          1593 => x"c0",
          1594 => x"52",
          1595 => x"87",
          1596 => x"08",
          1597 => x"2e",
          1598 => x"84",
          1599 => x"38",
          1600 => x"87",
          1601 => x"15",
          1602 => x"70",
          1603 => x"52",
          1604 => x"ff",
          1605 => x"39",
          1606 => x"81",
          1607 => x"80",
          1608 => x"52",
          1609 => x"90",
          1610 => x"80",
          1611 => x"71",
          1612 => x"7a",
          1613 => x"38",
          1614 => x"80",
          1615 => x"80",
          1616 => x"81",
          1617 => x"72",
          1618 => x"0c",
          1619 => x"04",
          1620 => x"7a",
          1621 => x"a3",
          1622 => x"88",
          1623 => x"33",
          1624 => x"56",
          1625 => x"3f",
          1626 => x"08",
          1627 => x"83",
          1628 => x"fe",
          1629 => x"87",
          1630 => x"0c",
          1631 => x"76",
          1632 => x"38",
          1633 => x"93",
          1634 => x"2b",
          1635 => x"8c",
          1636 => x"71",
          1637 => x"38",
          1638 => x"71",
          1639 => x"c6",
          1640 => x"39",
          1641 => x"81",
          1642 => x"06",
          1643 => x"71",
          1644 => x"38",
          1645 => x"8c",
          1646 => x"e8",
          1647 => x"98",
          1648 => x"71",
          1649 => x"73",
          1650 => x"92",
          1651 => x"72",
          1652 => x"06",
          1653 => x"f7",
          1654 => x"80",
          1655 => x"88",
          1656 => x"0c",
          1657 => x"80",
          1658 => x"56",
          1659 => x"56",
          1660 => x"81",
          1661 => x"88",
          1662 => x"fe",
          1663 => x"81",
          1664 => x"33",
          1665 => x"07",
          1666 => x"0c",
          1667 => x"3d",
          1668 => x"3d",
          1669 => x"11",
          1670 => x"33",
          1671 => x"71",
          1672 => x"81",
          1673 => x"72",
          1674 => x"75",
          1675 => x"81",
          1676 => x"52",
          1677 => x"54",
          1678 => x"0d",
          1679 => x"0d",
          1680 => x"05",
          1681 => x"52",
          1682 => x"70",
          1683 => x"34",
          1684 => x"51",
          1685 => x"83",
          1686 => x"ff",
          1687 => x"75",
          1688 => x"72",
          1689 => x"54",
          1690 => x"2a",
          1691 => x"70",
          1692 => x"34",
          1693 => x"51",
          1694 => x"81",
          1695 => x"70",
          1696 => x"70",
          1697 => x"3d",
          1698 => x"3d",
          1699 => x"77",
          1700 => x"70",
          1701 => x"38",
          1702 => x"05",
          1703 => x"70",
          1704 => x"34",
          1705 => x"eb",
          1706 => x"0d",
          1707 => x"0d",
          1708 => x"54",
          1709 => x"72",
          1710 => x"54",
          1711 => x"51",
          1712 => x"84",
          1713 => x"fc",
          1714 => x"77",
          1715 => x"53",
          1716 => x"05",
          1717 => x"70",
          1718 => x"33",
          1719 => x"ff",
          1720 => x"52",
          1721 => x"2e",
          1722 => x"80",
          1723 => x"71",
          1724 => x"0c",
          1725 => x"04",
          1726 => x"74",
          1727 => x"89",
          1728 => x"2e",
          1729 => x"11",
          1730 => x"52",
          1731 => x"70",
          1732 => x"e0",
          1733 => x"0d",
          1734 => x"81",
          1735 => x"04",
          1736 => x"ec",
          1737 => x"f7",
          1738 => x"56",
          1739 => x"17",
          1740 => x"74",
          1741 => x"d6",
          1742 => x"b0",
          1743 => x"b4",
          1744 => x"81",
          1745 => x"59",
          1746 => x"81",
          1747 => x"7a",
          1748 => x"06",
          1749 => x"ec",
          1750 => x"17",
          1751 => x"08",
          1752 => x"08",
          1753 => x"08",
          1754 => x"74",
          1755 => x"38",
          1756 => x"55",
          1757 => x"09",
          1758 => x"38",
          1759 => x"18",
          1760 => x"81",
          1761 => x"f9",
          1762 => x"39",
          1763 => x"81",
          1764 => x"8b",
          1765 => x"fa",
          1766 => x"7a",
          1767 => x"57",
          1768 => x"08",
          1769 => x"75",
          1770 => x"3f",
          1771 => x"08",
          1772 => x"e0",
          1773 => x"81",
          1774 => x"b4",
          1775 => x"16",
          1776 => x"be",
          1777 => x"e0",
          1778 => x"85",
          1779 => x"81",
          1780 => x"17",
          1781 => x"ec",
          1782 => x"3d",
          1783 => x"3d",
          1784 => x"52",
          1785 => x"3f",
          1786 => x"08",
          1787 => x"e0",
          1788 => x"38",
          1789 => x"74",
          1790 => x"81",
          1791 => x"38",
          1792 => x"59",
          1793 => x"09",
          1794 => x"e3",
          1795 => x"53",
          1796 => x"08",
          1797 => x"70",
          1798 => x"91",
          1799 => x"d5",
          1800 => x"17",
          1801 => x"3f",
          1802 => x"a4",
          1803 => x"51",
          1804 => x"86",
          1805 => x"f2",
          1806 => x"17",
          1807 => x"3f",
          1808 => x"52",
          1809 => x"51",
          1810 => x"8c",
          1811 => x"84",
          1812 => x"fc",
          1813 => x"17",
          1814 => x"70",
          1815 => x"79",
          1816 => x"52",
          1817 => x"51",
          1818 => x"77",
          1819 => x"80",
          1820 => x"81",
          1821 => x"f9",
          1822 => x"ec",
          1823 => x"2e",
          1824 => x"58",
          1825 => x"e0",
          1826 => x"0d",
          1827 => x"0d",
          1828 => x"98",
          1829 => x"05",
          1830 => x"80",
          1831 => x"27",
          1832 => x"14",
          1833 => x"29",
          1834 => x"05",
          1835 => x"81",
          1836 => x"87",
          1837 => x"f9",
          1838 => x"7a",
          1839 => x"54",
          1840 => x"27",
          1841 => x"76",
          1842 => x"27",
          1843 => x"ff",
          1844 => x"58",
          1845 => x"80",
          1846 => x"82",
          1847 => x"72",
          1848 => x"38",
          1849 => x"72",
          1850 => x"8e",
          1851 => x"39",
          1852 => x"17",
          1853 => x"a4",
          1854 => x"53",
          1855 => x"fd",
          1856 => x"ec",
          1857 => x"9f",
          1858 => x"ff",
          1859 => x"11",
          1860 => x"70",
          1861 => x"18",
          1862 => x"76",
          1863 => x"53",
          1864 => x"81",
          1865 => x"80",
          1866 => x"83",
          1867 => x"b4",
          1868 => x"88",
          1869 => x"79",
          1870 => x"84",
          1871 => x"58",
          1872 => x"80",
          1873 => x"9f",
          1874 => x"80",
          1875 => x"88",
          1876 => x"08",
          1877 => x"51",
          1878 => x"81",
          1879 => x"80",
          1880 => x"10",
          1881 => x"74",
          1882 => x"51",
          1883 => x"81",
          1884 => x"83",
          1885 => x"58",
          1886 => x"87",
          1887 => x"08",
          1888 => x"51",
          1889 => x"81",
          1890 => x"9b",
          1891 => x"2b",
          1892 => x"74",
          1893 => x"51",
          1894 => x"81",
          1895 => x"f0",
          1896 => x"83",
          1897 => x"77",
          1898 => x"0c",
          1899 => x"04",
          1900 => x"7a",
          1901 => x"58",
          1902 => x"81",
          1903 => x"9e",
          1904 => x"17",
          1905 => x"96",
          1906 => x"53",
          1907 => x"81",
          1908 => x"79",
          1909 => x"72",
          1910 => x"38",
          1911 => x"72",
          1912 => x"b8",
          1913 => x"39",
          1914 => x"17",
          1915 => x"a4",
          1916 => x"53",
          1917 => x"fb",
          1918 => x"ec",
          1919 => x"81",
          1920 => x"81",
          1921 => x"83",
          1922 => x"b4",
          1923 => x"78",
          1924 => x"56",
          1925 => x"76",
          1926 => x"38",
          1927 => x"9f",
          1928 => x"33",
          1929 => x"07",
          1930 => x"74",
          1931 => x"83",
          1932 => x"89",
          1933 => x"08",
          1934 => x"51",
          1935 => x"81",
          1936 => x"59",
          1937 => x"08",
          1938 => x"74",
          1939 => x"16",
          1940 => x"84",
          1941 => x"76",
          1942 => x"88",
          1943 => x"81",
          1944 => x"8f",
          1945 => x"53",
          1946 => x"80",
          1947 => x"88",
          1948 => x"08",
          1949 => x"51",
          1950 => x"81",
          1951 => x"59",
          1952 => x"08",
          1953 => x"77",
          1954 => x"06",
          1955 => x"83",
          1956 => x"05",
          1957 => x"f7",
          1958 => x"39",
          1959 => x"a4",
          1960 => x"52",
          1961 => x"ef",
          1962 => x"e0",
          1963 => x"ec",
          1964 => x"38",
          1965 => x"06",
          1966 => x"83",
          1967 => x"18",
          1968 => x"54",
          1969 => x"f6",
          1970 => x"ec",
          1971 => x"0a",
          1972 => x"52",
          1973 => x"83",
          1974 => x"83",
          1975 => x"81",
          1976 => x"8a",
          1977 => x"f8",
          1978 => x"7c",
          1979 => x"59",
          1980 => x"81",
          1981 => x"38",
          1982 => x"08",
          1983 => x"73",
          1984 => x"38",
          1985 => x"52",
          1986 => x"a4",
          1987 => x"e0",
          1988 => x"ec",
          1989 => x"f2",
          1990 => x"82",
          1991 => x"39",
          1992 => x"e6",
          1993 => x"e0",
          1994 => x"de",
          1995 => x"78",
          1996 => x"3f",
          1997 => x"08",
          1998 => x"e0",
          1999 => x"80",
          2000 => x"ec",
          2001 => x"2e",
          2002 => x"ec",
          2003 => x"2e",
          2004 => x"53",
          2005 => x"51",
          2006 => x"81",
          2007 => x"c5",
          2008 => x"08",
          2009 => x"18",
          2010 => x"57",
          2011 => x"90",
          2012 => x"90",
          2013 => x"16",
          2014 => x"54",
          2015 => x"34",
          2016 => x"78",
          2017 => x"38",
          2018 => x"81",
          2019 => x"8a",
          2020 => x"f6",
          2021 => x"7e",
          2022 => x"5b",
          2023 => x"38",
          2024 => x"58",
          2025 => x"88",
          2026 => x"08",
          2027 => x"38",
          2028 => x"39",
          2029 => x"51",
          2030 => x"81",
          2031 => x"ec",
          2032 => x"82",
          2033 => x"ec",
          2034 => x"81",
          2035 => x"ff",
          2036 => x"38",
          2037 => x"81",
          2038 => x"26",
          2039 => x"79",
          2040 => x"08",
          2041 => x"73",
          2042 => x"b9",
          2043 => x"2e",
          2044 => x"80",
          2045 => x"1a",
          2046 => x"08",
          2047 => x"38",
          2048 => x"52",
          2049 => x"af",
          2050 => x"81",
          2051 => x"81",
          2052 => x"06",
          2053 => x"ec",
          2054 => x"81",
          2055 => x"09",
          2056 => x"72",
          2057 => x"70",
          2058 => x"ec",
          2059 => x"51",
          2060 => x"73",
          2061 => x"81",
          2062 => x"80",
          2063 => x"8c",
          2064 => x"81",
          2065 => x"38",
          2066 => x"08",
          2067 => x"73",
          2068 => x"75",
          2069 => x"77",
          2070 => x"56",
          2071 => x"76",
          2072 => x"82",
          2073 => x"26",
          2074 => x"75",
          2075 => x"f8",
          2076 => x"ec",
          2077 => x"2e",
          2078 => x"59",
          2079 => x"08",
          2080 => x"81",
          2081 => x"81",
          2082 => x"59",
          2083 => x"08",
          2084 => x"70",
          2085 => x"25",
          2086 => x"51",
          2087 => x"73",
          2088 => x"75",
          2089 => x"81",
          2090 => x"38",
          2091 => x"f5",
          2092 => x"75",
          2093 => x"f9",
          2094 => x"ec",
          2095 => x"ec",
          2096 => x"70",
          2097 => x"08",
          2098 => x"51",
          2099 => x"80",
          2100 => x"73",
          2101 => x"38",
          2102 => x"52",
          2103 => x"d0",
          2104 => x"e0",
          2105 => x"a5",
          2106 => x"18",
          2107 => x"08",
          2108 => x"18",
          2109 => x"74",
          2110 => x"38",
          2111 => x"18",
          2112 => x"33",
          2113 => x"73",
          2114 => x"97",
          2115 => x"74",
          2116 => x"38",
          2117 => x"55",
          2118 => x"ec",
          2119 => x"85",
          2120 => x"75",
          2121 => x"ec",
          2122 => x"3d",
          2123 => x"3d",
          2124 => x"52",
          2125 => x"3f",
          2126 => x"08",
          2127 => x"81",
          2128 => x"80",
          2129 => x"52",
          2130 => x"c1",
          2131 => x"e0",
          2132 => x"e0",
          2133 => x"0c",
          2134 => x"53",
          2135 => x"15",
          2136 => x"f2",
          2137 => x"56",
          2138 => x"16",
          2139 => x"22",
          2140 => x"27",
          2141 => x"54",
          2142 => x"76",
          2143 => x"33",
          2144 => x"3f",
          2145 => x"08",
          2146 => x"38",
          2147 => x"76",
          2148 => x"70",
          2149 => x"9f",
          2150 => x"56",
          2151 => x"ec",
          2152 => x"3d",
          2153 => x"3d",
          2154 => x"71",
          2155 => x"57",
          2156 => x"0a",
          2157 => x"38",
          2158 => x"53",
          2159 => x"38",
          2160 => x"0c",
          2161 => x"54",
          2162 => x"75",
          2163 => x"73",
          2164 => x"a8",
          2165 => x"73",
          2166 => x"85",
          2167 => x"0b",
          2168 => x"5a",
          2169 => x"27",
          2170 => x"a8",
          2171 => x"18",
          2172 => x"39",
          2173 => x"70",
          2174 => x"58",
          2175 => x"b2",
          2176 => x"76",
          2177 => x"3f",
          2178 => x"08",
          2179 => x"e0",
          2180 => x"bd",
          2181 => x"81",
          2182 => x"27",
          2183 => x"16",
          2184 => x"e0",
          2185 => x"38",
          2186 => x"39",
          2187 => x"55",
          2188 => x"52",
          2189 => x"d5",
          2190 => x"e0",
          2191 => x"0c",
          2192 => x"0c",
          2193 => x"53",
          2194 => x"80",
          2195 => x"85",
          2196 => x"94",
          2197 => x"2a",
          2198 => x"0c",
          2199 => x"06",
          2200 => x"9c",
          2201 => x"58",
          2202 => x"e0",
          2203 => x"0d",
          2204 => x"0d",
          2205 => x"90",
          2206 => x"05",
          2207 => x"f0",
          2208 => x"27",
          2209 => x"0b",
          2210 => x"98",
          2211 => x"84",
          2212 => x"2e",
          2213 => x"76",
          2214 => x"58",
          2215 => x"38",
          2216 => x"15",
          2217 => x"08",
          2218 => x"38",
          2219 => x"88",
          2220 => x"53",
          2221 => x"81",
          2222 => x"c0",
          2223 => x"22",
          2224 => x"89",
          2225 => x"72",
          2226 => x"74",
          2227 => x"f3",
          2228 => x"ec",
          2229 => x"82",
          2230 => x"81",
          2231 => x"27",
          2232 => x"81",
          2233 => x"e0",
          2234 => x"80",
          2235 => x"16",
          2236 => x"e0",
          2237 => x"ca",
          2238 => x"38",
          2239 => x"0c",
          2240 => x"dd",
          2241 => x"08",
          2242 => x"f9",
          2243 => x"ec",
          2244 => x"87",
          2245 => x"e0",
          2246 => x"80",
          2247 => x"55",
          2248 => x"08",
          2249 => x"38",
          2250 => x"ec",
          2251 => x"2e",
          2252 => x"ec",
          2253 => x"75",
          2254 => x"3f",
          2255 => x"08",
          2256 => x"94",
          2257 => x"52",
          2258 => x"c1",
          2259 => x"e0",
          2260 => x"0c",
          2261 => x"0c",
          2262 => x"05",
          2263 => x"80",
          2264 => x"ec",
          2265 => x"3d",
          2266 => x"3d",
          2267 => x"71",
          2268 => x"57",
          2269 => x"51",
          2270 => x"81",
          2271 => x"54",
          2272 => x"08",
          2273 => x"81",
          2274 => x"56",
          2275 => x"52",
          2276 => x"83",
          2277 => x"e0",
          2278 => x"ec",
          2279 => x"d2",
          2280 => x"e0",
          2281 => x"08",
          2282 => x"54",
          2283 => x"e5",
          2284 => x"06",
          2285 => x"58",
          2286 => x"08",
          2287 => x"38",
          2288 => x"75",
          2289 => x"80",
          2290 => x"81",
          2291 => x"7a",
          2292 => x"06",
          2293 => x"39",
          2294 => x"08",
          2295 => x"76",
          2296 => x"3f",
          2297 => x"08",
          2298 => x"e0",
          2299 => x"ff",
          2300 => x"84",
          2301 => x"06",
          2302 => x"54",
          2303 => x"e0",
          2304 => x"0d",
          2305 => x"0d",
          2306 => x"52",
          2307 => x"3f",
          2308 => x"08",
          2309 => x"06",
          2310 => x"51",
          2311 => x"83",
          2312 => x"06",
          2313 => x"14",
          2314 => x"3f",
          2315 => x"08",
          2316 => x"07",
          2317 => x"ec",
          2318 => x"3d",
          2319 => x"3d",
          2320 => x"70",
          2321 => x"06",
          2322 => x"53",
          2323 => x"ed",
          2324 => x"33",
          2325 => x"83",
          2326 => x"06",
          2327 => x"90",
          2328 => x"15",
          2329 => x"3f",
          2330 => x"04",
          2331 => x"7b",
          2332 => x"84",
          2333 => x"58",
          2334 => x"80",
          2335 => x"38",
          2336 => x"52",
          2337 => x"8f",
          2338 => x"e0",
          2339 => x"ec",
          2340 => x"f5",
          2341 => x"08",
          2342 => x"53",
          2343 => x"84",
          2344 => x"39",
          2345 => x"70",
          2346 => x"81",
          2347 => x"51",
          2348 => x"16",
          2349 => x"e0",
          2350 => x"81",
          2351 => x"38",
          2352 => x"ae",
          2353 => x"81",
          2354 => x"54",
          2355 => x"2e",
          2356 => x"8f",
          2357 => x"81",
          2358 => x"76",
          2359 => x"54",
          2360 => x"09",
          2361 => x"38",
          2362 => x"7a",
          2363 => x"80",
          2364 => x"fa",
          2365 => x"ec",
          2366 => x"81",
          2367 => x"89",
          2368 => x"08",
          2369 => x"86",
          2370 => x"98",
          2371 => x"81",
          2372 => x"8b",
          2373 => x"fb",
          2374 => x"70",
          2375 => x"81",
          2376 => x"fc",
          2377 => x"ec",
          2378 => x"81",
          2379 => x"b4",
          2380 => x"08",
          2381 => x"ec",
          2382 => x"ec",
          2383 => x"81",
          2384 => x"a0",
          2385 => x"81",
          2386 => x"52",
          2387 => x"51",
          2388 => x"8b",
          2389 => x"52",
          2390 => x"51",
          2391 => x"81",
          2392 => x"34",
          2393 => x"e0",
          2394 => x"0d",
          2395 => x"0d",
          2396 => x"98",
          2397 => x"70",
          2398 => x"ec",
          2399 => x"ec",
          2400 => x"38",
          2401 => x"53",
          2402 => x"81",
          2403 => x"34",
          2404 => x"04",
          2405 => x"78",
          2406 => x"80",
          2407 => x"34",
          2408 => x"80",
          2409 => x"38",
          2410 => x"18",
          2411 => x"9c",
          2412 => x"70",
          2413 => x"56",
          2414 => x"a0",
          2415 => x"71",
          2416 => x"81",
          2417 => x"81",
          2418 => x"89",
          2419 => x"06",
          2420 => x"73",
          2421 => x"55",
          2422 => x"55",
          2423 => x"81",
          2424 => x"81",
          2425 => x"74",
          2426 => x"75",
          2427 => x"52",
          2428 => x"13",
          2429 => x"08",
          2430 => x"33",
          2431 => x"9c",
          2432 => x"11",
          2433 => x"8a",
          2434 => x"e0",
          2435 => x"96",
          2436 => x"e7",
          2437 => x"e0",
          2438 => x"23",
          2439 => x"e7",
          2440 => x"ec",
          2441 => x"17",
          2442 => x"0d",
          2443 => x"0d",
          2444 => x"5e",
          2445 => x"70",
          2446 => x"55",
          2447 => x"83",
          2448 => x"73",
          2449 => x"91",
          2450 => x"2e",
          2451 => x"1d",
          2452 => x"0c",
          2453 => x"15",
          2454 => x"70",
          2455 => x"56",
          2456 => x"09",
          2457 => x"38",
          2458 => x"80",
          2459 => x"30",
          2460 => x"78",
          2461 => x"54",
          2462 => x"73",
          2463 => x"60",
          2464 => x"54",
          2465 => x"96",
          2466 => x"0b",
          2467 => x"80",
          2468 => x"f6",
          2469 => x"ec",
          2470 => x"85",
          2471 => x"3d",
          2472 => x"5c",
          2473 => x"53",
          2474 => x"51",
          2475 => x"80",
          2476 => x"88",
          2477 => x"5c",
          2478 => x"09",
          2479 => x"d4",
          2480 => x"70",
          2481 => x"71",
          2482 => x"30",
          2483 => x"73",
          2484 => x"51",
          2485 => x"57",
          2486 => x"38",
          2487 => x"75",
          2488 => x"17",
          2489 => x"75",
          2490 => x"30",
          2491 => x"51",
          2492 => x"80",
          2493 => x"38",
          2494 => x"87",
          2495 => x"26",
          2496 => x"77",
          2497 => x"a4",
          2498 => x"27",
          2499 => x"a0",
          2500 => x"39",
          2501 => x"33",
          2502 => x"57",
          2503 => x"27",
          2504 => x"75",
          2505 => x"30",
          2506 => x"32",
          2507 => x"80",
          2508 => x"25",
          2509 => x"56",
          2510 => x"80",
          2511 => x"84",
          2512 => x"58",
          2513 => x"70",
          2514 => x"55",
          2515 => x"09",
          2516 => x"38",
          2517 => x"80",
          2518 => x"30",
          2519 => x"77",
          2520 => x"54",
          2521 => x"81",
          2522 => x"ae",
          2523 => x"06",
          2524 => x"54",
          2525 => x"74",
          2526 => x"80",
          2527 => x"7b",
          2528 => x"30",
          2529 => x"70",
          2530 => x"25",
          2531 => x"07",
          2532 => x"51",
          2533 => x"a7",
          2534 => x"8b",
          2535 => x"39",
          2536 => x"54",
          2537 => x"8c",
          2538 => x"ff",
          2539 => x"b0",
          2540 => x"54",
          2541 => x"e1",
          2542 => x"e0",
          2543 => x"b2",
          2544 => x"70",
          2545 => x"71",
          2546 => x"54",
          2547 => x"81",
          2548 => x"80",
          2549 => x"38",
          2550 => x"76",
          2551 => x"df",
          2552 => x"54",
          2553 => x"81",
          2554 => x"55",
          2555 => x"34",
          2556 => x"52",
          2557 => x"51",
          2558 => x"81",
          2559 => x"bf",
          2560 => x"16",
          2561 => x"26",
          2562 => x"16",
          2563 => x"06",
          2564 => x"17",
          2565 => x"34",
          2566 => x"fd",
          2567 => x"19",
          2568 => x"80",
          2569 => x"79",
          2570 => x"81",
          2571 => x"81",
          2572 => x"85",
          2573 => x"54",
          2574 => x"8f",
          2575 => x"86",
          2576 => x"39",
          2577 => x"f3",
          2578 => x"73",
          2579 => x"80",
          2580 => x"52",
          2581 => x"ce",
          2582 => x"e0",
          2583 => x"ec",
          2584 => x"d7",
          2585 => x"08",
          2586 => x"e6",
          2587 => x"ec",
          2588 => x"81",
          2589 => x"80",
          2590 => x"1b",
          2591 => x"55",
          2592 => x"2e",
          2593 => x"8b",
          2594 => x"06",
          2595 => x"1c",
          2596 => x"33",
          2597 => x"70",
          2598 => x"55",
          2599 => x"38",
          2600 => x"52",
          2601 => x"9f",
          2602 => x"e0",
          2603 => x"8b",
          2604 => x"7a",
          2605 => x"3f",
          2606 => x"75",
          2607 => x"57",
          2608 => x"2e",
          2609 => x"84",
          2610 => x"06",
          2611 => x"75",
          2612 => x"81",
          2613 => x"2a",
          2614 => x"73",
          2615 => x"38",
          2616 => x"54",
          2617 => x"fb",
          2618 => x"80",
          2619 => x"34",
          2620 => x"c1",
          2621 => x"06",
          2622 => x"38",
          2623 => x"39",
          2624 => x"70",
          2625 => x"54",
          2626 => x"86",
          2627 => x"84",
          2628 => x"06",
          2629 => x"73",
          2630 => x"38",
          2631 => x"83",
          2632 => x"b4",
          2633 => x"51",
          2634 => x"81",
          2635 => x"88",
          2636 => x"ea",
          2637 => x"ec",
          2638 => x"3d",
          2639 => x"3d",
          2640 => x"ff",
          2641 => x"71",
          2642 => x"5c",
          2643 => x"80",
          2644 => x"38",
          2645 => x"05",
          2646 => x"a0",
          2647 => x"71",
          2648 => x"38",
          2649 => x"71",
          2650 => x"81",
          2651 => x"38",
          2652 => x"11",
          2653 => x"06",
          2654 => x"70",
          2655 => x"38",
          2656 => x"81",
          2657 => x"05",
          2658 => x"76",
          2659 => x"38",
          2660 => x"dc",
          2661 => x"77",
          2662 => x"57",
          2663 => x"05",
          2664 => x"70",
          2665 => x"33",
          2666 => x"53",
          2667 => x"99",
          2668 => x"e0",
          2669 => x"ff",
          2670 => x"ff",
          2671 => x"70",
          2672 => x"38",
          2673 => x"81",
          2674 => x"51",
          2675 => x"9f",
          2676 => x"72",
          2677 => x"81",
          2678 => x"70",
          2679 => x"72",
          2680 => x"32",
          2681 => x"72",
          2682 => x"73",
          2683 => x"53",
          2684 => x"70",
          2685 => x"38",
          2686 => x"19",
          2687 => x"75",
          2688 => x"38",
          2689 => x"83",
          2690 => x"74",
          2691 => x"59",
          2692 => x"39",
          2693 => x"33",
          2694 => x"ec",
          2695 => x"3d",
          2696 => x"3d",
          2697 => x"80",
          2698 => x"34",
          2699 => x"17",
          2700 => x"75",
          2701 => x"3f",
          2702 => x"ec",
          2703 => x"80",
          2704 => x"16",
          2705 => x"3f",
          2706 => x"08",
          2707 => x"06",
          2708 => x"73",
          2709 => x"2e",
          2710 => x"80",
          2711 => x"0b",
          2712 => x"56",
          2713 => x"e9",
          2714 => x"06",
          2715 => x"57",
          2716 => x"32",
          2717 => x"80",
          2718 => x"51",
          2719 => x"8a",
          2720 => x"e8",
          2721 => x"06",
          2722 => x"53",
          2723 => x"52",
          2724 => x"51",
          2725 => x"81",
          2726 => x"55",
          2727 => x"08",
          2728 => x"38",
          2729 => x"db",
          2730 => x"86",
          2731 => x"97",
          2732 => x"e0",
          2733 => x"ec",
          2734 => x"2e",
          2735 => x"55",
          2736 => x"e0",
          2737 => x"0d",
          2738 => x"0d",
          2739 => x"05",
          2740 => x"33",
          2741 => x"75",
          2742 => x"fc",
          2743 => x"ec",
          2744 => x"8b",
          2745 => x"81",
          2746 => x"24",
          2747 => x"81",
          2748 => x"84",
          2749 => x"fc",
          2750 => x"55",
          2751 => x"73",
          2752 => x"e6",
          2753 => x"0c",
          2754 => x"06",
          2755 => x"57",
          2756 => x"ae",
          2757 => x"33",
          2758 => x"3f",
          2759 => x"08",
          2760 => x"70",
          2761 => x"55",
          2762 => x"76",
          2763 => x"b8",
          2764 => x"2a",
          2765 => x"51",
          2766 => x"72",
          2767 => x"86",
          2768 => x"74",
          2769 => x"15",
          2770 => x"81",
          2771 => x"d7",
          2772 => x"ec",
          2773 => x"ff",
          2774 => x"06",
          2775 => x"56",
          2776 => x"38",
          2777 => x"8f",
          2778 => x"2a",
          2779 => x"51",
          2780 => x"72",
          2781 => x"80",
          2782 => x"52",
          2783 => x"3f",
          2784 => x"08",
          2785 => x"57",
          2786 => x"09",
          2787 => x"e2",
          2788 => x"74",
          2789 => x"56",
          2790 => x"33",
          2791 => x"72",
          2792 => x"38",
          2793 => x"51",
          2794 => x"81",
          2795 => x"57",
          2796 => x"84",
          2797 => x"ff",
          2798 => x"56",
          2799 => x"25",
          2800 => x"0b",
          2801 => x"56",
          2802 => x"05",
          2803 => x"83",
          2804 => x"2e",
          2805 => x"52",
          2806 => x"c6",
          2807 => x"e0",
          2808 => x"06",
          2809 => x"27",
          2810 => x"16",
          2811 => x"27",
          2812 => x"56",
          2813 => x"84",
          2814 => x"56",
          2815 => x"84",
          2816 => x"14",
          2817 => x"3f",
          2818 => x"08",
          2819 => x"06",
          2820 => x"80",
          2821 => x"06",
          2822 => x"80",
          2823 => x"db",
          2824 => x"ec",
          2825 => x"ff",
          2826 => x"77",
          2827 => x"d8",
          2828 => x"de",
          2829 => x"e0",
          2830 => x"9c",
          2831 => x"c4",
          2832 => x"15",
          2833 => x"14",
          2834 => x"70",
          2835 => x"51",
          2836 => x"56",
          2837 => x"84",
          2838 => x"81",
          2839 => x"71",
          2840 => x"16",
          2841 => x"53",
          2842 => x"23",
          2843 => x"8b",
          2844 => x"73",
          2845 => x"80",
          2846 => x"8d",
          2847 => x"39",
          2848 => x"51",
          2849 => x"81",
          2850 => x"53",
          2851 => x"08",
          2852 => x"72",
          2853 => x"8d",
          2854 => x"ce",
          2855 => x"14",
          2856 => x"3f",
          2857 => x"08",
          2858 => x"06",
          2859 => x"38",
          2860 => x"51",
          2861 => x"81",
          2862 => x"55",
          2863 => x"51",
          2864 => x"81",
          2865 => x"83",
          2866 => x"53",
          2867 => x"80",
          2868 => x"38",
          2869 => x"78",
          2870 => x"2a",
          2871 => x"78",
          2872 => x"86",
          2873 => x"22",
          2874 => x"31",
          2875 => x"be",
          2876 => x"e0",
          2877 => x"ec",
          2878 => x"2e",
          2879 => x"81",
          2880 => x"80",
          2881 => x"f5",
          2882 => x"83",
          2883 => x"ff",
          2884 => x"38",
          2885 => x"9f",
          2886 => x"38",
          2887 => x"39",
          2888 => x"80",
          2889 => x"38",
          2890 => x"98",
          2891 => x"a0",
          2892 => x"1c",
          2893 => x"0c",
          2894 => x"17",
          2895 => x"76",
          2896 => x"81",
          2897 => x"80",
          2898 => x"d9",
          2899 => x"ec",
          2900 => x"ff",
          2901 => x"8d",
          2902 => x"8e",
          2903 => x"8a",
          2904 => x"14",
          2905 => x"3f",
          2906 => x"08",
          2907 => x"74",
          2908 => x"a2",
          2909 => x"79",
          2910 => x"ee",
          2911 => x"a8",
          2912 => x"15",
          2913 => x"2e",
          2914 => x"10",
          2915 => x"2a",
          2916 => x"05",
          2917 => x"ff",
          2918 => x"53",
          2919 => x"9c",
          2920 => x"81",
          2921 => x"0b",
          2922 => x"ff",
          2923 => x"0c",
          2924 => x"84",
          2925 => x"83",
          2926 => x"06",
          2927 => x"80",
          2928 => x"d8",
          2929 => x"ec",
          2930 => x"ff",
          2931 => x"72",
          2932 => x"81",
          2933 => x"38",
          2934 => x"73",
          2935 => x"3f",
          2936 => x"08",
          2937 => x"81",
          2938 => x"84",
          2939 => x"b2",
          2940 => x"87",
          2941 => x"e0",
          2942 => x"ff",
          2943 => x"82",
          2944 => x"09",
          2945 => x"c8",
          2946 => x"51",
          2947 => x"81",
          2948 => x"84",
          2949 => x"d2",
          2950 => x"06",
          2951 => x"98",
          2952 => x"ee",
          2953 => x"e0",
          2954 => x"85",
          2955 => x"09",
          2956 => x"38",
          2957 => x"51",
          2958 => x"81",
          2959 => x"90",
          2960 => x"a0",
          2961 => x"ca",
          2962 => x"e0",
          2963 => x"0c",
          2964 => x"81",
          2965 => x"81",
          2966 => x"81",
          2967 => x"72",
          2968 => x"80",
          2969 => x"0c",
          2970 => x"81",
          2971 => x"90",
          2972 => x"fb",
          2973 => x"54",
          2974 => x"80",
          2975 => x"73",
          2976 => x"80",
          2977 => x"72",
          2978 => x"80",
          2979 => x"86",
          2980 => x"15",
          2981 => x"71",
          2982 => x"81",
          2983 => x"81",
          2984 => x"d0",
          2985 => x"ec",
          2986 => x"06",
          2987 => x"38",
          2988 => x"54",
          2989 => x"80",
          2990 => x"71",
          2991 => x"81",
          2992 => x"87",
          2993 => x"fa",
          2994 => x"ab",
          2995 => x"58",
          2996 => x"05",
          2997 => x"e6",
          2998 => x"80",
          2999 => x"e0",
          3000 => x"38",
          3001 => x"08",
          3002 => x"ec",
          3003 => x"08",
          3004 => x"80",
          3005 => x"80",
          3006 => x"54",
          3007 => x"84",
          3008 => x"34",
          3009 => x"75",
          3010 => x"2e",
          3011 => x"53",
          3012 => x"53",
          3013 => x"f7",
          3014 => x"ec",
          3015 => x"73",
          3016 => x"0c",
          3017 => x"04",
          3018 => x"67",
          3019 => x"80",
          3020 => x"59",
          3021 => x"78",
          3022 => x"c8",
          3023 => x"06",
          3024 => x"3d",
          3025 => x"99",
          3026 => x"52",
          3027 => x"3f",
          3028 => x"08",
          3029 => x"e0",
          3030 => x"38",
          3031 => x"52",
          3032 => x"52",
          3033 => x"3f",
          3034 => x"08",
          3035 => x"e0",
          3036 => x"02",
          3037 => x"33",
          3038 => x"55",
          3039 => x"25",
          3040 => x"55",
          3041 => x"54",
          3042 => x"81",
          3043 => x"80",
          3044 => x"74",
          3045 => x"81",
          3046 => x"75",
          3047 => x"3f",
          3048 => x"08",
          3049 => x"02",
          3050 => x"91",
          3051 => x"81",
          3052 => x"82",
          3053 => x"06",
          3054 => x"80",
          3055 => x"88",
          3056 => x"39",
          3057 => x"58",
          3058 => x"38",
          3059 => x"70",
          3060 => x"54",
          3061 => x"81",
          3062 => x"52",
          3063 => x"a5",
          3064 => x"e0",
          3065 => x"88",
          3066 => x"62",
          3067 => x"d4",
          3068 => x"54",
          3069 => x"15",
          3070 => x"62",
          3071 => x"e8",
          3072 => x"52",
          3073 => x"51",
          3074 => x"7a",
          3075 => x"83",
          3076 => x"80",
          3077 => x"38",
          3078 => x"08",
          3079 => x"53",
          3080 => x"3d",
          3081 => x"dd",
          3082 => x"ec",
          3083 => x"81",
          3084 => x"82",
          3085 => x"39",
          3086 => x"38",
          3087 => x"33",
          3088 => x"70",
          3089 => x"55",
          3090 => x"2e",
          3091 => x"55",
          3092 => x"77",
          3093 => x"81",
          3094 => x"73",
          3095 => x"38",
          3096 => x"54",
          3097 => x"a0",
          3098 => x"82",
          3099 => x"52",
          3100 => x"a3",
          3101 => x"e0",
          3102 => x"18",
          3103 => x"55",
          3104 => x"e0",
          3105 => x"38",
          3106 => x"70",
          3107 => x"54",
          3108 => x"86",
          3109 => x"c0",
          3110 => x"b0",
          3111 => x"1b",
          3112 => x"1b",
          3113 => x"70",
          3114 => x"d9",
          3115 => x"e0",
          3116 => x"e0",
          3117 => x"0c",
          3118 => x"52",
          3119 => x"3f",
          3120 => x"08",
          3121 => x"08",
          3122 => x"77",
          3123 => x"86",
          3124 => x"1a",
          3125 => x"1a",
          3126 => x"91",
          3127 => x"0b",
          3128 => x"80",
          3129 => x"0c",
          3130 => x"70",
          3131 => x"54",
          3132 => x"81",
          3133 => x"ec",
          3134 => x"2e",
          3135 => x"81",
          3136 => x"94",
          3137 => x"17",
          3138 => x"2b",
          3139 => x"57",
          3140 => x"52",
          3141 => x"9f",
          3142 => x"e0",
          3143 => x"ec",
          3144 => x"26",
          3145 => x"55",
          3146 => x"08",
          3147 => x"81",
          3148 => x"79",
          3149 => x"31",
          3150 => x"70",
          3151 => x"25",
          3152 => x"76",
          3153 => x"81",
          3154 => x"55",
          3155 => x"38",
          3156 => x"0c",
          3157 => x"75",
          3158 => x"54",
          3159 => x"a2",
          3160 => x"7a",
          3161 => x"3f",
          3162 => x"08",
          3163 => x"55",
          3164 => x"89",
          3165 => x"e0",
          3166 => x"1a",
          3167 => x"80",
          3168 => x"54",
          3169 => x"e0",
          3170 => x"0d",
          3171 => x"0d",
          3172 => x"64",
          3173 => x"59",
          3174 => x"90",
          3175 => x"52",
          3176 => x"cf",
          3177 => x"e0",
          3178 => x"ec",
          3179 => x"38",
          3180 => x"55",
          3181 => x"86",
          3182 => x"82",
          3183 => x"19",
          3184 => x"55",
          3185 => x"80",
          3186 => x"38",
          3187 => x"0b",
          3188 => x"82",
          3189 => x"39",
          3190 => x"1a",
          3191 => x"82",
          3192 => x"19",
          3193 => x"08",
          3194 => x"7c",
          3195 => x"74",
          3196 => x"2e",
          3197 => x"94",
          3198 => x"83",
          3199 => x"56",
          3200 => x"38",
          3201 => x"22",
          3202 => x"89",
          3203 => x"55",
          3204 => x"75",
          3205 => x"19",
          3206 => x"39",
          3207 => x"52",
          3208 => x"93",
          3209 => x"e0",
          3210 => x"75",
          3211 => x"38",
          3212 => x"ff",
          3213 => x"98",
          3214 => x"19",
          3215 => x"51",
          3216 => x"81",
          3217 => x"80",
          3218 => x"38",
          3219 => x"08",
          3220 => x"2a",
          3221 => x"80",
          3222 => x"38",
          3223 => x"8a",
          3224 => x"5c",
          3225 => x"27",
          3226 => x"7a",
          3227 => x"54",
          3228 => x"52",
          3229 => x"51",
          3230 => x"81",
          3231 => x"fe",
          3232 => x"83",
          3233 => x"56",
          3234 => x"9f",
          3235 => x"08",
          3236 => x"74",
          3237 => x"38",
          3238 => x"b4",
          3239 => x"16",
          3240 => x"89",
          3241 => x"51",
          3242 => x"77",
          3243 => x"b9",
          3244 => x"1a",
          3245 => x"08",
          3246 => x"84",
          3247 => x"57",
          3248 => x"27",
          3249 => x"56",
          3250 => x"52",
          3251 => x"c7",
          3252 => x"e0",
          3253 => x"38",
          3254 => x"19",
          3255 => x"06",
          3256 => x"52",
          3257 => x"a2",
          3258 => x"31",
          3259 => x"7f",
          3260 => x"94",
          3261 => x"94",
          3262 => x"5c",
          3263 => x"80",
          3264 => x"ec",
          3265 => x"3d",
          3266 => x"3d",
          3267 => x"65",
          3268 => x"5d",
          3269 => x"0c",
          3270 => x"05",
          3271 => x"f6",
          3272 => x"ec",
          3273 => x"81",
          3274 => x"8a",
          3275 => x"33",
          3276 => x"2e",
          3277 => x"56",
          3278 => x"90",
          3279 => x"81",
          3280 => x"06",
          3281 => x"87",
          3282 => x"2e",
          3283 => x"95",
          3284 => x"91",
          3285 => x"56",
          3286 => x"81",
          3287 => x"34",
          3288 => x"8e",
          3289 => x"08",
          3290 => x"56",
          3291 => x"84",
          3292 => x"5c",
          3293 => x"82",
          3294 => x"18",
          3295 => x"ff",
          3296 => x"74",
          3297 => x"7e",
          3298 => x"ff",
          3299 => x"2a",
          3300 => x"7a",
          3301 => x"8c",
          3302 => x"08",
          3303 => x"38",
          3304 => x"39",
          3305 => x"52",
          3306 => x"e7",
          3307 => x"e0",
          3308 => x"ec",
          3309 => x"2e",
          3310 => x"74",
          3311 => x"91",
          3312 => x"2e",
          3313 => x"74",
          3314 => x"88",
          3315 => x"38",
          3316 => x"0c",
          3317 => x"15",
          3318 => x"08",
          3319 => x"06",
          3320 => x"51",
          3321 => x"81",
          3322 => x"fe",
          3323 => x"18",
          3324 => x"51",
          3325 => x"81",
          3326 => x"80",
          3327 => x"38",
          3328 => x"08",
          3329 => x"2a",
          3330 => x"80",
          3331 => x"38",
          3332 => x"8a",
          3333 => x"5b",
          3334 => x"27",
          3335 => x"7b",
          3336 => x"54",
          3337 => x"52",
          3338 => x"51",
          3339 => x"81",
          3340 => x"fe",
          3341 => x"b0",
          3342 => x"31",
          3343 => x"79",
          3344 => x"84",
          3345 => x"16",
          3346 => x"89",
          3347 => x"52",
          3348 => x"cc",
          3349 => x"55",
          3350 => x"16",
          3351 => x"2b",
          3352 => x"39",
          3353 => x"94",
          3354 => x"93",
          3355 => x"cd",
          3356 => x"ec",
          3357 => x"e3",
          3358 => x"b0",
          3359 => x"76",
          3360 => x"94",
          3361 => x"ff",
          3362 => x"71",
          3363 => x"7b",
          3364 => x"38",
          3365 => x"18",
          3366 => x"51",
          3367 => x"81",
          3368 => x"fd",
          3369 => x"53",
          3370 => x"18",
          3371 => x"06",
          3372 => x"51",
          3373 => x"7e",
          3374 => x"83",
          3375 => x"76",
          3376 => x"17",
          3377 => x"1e",
          3378 => x"18",
          3379 => x"0c",
          3380 => x"58",
          3381 => x"74",
          3382 => x"38",
          3383 => x"8c",
          3384 => x"90",
          3385 => x"33",
          3386 => x"55",
          3387 => x"34",
          3388 => x"81",
          3389 => x"90",
          3390 => x"f8",
          3391 => x"8b",
          3392 => x"53",
          3393 => x"f2",
          3394 => x"ec",
          3395 => x"81",
          3396 => x"80",
          3397 => x"16",
          3398 => x"2a",
          3399 => x"51",
          3400 => x"80",
          3401 => x"38",
          3402 => x"52",
          3403 => x"e7",
          3404 => x"e0",
          3405 => x"ec",
          3406 => x"d4",
          3407 => x"08",
          3408 => x"a0",
          3409 => x"73",
          3410 => x"88",
          3411 => x"74",
          3412 => x"51",
          3413 => x"8c",
          3414 => x"9c",
          3415 => x"fb",
          3416 => x"b2",
          3417 => x"15",
          3418 => x"3f",
          3419 => x"15",
          3420 => x"3f",
          3421 => x"0b",
          3422 => x"78",
          3423 => x"3f",
          3424 => x"08",
          3425 => x"81",
          3426 => x"57",
          3427 => x"34",
          3428 => x"e0",
          3429 => x"0d",
          3430 => x"0d",
          3431 => x"54",
          3432 => x"81",
          3433 => x"53",
          3434 => x"08",
          3435 => x"3d",
          3436 => x"73",
          3437 => x"3f",
          3438 => x"08",
          3439 => x"e0",
          3440 => x"81",
          3441 => x"74",
          3442 => x"ec",
          3443 => x"3d",
          3444 => x"3d",
          3445 => x"51",
          3446 => x"8b",
          3447 => x"81",
          3448 => x"24",
          3449 => x"ec",
          3450 => x"ed",
          3451 => x"52",
          3452 => x"e0",
          3453 => x"0d",
          3454 => x"0d",
          3455 => x"3d",
          3456 => x"94",
          3457 => x"c1",
          3458 => x"e0",
          3459 => x"ec",
          3460 => x"e0",
          3461 => x"63",
          3462 => x"d4",
          3463 => x"8d",
          3464 => x"e0",
          3465 => x"ec",
          3466 => x"38",
          3467 => x"05",
          3468 => x"2b",
          3469 => x"80",
          3470 => x"76",
          3471 => x"0c",
          3472 => x"02",
          3473 => x"70",
          3474 => x"81",
          3475 => x"56",
          3476 => x"9e",
          3477 => x"53",
          3478 => x"db",
          3479 => x"ec",
          3480 => x"15",
          3481 => x"81",
          3482 => x"84",
          3483 => x"06",
          3484 => x"55",
          3485 => x"e0",
          3486 => x"0d",
          3487 => x"0d",
          3488 => x"5b",
          3489 => x"80",
          3490 => x"ff",
          3491 => x"9f",
          3492 => x"b5",
          3493 => x"e0",
          3494 => x"ec",
          3495 => x"fc",
          3496 => x"7a",
          3497 => x"08",
          3498 => x"64",
          3499 => x"2e",
          3500 => x"a0",
          3501 => x"70",
          3502 => x"ea",
          3503 => x"e0",
          3504 => x"ec",
          3505 => x"d4",
          3506 => x"7b",
          3507 => x"3f",
          3508 => x"08",
          3509 => x"e0",
          3510 => x"38",
          3511 => x"51",
          3512 => x"81",
          3513 => x"45",
          3514 => x"51",
          3515 => x"81",
          3516 => x"57",
          3517 => x"08",
          3518 => x"80",
          3519 => x"da",
          3520 => x"ec",
          3521 => x"81",
          3522 => x"a4",
          3523 => x"7b",
          3524 => x"3f",
          3525 => x"e0",
          3526 => x"38",
          3527 => x"51",
          3528 => x"81",
          3529 => x"57",
          3530 => x"08",
          3531 => x"38",
          3532 => x"09",
          3533 => x"38",
          3534 => x"e0",
          3535 => x"dc",
          3536 => x"ff",
          3537 => x"74",
          3538 => x"3f",
          3539 => x"78",
          3540 => x"33",
          3541 => x"56",
          3542 => x"91",
          3543 => x"05",
          3544 => x"81",
          3545 => x"56",
          3546 => x"f5",
          3547 => x"54",
          3548 => x"81",
          3549 => x"80",
          3550 => x"78",
          3551 => x"55",
          3552 => x"11",
          3553 => x"18",
          3554 => x"58",
          3555 => x"34",
          3556 => x"ff",
          3557 => x"55",
          3558 => x"34",
          3559 => x"77",
          3560 => x"81",
          3561 => x"ff",
          3562 => x"55",
          3563 => x"34",
          3564 => x"ed",
          3565 => x"84",
          3566 => x"a0",
          3567 => x"70",
          3568 => x"56",
          3569 => x"76",
          3570 => x"81",
          3571 => x"70",
          3572 => x"56",
          3573 => x"82",
          3574 => x"78",
          3575 => x"80",
          3576 => x"27",
          3577 => x"19",
          3578 => x"7a",
          3579 => x"5c",
          3580 => x"55",
          3581 => x"7a",
          3582 => x"5c",
          3583 => x"2e",
          3584 => x"85",
          3585 => x"94",
          3586 => x"81",
          3587 => x"73",
          3588 => x"81",
          3589 => x"7a",
          3590 => x"38",
          3591 => x"76",
          3592 => x"0c",
          3593 => x"04",
          3594 => x"7b",
          3595 => x"fc",
          3596 => x"53",
          3597 => x"bb",
          3598 => x"e0",
          3599 => x"ec",
          3600 => x"fa",
          3601 => x"33",
          3602 => x"f2",
          3603 => x"08",
          3604 => x"27",
          3605 => x"15",
          3606 => x"2a",
          3607 => x"51",
          3608 => x"83",
          3609 => x"94",
          3610 => x"80",
          3611 => x"0c",
          3612 => x"2e",
          3613 => x"79",
          3614 => x"70",
          3615 => x"51",
          3616 => x"2e",
          3617 => x"52",
          3618 => x"ff",
          3619 => x"81",
          3620 => x"ff",
          3621 => x"70",
          3622 => x"ff",
          3623 => x"81",
          3624 => x"73",
          3625 => x"76",
          3626 => x"06",
          3627 => x"0c",
          3628 => x"98",
          3629 => x"58",
          3630 => x"39",
          3631 => x"54",
          3632 => x"73",
          3633 => x"cd",
          3634 => x"ec",
          3635 => x"81",
          3636 => x"81",
          3637 => x"38",
          3638 => x"08",
          3639 => x"9b",
          3640 => x"e0",
          3641 => x"0c",
          3642 => x"0c",
          3643 => x"81",
          3644 => x"76",
          3645 => x"38",
          3646 => x"94",
          3647 => x"94",
          3648 => x"16",
          3649 => x"2a",
          3650 => x"51",
          3651 => x"72",
          3652 => x"38",
          3653 => x"51",
          3654 => x"81",
          3655 => x"54",
          3656 => x"08",
          3657 => x"ec",
          3658 => x"a7",
          3659 => x"74",
          3660 => x"3f",
          3661 => x"08",
          3662 => x"2e",
          3663 => x"74",
          3664 => x"79",
          3665 => x"14",
          3666 => x"38",
          3667 => x"0c",
          3668 => x"94",
          3669 => x"94",
          3670 => x"83",
          3671 => x"72",
          3672 => x"38",
          3673 => x"51",
          3674 => x"81",
          3675 => x"94",
          3676 => x"91",
          3677 => x"53",
          3678 => x"81",
          3679 => x"34",
          3680 => x"39",
          3681 => x"81",
          3682 => x"05",
          3683 => x"08",
          3684 => x"08",
          3685 => x"38",
          3686 => x"0c",
          3687 => x"80",
          3688 => x"72",
          3689 => x"73",
          3690 => x"53",
          3691 => x"8c",
          3692 => x"16",
          3693 => x"38",
          3694 => x"0c",
          3695 => x"81",
          3696 => x"8b",
          3697 => x"f9",
          3698 => x"56",
          3699 => x"80",
          3700 => x"38",
          3701 => x"3d",
          3702 => x"8a",
          3703 => x"51",
          3704 => x"81",
          3705 => x"55",
          3706 => x"08",
          3707 => x"77",
          3708 => x"52",
          3709 => x"b5",
          3710 => x"e0",
          3711 => x"ec",
          3712 => x"c3",
          3713 => x"33",
          3714 => x"55",
          3715 => x"24",
          3716 => x"16",
          3717 => x"2a",
          3718 => x"51",
          3719 => x"80",
          3720 => x"9c",
          3721 => x"77",
          3722 => x"3f",
          3723 => x"08",
          3724 => x"77",
          3725 => x"22",
          3726 => x"74",
          3727 => x"ce",
          3728 => x"ec",
          3729 => x"74",
          3730 => x"81",
          3731 => x"85",
          3732 => x"74",
          3733 => x"38",
          3734 => x"74",
          3735 => x"ec",
          3736 => x"3d",
          3737 => x"3d",
          3738 => x"3d",
          3739 => x"70",
          3740 => x"ff",
          3741 => x"e0",
          3742 => x"81",
          3743 => x"73",
          3744 => x"0d",
          3745 => x"0d",
          3746 => x"3d",
          3747 => x"71",
          3748 => x"e7",
          3749 => x"ec",
          3750 => x"81",
          3751 => x"80",
          3752 => x"93",
          3753 => x"e0",
          3754 => x"51",
          3755 => x"81",
          3756 => x"53",
          3757 => x"81",
          3758 => x"52",
          3759 => x"ac",
          3760 => x"e0",
          3761 => x"ec",
          3762 => x"2e",
          3763 => x"85",
          3764 => x"87",
          3765 => x"e0",
          3766 => x"74",
          3767 => x"d5",
          3768 => x"52",
          3769 => x"89",
          3770 => x"e0",
          3771 => x"70",
          3772 => x"07",
          3773 => x"81",
          3774 => x"06",
          3775 => x"54",
          3776 => x"e0",
          3777 => x"0d",
          3778 => x"0d",
          3779 => x"53",
          3780 => x"53",
          3781 => x"56",
          3782 => x"81",
          3783 => x"55",
          3784 => x"08",
          3785 => x"52",
          3786 => x"81",
          3787 => x"e0",
          3788 => x"ec",
          3789 => x"38",
          3790 => x"05",
          3791 => x"2b",
          3792 => x"80",
          3793 => x"86",
          3794 => x"76",
          3795 => x"38",
          3796 => x"51",
          3797 => x"74",
          3798 => x"0c",
          3799 => x"04",
          3800 => x"63",
          3801 => x"80",
          3802 => x"ec",
          3803 => x"3d",
          3804 => x"3f",
          3805 => x"08",
          3806 => x"e0",
          3807 => x"38",
          3808 => x"73",
          3809 => x"08",
          3810 => x"13",
          3811 => x"58",
          3812 => x"26",
          3813 => x"7c",
          3814 => x"39",
          3815 => x"cc",
          3816 => x"81",
          3817 => x"ec",
          3818 => x"33",
          3819 => x"81",
          3820 => x"06",
          3821 => x"75",
          3822 => x"52",
          3823 => x"05",
          3824 => x"3f",
          3825 => x"08",
          3826 => x"38",
          3827 => x"08",
          3828 => x"38",
          3829 => x"08",
          3830 => x"ec",
          3831 => x"80",
          3832 => x"81",
          3833 => x"59",
          3834 => x"14",
          3835 => x"ca",
          3836 => x"39",
          3837 => x"81",
          3838 => x"57",
          3839 => x"38",
          3840 => x"18",
          3841 => x"ff",
          3842 => x"81",
          3843 => x"5b",
          3844 => x"08",
          3845 => x"7c",
          3846 => x"12",
          3847 => x"52",
          3848 => x"82",
          3849 => x"06",
          3850 => x"14",
          3851 => x"cb",
          3852 => x"e0",
          3853 => x"ff",
          3854 => x"70",
          3855 => x"82",
          3856 => x"51",
          3857 => x"b4",
          3858 => x"bb",
          3859 => x"ec",
          3860 => x"0a",
          3861 => x"70",
          3862 => x"84",
          3863 => x"51",
          3864 => x"ff",
          3865 => x"56",
          3866 => x"38",
          3867 => x"7c",
          3868 => x"0c",
          3869 => x"81",
          3870 => x"74",
          3871 => x"7a",
          3872 => x"0c",
          3873 => x"04",
          3874 => x"79",
          3875 => x"05",
          3876 => x"57",
          3877 => x"81",
          3878 => x"56",
          3879 => x"08",
          3880 => x"91",
          3881 => x"75",
          3882 => x"90",
          3883 => x"81",
          3884 => x"06",
          3885 => x"87",
          3886 => x"2e",
          3887 => x"94",
          3888 => x"73",
          3889 => x"27",
          3890 => x"73",
          3891 => x"ec",
          3892 => x"88",
          3893 => x"76",
          3894 => x"3f",
          3895 => x"08",
          3896 => x"0c",
          3897 => x"39",
          3898 => x"52",
          3899 => x"bf",
          3900 => x"ec",
          3901 => x"2e",
          3902 => x"83",
          3903 => x"81",
          3904 => x"81",
          3905 => x"06",
          3906 => x"56",
          3907 => x"a0",
          3908 => x"81",
          3909 => x"98",
          3910 => x"94",
          3911 => x"08",
          3912 => x"e0",
          3913 => x"51",
          3914 => x"81",
          3915 => x"56",
          3916 => x"8c",
          3917 => x"17",
          3918 => x"07",
          3919 => x"18",
          3920 => x"2e",
          3921 => x"91",
          3922 => x"55",
          3923 => x"e0",
          3924 => x"0d",
          3925 => x"0d",
          3926 => x"3d",
          3927 => x"52",
          3928 => x"da",
          3929 => x"ec",
          3930 => x"81",
          3931 => x"81",
          3932 => x"45",
          3933 => x"52",
          3934 => x"52",
          3935 => x"3f",
          3936 => x"08",
          3937 => x"e0",
          3938 => x"38",
          3939 => x"05",
          3940 => x"2a",
          3941 => x"51",
          3942 => x"55",
          3943 => x"38",
          3944 => x"54",
          3945 => x"81",
          3946 => x"80",
          3947 => x"70",
          3948 => x"54",
          3949 => x"81",
          3950 => x"52",
          3951 => x"c5",
          3952 => x"e0",
          3953 => x"2a",
          3954 => x"51",
          3955 => x"80",
          3956 => x"38",
          3957 => x"ec",
          3958 => x"15",
          3959 => x"86",
          3960 => x"81",
          3961 => x"5c",
          3962 => x"3d",
          3963 => x"c7",
          3964 => x"ec",
          3965 => x"81",
          3966 => x"80",
          3967 => x"ec",
          3968 => x"73",
          3969 => x"3f",
          3970 => x"08",
          3971 => x"e0",
          3972 => x"87",
          3973 => x"39",
          3974 => x"08",
          3975 => x"38",
          3976 => x"08",
          3977 => x"77",
          3978 => x"3f",
          3979 => x"08",
          3980 => x"08",
          3981 => x"ec",
          3982 => x"80",
          3983 => x"55",
          3984 => x"94",
          3985 => x"2e",
          3986 => x"53",
          3987 => x"51",
          3988 => x"81",
          3989 => x"55",
          3990 => x"78",
          3991 => x"fe",
          3992 => x"e0",
          3993 => x"81",
          3994 => x"a0",
          3995 => x"e9",
          3996 => x"53",
          3997 => x"05",
          3998 => x"51",
          3999 => x"81",
          4000 => x"54",
          4001 => x"08",
          4002 => x"78",
          4003 => x"8e",
          4004 => x"58",
          4005 => x"81",
          4006 => x"54",
          4007 => x"08",
          4008 => x"54",
          4009 => x"81",
          4010 => x"84",
          4011 => x"06",
          4012 => x"02",
          4013 => x"33",
          4014 => x"81",
          4015 => x"86",
          4016 => x"f6",
          4017 => x"74",
          4018 => x"70",
          4019 => x"c3",
          4020 => x"e0",
          4021 => x"56",
          4022 => x"08",
          4023 => x"54",
          4024 => x"08",
          4025 => x"81",
          4026 => x"82",
          4027 => x"e0",
          4028 => x"09",
          4029 => x"38",
          4030 => x"b4",
          4031 => x"b0",
          4032 => x"e0",
          4033 => x"51",
          4034 => x"81",
          4035 => x"54",
          4036 => x"08",
          4037 => x"8b",
          4038 => x"b4",
          4039 => x"b7",
          4040 => x"54",
          4041 => x"15",
          4042 => x"90",
          4043 => x"34",
          4044 => x"0a",
          4045 => x"19",
          4046 => x"9f",
          4047 => x"78",
          4048 => x"51",
          4049 => x"a0",
          4050 => x"11",
          4051 => x"05",
          4052 => x"b6",
          4053 => x"ae",
          4054 => x"15",
          4055 => x"78",
          4056 => x"53",
          4057 => x"3f",
          4058 => x"0b",
          4059 => x"77",
          4060 => x"3f",
          4061 => x"08",
          4062 => x"e0",
          4063 => x"82",
          4064 => x"52",
          4065 => x"51",
          4066 => x"3f",
          4067 => x"52",
          4068 => x"aa",
          4069 => x"90",
          4070 => x"34",
          4071 => x"0b",
          4072 => x"78",
          4073 => x"b6",
          4074 => x"e0",
          4075 => x"39",
          4076 => x"52",
          4077 => x"be",
          4078 => x"81",
          4079 => x"99",
          4080 => x"da",
          4081 => x"3d",
          4082 => x"d2",
          4083 => x"53",
          4084 => x"84",
          4085 => x"3d",
          4086 => x"3f",
          4087 => x"08",
          4088 => x"e0",
          4089 => x"38",
          4090 => x"3d",
          4091 => x"3d",
          4092 => x"cc",
          4093 => x"ec",
          4094 => x"81",
          4095 => x"82",
          4096 => x"81",
          4097 => x"81",
          4098 => x"86",
          4099 => x"aa",
          4100 => x"a4",
          4101 => x"a8",
          4102 => x"05",
          4103 => x"ea",
          4104 => x"77",
          4105 => x"70",
          4106 => x"b4",
          4107 => x"3d",
          4108 => x"51",
          4109 => x"81",
          4110 => x"55",
          4111 => x"08",
          4112 => x"6f",
          4113 => x"06",
          4114 => x"a2",
          4115 => x"92",
          4116 => x"81",
          4117 => x"ec",
          4118 => x"2e",
          4119 => x"81",
          4120 => x"51",
          4121 => x"81",
          4122 => x"55",
          4123 => x"08",
          4124 => x"68",
          4125 => x"a8",
          4126 => x"05",
          4127 => x"51",
          4128 => x"3f",
          4129 => x"33",
          4130 => x"8b",
          4131 => x"84",
          4132 => x"06",
          4133 => x"73",
          4134 => x"a0",
          4135 => x"8b",
          4136 => x"54",
          4137 => x"15",
          4138 => x"33",
          4139 => x"70",
          4140 => x"55",
          4141 => x"2e",
          4142 => x"6e",
          4143 => x"df",
          4144 => x"78",
          4145 => x"3f",
          4146 => x"08",
          4147 => x"ff",
          4148 => x"82",
          4149 => x"e0",
          4150 => x"80",
          4151 => x"ec",
          4152 => x"78",
          4153 => x"af",
          4154 => x"e0",
          4155 => x"d4",
          4156 => x"55",
          4157 => x"08",
          4158 => x"81",
          4159 => x"73",
          4160 => x"81",
          4161 => x"63",
          4162 => x"76",
          4163 => x"3f",
          4164 => x"0b",
          4165 => x"87",
          4166 => x"e0",
          4167 => x"77",
          4168 => x"3f",
          4169 => x"08",
          4170 => x"e0",
          4171 => x"78",
          4172 => x"aa",
          4173 => x"e0",
          4174 => x"81",
          4175 => x"a8",
          4176 => x"ed",
          4177 => x"80",
          4178 => x"02",
          4179 => x"df",
          4180 => x"57",
          4181 => x"3d",
          4182 => x"96",
          4183 => x"e9",
          4184 => x"e0",
          4185 => x"ec",
          4186 => x"cf",
          4187 => x"65",
          4188 => x"d4",
          4189 => x"b5",
          4190 => x"e0",
          4191 => x"ec",
          4192 => x"38",
          4193 => x"05",
          4194 => x"06",
          4195 => x"73",
          4196 => x"a7",
          4197 => x"09",
          4198 => x"71",
          4199 => x"06",
          4200 => x"55",
          4201 => x"15",
          4202 => x"81",
          4203 => x"34",
          4204 => x"b4",
          4205 => x"ec",
          4206 => x"74",
          4207 => x"0c",
          4208 => x"04",
          4209 => x"64",
          4210 => x"93",
          4211 => x"52",
          4212 => x"d1",
          4213 => x"ec",
          4214 => x"81",
          4215 => x"80",
          4216 => x"58",
          4217 => x"3d",
          4218 => x"c8",
          4219 => x"ec",
          4220 => x"81",
          4221 => x"b4",
          4222 => x"c7",
          4223 => x"a0",
          4224 => x"55",
          4225 => x"84",
          4226 => x"17",
          4227 => x"2b",
          4228 => x"96",
          4229 => x"b0",
          4230 => x"54",
          4231 => x"15",
          4232 => x"ff",
          4233 => x"81",
          4234 => x"55",
          4235 => x"e0",
          4236 => x"0d",
          4237 => x"0d",
          4238 => x"5a",
          4239 => x"3d",
          4240 => x"99",
          4241 => x"81",
          4242 => x"e0",
          4243 => x"e0",
          4244 => x"81",
          4245 => x"07",
          4246 => x"55",
          4247 => x"2e",
          4248 => x"81",
          4249 => x"55",
          4250 => x"2e",
          4251 => x"7b",
          4252 => x"80",
          4253 => x"70",
          4254 => x"be",
          4255 => x"ec",
          4256 => x"81",
          4257 => x"80",
          4258 => x"52",
          4259 => x"dc",
          4260 => x"e0",
          4261 => x"ec",
          4262 => x"38",
          4263 => x"08",
          4264 => x"08",
          4265 => x"56",
          4266 => x"19",
          4267 => x"59",
          4268 => x"74",
          4269 => x"56",
          4270 => x"ec",
          4271 => x"75",
          4272 => x"74",
          4273 => x"2e",
          4274 => x"16",
          4275 => x"33",
          4276 => x"73",
          4277 => x"38",
          4278 => x"84",
          4279 => x"06",
          4280 => x"7a",
          4281 => x"76",
          4282 => x"07",
          4283 => x"54",
          4284 => x"80",
          4285 => x"80",
          4286 => x"7b",
          4287 => x"53",
          4288 => x"93",
          4289 => x"e0",
          4290 => x"ec",
          4291 => x"38",
          4292 => x"55",
          4293 => x"56",
          4294 => x"8b",
          4295 => x"56",
          4296 => x"83",
          4297 => x"75",
          4298 => x"51",
          4299 => x"3f",
          4300 => x"08",
          4301 => x"81",
          4302 => x"98",
          4303 => x"e6",
          4304 => x"53",
          4305 => x"b8",
          4306 => x"3d",
          4307 => x"3f",
          4308 => x"08",
          4309 => x"08",
          4310 => x"ec",
          4311 => x"98",
          4312 => x"a0",
          4313 => x"70",
          4314 => x"ae",
          4315 => x"6d",
          4316 => x"81",
          4317 => x"57",
          4318 => x"74",
          4319 => x"38",
          4320 => x"81",
          4321 => x"81",
          4322 => x"52",
          4323 => x"89",
          4324 => x"e0",
          4325 => x"a5",
          4326 => x"33",
          4327 => x"54",
          4328 => x"3f",
          4329 => x"08",
          4330 => x"38",
          4331 => x"76",
          4332 => x"05",
          4333 => x"39",
          4334 => x"08",
          4335 => x"15",
          4336 => x"ff",
          4337 => x"73",
          4338 => x"38",
          4339 => x"83",
          4340 => x"56",
          4341 => x"75",
          4342 => x"81",
          4343 => x"33",
          4344 => x"2e",
          4345 => x"52",
          4346 => x"51",
          4347 => x"3f",
          4348 => x"08",
          4349 => x"ff",
          4350 => x"38",
          4351 => x"88",
          4352 => x"8a",
          4353 => x"38",
          4354 => x"ec",
          4355 => x"75",
          4356 => x"74",
          4357 => x"73",
          4358 => x"05",
          4359 => x"17",
          4360 => x"70",
          4361 => x"34",
          4362 => x"70",
          4363 => x"ff",
          4364 => x"55",
          4365 => x"26",
          4366 => x"8b",
          4367 => x"86",
          4368 => x"e5",
          4369 => x"38",
          4370 => x"99",
          4371 => x"05",
          4372 => x"70",
          4373 => x"73",
          4374 => x"81",
          4375 => x"ff",
          4376 => x"ed",
          4377 => x"80",
          4378 => x"91",
          4379 => x"55",
          4380 => x"3f",
          4381 => x"08",
          4382 => x"e0",
          4383 => x"38",
          4384 => x"51",
          4385 => x"3f",
          4386 => x"08",
          4387 => x"e0",
          4388 => x"76",
          4389 => x"67",
          4390 => x"34",
          4391 => x"81",
          4392 => x"84",
          4393 => x"06",
          4394 => x"80",
          4395 => x"2e",
          4396 => x"81",
          4397 => x"ff",
          4398 => x"81",
          4399 => x"54",
          4400 => x"08",
          4401 => x"53",
          4402 => x"08",
          4403 => x"ff",
          4404 => x"67",
          4405 => x"8b",
          4406 => x"53",
          4407 => x"51",
          4408 => x"3f",
          4409 => x"0b",
          4410 => x"79",
          4411 => x"ee",
          4412 => x"e0",
          4413 => x"55",
          4414 => x"e0",
          4415 => x"0d",
          4416 => x"0d",
          4417 => x"88",
          4418 => x"05",
          4419 => x"fc",
          4420 => x"54",
          4421 => x"d2",
          4422 => x"ec",
          4423 => x"81",
          4424 => x"82",
          4425 => x"1a",
          4426 => x"82",
          4427 => x"80",
          4428 => x"8c",
          4429 => x"78",
          4430 => x"1a",
          4431 => x"2a",
          4432 => x"51",
          4433 => x"90",
          4434 => x"82",
          4435 => x"58",
          4436 => x"81",
          4437 => x"39",
          4438 => x"22",
          4439 => x"70",
          4440 => x"56",
          4441 => x"ff",
          4442 => x"14",
          4443 => x"30",
          4444 => x"9f",
          4445 => x"e0",
          4446 => x"19",
          4447 => x"5a",
          4448 => x"81",
          4449 => x"38",
          4450 => x"77",
          4451 => x"82",
          4452 => x"56",
          4453 => x"74",
          4454 => x"ff",
          4455 => x"81",
          4456 => x"55",
          4457 => x"75",
          4458 => x"82",
          4459 => x"e0",
          4460 => x"ff",
          4461 => x"ec",
          4462 => x"2e",
          4463 => x"81",
          4464 => x"8e",
          4465 => x"56",
          4466 => x"09",
          4467 => x"38",
          4468 => x"59",
          4469 => x"77",
          4470 => x"06",
          4471 => x"87",
          4472 => x"39",
          4473 => x"ba",
          4474 => x"55",
          4475 => x"2e",
          4476 => x"15",
          4477 => x"2e",
          4478 => x"83",
          4479 => x"75",
          4480 => x"7e",
          4481 => x"a8",
          4482 => x"e0",
          4483 => x"ec",
          4484 => x"ce",
          4485 => x"16",
          4486 => x"56",
          4487 => x"38",
          4488 => x"19",
          4489 => x"8c",
          4490 => x"7d",
          4491 => x"38",
          4492 => x"0c",
          4493 => x"0c",
          4494 => x"80",
          4495 => x"73",
          4496 => x"98",
          4497 => x"05",
          4498 => x"57",
          4499 => x"26",
          4500 => x"7b",
          4501 => x"0c",
          4502 => x"81",
          4503 => x"84",
          4504 => x"54",
          4505 => x"e0",
          4506 => x"0d",
          4507 => x"0d",
          4508 => x"88",
          4509 => x"05",
          4510 => x"54",
          4511 => x"c5",
          4512 => x"56",
          4513 => x"ec",
          4514 => x"8b",
          4515 => x"ec",
          4516 => x"29",
          4517 => x"05",
          4518 => x"55",
          4519 => x"84",
          4520 => x"34",
          4521 => x"08",
          4522 => x"5f",
          4523 => x"51",
          4524 => x"3f",
          4525 => x"08",
          4526 => x"70",
          4527 => x"57",
          4528 => x"8b",
          4529 => x"82",
          4530 => x"06",
          4531 => x"56",
          4532 => x"38",
          4533 => x"05",
          4534 => x"7e",
          4535 => x"f0",
          4536 => x"e0",
          4537 => x"67",
          4538 => x"2e",
          4539 => x"82",
          4540 => x"8b",
          4541 => x"75",
          4542 => x"80",
          4543 => x"81",
          4544 => x"2e",
          4545 => x"80",
          4546 => x"38",
          4547 => x"0a",
          4548 => x"ff",
          4549 => x"55",
          4550 => x"86",
          4551 => x"8a",
          4552 => x"89",
          4553 => x"2a",
          4554 => x"77",
          4555 => x"59",
          4556 => x"81",
          4557 => x"70",
          4558 => x"07",
          4559 => x"56",
          4560 => x"38",
          4561 => x"05",
          4562 => x"7e",
          4563 => x"80",
          4564 => x"81",
          4565 => x"8a",
          4566 => x"83",
          4567 => x"06",
          4568 => x"08",
          4569 => x"74",
          4570 => x"41",
          4571 => x"56",
          4572 => x"8a",
          4573 => x"61",
          4574 => x"55",
          4575 => x"27",
          4576 => x"93",
          4577 => x"80",
          4578 => x"38",
          4579 => x"70",
          4580 => x"43",
          4581 => x"95",
          4582 => x"06",
          4583 => x"2e",
          4584 => x"77",
          4585 => x"74",
          4586 => x"83",
          4587 => x"06",
          4588 => x"82",
          4589 => x"2e",
          4590 => x"78",
          4591 => x"2e",
          4592 => x"80",
          4593 => x"ae",
          4594 => x"2a",
          4595 => x"81",
          4596 => x"56",
          4597 => x"2e",
          4598 => x"77",
          4599 => x"81",
          4600 => x"79",
          4601 => x"70",
          4602 => x"5a",
          4603 => x"86",
          4604 => x"27",
          4605 => x"52",
          4606 => x"fa",
          4607 => x"ec",
          4608 => x"29",
          4609 => x"70",
          4610 => x"55",
          4611 => x"0b",
          4612 => x"08",
          4613 => x"05",
          4614 => x"ff",
          4615 => x"27",
          4616 => x"88",
          4617 => x"ae",
          4618 => x"2a",
          4619 => x"81",
          4620 => x"56",
          4621 => x"2e",
          4622 => x"77",
          4623 => x"81",
          4624 => x"79",
          4625 => x"70",
          4626 => x"5a",
          4627 => x"86",
          4628 => x"27",
          4629 => x"52",
          4630 => x"f9",
          4631 => x"ec",
          4632 => x"84",
          4633 => x"ec",
          4634 => x"f5",
          4635 => x"81",
          4636 => x"e0",
          4637 => x"ec",
          4638 => x"71",
          4639 => x"83",
          4640 => x"5e",
          4641 => x"89",
          4642 => x"5c",
          4643 => x"1c",
          4644 => x"05",
          4645 => x"ff",
          4646 => x"70",
          4647 => x"31",
          4648 => x"57",
          4649 => x"83",
          4650 => x"06",
          4651 => x"1c",
          4652 => x"5c",
          4653 => x"1d",
          4654 => x"29",
          4655 => x"31",
          4656 => x"55",
          4657 => x"87",
          4658 => x"7c",
          4659 => x"7a",
          4660 => x"31",
          4661 => x"f8",
          4662 => x"ec",
          4663 => x"7d",
          4664 => x"81",
          4665 => x"81",
          4666 => x"83",
          4667 => x"80",
          4668 => x"87",
          4669 => x"81",
          4670 => x"fd",
          4671 => x"f8",
          4672 => x"2e",
          4673 => x"80",
          4674 => x"ff",
          4675 => x"ec",
          4676 => x"a0",
          4677 => x"38",
          4678 => x"74",
          4679 => x"86",
          4680 => x"fd",
          4681 => x"81",
          4682 => x"80",
          4683 => x"83",
          4684 => x"39",
          4685 => x"08",
          4686 => x"92",
          4687 => x"b8",
          4688 => x"59",
          4689 => x"27",
          4690 => x"86",
          4691 => x"55",
          4692 => x"09",
          4693 => x"38",
          4694 => x"f5",
          4695 => x"38",
          4696 => x"55",
          4697 => x"86",
          4698 => x"80",
          4699 => x"7a",
          4700 => x"b9",
          4701 => x"81",
          4702 => x"7a",
          4703 => x"8a",
          4704 => x"52",
          4705 => x"ff",
          4706 => x"79",
          4707 => x"7b",
          4708 => x"06",
          4709 => x"51",
          4710 => x"3f",
          4711 => x"1c",
          4712 => x"32",
          4713 => x"96",
          4714 => x"06",
          4715 => x"91",
          4716 => x"a1",
          4717 => x"55",
          4718 => x"ff",
          4719 => x"74",
          4720 => x"06",
          4721 => x"51",
          4722 => x"3f",
          4723 => x"52",
          4724 => x"ff",
          4725 => x"f8",
          4726 => x"34",
          4727 => x"1b",
          4728 => x"d9",
          4729 => x"52",
          4730 => x"ff",
          4731 => x"60",
          4732 => x"51",
          4733 => x"3f",
          4734 => x"09",
          4735 => x"cb",
          4736 => x"b2",
          4737 => x"c3",
          4738 => x"a0",
          4739 => x"52",
          4740 => x"ff",
          4741 => x"82",
          4742 => x"51",
          4743 => x"3f",
          4744 => x"1b",
          4745 => x"95",
          4746 => x"b2",
          4747 => x"a0",
          4748 => x"80",
          4749 => x"1c",
          4750 => x"80",
          4751 => x"93",
          4752 => x"f8",
          4753 => x"1b",
          4754 => x"82",
          4755 => x"52",
          4756 => x"ff",
          4757 => x"7c",
          4758 => x"06",
          4759 => x"51",
          4760 => x"3f",
          4761 => x"a4",
          4762 => x"0b",
          4763 => x"93",
          4764 => x"8c",
          4765 => x"51",
          4766 => x"3f",
          4767 => x"52",
          4768 => x"70",
          4769 => x"9f",
          4770 => x"54",
          4771 => x"52",
          4772 => x"9b",
          4773 => x"56",
          4774 => x"08",
          4775 => x"7d",
          4776 => x"81",
          4777 => x"38",
          4778 => x"86",
          4779 => x"52",
          4780 => x"9b",
          4781 => x"80",
          4782 => x"7a",
          4783 => x"ed",
          4784 => x"85",
          4785 => x"7a",
          4786 => x"8f",
          4787 => x"85",
          4788 => x"83",
          4789 => x"ff",
          4790 => x"ff",
          4791 => x"e8",
          4792 => x"9e",
          4793 => x"52",
          4794 => x"51",
          4795 => x"3f",
          4796 => x"52",
          4797 => x"9e",
          4798 => x"54",
          4799 => x"53",
          4800 => x"51",
          4801 => x"3f",
          4802 => x"16",
          4803 => x"7e",
          4804 => x"d8",
          4805 => x"80",
          4806 => x"ff",
          4807 => x"7f",
          4808 => x"7d",
          4809 => x"81",
          4810 => x"f8",
          4811 => x"ff",
          4812 => x"ff",
          4813 => x"51",
          4814 => x"3f",
          4815 => x"88",
          4816 => x"39",
          4817 => x"f8",
          4818 => x"2e",
          4819 => x"55",
          4820 => x"51",
          4821 => x"3f",
          4822 => x"57",
          4823 => x"83",
          4824 => x"76",
          4825 => x"7a",
          4826 => x"ff",
          4827 => x"81",
          4828 => x"82",
          4829 => x"80",
          4830 => x"e0",
          4831 => x"51",
          4832 => x"3f",
          4833 => x"78",
          4834 => x"74",
          4835 => x"18",
          4836 => x"2e",
          4837 => x"79",
          4838 => x"2e",
          4839 => x"55",
          4840 => x"62",
          4841 => x"74",
          4842 => x"75",
          4843 => x"7e",
          4844 => x"b8",
          4845 => x"e0",
          4846 => x"38",
          4847 => x"78",
          4848 => x"74",
          4849 => x"56",
          4850 => x"93",
          4851 => x"66",
          4852 => x"26",
          4853 => x"56",
          4854 => x"83",
          4855 => x"64",
          4856 => x"77",
          4857 => x"84",
          4858 => x"52",
          4859 => x"9d",
          4860 => x"d4",
          4861 => x"51",
          4862 => x"3f",
          4863 => x"55",
          4864 => x"81",
          4865 => x"34",
          4866 => x"16",
          4867 => x"16",
          4868 => x"16",
          4869 => x"05",
          4870 => x"c1",
          4871 => x"fe",
          4872 => x"fe",
          4873 => x"34",
          4874 => x"08",
          4875 => x"07",
          4876 => x"16",
          4877 => x"e0",
          4878 => x"34",
          4879 => x"c6",
          4880 => x"9c",
          4881 => x"52",
          4882 => x"51",
          4883 => x"3f",
          4884 => x"53",
          4885 => x"51",
          4886 => x"3f",
          4887 => x"ec",
          4888 => x"38",
          4889 => x"52",
          4890 => x"99",
          4891 => x"56",
          4892 => x"08",
          4893 => x"39",
          4894 => x"39",
          4895 => x"39",
          4896 => x"08",
          4897 => x"ec",
          4898 => x"3d",
          4899 => x"3d",
          4900 => x"5b",
          4901 => x"60",
          4902 => x"57",
          4903 => x"25",
          4904 => x"3d",
          4905 => x"55",
          4906 => x"15",
          4907 => x"c9",
          4908 => x"81",
          4909 => x"06",
          4910 => x"3d",
          4911 => x"8d",
          4912 => x"74",
          4913 => x"05",
          4914 => x"17",
          4915 => x"2e",
          4916 => x"c9",
          4917 => x"34",
          4918 => x"83",
          4919 => x"74",
          4920 => x"0c",
          4921 => x"04",
          4922 => x"78",
          4923 => x"55",
          4924 => x"80",
          4925 => x"38",
          4926 => x"77",
          4927 => x"33",
          4928 => x"39",
          4929 => x"80",
          4930 => x"56",
          4931 => x"83",
          4932 => x"73",
          4933 => x"2a",
          4934 => x"53",
          4935 => x"73",
          4936 => x"81",
          4937 => x"72",
          4938 => x"05",
          4939 => x"56",
          4940 => x"81",
          4941 => x"77",
          4942 => x"08",
          4943 => x"f3",
          4944 => x"ec",
          4945 => x"38",
          4946 => x"53",
          4947 => x"ff",
          4948 => x"16",
          4949 => x"06",
          4950 => x"76",
          4951 => x"ff",
          4952 => x"ec",
          4953 => x"3d",
          4954 => x"3d",
          4955 => x"71",
          4956 => x"8e",
          4957 => x"29",
          4958 => x"05",
          4959 => x"04",
          4960 => x"51",
          4961 => x"81",
          4962 => x"80",
          4963 => x"df",
          4964 => x"f2",
          4965 => x"b0",
          4966 => x"39",
          4967 => x"51",
          4968 => x"81",
          4969 => x"80",
          4970 => x"df",
          4971 => x"d6",
          4972 => x"f4",
          4973 => x"39",
          4974 => x"51",
          4975 => x"81",
          4976 => x"80",
          4977 => x"e0",
          4978 => x"39",
          4979 => x"51",
          4980 => x"e0",
          4981 => x"39",
          4982 => x"51",
          4983 => x"e1",
          4984 => x"39",
          4985 => x"51",
          4986 => x"e1",
          4987 => x"39",
          4988 => x"51",
          4989 => x"e2",
          4990 => x"39",
          4991 => x"51",
          4992 => x"e2",
          4993 => x"86",
          4994 => x"3d",
          4995 => x"3d",
          4996 => x"56",
          4997 => x"e7",
          4998 => x"74",
          4999 => x"e8",
          5000 => x"39",
          5001 => x"74",
          5002 => x"82",
          5003 => x"e0",
          5004 => x"51",
          5005 => x"3f",
          5006 => x"08",
          5007 => x"75",
          5008 => x"c4",
          5009 => x"c4",
          5010 => x"0d",
          5011 => x"0d",
          5012 => x"05",
          5013 => x"33",
          5014 => x"68",
          5015 => x"7a",
          5016 => x"51",
          5017 => x"78",
          5018 => x"ff",
          5019 => x"81",
          5020 => x"07",
          5021 => x"06",
          5022 => x"56",
          5023 => x"38",
          5024 => x"52",
          5025 => x"52",
          5026 => x"3f",
          5027 => x"08",
          5028 => x"e0",
          5029 => x"81",
          5030 => x"87",
          5031 => x"0c",
          5032 => x"08",
          5033 => x"d4",
          5034 => x"80",
          5035 => x"75",
          5036 => x"3f",
          5037 => x"08",
          5038 => x"e0",
          5039 => x"7a",
          5040 => x"2e",
          5041 => x"19",
          5042 => x"59",
          5043 => x"3d",
          5044 => x"cd",
          5045 => x"30",
          5046 => x"80",
          5047 => x"70",
          5048 => x"06",
          5049 => x"56",
          5050 => x"90",
          5051 => x"e8",
          5052 => x"98",
          5053 => x"78",
          5054 => x"3f",
          5055 => x"81",
          5056 => x"96",
          5057 => x"f9",
          5058 => x"02",
          5059 => x"05",
          5060 => x"ff",
          5061 => x"7a",
          5062 => x"fe",
          5063 => x"ec",
          5064 => x"38",
          5065 => x"88",
          5066 => x"2e",
          5067 => x"39",
          5068 => x"54",
          5069 => x"53",
          5070 => x"51",
          5071 => x"ec",
          5072 => x"83",
          5073 => x"76",
          5074 => x"0c",
          5075 => x"04",
          5076 => x"7f",
          5077 => x"8c",
          5078 => x"05",
          5079 => x"15",
          5080 => x"5c",
          5081 => x"5e",
          5082 => x"e2",
          5083 => x"89",
          5084 => x"e2",
          5085 => x"83",
          5086 => x"55",
          5087 => x"80",
          5088 => x"90",
          5089 => x"7b",
          5090 => x"38",
          5091 => x"74",
          5092 => x"7a",
          5093 => x"72",
          5094 => x"e2",
          5095 => x"88",
          5096 => x"39",
          5097 => x"51",
          5098 => x"3f",
          5099 => x"80",
          5100 => x"18",
          5101 => x"27",
          5102 => x"08",
          5103 => x"f0",
          5104 => x"c8",
          5105 => x"81",
          5106 => x"ff",
          5107 => x"84",
          5108 => x"39",
          5109 => x"72",
          5110 => x"38",
          5111 => x"81",
          5112 => x"ff",
          5113 => x"89",
          5114 => x"98",
          5115 => x"b8",
          5116 => x"55",
          5117 => x"81",
          5118 => x"80",
          5119 => x"9c",
          5120 => x"a4",
          5121 => x"74",
          5122 => x"38",
          5123 => x"33",
          5124 => x"56",
          5125 => x"83",
          5126 => x"80",
          5127 => x"27",
          5128 => x"53",
          5129 => x"70",
          5130 => x"51",
          5131 => x"2e",
          5132 => x"80",
          5133 => x"38",
          5134 => x"39",
          5135 => x"81",
          5136 => x"15",
          5137 => x"81",
          5138 => x"ff",
          5139 => x"78",
          5140 => x"5c",
          5141 => x"dc",
          5142 => x"e0",
          5143 => x"70",
          5144 => x"57",
          5145 => x"09",
          5146 => x"38",
          5147 => x"3f",
          5148 => x"08",
          5149 => x"98",
          5150 => x"32",
          5151 => x"9b",
          5152 => x"70",
          5153 => x"75",
          5154 => x"58",
          5155 => x"51",
          5156 => x"24",
          5157 => x"9b",
          5158 => x"06",
          5159 => x"53",
          5160 => x"1e",
          5161 => x"26",
          5162 => x"ff",
          5163 => x"ec",
          5164 => x"3d",
          5165 => x"3d",
          5166 => x"05",
          5167 => x"a4",
          5168 => x"a8",
          5169 => x"86",
          5170 => x"e9",
          5171 => x"fe",
          5172 => x"81",
          5173 => x"81",
          5174 => x"81",
          5175 => x"52",
          5176 => x"51",
          5177 => x"3f",
          5178 => x"85",
          5179 => x"e8",
          5180 => x"0d",
          5181 => x"0d",
          5182 => x"80",
          5183 => x"ff",
          5184 => x"51",
          5185 => x"3f",
          5186 => x"51",
          5187 => x"3f",
          5188 => x"f1",
          5189 => x"81",
          5190 => x"06",
          5191 => x"80",
          5192 => x"81",
          5193 => x"a0",
          5194 => x"fc",
          5195 => x"98",
          5196 => x"fe",
          5197 => x"72",
          5198 => x"81",
          5199 => x"71",
          5200 => x"38",
          5201 => x"f0",
          5202 => x"e4",
          5203 => x"f2",
          5204 => x"51",
          5205 => x"3f",
          5206 => x"70",
          5207 => x"52",
          5208 => x"95",
          5209 => x"fe",
          5210 => x"81",
          5211 => x"fe",
          5212 => x"80",
          5213 => x"d0",
          5214 => x"2a",
          5215 => x"51",
          5216 => x"2e",
          5217 => x"51",
          5218 => x"3f",
          5219 => x"51",
          5220 => x"3f",
          5221 => x"f0",
          5222 => x"85",
          5223 => x"06",
          5224 => x"80",
          5225 => x"81",
          5226 => x"9c",
          5227 => x"c8",
          5228 => x"94",
          5229 => x"fe",
          5230 => x"72",
          5231 => x"81",
          5232 => x"71",
          5233 => x"38",
          5234 => x"ef",
          5235 => x"e4",
          5236 => x"f1",
          5237 => x"51",
          5238 => x"3f",
          5239 => x"70",
          5240 => x"52",
          5241 => x"95",
          5242 => x"fe",
          5243 => x"81",
          5244 => x"fe",
          5245 => x"80",
          5246 => x"cc",
          5247 => x"2a",
          5248 => x"51",
          5249 => x"2e",
          5250 => x"51",
          5251 => x"3f",
          5252 => x"51",
          5253 => x"3f",
          5254 => x"ef",
          5255 => x"fd",
          5256 => x"3d",
          5257 => x"3d",
          5258 => x"70",
          5259 => x"80",
          5260 => x"fe",
          5261 => x"81",
          5262 => x"54",
          5263 => x"81",
          5264 => x"c4",
          5265 => x"e4",
          5266 => x"dc",
          5267 => x"e0",
          5268 => x"81",
          5269 => x"07",
          5270 => x"71",
          5271 => x"54",
          5272 => x"ec",
          5273 => x"ec",
          5274 => x"81",
          5275 => x"06",
          5276 => x"83",
          5277 => x"52",
          5278 => x"92",
          5279 => x"e0",
          5280 => x"8c",
          5281 => x"e0",
          5282 => x"fd",
          5283 => x"39",
          5284 => x"51",
          5285 => x"82",
          5286 => x"ec",
          5287 => x"ec",
          5288 => x"82",
          5289 => x"06",
          5290 => x"52",
          5291 => x"83",
          5292 => x"0b",
          5293 => x"0c",
          5294 => x"04",
          5295 => x"80",
          5296 => x"83",
          5297 => x"5d",
          5298 => x"51",
          5299 => x"3f",
          5300 => x"08",
          5301 => x"59",
          5302 => x"09",
          5303 => x"38",
          5304 => x"52",
          5305 => x"52",
          5306 => x"b6",
          5307 => x"78",
          5308 => x"90",
          5309 => x"cf",
          5310 => x"e0",
          5311 => x"88",
          5312 => x"d8",
          5313 => x"39",
          5314 => x"5d",
          5315 => x"51",
          5316 => x"3f",
          5317 => x"46",
          5318 => x"52",
          5319 => x"86",
          5320 => x"ff",
          5321 => x"f3",
          5322 => x"ec",
          5323 => x"2b",
          5324 => x"51",
          5325 => x"c2",
          5326 => x"38",
          5327 => x"24",
          5328 => x"bd",
          5329 => x"38",
          5330 => x"90",
          5331 => x"2e",
          5332 => x"78",
          5333 => x"da",
          5334 => x"39",
          5335 => x"2e",
          5336 => x"78",
          5337 => x"85",
          5338 => x"bf",
          5339 => x"38",
          5340 => x"78",
          5341 => x"89",
          5342 => x"80",
          5343 => x"38",
          5344 => x"2e",
          5345 => x"78",
          5346 => x"89",
          5347 => x"b4",
          5348 => x"83",
          5349 => x"38",
          5350 => x"24",
          5351 => x"81",
          5352 => x"fd",
          5353 => x"39",
          5354 => x"2e",
          5355 => x"8a",
          5356 => x"3d",
          5357 => x"53",
          5358 => x"51",
          5359 => x"3f",
          5360 => x"08",
          5361 => x"c4",
          5362 => x"fe",
          5363 => x"ff",
          5364 => x"ff",
          5365 => x"81",
          5366 => x"80",
          5367 => x"38",
          5368 => x"f8",
          5369 => x"84",
          5370 => x"82",
          5371 => x"ec",
          5372 => x"38",
          5373 => x"08",
          5374 => x"94",
          5375 => x"a8",
          5376 => x"5c",
          5377 => x"27",
          5378 => x"61",
          5379 => x"70",
          5380 => x"0c",
          5381 => x"f5",
          5382 => x"39",
          5383 => x"80",
          5384 => x"84",
          5385 => x"81",
          5386 => x"ec",
          5387 => x"2e",
          5388 => x"b4",
          5389 => x"11",
          5390 => x"05",
          5391 => x"c1",
          5392 => x"e0",
          5393 => x"fd",
          5394 => x"3d",
          5395 => x"53",
          5396 => x"51",
          5397 => x"3f",
          5398 => x"08",
          5399 => x"ac",
          5400 => x"a4",
          5401 => x"c0",
          5402 => x"79",
          5403 => x"8c",
          5404 => x"79",
          5405 => x"5b",
          5406 => x"61",
          5407 => x"eb",
          5408 => x"ff",
          5409 => x"ff",
          5410 => x"ff",
          5411 => x"81",
          5412 => x"80",
          5413 => x"38",
          5414 => x"fc",
          5415 => x"84",
          5416 => x"80",
          5417 => x"ec",
          5418 => x"2e",
          5419 => x"b4",
          5420 => x"11",
          5421 => x"05",
          5422 => x"c5",
          5423 => x"e0",
          5424 => x"fc",
          5425 => x"e6",
          5426 => x"f8",
          5427 => x"5a",
          5428 => x"a8",
          5429 => x"33",
          5430 => x"5a",
          5431 => x"2e",
          5432 => x"55",
          5433 => x"33",
          5434 => x"81",
          5435 => x"fe",
          5436 => x"81",
          5437 => x"05",
          5438 => x"39",
          5439 => x"51",
          5440 => x"b4",
          5441 => x"11",
          5442 => x"05",
          5443 => x"f1",
          5444 => x"e0",
          5445 => x"38",
          5446 => x"33",
          5447 => x"2e",
          5448 => x"e9",
          5449 => x"80",
          5450 => x"e9",
          5451 => x"78",
          5452 => x"38",
          5453 => x"08",
          5454 => x"81",
          5455 => x"59",
          5456 => x"88",
          5457 => x"9c",
          5458 => x"39",
          5459 => x"33",
          5460 => x"2e",
          5461 => x"e9",
          5462 => x"9a",
          5463 => x"d2",
          5464 => x"80",
          5465 => x"81",
          5466 => x"44",
          5467 => x"e9",
          5468 => x"80",
          5469 => x"3d",
          5470 => x"53",
          5471 => x"51",
          5472 => x"3f",
          5473 => x"08",
          5474 => x"81",
          5475 => x"59",
          5476 => x"89",
          5477 => x"90",
          5478 => x"cc",
          5479 => x"d5",
          5480 => x"80",
          5481 => x"81",
          5482 => x"43",
          5483 => x"e9",
          5484 => x"78",
          5485 => x"38",
          5486 => x"08",
          5487 => x"81",
          5488 => x"59",
          5489 => x"88",
          5490 => x"a8",
          5491 => x"39",
          5492 => x"33",
          5493 => x"2e",
          5494 => x"e9",
          5495 => x"88",
          5496 => x"bc",
          5497 => x"43",
          5498 => x"f8",
          5499 => x"84",
          5500 => x"fe",
          5501 => x"ec",
          5502 => x"2e",
          5503 => x"62",
          5504 => x"88",
          5505 => x"81",
          5506 => x"32",
          5507 => x"72",
          5508 => x"70",
          5509 => x"51",
          5510 => x"80",
          5511 => x"7a",
          5512 => x"38",
          5513 => x"e6",
          5514 => x"f5",
          5515 => x"55",
          5516 => x"53",
          5517 => x"51",
          5518 => x"81",
          5519 => x"fe",
          5520 => x"f9",
          5521 => x"3d",
          5522 => x"53",
          5523 => x"51",
          5524 => x"3f",
          5525 => x"08",
          5526 => x"b0",
          5527 => x"fe",
          5528 => x"ff",
          5529 => x"fe",
          5530 => x"81",
          5531 => x"80",
          5532 => x"63",
          5533 => x"cb",
          5534 => x"34",
          5535 => x"44",
          5536 => x"fc",
          5537 => x"84",
          5538 => x"fc",
          5539 => x"ec",
          5540 => x"38",
          5541 => x"63",
          5542 => x"52",
          5543 => x"51",
          5544 => x"3f",
          5545 => x"79",
          5546 => x"ba",
          5547 => x"79",
          5548 => x"ae",
          5549 => x"38",
          5550 => x"a0",
          5551 => x"fe",
          5552 => x"ff",
          5553 => x"fe",
          5554 => x"81",
          5555 => x"80",
          5556 => x"63",
          5557 => x"cb",
          5558 => x"34",
          5559 => x"44",
          5560 => x"81",
          5561 => x"fe",
          5562 => x"ff",
          5563 => x"3d",
          5564 => x"53",
          5565 => x"51",
          5566 => x"3f",
          5567 => x"08",
          5568 => x"88",
          5569 => x"fe",
          5570 => x"ff",
          5571 => x"fe",
          5572 => x"81",
          5573 => x"80",
          5574 => x"60",
          5575 => x"05",
          5576 => x"82",
          5577 => x"78",
          5578 => x"fe",
          5579 => x"ff",
          5580 => x"fe",
          5581 => x"81",
          5582 => x"df",
          5583 => x"39",
          5584 => x"54",
          5585 => x"8c",
          5586 => x"c0",
          5587 => x"52",
          5588 => x"fa",
          5589 => x"45",
          5590 => x"78",
          5591 => x"ac",
          5592 => x"26",
          5593 => x"82",
          5594 => x"39",
          5595 => x"f0",
          5596 => x"84",
          5597 => x"fc",
          5598 => x"ec",
          5599 => x"2e",
          5600 => x"59",
          5601 => x"22",
          5602 => x"05",
          5603 => x"41",
          5604 => x"81",
          5605 => x"fe",
          5606 => x"ff",
          5607 => x"3d",
          5608 => x"53",
          5609 => x"51",
          5610 => x"3f",
          5611 => x"08",
          5612 => x"d8",
          5613 => x"fe",
          5614 => x"ff",
          5615 => x"fe",
          5616 => x"81",
          5617 => x"80",
          5618 => x"60",
          5619 => x"59",
          5620 => x"41",
          5621 => x"f0",
          5622 => x"84",
          5623 => x"fc",
          5624 => x"ec",
          5625 => x"38",
          5626 => x"60",
          5627 => x"52",
          5628 => x"51",
          5629 => x"3f",
          5630 => x"79",
          5631 => x"e6",
          5632 => x"79",
          5633 => x"ae",
          5634 => x"38",
          5635 => x"9c",
          5636 => x"fe",
          5637 => x"ff",
          5638 => x"fe",
          5639 => x"81",
          5640 => x"80",
          5641 => x"60",
          5642 => x"59",
          5643 => x"41",
          5644 => x"81",
          5645 => x"fe",
          5646 => x"ff",
          5647 => x"3d",
          5648 => x"53",
          5649 => x"51",
          5650 => x"3f",
          5651 => x"08",
          5652 => x"b8",
          5653 => x"81",
          5654 => x"fe",
          5655 => x"63",
          5656 => x"b4",
          5657 => x"11",
          5658 => x"05",
          5659 => x"91",
          5660 => x"e0",
          5661 => x"f5",
          5662 => x"52",
          5663 => x"51",
          5664 => x"3f",
          5665 => x"2d",
          5666 => x"08",
          5667 => x"fc",
          5668 => x"e0",
          5669 => x"e7",
          5670 => x"f6",
          5671 => x"ec",
          5672 => x"f8",
          5673 => x"80",
          5674 => x"e2",
          5675 => x"39",
          5676 => x"51",
          5677 => x"3f",
          5678 => x"a5",
          5679 => x"98",
          5680 => x"39",
          5681 => x"51",
          5682 => x"2e",
          5683 => x"7d",
          5684 => x"78",
          5685 => x"d8",
          5686 => x"ff",
          5687 => x"fe",
          5688 => x"81",
          5689 => x"5c",
          5690 => x"82",
          5691 => x"7a",
          5692 => x"38",
          5693 => x"8c",
          5694 => x"39",
          5695 => x"b0",
          5696 => x"39",
          5697 => x"56",
          5698 => x"e8",
          5699 => x"53",
          5700 => x"52",
          5701 => x"b0",
          5702 => x"f6",
          5703 => x"39",
          5704 => x"52",
          5705 => x"b0",
          5706 => x"f5",
          5707 => x"39",
          5708 => x"e8",
          5709 => x"53",
          5710 => x"52",
          5711 => x"b0",
          5712 => x"f5",
          5713 => x"39",
          5714 => x"53",
          5715 => x"52",
          5716 => x"b0",
          5717 => x"f5",
          5718 => x"e9",
          5719 => x"ed",
          5720 => x"56",
          5721 => x"46",
          5722 => x"80",
          5723 => x"80",
          5724 => x"80",
          5725 => x"ff",
          5726 => x"eb",
          5727 => x"ec",
          5728 => x"ec",
          5729 => x"70",
          5730 => x"07",
          5731 => x"5b",
          5732 => x"5a",
          5733 => x"83",
          5734 => x"78",
          5735 => x"78",
          5736 => x"38",
          5737 => x"81",
          5738 => x"59",
          5739 => x"38",
          5740 => x"7d",
          5741 => x"59",
          5742 => x"7e",
          5743 => x"81",
          5744 => x"38",
          5745 => x"51",
          5746 => x"3f",
          5747 => x"fc",
          5748 => x"0b",
          5749 => x"34",
          5750 => x"8c",
          5751 => x"55",
          5752 => x"52",
          5753 => x"d6",
          5754 => x"ec",
          5755 => x"2b",
          5756 => x"53",
          5757 => x"52",
          5758 => x"d6",
          5759 => x"81",
          5760 => x"07",
          5761 => x"c0",
          5762 => x"08",
          5763 => x"84",
          5764 => x"51",
          5765 => x"3f",
          5766 => x"08",
          5767 => x"08",
          5768 => x"84",
          5769 => x"51",
          5770 => x"3f",
          5771 => x"e0",
          5772 => x"0c",
          5773 => x"0b",
          5774 => x"84",
          5775 => x"83",
          5776 => x"94",
          5777 => x"df",
          5778 => x"f0",
          5779 => x"0b",
          5780 => x"0c",
          5781 => x"3f",
          5782 => x"3f",
          5783 => x"51",
          5784 => x"3f",
          5785 => x"51",
          5786 => x"3f",
          5787 => x"51",
          5788 => x"3f",
          5789 => x"be",
          5790 => x"3f",
          5791 => x"00",
          5792 => x"00",
          5793 => x"00",
          5794 => x"00",
          5795 => x"00",
          5796 => x"00",
          5797 => x"00",
          5798 => x"00",
          5799 => x"00",
          5800 => x"00",
          5801 => x"00",
          5802 => x"00",
          5803 => x"00",
          5804 => x"00",
          5805 => x"00",
          5806 => x"00",
          5807 => x"00",
          5808 => x"00",
          5809 => x"00",
          5810 => x"00",
          5811 => x"00",
          5812 => x"00",
          5813 => x"00",
          5814 => x"00",
          5815 => x"00",
          5816 => x"25",
          5817 => x"64",
          5818 => x"20",
          5819 => x"25",
          5820 => x"64",
          5821 => x"25",
          5822 => x"53",
          5823 => x"43",
          5824 => x"69",
          5825 => x"61",
          5826 => x"6e",
          5827 => x"20",
          5828 => x"6f",
          5829 => x"6f",
          5830 => x"6f",
          5831 => x"67",
          5832 => x"3a",
          5833 => x"76",
          5834 => x"73",
          5835 => x"70",
          5836 => x"65",
          5837 => x"64",
          5838 => x"20",
          5839 => x"57",
          5840 => x"44",
          5841 => x"20",
          5842 => x"30",
          5843 => x"25",
          5844 => x"29",
          5845 => x"20",
          5846 => x"53",
          5847 => x"4d",
          5848 => x"20",
          5849 => x"30",
          5850 => x"25",
          5851 => x"29",
          5852 => x"20",
          5853 => x"49",
          5854 => x"20",
          5855 => x"4d",
          5856 => x"30",
          5857 => x"25",
          5858 => x"29",
          5859 => x"20",
          5860 => x"42",
          5861 => x"20",
          5862 => x"20",
          5863 => x"30",
          5864 => x"25",
          5865 => x"29",
          5866 => x"20",
          5867 => x"52",
          5868 => x"20",
          5869 => x"20",
          5870 => x"30",
          5871 => x"25",
          5872 => x"29",
          5873 => x"20",
          5874 => x"53",
          5875 => x"41",
          5876 => x"20",
          5877 => x"65",
          5878 => x"65",
          5879 => x"25",
          5880 => x"29",
          5881 => x"20",
          5882 => x"54",
          5883 => x"52",
          5884 => x"20",
          5885 => x"69",
          5886 => x"73",
          5887 => x"25",
          5888 => x"29",
          5889 => x"20",
          5890 => x"49",
          5891 => x"20",
          5892 => x"4c",
          5893 => x"68",
          5894 => x"65",
          5895 => x"25",
          5896 => x"29",
          5897 => x"20",
          5898 => x"57",
          5899 => x"42",
          5900 => x"20",
          5901 => x"0a",
          5902 => x"20",
          5903 => x"57",
          5904 => x"32",
          5905 => x"20",
          5906 => x"49",
          5907 => x"4c",
          5908 => x"20",
          5909 => x"50",
          5910 => x"00",
          5911 => x"20",
          5912 => x"53",
          5913 => x"00",
          5914 => x"41",
          5915 => x"65",
          5916 => x"73",
          5917 => x"20",
          5918 => x"43",
          5919 => x"52",
          5920 => x"74",
          5921 => x"63",
          5922 => x"20",
          5923 => x"72",
          5924 => x"20",
          5925 => x"30",
          5926 => x"00",
          5927 => x"20",
          5928 => x"43",
          5929 => x"4d",
          5930 => x"72",
          5931 => x"74",
          5932 => x"20",
          5933 => x"72",
          5934 => x"20",
          5935 => x"30",
          5936 => x"00",
          5937 => x"20",
          5938 => x"53",
          5939 => x"6b",
          5940 => x"61",
          5941 => x"41",
          5942 => x"65",
          5943 => x"20",
          5944 => x"20",
          5945 => x"30",
          5946 => x"00",
          5947 => x"4d",
          5948 => x"3a",
          5949 => x"20",
          5950 => x"5a",
          5951 => x"49",
          5952 => x"20",
          5953 => x"20",
          5954 => x"20",
          5955 => x"20",
          5956 => x"20",
          5957 => x"30",
          5958 => x"00",
          5959 => x"20",
          5960 => x"53",
          5961 => x"65",
          5962 => x"6c",
          5963 => x"20",
          5964 => x"71",
          5965 => x"20",
          5966 => x"20",
          5967 => x"64",
          5968 => x"34",
          5969 => x"7a",
          5970 => x"20",
          5971 => x"53",
          5972 => x"4d",
          5973 => x"6f",
          5974 => x"46",
          5975 => x"20",
          5976 => x"20",
          5977 => x"20",
          5978 => x"64",
          5979 => x"34",
          5980 => x"7a",
          5981 => x"20",
          5982 => x"57",
          5983 => x"62",
          5984 => x"20",
          5985 => x"41",
          5986 => x"6c",
          5987 => x"20",
          5988 => x"71",
          5989 => x"64",
          5990 => x"34",
          5991 => x"7a",
          5992 => x"53",
          5993 => x"6c",
          5994 => x"4d",
          5995 => x"75",
          5996 => x"46",
          5997 => x"00",
          5998 => x"45",
          5999 => x"45",
          6000 => x"69",
          6001 => x"55",
          6002 => x"6f",
          6003 => x"53",
          6004 => x"22",
          6005 => x"3a",
          6006 => x"3e",
          6007 => x"7c",
          6008 => x"46",
          6009 => x"46",
          6010 => x"32",
          6011 => x"eb",
          6012 => x"53",
          6013 => x"35",
          6014 => x"4e",
          6015 => x"41",
          6016 => x"20",
          6017 => x"41",
          6018 => x"20",
          6019 => x"4e",
          6020 => x"41",
          6021 => x"20",
          6022 => x"41",
          6023 => x"20",
          6024 => x"00",
          6025 => x"00",
          6026 => x"00",
          6027 => x"00",
          6028 => x"80",
          6029 => x"8e",
          6030 => x"45",
          6031 => x"49",
          6032 => x"90",
          6033 => x"99",
          6034 => x"59",
          6035 => x"9c",
          6036 => x"41",
          6037 => x"a5",
          6038 => x"a8",
          6039 => x"ac",
          6040 => x"b0",
          6041 => x"b4",
          6042 => x"b8",
          6043 => x"bc",
          6044 => x"c0",
          6045 => x"c4",
          6046 => x"c8",
          6047 => x"cc",
          6048 => x"d0",
          6049 => x"d4",
          6050 => x"d8",
          6051 => x"dc",
          6052 => x"e0",
          6053 => x"e4",
          6054 => x"e8",
          6055 => x"ec",
          6056 => x"f0",
          6057 => x"f4",
          6058 => x"f8",
          6059 => x"fc",
          6060 => x"2b",
          6061 => x"3d",
          6062 => x"5c",
          6063 => x"3c",
          6064 => x"7f",
          6065 => x"00",
          6066 => x"00",
          6067 => x"01",
          6068 => x"00",
          6069 => x"00",
          6070 => x"00",
          6071 => x"00",
          6072 => x"00",
          6073 => x"64",
          6074 => x"74",
          6075 => x"64",
          6076 => x"74",
          6077 => x"66",
          6078 => x"74",
          6079 => x"66",
          6080 => x"64",
          6081 => x"66",
          6082 => x"63",
          6083 => x"6d",
          6084 => x"61",
          6085 => x"6d",
          6086 => x"79",
          6087 => x"6d",
          6088 => x"66",
          6089 => x"6d",
          6090 => x"70",
          6091 => x"6d",
          6092 => x"6d",
          6093 => x"6d",
          6094 => x"68",
          6095 => x"68",
          6096 => x"68",
          6097 => x"68",
          6098 => x"63",
          6099 => x"00",
          6100 => x"6a",
          6101 => x"72",
          6102 => x"61",
          6103 => x"72",
          6104 => x"74",
          6105 => x"69",
          6106 => x"00",
          6107 => x"74",
          6108 => x"00",
          6109 => x"74",
          6110 => x"69",
          6111 => x"44",
          6112 => x"20",
          6113 => x"6f",
          6114 => x"49",
          6115 => x"72",
          6116 => x"20",
          6117 => x"6f",
          6118 => x"00",
          6119 => x"44",
          6120 => x"20",
          6121 => x"20",
          6122 => x"64",
          6123 => x"00",
          6124 => x"4e",
          6125 => x"69",
          6126 => x"66",
          6127 => x"64",
          6128 => x"4e",
          6129 => x"61",
          6130 => x"66",
          6131 => x"64",
          6132 => x"49",
          6133 => x"6c",
          6134 => x"66",
          6135 => x"6e",
          6136 => x"2e",
          6137 => x"41",
          6138 => x"73",
          6139 => x"65",
          6140 => x"64",
          6141 => x"46",
          6142 => x"20",
          6143 => x"65",
          6144 => x"20",
          6145 => x"73",
          6146 => x"0a",
          6147 => x"46",
          6148 => x"20",
          6149 => x"64",
          6150 => x"69",
          6151 => x"6c",
          6152 => x"0a",
          6153 => x"53",
          6154 => x"73",
          6155 => x"69",
          6156 => x"70",
          6157 => x"65",
          6158 => x"64",
          6159 => x"44",
          6160 => x"65",
          6161 => x"6d",
          6162 => x"20",
          6163 => x"69",
          6164 => x"6c",
          6165 => x"0a",
          6166 => x"44",
          6167 => x"20",
          6168 => x"20",
          6169 => x"62",
          6170 => x"2e",
          6171 => x"4e",
          6172 => x"6f",
          6173 => x"74",
          6174 => x"65",
          6175 => x"6c",
          6176 => x"73",
          6177 => x"20",
          6178 => x"6e",
          6179 => x"6e",
          6180 => x"73",
          6181 => x"00",
          6182 => x"46",
          6183 => x"61",
          6184 => x"62",
          6185 => x"65",
          6186 => x"00",
          6187 => x"54",
          6188 => x"6f",
          6189 => x"20",
          6190 => x"72",
          6191 => x"6f",
          6192 => x"61",
          6193 => x"6c",
          6194 => x"2e",
          6195 => x"46",
          6196 => x"20",
          6197 => x"6c",
          6198 => x"65",
          6199 => x"00",
          6200 => x"49",
          6201 => x"66",
          6202 => x"69",
          6203 => x"20",
          6204 => x"6f",
          6205 => x"0a",
          6206 => x"54",
          6207 => x"6d",
          6208 => x"20",
          6209 => x"6e",
          6210 => x"6c",
          6211 => x"0a",
          6212 => x"50",
          6213 => x"6d",
          6214 => x"72",
          6215 => x"6e",
          6216 => x"72",
          6217 => x"2e",
          6218 => x"53",
          6219 => x"65",
          6220 => x"0a",
          6221 => x"55",
          6222 => x"6f",
          6223 => x"65",
          6224 => x"72",
          6225 => x"0a",
          6226 => x"20",
          6227 => x"65",
          6228 => x"73",
          6229 => x"20",
          6230 => x"20",
          6231 => x"65",
          6232 => x"65",
          6233 => x"00",
          6234 => x"72",
          6235 => x"00",
          6236 => x"25",
          6237 => x"00",
          6238 => x"3a",
          6239 => x"25",
          6240 => x"00",
          6241 => x"20",
          6242 => x"20",
          6243 => x"00",
          6244 => x"25",
          6245 => x"00",
          6246 => x"20",
          6247 => x"20",
          6248 => x"7c",
          6249 => x"7a",
          6250 => x"0a",
          6251 => x"25",
          6252 => x"00",
          6253 => x"31",
          6254 => x"34",
          6255 => x"32",
          6256 => x"76",
          6257 => x"00",
          6258 => x"20",
          6259 => x"2c",
          6260 => x"76",
          6261 => x"32",
          6262 => x"25",
          6263 => x"73",
          6264 => x"0a",
          6265 => x"5a",
          6266 => x"49",
          6267 => x"72",
          6268 => x"74",
          6269 => x"6e",
          6270 => x"72",
          6271 => x"54",
          6272 => x"72",
          6273 => x"74",
          6274 => x"75",
          6275 => x"00",
          6276 => x"50",
          6277 => x"69",
          6278 => x"72",
          6279 => x"74",
          6280 => x"49",
          6281 => x"4c",
          6282 => x"20",
          6283 => x"65",
          6284 => x"70",
          6285 => x"49",
          6286 => x"4c",
          6287 => x"20",
          6288 => x"65",
          6289 => x"70",
          6290 => x"55",
          6291 => x"30",
          6292 => x"20",
          6293 => x"65",
          6294 => x"70",
          6295 => x"55",
          6296 => x"30",
          6297 => x"20",
          6298 => x"65",
          6299 => x"70",
          6300 => x"55",
          6301 => x"31",
          6302 => x"20",
          6303 => x"65",
          6304 => x"70",
          6305 => x"55",
          6306 => x"31",
          6307 => x"20",
          6308 => x"65",
          6309 => x"70",
          6310 => x"53",
          6311 => x"69",
          6312 => x"75",
          6313 => x"69",
          6314 => x"2e",
          6315 => x"00",
          6316 => x"45",
          6317 => x"6c",
          6318 => x"20",
          6319 => x"65",
          6320 => x"2e",
          6321 => x"61",
          6322 => x"65",
          6323 => x"2e",
          6324 => x"00",
          6325 => x"30",
          6326 => x"46",
          6327 => x"65",
          6328 => x"6f",
          6329 => x"69",
          6330 => x"6c",
          6331 => x"20",
          6332 => x"63",
          6333 => x"20",
          6334 => x"70",
          6335 => x"73",
          6336 => x"6e",
          6337 => x"6d",
          6338 => x"61",
          6339 => x"2e",
          6340 => x"2a",
          6341 => x"43",
          6342 => x"72",
          6343 => x"2e",
          6344 => x"00",
          6345 => x"43",
          6346 => x"69",
          6347 => x"2e",
          6348 => x"43",
          6349 => x"61",
          6350 => x"67",
          6351 => x"00",
          6352 => x"25",
          6353 => x"78",
          6354 => x"38",
          6355 => x"3e",
          6356 => x"6c",
          6357 => x"30",
          6358 => x"0a",
          6359 => x"44",
          6360 => x"20",
          6361 => x"6f",
          6362 => x"00",
          6363 => x"0a",
          6364 => x"70",
          6365 => x"65",
          6366 => x"25",
          6367 => x"20",
          6368 => x"58",
          6369 => x"3f",
          6370 => x"00",
          6371 => x"25",
          6372 => x"20",
          6373 => x"58",
          6374 => x"25",
          6375 => x"20",
          6376 => x"58",
          6377 => x"45",
          6378 => x"75",
          6379 => x"67",
          6380 => x"64",
          6381 => x"20",
          6382 => x"78",
          6383 => x"2e",
          6384 => x"43",
          6385 => x"69",
          6386 => x"63",
          6387 => x"20",
          6388 => x"30",
          6389 => x"2e",
          6390 => x"00",
          6391 => x"43",
          6392 => x"20",
          6393 => x"75",
          6394 => x"64",
          6395 => x"64",
          6396 => x"25",
          6397 => x"0a",
          6398 => x"52",
          6399 => x"61",
          6400 => x"6e",
          6401 => x"70",
          6402 => x"63",
          6403 => x"6f",
          6404 => x"2e",
          6405 => x"43",
          6406 => x"20",
          6407 => x"6f",
          6408 => x"6e",
          6409 => x"2e",
          6410 => x"5a",
          6411 => x"62",
          6412 => x"25",
          6413 => x"25",
          6414 => x"73",
          6415 => x"00",
          6416 => x"25",
          6417 => x"25",
          6418 => x"73",
          6419 => x"25",
          6420 => x"25",
          6421 => x"42",
          6422 => x"63",
          6423 => x"61",
          6424 => x"0a",
          6425 => x"52",
          6426 => x"69",
          6427 => x"2e",
          6428 => x"45",
          6429 => x"6c",
          6430 => x"20",
          6431 => x"65",
          6432 => x"70",
          6433 => x"2e",
          6434 => x"00",
          6435 => x"00",
          6436 => x"00",
          6437 => x"00",
          6438 => x"00",
          6439 => x"00",
          6440 => x"00",
          6441 => x"00",
          6442 => x"00",
          6443 => x"01",
          6444 => x"01",
          6445 => x"00",
          6446 => x"00",
          6447 => x"00",
          6448 => x"00",
          6449 => x"05",
          6450 => x"05",
          6451 => x"05",
          6452 => x"00",
          6453 => x"01",
          6454 => x"01",
          6455 => x"01",
          6456 => x"01",
          6457 => x"00",
          6458 => x"01",
          6459 => x"00",
          6460 => x"00",
          6461 => x"01",
          6462 => x"00",
          6463 => x"00",
          6464 => x"00",
          6465 => x"01",
          6466 => x"00",
          6467 => x"00",
          6468 => x"00",
          6469 => x"01",
          6470 => x"00",
          6471 => x"00",
          6472 => x"00",
          6473 => x"01",
          6474 => x"00",
          6475 => x"00",
          6476 => x"00",
          6477 => x"01",
          6478 => x"00",
          6479 => x"00",
          6480 => x"00",
          6481 => x"01",
          6482 => x"00",
          6483 => x"00",
          6484 => x"00",
          6485 => x"01",
          6486 => x"00",
          6487 => x"00",
          6488 => x"00",
          6489 => x"01",
          6490 => x"00",
          6491 => x"00",
          6492 => x"00",
          6493 => x"01",
          6494 => x"00",
          6495 => x"00",
          6496 => x"00",
          6497 => x"01",
          6498 => x"00",
          6499 => x"00",
          6500 => x"00",
          6501 => x"01",
          6502 => x"00",
          6503 => x"00",
          6504 => x"00",
          6505 => x"01",
          6506 => x"00",
          6507 => x"00",
          6508 => x"00",
          6509 => x"01",
          6510 => x"00",
          6511 => x"00",
          6512 => x"00",
          6513 => x"01",
          6514 => x"00",
          6515 => x"00",
          6516 => x"00",
          6517 => x"01",
          6518 => x"00",
          6519 => x"00",
          6520 => x"00",
          6521 => x"01",
          6522 => x"00",
          6523 => x"00",
          6524 => x"00",
          6525 => x"01",
          6526 => x"00",
          6527 => x"00",
          6528 => x"00",
          6529 => x"01",
          6530 => x"00",
          6531 => x"00",
          6532 => x"00",
          6533 => x"01",
          6534 => x"00",
          6535 => x"00",
          6536 => x"00",
          6537 => x"01",
          6538 => x"00",
          6539 => x"00",
          6540 => x"00",
          6541 => x"01",
          6542 => x"00",
          6543 => x"00",
          6544 => x"00",
          6545 => x"01",
          6546 => x"00",
          6547 => x"00",
          6548 => x"00",
          6549 => x"01",
          6550 => x"00",
          6551 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
