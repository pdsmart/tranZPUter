-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b92",
             1 => x"d8040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b92",
            73 => x"bc040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b929f",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b81c5",
           162 => x"f0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"92a40400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b93",
           171 => x"dd2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b95",
           179 => x"c92d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"94040b0b",
           269 => x"0b8ca304",
           270 => x"0b0b0b8c",
           271 => x"b2040b0b",
           272 => x"0b8cc104",
           273 => x"0b0b0b8c",
           274 => x"d0040b0b",
           275 => x"0b8cdf04",
           276 => x"0b0b0b8c",
           277 => x"ee040b0b",
           278 => x"0b8cfd04",
           279 => x"0b0b0b8d",
           280 => x"8c040b0b",
           281 => x"0b8d9b04",
           282 => x"0b0b0b8d",
           283 => x"aa040b0b",
           284 => x"0b8db904",
           285 => x"0b0b0b8d",
           286 => x"c8040b0b",
           287 => x"0b8dd704",
           288 => x"0b0b0b8d",
           289 => x"e6040b0b",
           290 => x"0b8df504",
           291 => x"0b0b0b8e",
           292 => x"84040b0b",
           293 => x"0b8e9404",
           294 => x"0b0b0b8e",
           295 => x"a4040b0b",
           296 => x"0b8eb404",
           297 => x"0b0b0b8e",
           298 => x"c4040b0b",
           299 => x"0b8ed404",
           300 => x"0b0b0b8e",
           301 => x"e4040b0b",
           302 => x"0b8ef404",
           303 => x"0b0b0b8f",
           304 => x"84040b0b",
           305 => x"0b8f9404",
           306 => x"0b0b0b8f",
           307 => x"a4040b0b",
           308 => x"0b8fb404",
           309 => x"0b0b0b8f",
           310 => x"c4040b0b",
           311 => x"0b8fd404",
           312 => x"0b0b0b8f",
           313 => x"e4040b0b",
           314 => x"0b8ff404",
           315 => x"0b0b0b90",
           316 => x"84040b0b",
           317 => x"0b909404",
           318 => x"0b0b0b90",
           319 => x"a4040b0b",
           320 => x"0b90b404",
           321 => x"0b0b0b90",
           322 => x"c4040b0b",
           323 => x"0b90d404",
           324 => x"0b0b0b90",
           325 => x"e4040b0b",
           326 => x"0b90f404",
           327 => x"0b0b0b91",
           328 => x"84040b0b",
           329 => x"0b919404",
           330 => x"0b0b0b91",
           331 => x"a3040b0b",
           332 => x"0b91b204",
           333 => x"0b0b0b91",
           334 => x"c1040b0b",
           335 => x"0b91d004",
           336 => x"0b0b0b91",
           337 => x"df040b0b",
           338 => x"0b91ee04",
           339 => x"ffffffff",
           340 => x"ffffffff",
           341 => x"ffffffff",
           342 => x"ffffffff",
           343 => x"ffffffff",
           344 => x"ffffffff",
           345 => x"ffffffff",
           346 => x"ffffffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0481decc",
           386 => x"0ca0ae2d",
           387 => x"81decc08",
           388 => x"82809004",
           389 => x"81decc0c",
           390 => x"ade22d81",
           391 => x"decc0882",
           392 => x"80900481",
           393 => x"decc0cae",
           394 => x"a12d81de",
           395 => x"cc088280",
           396 => x"900481de",
           397 => x"cc0caebf",
           398 => x"2d81decc",
           399 => x"08828090",
           400 => x"0481decc",
           401 => x"0cb4fd2d",
           402 => x"81decc08",
           403 => x"82809004",
           404 => x"81decc0c",
           405 => x"b5fb2d81",
           406 => x"decc0882",
           407 => x"80900481",
           408 => x"decc0cae",
           409 => x"e22d81de",
           410 => x"cc088280",
           411 => x"900481de",
           412 => x"cc0cb698",
           413 => x"2d81decc",
           414 => x"08828090",
           415 => x"0481decc",
           416 => x"0cb88a2d",
           417 => x"81decc08",
           418 => x"82809004",
           419 => x"81decc0c",
           420 => x"b4a32d81",
           421 => x"decc0882",
           422 => x"80900481",
           423 => x"decc0cb4",
           424 => x"b92d81de",
           425 => x"cc088280",
           426 => x"900481de",
           427 => x"cc0cb4dd",
           428 => x"2d81decc",
           429 => x"08828090",
           430 => x"0481decc",
           431 => x"0ca2bb2d",
           432 => x"81decc08",
           433 => x"82809004",
           434 => x"81decc0c",
           435 => x"a38c2d81",
           436 => x"decc0882",
           437 => x"80900481",
           438 => x"decc0c9b",
           439 => x"a82d81de",
           440 => x"cc088280",
           441 => x"900481de",
           442 => x"cc0c9cdd",
           443 => x"2d81decc",
           444 => x"08828090",
           445 => x"0481decc",
           446 => x"0c9e902d",
           447 => x"81decc08",
           448 => x"82809004",
           449 => x"81decc0c",
           450 => x"80eabf2d",
           451 => x"81decc08",
           452 => x"82809004",
           453 => x"81decc0c",
           454 => x"80f7b02d",
           455 => x"81decc08",
           456 => x"82809004",
           457 => x"81decc0c",
           458 => x"80efa42d",
           459 => x"81decc08",
           460 => x"82809004",
           461 => x"81decc0c",
           462 => x"80f2a12d",
           463 => x"81decc08",
           464 => x"82809004",
           465 => x"81decc0c",
           466 => x"80fcbf2d",
           467 => x"81decc08",
           468 => x"82809004",
           469 => x"81decc0c",
           470 => x"81859f2d",
           471 => x"81decc08",
           472 => x"82809004",
           473 => x"81decc0c",
           474 => x"80f6922d",
           475 => x"81decc08",
           476 => x"82809004",
           477 => x"81decc0c",
           478 => x"80ffde2d",
           479 => x"81decc08",
           480 => x"82809004",
           481 => x"81decc0c",
           482 => x"8180fd2d",
           483 => x"81decc08",
           484 => x"82809004",
           485 => x"81decc0c",
           486 => x"81819c2d",
           487 => x"81decc08",
           488 => x"82809004",
           489 => x"81decc0c",
           490 => x"8189862d",
           491 => x"81decc08",
           492 => x"82809004",
           493 => x"81decc0c",
           494 => x"8186ec2d",
           495 => x"81decc08",
           496 => x"82809004",
           497 => x"81decc0c",
           498 => x"818bda2d",
           499 => x"81decc08",
           500 => x"82809004",
           501 => x"81decc0c",
           502 => x"8182a02d",
           503 => x"81decc08",
           504 => x"82809004",
           505 => x"81decc0c",
           506 => x"818eda2d",
           507 => x"81decc08",
           508 => x"82809004",
           509 => x"81decc0c",
           510 => x"818fdb2d",
           511 => x"81decc08",
           512 => x"82809004",
           513 => x"81decc0c",
           514 => x"80f8902d",
           515 => x"81decc08",
           516 => x"82809004",
           517 => x"81decc0c",
           518 => x"80f7e92d",
           519 => x"81decc08",
           520 => x"82809004",
           521 => x"81decc0c",
           522 => x"80f9942d",
           523 => x"81decc08",
           524 => x"82809004",
           525 => x"81decc0c",
           526 => x"8182f72d",
           527 => x"81decc08",
           528 => x"82809004",
           529 => x"81decc0c",
           530 => x"8190cc2d",
           531 => x"81decc08",
           532 => x"82809004",
           533 => x"81decc0c",
           534 => x"8192d62d",
           535 => x"81decc08",
           536 => x"82809004",
           537 => x"81decc0c",
           538 => x"8196982d",
           539 => x"81decc08",
           540 => x"82809004",
           541 => x"81decc0c",
           542 => x"80e9de2d",
           543 => x"81decc08",
           544 => x"82809004",
           545 => x"81decc0c",
           546 => x"8199842d",
           547 => x"81decc08",
           548 => x"82809004",
           549 => x"81decc0c",
           550 => x"bb992d81",
           551 => x"decc0882",
           552 => x"80900481",
           553 => x"decc0cbd",
           554 => x"832d81de",
           555 => x"cc088280",
           556 => x"900481de",
           557 => x"cc0cbee7",
           558 => x"2d81decc",
           559 => x"08828090",
           560 => x"0481decc",
           561 => x"0c9bd12d",
           562 => x"81decc08",
           563 => x"82809004",
           564 => x"81decc0c",
           565 => x"9cb32d81",
           566 => x"decc0882",
           567 => x"80900481",
           568 => x"decc0c9f",
           569 => x"a02d81de",
           570 => x"cc088280",
           571 => x"900481de",
           572 => x"cc0c81a5",
           573 => x"ff2d81de",
           574 => x"cc088280",
           575 => x"90043c04",
           576 => x"10101010",
           577 => x"10101010",
           578 => x"10101010",
           579 => x"10101010",
           580 => x"10101010",
           581 => x"10101010",
           582 => x"10101010",
           583 => x"10101053",
           584 => x"51040000",
           585 => x"7381ff06",
           586 => x"73830609",
           587 => x"81058305",
           588 => x"1010102b",
           589 => x"0772fc06",
           590 => x"0c515104",
           591 => x"72728072",
           592 => x"8106ff05",
           593 => x"09720605",
           594 => x"71105272",
           595 => x"0a100a53",
           596 => x"72ed3851",
           597 => x"51535104",
           598 => x"81dec070",
           599 => x"81f5ec27",
           600 => x"8e388071",
           601 => x"70840553",
           602 => x"0c0b0b0b",
           603 => x"92db048c",
           604 => x"815181c4",
           605 => x"be040081",
           606 => x"decc0802",
           607 => x"81decc0c",
           608 => x"fd3d0d80",
           609 => x"5381decc",
           610 => x"088c0508",
           611 => x"5281decc",
           612 => x"08880508",
           613 => x"5183d43f",
           614 => x"81dec008",
           615 => x"7081dec0",
           616 => x"0c54853d",
           617 => x"0d81decc",
           618 => x"0c0481de",
           619 => x"cc080281",
           620 => x"decc0cfd",
           621 => x"3d0d8153",
           622 => x"81decc08",
           623 => x"8c050852",
           624 => x"81decc08",
           625 => x"88050851",
           626 => x"83a13f81",
           627 => x"dec00870",
           628 => x"81dec00c",
           629 => x"54853d0d",
           630 => x"81decc0c",
           631 => x"0481decc",
           632 => x"080281de",
           633 => x"cc0cf93d",
           634 => x"0d800b81",
           635 => x"decc08fc",
           636 => x"050c81de",
           637 => x"cc088805",
           638 => x"088025b9",
           639 => x"3881decc",
           640 => x"08880508",
           641 => x"3081decc",
           642 => x"0888050c",
           643 => x"800b81de",
           644 => x"cc08f405",
           645 => x"0c81decc",
           646 => x"08fc0508",
           647 => x"8a38810b",
           648 => x"81decc08",
           649 => x"f4050c81",
           650 => x"decc08f4",
           651 => x"050881de",
           652 => x"cc08fc05",
           653 => x"0c81decc",
           654 => x"088c0508",
           655 => x"8025b938",
           656 => x"81decc08",
           657 => x"8c050830",
           658 => x"81decc08",
           659 => x"8c050c80",
           660 => x"0b81decc",
           661 => x"08f0050c",
           662 => x"81decc08",
           663 => x"fc05088a",
           664 => x"38810b81",
           665 => x"decc08f0",
           666 => x"050c81de",
           667 => x"cc08f005",
           668 => x"0881decc",
           669 => x"08fc050c",
           670 => x"805381de",
           671 => x"cc088c05",
           672 => x"085281de",
           673 => x"cc088805",
           674 => x"085181df",
           675 => x"3f81dec0",
           676 => x"087081de",
           677 => x"cc08f805",
           678 => x"0c5481de",
           679 => x"cc08fc05",
           680 => x"08802e90",
           681 => x"3881decc",
           682 => x"08f80508",
           683 => x"3081decc",
           684 => x"08f8050c",
           685 => x"81decc08",
           686 => x"f8050870",
           687 => x"81dec00c",
           688 => x"54893d0d",
           689 => x"81decc0c",
           690 => x"0481decc",
           691 => x"080281de",
           692 => x"cc0cfb3d",
           693 => x"0d800b81",
           694 => x"decc08fc",
           695 => x"050c81de",
           696 => x"cc088805",
           697 => x"08802599",
           698 => x"3881decc",
           699 => x"08880508",
           700 => x"3081decc",
           701 => x"0888050c",
           702 => x"810b81de",
           703 => x"cc08fc05",
           704 => x"0c81decc",
           705 => x"088c0508",
           706 => x"80259038",
           707 => x"81decc08",
           708 => x"8c050830",
           709 => x"81decc08",
           710 => x"8c050c81",
           711 => x"5381decc",
           712 => x"088c0508",
           713 => x"5281decc",
           714 => x"08880508",
           715 => x"51bd3f81",
           716 => x"dec00870",
           717 => x"81decc08",
           718 => x"f8050c54",
           719 => x"81decc08",
           720 => x"fc050880",
           721 => x"2e903881",
           722 => x"decc08f8",
           723 => x"05083081",
           724 => x"decc08f8",
           725 => x"050c81de",
           726 => x"cc08f805",
           727 => x"087081de",
           728 => x"c00c5487",
           729 => x"3d0d81de",
           730 => x"cc0c0481",
           731 => x"decc0802",
           732 => x"81decc0c",
           733 => x"fd3d0d81",
           734 => x"0b81decc",
           735 => x"08fc050c",
           736 => x"800b81de",
           737 => x"cc08f805",
           738 => x"0c81decc",
           739 => x"088c0508",
           740 => x"81decc08",
           741 => x"88050827",
           742 => x"b93881de",
           743 => x"cc08fc05",
           744 => x"08802eae",
           745 => x"38800b81",
           746 => x"decc088c",
           747 => x"050824a2",
           748 => x"3881decc",
           749 => x"088c0508",
           750 => x"1081decc",
           751 => x"088c050c",
           752 => x"81decc08",
           753 => x"fc050810",
           754 => x"81decc08",
           755 => x"fc050cff",
           756 => x"b83981de",
           757 => x"cc08fc05",
           758 => x"08802e80",
           759 => x"e13881de",
           760 => x"cc088c05",
           761 => x"0881decc",
           762 => x"08880508",
           763 => x"26ad3881",
           764 => x"decc0888",
           765 => x"050881de",
           766 => x"cc088c05",
           767 => x"083181de",
           768 => x"cc088805",
           769 => x"0c81decc",
           770 => x"08f80508",
           771 => x"81decc08",
           772 => x"fc050807",
           773 => x"81decc08",
           774 => x"f8050c81",
           775 => x"decc08fc",
           776 => x"0508812a",
           777 => x"81decc08",
           778 => x"fc050c81",
           779 => x"decc088c",
           780 => x"0508812a",
           781 => x"81decc08",
           782 => x"8c050cff",
           783 => x"953981de",
           784 => x"cc089005",
           785 => x"08802e93",
           786 => x"3881decc",
           787 => x"08880508",
           788 => x"7081decc",
           789 => x"08f4050c",
           790 => x"51913981",
           791 => x"decc08f8",
           792 => x"05087081",
           793 => x"decc08f4",
           794 => x"050c5181",
           795 => x"decc08f4",
           796 => x"050881de",
           797 => x"c00c853d",
           798 => x"0d81decc",
           799 => x"0c04fc3d",
           800 => x"0d767971",
           801 => x"028c059f",
           802 => x"05335755",
           803 => x"53558372",
           804 => x"278a3874",
           805 => x"83065170",
           806 => x"802ea438",
           807 => x"ff125271",
           808 => x"ff2e9338",
           809 => x"73737081",
           810 => x"055534ff",
           811 => x"125271ff",
           812 => x"2e098106",
           813 => x"ef387481",
           814 => x"dec00c86",
           815 => x"3d0d0474",
           816 => x"74882b75",
           817 => x"07707190",
           818 => x"2b075154",
           819 => x"518f7227",
           820 => x"a5387271",
           821 => x"70840553",
           822 => x"0c727170",
           823 => x"8405530c",
           824 => x"72717084",
           825 => x"05530c72",
           826 => x"71708405",
           827 => x"530cf012",
           828 => x"52718f26",
           829 => x"dd388372",
           830 => x"27903872",
           831 => x"71708405",
           832 => x"530cfc12",
           833 => x"52718326",
           834 => x"f2387053",
           835 => x"ff8e39fb",
           836 => x"3d0d7779",
           837 => x"70720783",
           838 => x"06535452",
           839 => x"70933871",
           840 => x"73730854",
           841 => x"56547173",
           842 => x"082e80c6",
           843 => x"38737554",
           844 => x"52713370",
           845 => x"81ff0652",
           846 => x"5470802e",
           847 => x"9d387233",
           848 => x"5570752e",
           849 => x"09810695",
           850 => x"38811281",
           851 => x"14713370",
           852 => x"81ff0654",
           853 => x"56545270",
           854 => x"e5387233",
           855 => x"557381ff",
           856 => x"067581ff",
           857 => x"06717131",
           858 => x"81dec00c",
           859 => x"5252873d",
           860 => x"0d047109",
           861 => x"70f7fbfd",
           862 => x"ff140670",
           863 => x"f8848281",
           864 => x"80065151",
           865 => x"51709738",
           866 => x"84148416",
           867 => x"71085456",
           868 => x"54717508",
           869 => x"2edc3873",
           870 => x"755452ff",
           871 => x"9439800b",
           872 => x"81dec00c",
           873 => x"873d0d04",
           874 => x"fe3d0d80",
           875 => x"52835371",
           876 => x"882b5287",
           877 => x"863f81de",
           878 => x"c00881ff",
           879 => x"067207ff",
           880 => x"14545272",
           881 => x"8025e838",
           882 => x"7181dec0",
           883 => x"0c843d0d",
           884 => x"04fb3d0d",
           885 => x"77700870",
           886 => x"53535671",
           887 => x"802e80ca",
           888 => x"38713351",
           889 => x"70a02e09",
           890 => x"81068638",
           891 => x"811252f1",
           892 => x"39715384",
           893 => x"39811353",
           894 => x"80733370",
           895 => x"81ff0653",
           896 => x"555570a0",
           897 => x"2e833881",
           898 => x"5570802e",
           899 => x"843874e5",
           900 => x"387381ff",
           901 => x"065170a0",
           902 => x"2e098106",
           903 => x"88388073",
           904 => x"70810555",
           905 => x"3472760c",
           906 => x"71517081",
           907 => x"dec00c87",
           908 => x"3d0d04fc",
           909 => x"3d0d7653",
           910 => x"7208802e",
           911 => x"9138863d",
           912 => x"fc055272",
           913 => x"519bc33f",
           914 => x"81dec008",
           915 => x"85388053",
           916 => x"83397453",
           917 => x"7281dec0",
           918 => x"0c863d0d",
           919 => x"04fc3d0d",
           920 => x"76821133",
           921 => x"ff055253",
           922 => x"8152708b",
           923 => x"26819838",
           924 => x"831333ff",
           925 => x"05518252",
           926 => x"709e2681",
           927 => x"8a388413",
           928 => x"33518352",
           929 => x"70972680",
           930 => x"fe388513",
           931 => x"33518452",
           932 => x"70bb2680",
           933 => x"f2388613",
           934 => x"33518552",
           935 => x"70bb2680",
           936 => x"e6388813",
           937 => x"22558652",
           938 => x"7487e726",
           939 => x"80d9388a",
           940 => x"13225487",
           941 => x"527387e7",
           942 => x"2680cc38",
           943 => x"810b87c0",
           944 => x"989c0c72",
           945 => x"2287c098",
           946 => x"bc0c8213",
           947 => x"3387c098",
           948 => x"b80c8313",
           949 => x"3387c098",
           950 => x"b40c8413",
           951 => x"3387c098",
           952 => x"b00c8513",
           953 => x"3387c098",
           954 => x"ac0c8613",
           955 => x"3387c098",
           956 => x"a80c7487",
           957 => x"c098a40c",
           958 => x"7387c098",
           959 => x"a00c800b",
           960 => x"87c0989c",
           961 => x"0c805271",
           962 => x"81dec00c",
           963 => x"863d0d04",
           964 => x"f33d0d7f",
           965 => x"5b87c098",
           966 => x"9c5d817d",
           967 => x"0c87c098",
           968 => x"bc085e7d",
           969 => x"7b2387c0",
           970 => x"98b8085a",
           971 => x"79821c34",
           972 => x"87c098b4",
           973 => x"085a7983",
           974 => x"1c3487c0",
           975 => x"98b0085a",
           976 => x"79841c34",
           977 => x"87c098ac",
           978 => x"085a7985",
           979 => x"1c3487c0",
           980 => x"98a8085a",
           981 => x"79861c34",
           982 => x"87c098a4",
           983 => x"085c7b88",
           984 => x"1c2387c0",
           985 => x"98a0085a",
           986 => x"798a1c23",
           987 => x"807d0c79",
           988 => x"83ffff06",
           989 => x"597b83ff",
           990 => x"ff065886",
           991 => x"1b335785",
           992 => x"1b335684",
           993 => x"1b335583",
           994 => x"1b335482",
           995 => x"1b33537d",
           996 => x"83ffff06",
           997 => x"5281c6e4",
           998 => x"5195883f",
           999 => x"8f3d0d04",
          1000 => x"ff3d0d02",
          1001 => x"8f053370",
          1002 => x"30709f2a",
          1003 => x"51525270",
          1004 => x"0b0b81db",
          1005 => x"8834833d",
          1006 => x"0d04fb3d",
          1007 => x"0d770b0b",
          1008 => x"81db8833",
          1009 => x"7081ff06",
          1010 => x"57555687",
          1011 => x"c0948451",
          1012 => x"74802e86",
          1013 => x"3887c094",
          1014 => x"94517008",
          1015 => x"70962a70",
          1016 => x"81065354",
          1017 => x"5270802e",
          1018 => x"8c387191",
          1019 => x"2a708106",
          1020 => x"515170d7",
          1021 => x"38728132",
          1022 => x"70810651",
          1023 => x"5170802e",
          1024 => x"8d387193",
          1025 => x"2a708106",
          1026 => x"515170ff",
          1027 => x"be387381",
          1028 => x"ff065187",
          1029 => x"c0948052",
          1030 => x"70802e86",
          1031 => x"3887c094",
          1032 => x"90527572",
          1033 => x"0c7581de",
          1034 => x"c00c873d",
          1035 => x"0d04fb3d",
          1036 => x"0d029f05",
          1037 => x"330b0b81",
          1038 => x"db883370",
          1039 => x"81ff0657",
          1040 => x"555687c0",
          1041 => x"94845174",
          1042 => x"802e8638",
          1043 => x"87c09494",
          1044 => x"51700870",
          1045 => x"962a7081",
          1046 => x"06535452",
          1047 => x"70802e8c",
          1048 => x"3871912a",
          1049 => x"70810651",
          1050 => x"5170d738",
          1051 => x"72813270",
          1052 => x"81065151",
          1053 => x"70802e8d",
          1054 => x"3871932a",
          1055 => x"70810651",
          1056 => x"5170ffbe",
          1057 => x"387381ff",
          1058 => x"065187c0",
          1059 => x"94805270",
          1060 => x"802e8638",
          1061 => x"87c09490",
          1062 => x"5275720c",
          1063 => x"873d0d04",
          1064 => x"f93d0d79",
          1065 => x"54807433",
          1066 => x"7081ff06",
          1067 => x"53535770",
          1068 => x"772e80fe",
          1069 => x"387181ff",
          1070 => x"0681150b",
          1071 => x"0b81db88",
          1072 => x"337081ff",
          1073 => x"06595755",
          1074 => x"5887c094",
          1075 => x"84517580",
          1076 => x"2e863887",
          1077 => x"c0949451",
          1078 => x"70087096",
          1079 => x"2a708106",
          1080 => x"53545270",
          1081 => x"802e8c38",
          1082 => x"71912a70",
          1083 => x"81065151",
          1084 => x"70d73872",
          1085 => x"81327081",
          1086 => x"06515170",
          1087 => x"802e8d38",
          1088 => x"71932a70",
          1089 => x"81065151",
          1090 => x"70ffbe38",
          1091 => x"7481ff06",
          1092 => x"5187c094",
          1093 => x"80527080",
          1094 => x"2e863887",
          1095 => x"c0949052",
          1096 => x"77720c81",
          1097 => x"17743370",
          1098 => x"81ff0653",
          1099 => x"535770ff",
          1100 => x"84387681",
          1101 => x"dec00c89",
          1102 => x"3d0d04fe",
          1103 => x"3d0d0b0b",
          1104 => x"81db8833",
          1105 => x"7081ff06",
          1106 => x"545287c0",
          1107 => x"94845172",
          1108 => x"802e8638",
          1109 => x"87c09494",
          1110 => x"51700870",
          1111 => x"822a7081",
          1112 => x"06515151",
          1113 => x"70802ee2",
          1114 => x"387181ff",
          1115 => x"065187c0",
          1116 => x"94805270",
          1117 => x"802e8638",
          1118 => x"87c09490",
          1119 => x"52710870",
          1120 => x"81ff0681",
          1121 => x"dec00c51",
          1122 => x"843d0d04",
          1123 => x"fe3d0d0b",
          1124 => x"0b81db88",
          1125 => x"337081ff",
          1126 => x"06525387",
          1127 => x"c0948452",
          1128 => x"70802e86",
          1129 => x"3887c094",
          1130 => x"94527108",
          1131 => x"70822a70",
          1132 => x"81065151",
          1133 => x"51ff5270",
          1134 => x"802ea038",
          1135 => x"7281ff06",
          1136 => x"5187c094",
          1137 => x"80527080",
          1138 => x"2e863887",
          1139 => x"c0949052",
          1140 => x"71087098",
          1141 => x"2b70982c",
          1142 => x"51535171",
          1143 => x"81dec00c",
          1144 => x"843d0d04",
          1145 => x"ff3d0d87",
          1146 => x"c09e8008",
          1147 => x"709c2a8a",
          1148 => x"06515170",
          1149 => x"802e84b4",
          1150 => x"3887c09e",
          1151 => x"a40881db",
          1152 => x"8c0c87c0",
          1153 => x"9ea80881",
          1154 => x"db900c87",
          1155 => x"c09e9408",
          1156 => x"81db940c",
          1157 => x"87c09e98",
          1158 => x"0881db98",
          1159 => x"0c87c09e",
          1160 => x"9c0881db",
          1161 => x"9c0c87c0",
          1162 => x"9ea00881",
          1163 => x"dba00c87",
          1164 => x"c09eac08",
          1165 => x"81dba40c",
          1166 => x"87c09eb0",
          1167 => x"0881dba8",
          1168 => x"0c87c09e",
          1169 => x"b40881db",
          1170 => x"ac0c87c0",
          1171 => x"9eb80881",
          1172 => x"dbb00c87",
          1173 => x"c09ebc08",
          1174 => x"81dbb40c",
          1175 => x"87c09ec0",
          1176 => x"0881dbb8",
          1177 => x"0c87c09e",
          1178 => x"c40881db",
          1179 => x"bc0c87c0",
          1180 => x"9e800851",
          1181 => x"7081dbc0",
          1182 => x"2387c09e",
          1183 => x"840881db",
          1184 => x"c40c87c0",
          1185 => x"9e880881",
          1186 => x"dbc80c87",
          1187 => x"c09e8c08",
          1188 => x"81dbcc0c",
          1189 => x"810b81db",
          1190 => x"d034800b",
          1191 => x"87c09e90",
          1192 => x"08708480",
          1193 => x"0a065152",
          1194 => x"5270802e",
          1195 => x"83388152",
          1196 => x"7181dbd1",
          1197 => x"34800b87",
          1198 => x"c09e9008",
          1199 => x"7088800a",
          1200 => x"06515252",
          1201 => x"70802e83",
          1202 => x"38815271",
          1203 => x"81dbd234",
          1204 => x"800b87c0",
          1205 => x"9e900870",
          1206 => x"90800a06",
          1207 => x"51525270",
          1208 => x"802e8338",
          1209 => x"81527181",
          1210 => x"dbd33480",
          1211 => x"0b87c09e",
          1212 => x"90087088",
          1213 => x"80800651",
          1214 => x"52527080",
          1215 => x"2e833881",
          1216 => x"527181db",
          1217 => x"d434800b",
          1218 => x"87c09e90",
          1219 => x"0870a080",
          1220 => x"80065152",
          1221 => x"5270802e",
          1222 => x"83388152",
          1223 => x"7181dbd5",
          1224 => x"34800b87",
          1225 => x"c09e9008",
          1226 => x"70908080",
          1227 => x"06515252",
          1228 => x"70802e83",
          1229 => x"38815271",
          1230 => x"81dbd634",
          1231 => x"800b87c0",
          1232 => x"9e900870",
          1233 => x"84808006",
          1234 => x"51525270",
          1235 => x"802e8338",
          1236 => x"81527181",
          1237 => x"dbd73480",
          1238 => x"0b87c09e",
          1239 => x"90087082",
          1240 => x"80800651",
          1241 => x"52527080",
          1242 => x"2e833881",
          1243 => x"527181db",
          1244 => x"d834800b",
          1245 => x"87c09e90",
          1246 => x"08708180",
          1247 => x"80065152",
          1248 => x"5270802e",
          1249 => x"83388152",
          1250 => x"7181dbd9",
          1251 => x"34800b87",
          1252 => x"c09e9008",
          1253 => x"7080c080",
          1254 => x"06515252",
          1255 => x"70802e83",
          1256 => x"38815271",
          1257 => x"81dbda34",
          1258 => x"800b87c0",
          1259 => x"9e900870",
          1260 => x"a0800651",
          1261 => x"52527080",
          1262 => x"2e833881",
          1263 => x"527181db",
          1264 => x"db3487c0",
          1265 => x"9e900870",
          1266 => x"98800670",
          1267 => x"8a2a5151",
          1268 => x"517081db",
          1269 => x"dc34800b",
          1270 => x"87c09e90",
          1271 => x"08708480",
          1272 => x"06515252",
          1273 => x"70802e83",
          1274 => x"38815271",
          1275 => x"81dbdd34",
          1276 => x"87c09e90",
          1277 => x"087083f0",
          1278 => x"0670842a",
          1279 => x"51515170",
          1280 => x"81dbde34",
          1281 => x"800b87c0",
          1282 => x"9e900870",
          1283 => x"88065152",
          1284 => x"5270802e",
          1285 => x"83388152",
          1286 => x"7181dbdf",
          1287 => x"3487c09e",
          1288 => x"90087087",
          1289 => x"06515170",
          1290 => x"81dbe034",
          1291 => x"833d0d04",
          1292 => x"fb3d0d81",
          1293 => x"c6fc5186",
          1294 => x"863f81db",
          1295 => x"d0335473",
          1296 => x"802e8838",
          1297 => x"81c79051",
          1298 => x"85f53f81",
          1299 => x"c7a45185",
          1300 => x"ee3f81db",
          1301 => x"d2335473",
          1302 => x"802e9338",
          1303 => x"81dbac08",
          1304 => x"81dbb008",
          1305 => x"11545281",
          1306 => x"c7bc518b",
          1307 => x"b63f81db",
          1308 => x"d7335473",
          1309 => x"802e9338",
          1310 => x"81dba408",
          1311 => x"81dba808",
          1312 => x"11545281",
          1313 => x"c7d8518b",
          1314 => x"9a3f81db",
          1315 => x"d4335473",
          1316 => x"802e9338",
          1317 => x"81db8c08",
          1318 => x"81db9008",
          1319 => x"11545281",
          1320 => x"c7f4518a",
          1321 => x"fe3f81db",
          1322 => x"d5335473",
          1323 => x"802e9338",
          1324 => x"81db9408",
          1325 => x"81db9808",
          1326 => x"11545281",
          1327 => x"c890518a",
          1328 => x"e23f81db",
          1329 => x"d6335473",
          1330 => x"802e9338",
          1331 => x"81db9c08",
          1332 => x"81dba008",
          1333 => x"11545281",
          1334 => x"c8ac518a",
          1335 => x"c63f81db",
          1336 => x"db335473",
          1337 => x"802e8d38",
          1338 => x"81dbdc33",
          1339 => x"5281c8c8",
          1340 => x"518ab03f",
          1341 => x"81dbdf33",
          1342 => x"5473802e",
          1343 => x"8d3881db",
          1344 => x"e0335281",
          1345 => x"c8e8518a",
          1346 => x"9a3f81db",
          1347 => x"dd335473",
          1348 => x"802e8d38",
          1349 => x"81dbde33",
          1350 => x"5281c988",
          1351 => x"518a843f",
          1352 => x"81dbd133",
          1353 => x"5473802e",
          1354 => x"883881c9",
          1355 => x"a851848f",
          1356 => x"3f81dbd3",
          1357 => x"33547380",
          1358 => x"2e883881",
          1359 => x"c9bc5183",
          1360 => x"fe3f81db",
          1361 => x"d8335473",
          1362 => x"802e8838",
          1363 => x"81c9c851",
          1364 => x"83ed3f81",
          1365 => x"dbd93354",
          1366 => x"73802e88",
          1367 => x"3881c9d4",
          1368 => x"5183dc3f",
          1369 => x"81dbda33",
          1370 => x"5473802e",
          1371 => x"883881c9",
          1372 => x"e05183cb",
          1373 => x"3f81c9ec",
          1374 => x"5183c43f",
          1375 => x"81dbb408",
          1376 => x"5281c9f8",
          1377 => x"51899c3f",
          1378 => x"81dbb808",
          1379 => x"5281caa0",
          1380 => x"5189903f",
          1381 => x"81dbbc08",
          1382 => x"5281cac8",
          1383 => x"5189843f",
          1384 => x"81caf051",
          1385 => x"f5fa3f81",
          1386 => x"dbc02252",
          1387 => x"81caf851",
          1388 => x"88f13f81",
          1389 => x"dbc40856",
          1390 => x"bd84c052",
          1391 => x"7551e7b7",
          1392 => x"3f81dec0",
          1393 => x"08bd84c0",
          1394 => x"29767131",
          1395 => x"545481de",
          1396 => x"c0085281",
          1397 => x"cba05188",
          1398 => x"ca3f81db",
          1399 => x"d7335473",
          1400 => x"802ea838",
          1401 => x"81dbc808",
          1402 => x"56bd84c0",
          1403 => x"527551e7",
          1404 => x"863f81de",
          1405 => x"c008bd84",
          1406 => x"c0297671",
          1407 => x"31545481",
          1408 => x"dec00852",
          1409 => x"81cbcc51",
          1410 => x"88993f81",
          1411 => x"dbd23354",
          1412 => x"73802ea8",
          1413 => x"3881dbcc",
          1414 => x"0856bd84",
          1415 => x"c0527551",
          1416 => x"e6d53f81",
          1417 => x"dec008bd",
          1418 => x"84c02976",
          1419 => x"71315454",
          1420 => x"81dec008",
          1421 => x"5281cbf8",
          1422 => x"5187e83f",
          1423 => x"81d79c51",
          1424 => x"81fd3f87",
          1425 => x"3d0d04fe",
          1426 => x"3d0d0292",
          1427 => x"0533ff05",
          1428 => x"52718426",
          1429 => x"aa387184",
          1430 => x"2981c680",
          1431 => x"05527108",
          1432 => x"0481cca4",
          1433 => x"519d3981",
          1434 => x"ccac5197",
          1435 => x"3981ccb4",
          1436 => x"51913981",
          1437 => x"ccbc518b",
          1438 => x"3981ccc0",
          1439 => x"51853981",
          1440 => x"ccc851f4",
          1441 => x"9b3f843d",
          1442 => x"0d047188",
          1443 => x"800c0480",
          1444 => x"0b87c096",
          1445 => x"840c04ff",
          1446 => x"3d0d87c0",
          1447 => x"96847008",
          1448 => x"52528072",
          1449 => x"0c707407",
          1450 => x"7081dbe4",
          1451 => x"0c720c83",
          1452 => x"3d0d04ff",
          1453 => x"3d0d87c0",
          1454 => x"96847008",
          1455 => x"81dbe40c",
          1456 => x"5280720c",
          1457 => x"73097081",
          1458 => x"dbe40806",
          1459 => x"7081dbe4",
          1460 => x"0c730c51",
          1461 => x"833d0d04",
          1462 => x"81dbe408",
          1463 => x"87c09684",
          1464 => x"0c04fe3d",
          1465 => x"0d029305",
          1466 => x"3353728a",
          1467 => x"2e098106",
          1468 => x"85388d51",
          1469 => x"ed3f81de",
          1470 => x"d8085271",
          1471 => x"802e9038",
          1472 => x"72723481",
          1473 => x"ded80881",
          1474 => x"0581ded8",
          1475 => x"0c8f3981",
          1476 => x"ded00852",
          1477 => x"71802e85",
          1478 => x"38725171",
          1479 => x"2d843d0d",
          1480 => x"04fe3d0d",
          1481 => x"02970533",
          1482 => x"81ded008",
          1483 => x"7681ded0",
          1484 => x"0c5451ff",
          1485 => x"ad3f7281",
          1486 => x"ded00c84",
          1487 => x"3d0d04fd",
          1488 => x"3d0d7554",
          1489 => x"73337081",
          1490 => x"ff065353",
          1491 => x"71802e8e",
          1492 => x"387281ff",
          1493 => x"06518114",
          1494 => x"54ff873f",
          1495 => x"e739853d",
          1496 => x"0d04fc3d",
          1497 => x"0d7781de",
          1498 => x"d0087881",
          1499 => x"ded00c56",
          1500 => x"54733370",
          1501 => x"81ff0653",
          1502 => x"5371802e",
          1503 => x"8e387281",
          1504 => x"ff065181",
          1505 => x"1454feda",
          1506 => x"3fe73974",
          1507 => x"81ded00c",
          1508 => x"863d0d04",
          1509 => x"ec3d0d66",
          1510 => x"68595978",
          1511 => x"7081055a",
          1512 => x"33567580",
          1513 => x"2e84f838",
          1514 => x"75a52e09",
          1515 => x"810682de",
          1516 => x"3880707a",
          1517 => x"7081055c",
          1518 => x"33585b5b",
          1519 => x"75b02e09",
          1520 => x"81068538",
          1521 => x"815a8b39",
          1522 => x"75ad2e09",
          1523 => x"81068a38",
          1524 => x"825a7870",
          1525 => x"81055a33",
          1526 => x"5675aa2e",
          1527 => x"09810692",
          1528 => x"38778419",
          1529 => x"71087b70",
          1530 => x"81055d33",
          1531 => x"595d5953",
          1532 => x"9d39d016",
          1533 => x"53728926",
          1534 => x"95387a88",
          1535 => x"297b1005",
          1536 => x"7605d005",
          1537 => x"79708105",
          1538 => x"5b33575b",
          1539 => x"e5397580",
          1540 => x"ec327030",
          1541 => x"70720780",
          1542 => x"257880cc",
          1543 => x"32703070",
          1544 => x"72078025",
          1545 => x"73075354",
          1546 => x"58515553",
          1547 => x"73802e8c",
          1548 => x"38798407",
          1549 => x"79708105",
          1550 => x"5b33575a",
          1551 => x"75802e83",
          1552 => x"de387554",
          1553 => x"80e07627",
          1554 => x"8938e016",
          1555 => x"7081ff06",
          1556 => x"55537380",
          1557 => x"cf2e81aa",
          1558 => x"387380cf",
          1559 => x"24a23873",
          1560 => x"80c32e81",
          1561 => x"8e387380",
          1562 => x"c3248b38",
          1563 => x"7380c22e",
          1564 => x"818c3881",
          1565 => x"99397380",
          1566 => x"c42e818a",
          1567 => x"38818f39",
          1568 => x"7380d52e",
          1569 => x"81803873",
          1570 => x"80d5248a",
          1571 => x"387380d3",
          1572 => x"2e8e3880",
          1573 => x"f9397380",
          1574 => x"d82e80ee",
          1575 => x"3880ef39",
          1576 => x"77841971",
          1577 => x"08565953",
          1578 => x"80743354",
          1579 => x"5572752e",
          1580 => x"8d388115",
          1581 => x"70157033",
          1582 => x"51545572",
          1583 => x"f5387981",
          1584 => x"2a569039",
          1585 => x"74811656",
          1586 => x"53727b27",
          1587 => x"8f38a051",
          1588 => x"fc903f75",
          1589 => x"81065372",
          1590 => x"802ee938",
          1591 => x"7351fcdf",
          1592 => x"3f748116",
          1593 => x"5653727b",
          1594 => x"27fdb038",
          1595 => x"a051fbf2",
          1596 => x"3fef3977",
          1597 => x"84198312",
          1598 => x"33535953",
          1599 => x"9339825c",
          1600 => x"9539885c",
          1601 => x"91398a5c",
          1602 => x"8d39905c",
          1603 => x"89397551",
          1604 => x"fbd03ffd",
          1605 => x"86397982",
          1606 => x"2a708106",
          1607 => x"51537280",
          1608 => x"2e883877",
          1609 => x"84195953",
          1610 => x"86398418",
          1611 => x"78545872",
          1612 => x"087480c4",
          1613 => x"32703070",
          1614 => x"72078025",
          1615 => x"51555555",
          1616 => x"7480258d",
          1617 => x"3872802e",
          1618 => x"88387430",
          1619 => x"7a90075b",
          1620 => x"55800b8f",
          1621 => x"3d5e577b",
          1622 => x"527451e0",
          1623 => x"cd3f81de",
          1624 => x"c00881ff",
          1625 => x"067c5375",
          1626 => x"5254e08b",
          1627 => x"3f81dec0",
          1628 => x"08558974",
          1629 => x"279238a7",
          1630 => x"14537580",
          1631 => x"f82e8438",
          1632 => x"87145372",
          1633 => x"81ff0654",
          1634 => x"b0145372",
          1635 => x"7d708105",
          1636 => x"5f348117",
          1637 => x"75307077",
          1638 => x"079f2a51",
          1639 => x"5457769f",
          1640 => x"26853872",
          1641 => x"ffb13879",
          1642 => x"842a7081",
          1643 => x"06515372",
          1644 => x"802e8e38",
          1645 => x"963d7705",
          1646 => x"e00553ad",
          1647 => x"73348117",
          1648 => x"57767a81",
          1649 => x"065455b0",
          1650 => x"54728338",
          1651 => x"a0547981",
          1652 => x"2a708106",
          1653 => x"5456729f",
          1654 => x"38811755",
          1655 => x"767b2797",
          1656 => x"387351f9",
          1657 => x"fd3f7581",
          1658 => x"0653728b",
          1659 => x"38748116",
          1660 => x"56537a73",
          1661 => x"26eb3896",
          1662 => x"3d7705e0",
          1663 => x"0553ff17",
          1664 => x"ff147033",
          1665 => x"535457f9",
          1666 => x"d93f76f2",
          1667 => x"38748116",
          1668 => x"5653727b",
          1669 => x"27fb8438",
          1670 => x"a051f9c6",
          1671 => x"3fef3996",
          1672 => x"3d0d04fd",
          1673 => x"3d0d863d",
          1674 => x"70708405",
          1675 => x"52085552",
          1676 => x"7351fae0",
          1677 => x"3f853d0d",
          1678 => x"04fe3d0d",
          1679 => x"7481ded8",
          1680 => x"0c853d88",
          1681 => x"05527551",
          1682 => x"faca3f81",
          1683 => x"ded80853",
          1684 => x"80733480",
          1685 => x"0b81ded8",
          1686 => x"0c843d0d",
          1687 => x"04fd3d0d",
          1688 => x"81ded008",
          1689 => x"7681ded0",
          1690 => x"0c873d88",
          1691 => x"05537752",
          1692 => x"53faa13f",
          1693 => x"7281ded0",
          1694 => x"0c853d0d",
          1695 => x"04fb3d0d",
          1696 => x"777981de",
          1697 => x"d4087056",
          1698 => x"54575580",
          1699 => x"5471802e",
          1700 => x"80e03881",
          1701 => x"ded40852",
          1702 => x"712d81de",
          1703 => x"c00881ff",
          1704 => x"06537280",
          1705 => x"2e80cb38",
          1706 => x"728d2eb9",
          1707 => x"38728832",
          1708 => x"70307080",
          1709 => x"25515152",
          1710 => x"73802e8b",
          1711 => x"3871802e",
          1712 => x"8638ff14",
          1713 => x"5497399f",
          1714 => x"7325c838",
          1715 => x"ff165273",
          1716 => x"7225c038",
          1717 => x"74145272",
          1718 => x"72348114",
          1719 => x"547251f8",
          1720 => x"813fffaf",
          1721 => x"39731552",
          1722 => x"8072348a",
          1723 => x"51f7f33f",
          1724 => x"81537281",
          1725 => x"dec00c87",
          1726 => x"3d0d04fe",
          1727 => x"3d0d81de",
          1728 => x"d4087581",
          1729 => x"ded40c77",
          1730 => x"53765253",
          1731 => x"feef3f72",
          1732 => x"81ded40c",
          1733 => x"843d0d04",
          1734 => x"f83d0d7a",
          1735 => x"7c5a5680",
          1736 => x"707a0c58",
          1737 => x"75087033",
          1738 => x"555373a0",
          1739 => x"2e098106",
          1740 => x"87388113",
          1741 => x"760ced39",
          1742 => x"73ad2e09",
          1743 => x"81068e38",
          1744 => x"81760811",
          1745 => x"770c7608",
          1746 => x"70335654",
          1747 => x"5873b02e",
          1748 => x"09810680",
          1749 => x"c2387508",
          1750 => x"8105760c",
          1751 => x"75087033",
          1752 => x"55537380",
          1753 => x"e22e8b38",
          1754 => x"90577380",
          1755 => x"f82e8538",
          1756 => x"8f398257",
          1757 => x"8113760c",
          1758 => x"75087033",
          1759 => x"5553ac39",
          1760 => x"8155a074",
          1761 => x"2780fa38",
          1762 => x"d0145380",
          1763 => x"55885789",
          1764 => x"73279838",
          1765 => x"80eb39d0",
          1766 => x"14538055",
          1767 => x"72892680",
          1768 => x"e0388639",
          1769 => x"805580d9",
          1770 => x"398a5780",
          1771 => x"55a07427",
          1772 => x"80c23880",
          1773 => x"e0742789",
          1774 => x"38e01470",
          1775 => x"81ff0655",
          1776 => x"53d01470",
          1777 => x"81ff0655",
          1778 => x"53907427",
          1779 => x"8e38f914",
          1780 => x"7081ff06",
          1781 => x"55538974",
          1782 => x"27ca3873",
          1783 => x"7727c538",
          1784 => x"74772914",
          1785 => x"76088105",
          1786 => x"770c7608",
          1787 => x"70335654",
          1788 => x"55ffba39",
          1789 => x"77802e84",
          1790 => x"38743055",
          1791 => x"74790c81",
          1792 => x"557481de",
          1793 => x"c00c8a3d",
          1794 => x"0d04f83d",
          1795 => x"0d7a7c5a",
          1796 => x"5680707a",
          1797 => x"0c587508",
          1798 => x"70335553",
          1799 => x"73a02e09",
          1800 => x"81068738",
          1801 => x"8113760c",
          1802 => x"ed3973ad",
          1803 => x"2e098106",
          1804 => x"8e388176",
          1805 => x"0811770c",
          1806 => x"76087033",
          1807 => x"56545873",
          1808 => x"b02e0981",
          1809 => x"0680c238",
          1810 => x"75088105",
          1811 => x"760c7508",
          1812 => x"70335553",
          1813 => x"7380e22e",
          1814 => x"8b389057",
          1815 => x"7380f82e",
          1816 => x"85388f39",
          1817 => x"82578113",
          1818 => x"760c7508",
          1819 => x"70335553",
          1820 => x"ac398155",
          1821 => x"a0742780",
          1822 => x"fa38d014",
          1823 => x"53805588",
          1824 => x"57897327",
          1825 => x"983880eb",
          1826 => x"39d01453",
          1827 => x"80557289",
          1828 => x"2680e038",
          1829 => x"86398055",
          1830 => x"80d9398a",
          1831 => x"578055a0",
          1832 => x"742780c2",
          1833 => x"3880e074",
          1834 => x"278938e0",
          1835 => x"147081ff",
          1836 => x"065553d0",
          1837 => x"147081ff",
          1838 => x"06555390",
          1839 => x"74278e38",
          1840 => x"f9147081",
          1841 => x"ff065553",
          1842 => x"897427ca",
          1843 => x"38737727",
          1844 => x"c5387477",
          1845 => x"29147608",
          1846 => x"8105770c",
          1847 => x"76087033",
          1848 => x"565455ff",
          1849 => x"ba397780",
          1850 => x"2e843874",
          1851 => x"30557479",
          1852 => x"0c815574",
          1853 => x"81dec00c",
          1854 => x"8a3d0d04",
          1855 => x"ff3d0d02",
          1856 => x"8f053351",
          1857 => x"81527072",
          1858 => x"26873881",
          1859 => x"dbe81133",
          1860 => x"527181de",
          1861 => x"c00c833d",
          1862 => x"0d04fc3d",
          1863 => x"0d029b05",
          1864 => x"33028405",
          1865 => x"9f053356",
          1866 => x"53835172",
          1867 => x"812680e0",
          1868 => x"3872842b",
          1869 => x"87c0928c",
          1870 => x"11535188",
          1871 => x"5474802e",
          1872 => x"84388188",
          1873 => x"5473720c",
          1874 => x"87c0928c",
          1875 => x"11518171",
          1876 => x"0c850b87",
          1877 => x"c0988c0c",
          1878 => x"70527108",
          1879 => x"70820651",
          1880 => x"5170802e",
          1881 => x"8a3887c0",
          1882 => x"988c0851",
          1883 => x"70ec3871",
          1884 => x"08fc8080",
          1885 => x"06527192",
          1886 => x"3887c098",
          1887 => x"8c085170",
          1888 => x"802e8738",
          1889 => x"7181dbe8",
          1890 => x"143481db",
          1891 => x"e8133351",
          1892 => x"7081dec0",
          1893 => x"0c863d0d",
          1894 => x"04f33d0d",
          1895 => x"60626402",
          1896 => x"8c05bf05",
          1897 => x"33574058",
          1898 => x"5b837452",
          1899 => x"5afecd3f",
          1900 => x"81dec008",
          1901 => x"81067a54",
          1902 => x"527181be",
          1903 => x"38717275",
          1904 => x"842b87c0",
          1905 => x"92801187",
          1906 => x"c0928c12",
          1907 => x"87c09284",
          1908 => x"13415a40",
          1909 => x"575a5885",
          1910 => x"0b87c098",
          1911 => x"8c0c767d",
          1912 => x"0c84760c",
          1913 => x"75087085",
          1914 => x"2a708106",
          1915 => x"51535471",
          1916 => x"802e8e38",
          1917 => x"7b085271",
          1918 => x"7b708105",
          1919 => x"5d348119",
          1920 => x"598074a2",
          1921 => x"06535371",
          1922 => x"732e8338",
          1923 => x"81537883",
          1924 => x"ff268f38",
          1925 => x"72802e8a",
          1926 => x"3887c098",
          1927 => x"8c085271",
          1928 => x"c33887c0",
          1929 => x"988c0852",
          1930 => x"71802e87",
          1931 => x"38788480",
          1932 => x"2e993881",
          1933 => x"760c87c0",
          1934 => x"928c1553",
          1935 => x"72087082",
          1936 => x"06515271",
          1937 => x"f738ff1a",
          1938 => x"5a8d3984",
          1939 => x"80178119",
          1940 => x"7081ff06",
          1941 => x"5a535779",
          1942 => x"802e9038",
          1943 => x"73fc8080",
          1944 => x"06527187",
          1945 => x"387d7826",
          1946 => x"feed3873",
          1947 => x"fc808006",
          1948 => x"5271802e",
          1949 => x"83388152",
          1950 => x"71537281",
          1951 => x"dec00c8f",
          1952 => x"3d0d04f3",
          1953 => x"3d0d6062",
          1954 => x"64028c05",
          1955 => x"bf053357",
          1956 => x"40585b83",
          1957 => x"59807452",
          1958 => x"58fce13f",
          1959 => x"81dec008",
          1960 => x"81067954",
          1961 => x"5271782e",
          1962 => x"09810681",
          1963 => x"b1387774",
          1964 => x"842b87c0",
          1965 => x"92801187",
          1966 => x"c0928c12",
          1967 => x"87c09284",
          1968 => x"1340595f",
          1969 => x"565a850b",
          1970 => x"87c0988c",
          1971 => x"0c767d0c",
          1972 => x"82760c80",
          1973 => x"58750870",
          1974 => x"842a7081",
          1975 => x"06515354",
          1976 => x"71802e8c",
          1977 => x"387a7081",
          1978 => x"055c337c",
          1979 => x"0c811858",
          1980 => x"73812a70",
          1981 => x"81065152",
          1982 => x"71802e8a",
          1983 => x"3887c098",
          1984 => x"8c085271",
          1985 => x"d03887c0",
          1986 => x"988c0852",
          1987 => x"71802e87",
          1988 => x"38778480",
          1989 => x"2e993881",
          1990 => x"760c87c0",
          1991 => x"928c1553",
          1992 => x"72087082",
          1993 => x"06515271",
          1994 => x"f738ff19",
          1995 => x"598d3981",
          1996 => x"1a7081ff",
          1997 => x"06848019",
          1998 => x"595b5278",
          1999 => x"802e9038",
          2000 => x"73fc8080",
          2001 => x"06527187",
          2002 => x"387d7a26",
          2003 => x"fef83873",
          2004 => x"fc808006",
          2005 => x"5271802e",
          2006 => x"83388152",
          2007 => x"71537281",
          2008 => x"dec00c8f",
          2009 => x"3d0d04f6",
          2010 => x"3d0d7e02",
          2011 => x"8405b305",
          2012 => x"33028805",
          2013 => x"b7053371",
          2014 => x"54545657",
          2015 => x"fafe3f81",
          2016 => x"dec00881",
          2017 => x"06538354",
          2018 => x"7280fe38",
          2019 => x"850b87c0",
          2020 => x"988c0c81",
          2021 => x"5671762e",
          2022 => x"80dc3871",
          2023 => x"76249338",
          2024 => x"74842b87",
          2025 => x"c0928c11",
          2026 => x"54547180",
          2027 => x"2e8d3880",
          2028 => x"d4397183",
          2029 => x"2e80c638",
          2030 => x"80cb3972",
          2031 => x"0870812a",
          2032 => x"70810651",
          2033 => x"51527180",
          2034 => x"2e8a3887",
          2035 => x"c0988c08",
          2036 => x"5271e838",
          2037 => x"87c0988c",
          2038 => x"08527196",
          2039 => x"3881730c",
          2040 => x"87c0928c",
          2041 => x"14537208",
          2042 => x"70820651",
          2043 => x"5271f738",
          2044 => x"96398056",
          2045 => x"92398880",
          2046 => x"0a770c85",
          2047 => x"39818077",
          2048 => x"0c725683",
          2049 => x"39845675",
          2050 => x"547381de",
          2051 => x"c00c8c3d",
          2052 => x"0d04fe3d",
          2053 => x"0d748111",
          2054 => x"33713371",
          2055 => x"882b0781",
          2056 => x"dec00c53",
          2057 => x"51843d0d",
          2058 => x"04fd3d0d",
          2059 => x"75831133",
          2060 => x"82123371",
          2061 => x"902b7188",
          2062 => x"2b078114",
          2063 => x"33707207",
          2064 => x"882b7533",
          2065 => x"710781de",
          2066 => x"c00c5253",
          2067 => x"54565452",
          2068 => x"853d0d04",
          2069 => x"ff3d0d73",
          2070 => x"02840592",
          2071 => x"05225252",
          2072 => x"70727081",
          2073 => x"05543470",
          2074 => x"882a5170",
          2075 => x"7234833d",
          2076 => x"0d04ff3d",
          2077 => x"0d737552",
          2078 => x"52707270",
          2079 => x"81055434",
          2080 => x"70882a51",
          2081 => x"70727081",
          2082 => x"05543470",
          2083 => x"882a5170",
          2084 => x"72708105",
          2085 => x"54347088",
          2086 => x"2a517072",
          2087 => x"34833d0d",
          2088 => x"04fe3d0d",
          2089 => x"76757754",
          2090 => x"54517080",
          2091 => x"2e923871",
          2092 => x"70810553",
          2093 => x"33737081",
          2094 => x"055534ff",
          2095 => x"1151eb39",
          2096 => x"843d0d04",
          2097 => x"fe3d0d75",
          2098 => x"77765452",
          2099 => x"53727270",
          2100 => x"81055434",
          2101 => x"ff115170",
          2102 => x"f438843d",
          2103 => x"0d04fc3d",
          2104 => x"0d787779",
          2105 => x"56565374",
          2106 => x"70810556",
          2107 => x"33747081",
          2108 => x"05563371",
          2109 => x"7131ff16",
          2110 => x"56525252",
          2111 => x"72802e86",
          2112 => x"3871802e",
          2113 => x"e2387181",
          2114 => x"dec00c86",
          2115 => x"3d0d04fe",
          2116 => x"3d0d7476",
          2117 => x"54518939",
          2118 => x"71732e8a",
          2119 => x"38811151",
          2120 => x"70335271",
          2121 => x"f3387033",
          2122 => x"81dec00c",
          2123 => x"843d0d04",
          2124 => x"800b81de",
          2125 => x"c00c0480",
          2126 => x"0b81dec0",
          2127 => x"0c04f73d",
          2128 => x"0d7b5680",
          2129 => x"0b831733",
          2130 => x"565a747a",
          2131 => x"2e80d638",
          2132 => x"8154b016",
          2133 => x"0853b416",
          2134 => x"70538117",
          2135 => x"335259fa",
          2136 => x"a23f81de",
          2137 => x"c0087a2e",
          2138 => x"098106b7",
          2139 => x"3881dec0",
          2140 => x"08831734",
          2141 => x"b0160870",
          2142 => x"a4180831",
          2143 => x"9c180859",
          2144 => x"56587477",
          2145 => x"279f3882",
          2146 => x"16335574",
          2147 => x"822e0981",
          2148 => x"06933881",
          2149 => x"54761853",
          2150 => x"78528116",
          2151 => x"3351f9e3",
          2152 => x"3f833981",
          2153 => x"5a7981de",
          2154 => x"c00c8b3d",
          2155 => x"0d04fa3d",
          2156 => x"0d787a56",
          2157 => x"56805774",
          2158 => x"b017082e",
          2159 => x"af387551",
          2160 => x"fefc3f81",
          2161 => x"dec00857",
          2162 => x"81dec008",
          2163 => x"9f388154",
          2164 => x"7453b416",
          2165 => x"52811633",
          2166 => x"51f7be3f",
          2167 => x"81dec008",
          2168 => x"802e8538",
          2169 => x"ff558157",
          2170 => x"74b0170c",
          2171 => x"7681dec0",
          2172 => x"0c883d0d",
          2173 => x"04f83d0d",
          2174 => x"7a705257",
          2175 => x"fec03f81",
          2176 => x"dec00858",
          2177 => x"81dec008",
          2178 => x"81913876",
          2179 => x"33557483",
          2180 => x"2e098106",
          2181 => x"80f03884",
          2182 => x"17335978",
          2183 => x"812e0981",
          2184 => x"0680e338",
          2185 => x"84805381",
          2186 => x"dec00852",
          2187 => x"b4177052",
          2188 => x"56fd913f",
          2189 => x"82d4d552",
          2190 => x"84b21751",
          2191 => x"fc963f84",
          2192 => x"8b85a4d2",
          2193 => x"527551fc",
          2194 => x"a93f868a",
          2195 => x"85e4f252",
          2196 => x"84981751",
          2197 => x"fc9c3f90",
          2198 => x"17085284",
          2199 => x"9c1751fc",
          2200 => x"913f8c17",
          2201 => x"085284a0",
          2202 => x"1751fc86",
          2203 => x"3fa01708",
          2204 => x"810570b0",
          2205 => x"190c7955",
          2206 => x"53755281",
          2207 => x"173351f8",
          2208 => x"823f7784",
          2209 => x"18348053",
          2210 => x"80528117",
          2211 => x"3351f9d7",
          2212 => x"3f81dec0",
          2213 => x"08802e83",
          2214 => x"38815877",
          2215 => x"81dec00c",
          2216 => x"8a3d0d04",
          2217 => x"fb3d0d77",
          2218 => x"fe1a9812",
          2219 => x"08fe0555",
          2220 => x"56548056",
          2221 => x"7473278d",
          2222 => x"388a1422",
          2223 => x"757129ac",
          2224 => x"16080557",
          2225 => x"537581de",
          2226 => x"c00c873d",
          2227 => x"0d04f93d",
          2228 => x"0d7a7a70",
          2229 => x"08565457",
          2230 => x"81772781",
          2231 => x"df387698",
          2232 => x"15082781",
          2233 => x"d738ff74",
          2234 => x"33545872",
          2235 => x"822e80f5",
          2236 => x"38728224",
          2237 => x"89387281",
          2238 => x"2e8d3881",
          2239 => x"bf397283",
          2240 => x"2e818e38",
          2241 => x"81b63976",
          2242 => x"812a1770",
          2243 => x"892aa416",
          2244 => x"08055374",
          2245 => x"5255fd96",
          2246 => x"3f81dec0",
          2247 => x"08819f38",
          2248 => x"7483ff06",
          2249 => x"14b41133",
          2250 => x"81177089",
          2251 => x"2aa41808",
          2252 => x"05557654",
          2253 => x"575753fc",
          2254 => x"f53f81de",
          2255 => x"c00880fe",
          2256 => x"387483ff",
          2257 => x"0614b411",
          2258 => x"3370882b",
          2259 => x"78077981",
          2260 => x"0671842a",
          2261 => x"5c525851",
          2262 => x"537280e2",
          2263 => x"38759fff",
          2264 => x"065880da",
          2265 => x"3976882a",
          2266 => x"a4150805",
          2267 => x"527351fc",
          2268 => x"bd3f81de",
          2269 => x"c00880c6",
          2270 => x"38761083",
          2271 => x"fe067405",
          2272 => x"b40551f9",
          2273 => x"8d3f81de",
          2274 => x"c00883ff",
          2275 => x"ff0658ae",
          2276 => x"3976872a",
          2277 => x"a4150805",
          2278 => x"527351fc",
          2279 => x"913f81de",
          2280 => x"c0089b38",
          2281 => x"76822b83",
          2282 => x"fc067405",
          2283 => x"b40551f8",
          2284 => x"f83f81de",
          2285 => x"c008f00a",
          2286 => x"06588339",
          2287 => x"81587781",
          2288 => x"dec00c89",
          2289 => x"3d0d04f8",
          2290 => x"3d0d7a7c",
          2291 => x"7e5a5856",
          2292 => x"82598177",
          2293 => x"27829e38",
          2294 => x"76981708",
          2295 => x"27829638",
          2296 => x"75335372",
          2297 => x"792e819d",
          2298 => x"38727924",
          2299 => x"89387281",
          2300 => x"2e8d3882",
          2301 => x"80397283",
          2302 => x"2e81b838",
          2303 => x"81f73976",
          2304 => x"812a1770",
          2305 => x"892aa418",
          2306 => x"08055376",
          2307 => x"5255fb9e",
          2308 => x"3f81dec0",
          2309 => x"085981de",
          2310 => x"c00881d9",
          2311 => x"387483ff",
          2312 => x"0616b405",
          2313 => x"81167881",
          2314 => x"06595654",
          2315 => x"77537680",
          2316 => x"2e8f3877",
          2317 => x"842b9ff0",
          2318 => x"0674338f",
          2319 => x"06710751",
          2320 => x"53727434",
          2321 => x"810b8317",
          2322 => x"3474892a",
          2323 => x"a4170805",
          2324 => x"527551fa",
          2325 => x"d93f81de",
          2326 => x"c0085981",
          2327 => x"dec00881",
          2328 => x"94387483",
          2329 => x"ff0616b4",
          2330 => x"0578842a",
          2331 => x"5454768f",
          2332 => x"3877882a",
          2333 => x"743381f0",
          2334 => x"06718f06",
          2335 => x"07515372",
          2336 => x"743480ec",
          2337 => x"3976882a",
          2338 => x"a4170805",
          2339 => x"527551fa",
          2340 => x"9d3f81de",
          2341 => x"c0085981",
          2342 => x"dec00880",
          2343 => x"d8387783",
          2344 => x"ffff0652",
          2345 => x"761083fe",
          2346 => x"067605b4",
          2347 => x"0551f7a4",
          2348 => x"3fbe3976",
          2349 => x"872aa417",
          2350 => x"08055275",
          2351 => x"51f9ef3f",
          2352 => x"81dec008",
          2353 => x"5981dec0",
          2354 => x"08ab3877",
          2355 => x"f00a0677",
          2356 => x"822b83fc",
          2357 => x"067018b4",
          2358 => x"05705451",
          2359 => x"5454f6c9",
          2360 => x"3f81dec0",
          2361 => x"088f0a06",
          2362 => x"74075272",
          2363 => x"51f7833f",
          2364 => x"810b8317",
          2365 => x"347881de",
          2366 => x"c00c8a3d",
          2367 => x"0d04f83d",
          2368 => x"0d7a7c7e",
          2369 => x"72085956",
          2370 => x"56598175",
          2371 => x"27a43874",
          2372 => x"98170827",
          2373 => x"9d387380",
          2374 => x"2eaa38ff",
          2375 => x"53735275",
          2376 => x"51fda43f",
          2377 => x"81dec008",
          2378 => x"5481dec0",
          2379 => x"0880f238",
          2380 => x"93398254",
          2381 => x"80eb3981",
          2382 => x"5480e639",
          2383 => x"81dec008",
          2384 => x"5480de39",
          2385 => x"74527851",
          2386 => x"fb843f81",
          2387 => x"dec00858",
          2388 => x"81dec008",
          2389 => x"802e80c7",
          2390 => x"3881dec0",
          2391 => x"08812ed2",
          2392 => x"3881dec0",
          2393 => x"08ff2ecf",
          2394 => x"38805374",
          2395 => x"527551fc",
          2396 => x"d63f81de",
          2397 => x"c008c538",
          2398 => x"981608fe",
          2399 => x"11901808",
          2400 => x"57555774",
          2401 => x"74279038",
          2402 => x"81159017",
          2403 => x"0c841633",
          2404 => x"81075473",
          2405 => x"84173477",
          2406 => x"55767826",
          2407 => x"ffa63880",
          2408 => x"547381de",
          2409 => x"c00c8a3d",
          2410 => x"0d04f63d",
          2411 => x"0d7c7e71",
          2412 => x"08595b5b",
          2413 => x"7995388c",
          2414 => x"17085877",
          2415 => x"802e8838",
          2416 => x"98170878",
          2417 => x"26b23881",
          2418 => x"58ae3979",
          2419 => x"527a51f9",
          2420 => x"fd3f8155",
          2421 => x"7481dec0",
          2422 => x"082782e0",
          2423 => x"3881dec0",
          2424 => x"085581de",
          2425 => x"c008ff2e",
          2426 => x"82d23898",
          2427 => x"170881de",
          2428 => x"c0082682",
          2429 => x"c7387958",
          2430 => x"90170870",
          2431 => x"56547380",
          2432 => x"2e82b938",
          2433 => x"777a2e09",
          2434 => x"810680e2",
          2435 => x"38811a56",
          2436 => x"98170876",
          2437 => x"26833882",
          2438 => x"5675527a",
          2439 => x"51f9af3f",
          2440 => x"805981de",
          2441 => x"c008812e",
          2442 => x"09810686",
          2443 => x"3881dec0",
          2444 => x"085981de",
          2445 => x"c0080970",
          2446 => x"30707207",
          2447 => x"8025707c",
          2448 => x"0781dec0",
          2449 => x"08545151",
          2450 => x"55557381",
          2451 => x"ef3881de",
          2452 => x"c008802e",
          2453 => x"95388c17",
          2454 => x"08548174",
          2455 => x"27903873",
          2456 => x"98180827",
          2457 => x"89387358",
          2458 => x"85397580",
          2459 => x"db387756",
          2460 => x"81165698",
          2461 => x"17087626",
          2462 => x"89388256",
          2463 => x"75782681",
          2464 => x"ac387552",
          2465 => x"7a51f8c6",
          2466 => x"3f81dec0",
          2467 => x"08802eb8",
          2468 => x"38805981",
          2469 => x"dec00881",
          2470 => x"2e098106",
          2471 => x"863881de",
          2472 => x"c0085981",
          2473 => x"dec00809",
          2474 => x"70307072",
          2475 => x"07802570",
          2476 => x"7c075151",
          2477 => x"55557380",
          2478 => x"f8387578",
          2479 => x"2e098106",
          2480 => x"ffae3873",
          2481 => x"5580f539",
          2482 => x"ff537552",
          2483 => x"7651f9f7",
          2484 => x"3f81dec0",
          2485 => x"0881dec0",
          2486 => x"08307081",
          2487 => x"dec00807",
          2488 => x"80255155",
          2489 => x"5579802e",
          2490 => x"94387380",
          2491 => x"2e8f3875",
          2492 => x"53795276",
          2493 => x"51f9d03f",
          2494 => x"81dec008",
          2495 => x"5574a538",
          2496 => x"758c180c",
          2497 => x"981708fe",
          2498 => x"05901808",
          2499 => x"56547474",
          2500 => x"268638ff",
          2501 => x"1590180c",
          2502 => x"84173381",
          2503 => x"07547384",
          2504 => x"18349739",
          2505 => x"ff567481",
          2506 => x"2e90388c",
          2507 => x"3980558c",
          2508 => x"3981dec0",
          2509 => x"08558539",
          2510 => x"81567555",
          2511 => x"7481dec0",
          2512 => x"0c8c3d0d",
          2513 => x"04f83d0d",
          2514 => x"7a705255",
          2515 => x"f3f03f81",
          2516 => x"dec00858",
          2517 => x"815681de",
          2518 => x"c00880d8",
          2519 => x"387b5274",
          2520 => x"51f6c13f",
          2521 => x"81dec008",
          2522 => x"81dec008",
          2523 => x"b0170c59",
          2524 => x"84805377",
          2525 => x"52b41570",
          2526 => x"5257f2c8",
          2527 => x"3f775684",
          2528 => x"39811656",
          2529 => x"8a152258",
          2530 => x"75782797",
          2531 => x"38815475",
          2532 => x"19537652",
          2533 => x"81153351",
          2534 => x"ede93f81",
          2535 => x"dec00880",
          2536 => x"2edf388a",
          2537 => x"15227632",
          2538 => x"70307072",
          2539 => x"07709f2a",
          2540 => x"53515656",
          2541 => x"7581dec0",
          2542 => x"0c8a3d0d",
          2543 => x"04f83d0d",
          2544 => x"7a7c7108",
          2545 => x"58565774",
          2546 => x"f0800a26",
          2547 => x"80f13874",
          2548 => x"9f065372",
          2549 => x"80e93874",
          2550 => x"90180c88",
          2551 => x"17085473",
          2552 => x"aa387533",
          2553 => x"53827327",
          2554 => x"8838a816",
          2555 => x"0854739b",
          2556 => x"3874852a",
          2557 => x"53820b88",
          2558 => x"17225a58",
          2559 => x"72792780",
          2560 => x"fe38a816",
          2561 => x"0898180c",
          2562 => x"80cd398a",
          2563 => x"16227089",
          2564 => x"2b545872",
          2565 => x"7526b238",
          2566 => x"73527651",
          2567 => x"f5b03f81",
          2568 => x"dec00854",
          2569 => x"81dec008",
          2570 => x"ff2ebd38",
          2571 => x"810b81de",
          2572 => x"c008278b",
          2573 => x"38981608",
          2574 => x"81dec008",
          2575 => x"26853882",
          2576 => x"58bd3974",
          2577 => x"733155cb",
          2578 => x"39735275",
          2579 => x"51f4d53f",
          2580 => x"81dec008",
          2581 => x"98180c73",
          2582 => x"94180c98",
          2583 => x"17085382",
          2584 => x"5872802e",
          2585 => x"9a388539",
          2586 => x"81589439",
          2587 => x"74892a13",
          2588 => x"98180c74",
          2589 => x"83ff0616",
          2590 => x"b4059c18",
          2591 => x"0c805877",
          2592 => x"81dec00c",
          2593 => x"8a3d0d04",
          2594 => x"f83d0d7a",
          2595 => x"70089012",
          2596 => x"08a00559",
          2597 => x"5754f080",
          2598 => x"0a772786",
          2599 => x"38800b98",
          2600 => x"150c9814",
          2601 => x"08538455",
          2602 => x"72802e81",
          2603 => x"cb387683",
          2604 => x"ff065877",
          2605 => x"81b53881",
          2606 => x"1398150c",
          2607 => x"94140855",
          2608 => x"74923876",
          2609 => x"852a8817",
          2610 => x"22565374",
          2611 => x"7326819b",
          2612 => x"3880c039",
          2613 => x"8a1622ff",
          2614 => x"0577892a",
          2615 => x"06537281",
          2616 => x"8a387452",
          2617 => x"7351f3e6",
          2618 => x"3f81dec0",
          2619 => x"08538255",
          2620 => x"810b81de",
          2621 => x"c0082780",
          2622 => x"ff388155",
          2623 => x"81dec008",
          2624 => x"ff2e80f4",
          2625 => x"38981608",
          2626 => x"81dec008",
          2627 => x"2680ca38",
          2628 => x"7b8a3877",
          2629 => x"98150c84",
          2630 => x"5580dd39",
          2631 => x"94140852",
          2632 => x"7351f986",
          2633 => x"3f81dec0",
          2634 => x"08538755",
          2635 => x"81dec008",
          2636 => x"802e80c4",
          2637 => x"38825581",
          2638 => x"dec00881",
          2639 => x"2eba3881",
          2640 => x"5581dec0",
          2641 => x"08ff2eb0",
          2642 => x"3881dec0",
          2643 => x"08527551",
          2644 => x"fbf33f81",
          2645 => x"dec008a0",
          2646 => x"38729415",
          2647 => x"0c725275",
          2648 => x"51f2c13f",
          2649 => x"81dec008",
          2650 => x"98150c76",
          2651 => x"90150c77",
          2652 => x"16b4059c",
          2653 => x"150c8055",
          2654 => x"7481dec0",
          2655 => x"0c8a3d0d",
          2656 => x"04f73d0d",
          2657 => x"7b7d7108",
          2658 => x"5b5b5780",
          2659 => x"527651fc",
          2660 => x"ac3f81de",
          2661 => x"c0085481",
          2662 => x"dec00880",
          2663 => x"ec3881de",
          2664 => x"c0085698",
          2665 => x"17085278",
          2666 => x"51f0833f",
          2667 => x"81dec008",
          2668 => x"5481dec0",
          2669 => x"0880d238",
          2670 => x"81dec008",
          2671 => x"9c180870",
          2672 => x"33515458",
          2673 => x"7281e52e",
          2674 => x"09810683",
          2675 => x"38815881",
          2676 => x"dec00855",
          2677 => x"72833881",
          2678 => x"55777507",
          2679 => x"5372802e",
          2680 => x"8e388116",
          2681 => x"56757a2e",
          2682 => x"09810688",
          2683 => x"38a53981",
          2684 => x"dec00856",
          2685 => x"81527651",
          2686 => x"fd8e3f81",
          2687 => x"dec00854",
          2688 => x"81dec008",
          2689 => x"802eff9b",
          2690 => x"3873842e",
          2691 => x"09810683",
          2692 => x"38875473",
          2693 => x"81dec00c",
          2694 => x"8b3d0d04",
          2695 => x"fd3d0d76",
          2696 => x"9a115254",
          2697 => x"ebec3f81",
          2698 => x"dec00883",
          2699 => x"ffff0676",
          2700 => x"70335153",
          2701 => x"5371832e",
          2702 => x"09810690",
          2703 => x"38941451",
          2704 => x"ebd03f81",
          2705 => x"dec00890",
          2706 => x"2b730753",
          2707 => x"7281dec0",
          2708 => x"0c853d0d",
          2709 => x"04fc3d0d",
          2710 => x"77797083",
          2711 => x"ffff0654",
          2712 => x"9a125355",
          2713 => x"55ebed3f",
          2714 => x"76703351",
          2715 => x"5372832e",
          2716 => x"0981068b",
          2717 => x"3873902a",
          2718 => x"52941551",
          2719 => x"ebd63f86",
          2720 => x"3d0d04f7",
          2721 => x"3d0d7b7d",
          2722 => x"5b558475",
          2723 => x"085a5898",
          2724 => x"1508802e",
          2725 => x"818a3898",
          2726 => x"15085278",
          2727 => x"51ee8f3f",
          2728 => x"81dec008",
          2729 => x"5881dec0",
          2730 => x"0880f538",
          2731 => x"9c150870",
          2732 => x"33555373",
          2733 => x"86388458",
          2734 => x"80e6398b",
          2735 => x"133370bf",
          2736 => x"067081ff",
          2737 => x"06585153",
          2738 => x"72861634",
          2739 => x"81dec008",
          2740 => x"537381e5",
          2741 => x"2e833881",
          2742 => x"5373ae2e",
          2743 => x"a9388170",
          2744 => x"74065457",
          2745 => x"72802e9e",
          2746 => x"38758f2e",
          2747 => x"993881de",
          2748 => x"c00876df",
          2749 => x"06545472",
          2750 => x"882e0981",
          2751 => x"06833876",
          2752 => x"54737a2e",
          2753 => x"a0388052",
          2754 => x"7451fafc",
          2755 => x"3f81dec0",
          2756 => x"085881de",
          2757 => x"c0088938",
          2758 => x"981508fe",
          2759 => x"fa388639",
          2760 => x"800b9816",
          2761 => x"0c7781de",
          2762 => x"c00c8b3d",
          2763 => x"0d04fb3d",
          2764 => x"0d777008",
          2765 => x"57548152",
          2766 => x"7351fcc5",
          2767 => x"3f81dec0",
          2768 => x"085581de",
          2769 => x"c008b438",
          2770 => x"98140852",
          2771 => x"7551ecde",
          2772 => x"3f81dec0",
          2773 => x"085581de",
          2774 => x"c008a038",
          2775 => x"a05381de",
          2776 => x"c008529c",
          2777 => x"140851ea",
          2778 => x"db3f8b53",
          2779 => x"a014529c",
          2780 => x"140851ea",
          2781 => x"ac3f810b",
          2782 => x"83173474",
          2783 => x"81dec00c",
          2784 => x"873d0d04",
          2785 => x"fd3d0d75",
          2786 => x"70089812",
          2787 => x"08547053",
          2788 => x"5553ec9a",
          2789 => x"3f81dec0",
          2790 => x"088d389c",
          2791 => x"130853e5",
          2792 => x"7334810b",
          2793 => x"83153485",
          2794 => x"3d0d04fa",
          2795 => x"3d0d787a",
          2796 => x"5757800b",
          2797 => x"89173498",
          2798 => x"1708802e",
          2799 => x"81823880",
          2800 => x"70891855",
          2801 => x"55559c17",
          2802 => x"08147033",
          2803 => x"81165651",
          2804 => x"5271a02e",
          2805 => x"a8387185",
          2806 => x"2e098106",
          2807 => x"843881e5",
          2808 => x"5273892e",
          2809 => x"0981068b",
          2810 => x"38ae7370",
          2811 => x"81055534",
          2812 => x"81155571",
          2813 => x"73708105",
          2814 => x"55348115",
          2815 => x"558a7427",
          2816 => x"c5387515",
          2817 => x"88055280",
          2818 => x"0b811334",
          2819 => x"9c170852",
          2820 => x"8b123388",
          2821 => x"17349c17",
          2822 => x"089c1152",
          2823 => x"52e88a3f",
          2824 => x"81dec008",
          2825 => x"760c9612",
          2826 => x"51e7e73f",
          2827 => x"81dec008",
          2828 => x"86172398",
          2829 => x"1251e7da",
          2830 => x"3f81dec0",
          2831 => x"08841723",
          2832 => x"883d0d04",
          2833 => x"f33d0d7f",
          2834 => x"70085e5b",
          2835 => x"80617033",
          2836 => x"51555573",
          2837 => x"af2e8338",
          2838 => x"81557380",
          2839 => x"dc2e9138",
          2840 => x"74802e8c",
          2841 => x"38941d08",
          2842 => x"881c0caa",
          2843 => x"39811541",
          2844 => x"80617033",
          2845 => x"56565673",
          2846 => x"af2e0981",
          2847 => x"06833881",
          2848 => x"567380dc",
          2849 => x"32703070",
          2850 => x"80257807",
          2851 => x"51515473",
          2852 => x"dc387388",
          2853 => x"1c0c6070",
          2854 => x"33515473",
          2855 => x"9f269638",
          2856 => x"ff800bab",
          2857 => x"1c348052",
          2858 => x"7a51f691",
          2859 => x"3f81dec0",
          2860 => x"08558598",
          2861 => x"39913d61",
          2862 => x"a01d5c5a",
          2863 => x"5e8b53a0",
          2864 => x"527951e7",
          2865 => x"ff3f8070",
          2866 => x"59578879",
          2867 => x"33555c73",
          2868 => x"ae2e0981",
          2869 => x"0680d438",
          2870 => x"78187033",
          2871 => x"811a71ae",
          2872 => x"32703070",
          2873 => x"9f2a7382",
          2874 => x"26075151",
          2875 => x"535a5754",
          2876 => x"738c3879",
          2877 => x"17547574",
          2878 => x"34811757",
          2879 => x"db3975af",
          2880 => x"32703070",
          2881 => x"9f2a5151",
          2882 => x"547580dc",
          2883 => x"2e8c3873",
          2884 => x"802e8738",
          2885 => x"75a02682",
          2886 => x"bd387719",
          2887 => x"7e0ca454",
          2888 => x"a0762782",
          2889 => x"bd38a054",
          2890 => x"82b83978",
          2891 => x"18703381",
          2892 => x"1a5a5754",
          2893 => x"a0762781",
          2894 => x"fc3875af",
          2895 => x"32703077",
          2896 => x"80dc3270",
          2897 => x"30728025",
          2898 => x"71802507",
          2899 => x"51515651",
          2900 => x"5573802e",
          2901 => x"ac388439",
          2902 => x"81185880",
          2903 => x"781a7033",
          2904 => x"51555573",
          2905 => x"af2e0981",
          2906 => x"06833881",
          2907 => x"557380dc",
          2908 => x"32703070",
          2909 => x"80257707",
          2910 => x"51515473",
          2911 => x"db3881b5",
          2912 => x"3975ae2e",
          2913 => x"09810683",
          2914 => x"38815476",
          2915 => x"7c277407",
          2916 => x"5473802e",
          2917 => x"a2387b8b",
          2918 => x"32703077",
          2919 => x"ae327030",
          2920 => x"72802571",
          2921 => x"9f2a0753",
          2922 => x"51565155",
          2923 => x"7481a738",
          2924 => x"88578b5c",
          2925 => x"fef53975",
          2926 => x"982b5473",
          2927 => x"80258c38",
          2928 => x"7580ff06",
          2929 => x"81cdb411",
          2930 => x"33575475",
          2931 => x"51e6e13f",
          2932 => x"81dec008",
          2933 => x"802eb238",
          2934 => x"78187033",
          2935 => x"811a7154",
          2936 => x"5a5654e6",
          2937 => x"d23f81de",
          2938 => x"c008802e",
          2939 => x"80e838ff",
          2940 => x"1c547674",
          2941 => x"2780df38",
          2942 => x"79175475",
          2943 => x"74348117",
          2944 => x"7a115557",
          2945 => x"747434a7",
          2946 => x"39755281",
          2947 => x"ccd451e5",
          2948 => x"fe3f81de",
          2949 => x"c008bf38",
          2950 => x"ff9f1654",
          2951 => x"73992689",
          2952 => x"38e01670",
          2953 => x"81ff0657",
          2954 => x"54791754",
          2955 => x"75743481",
          2956 => x"1757fdf7",
          2957 => x"3977197e",
          2958 => x"0c76802e",
          2959 => x"99387933",
          2960 => x"547381e5",
          2961 => x"2e098106",
          2962 => x"8438857a",
          2963 => x"348454a0",
          2964 => x"76278f38",
          2965 => x"8b398655",
          2966 => x"81f23984",
          2967 => x"5680f339",
          2968 => x"8054738b",
          2969 => x"1b34807b",
          2970 => x"0858527a",
          2971 => x"51f2ce3f",
          2972 => x"81dec008",
          2973 => x"5681dec0",
          2974 => x"0880d738",
          2975 => x"981b0852",
          2976 => x"7651e6aa",
          2977 => x"3f81dec0",
          2978 => x"085681de",
          2979 => x"c00880c2",
          2980 => x"389c1b08",
          2981 => x"70335555",
          2982 => x"73802eff",
          2983 => x"be388b15",
          2984 => x"33bf0654",
          2985 => x"73861c34",
          2986 => x"8b153370",
          2987 => x"832a7081",
          2988 => x"06515558",
          2989 => x"7392388b",
          2990 => x"53795274",
          2991 => x"51e49f3f",
          2992 => x"81dec008",
          2993 => x"802e8b38",
          2994 => x"75527a51",
          2995 => x"f3ba3fff",
          2996 => x"9f3975ab",
          2997 => x"1c335755",
          2998 => x"74802ebb",
          2999 => x"3874842e",
          3000 => x"09810680",
          3001 => x"e7387585",
          3002 => x"2a708106",
          3003 => x"77822a58",
          3004 => x"51547380",
          3005 => x"2e963875",
          3006 => x"81065473",
          3007 => x"802efbb5",
          3008 => x"38ff800b",
          3009 => x"ab1c3480",
          3010 => x"5580c139",
          3011 => x"75810654",
          3012 => x"73ba3885",
          3013 => x"55b63975",
          3014 => x"822a7081",
          3015 => x"06515473",
          3016 => x"ab38861b",
          3017 => x"3370842a",
          3018 => x"70810651",
          3019 => x"55557380",
          3020 => x"2ee13890",
          3021 => x"1b0883ff",
          3022 => x"061db405",
          3023 => x"527c51f5",
          3024 => x"db3f81de",
          3025 => x"c008881c",
          3026 => x"0cfaea39",
          3027 => x"7481dec0",
          3028 => x"0c8f3d0d",
          3029 => x"04f63d0d",
          3030 => x"7c5bff7b",
          3031 => x"08707173",
          3032 => x"55595c55",
          3033 => x"5973802e",
          3034 => x"81c63875",
          3035 => x"70810557",
          3036 => x"3370a026",
          3037 => x"525271ba",
          3038 => x"2e8d3870",
          3039 => x"ee3871ba",
          3040 => x"2e098106",
          3041 => x"81a53873",
          3042 => x"33d01170",
          3043 => x"81ff0651",
          3044 => x"52537089",
          3045 => x"26913882",
          3046 => x"147381ff",
          3047 => x"06d00556",
          3048 => x"5271762e",
          3049 => x"80f73880",
          3050 => x"0b81cda4",
          3051 => x"59557708",
          3052 => x"7a555776",
          3053 => x"70810558",
          3054 => x"33747081",
          3055 => x"055633ff",
          3056 => x"9f125353",
          3057 => x"53709926",
          3058 => x"8938e013",
          3059 => x"7081ff06",
          3060 => x"5451ff9f",
          3061 => x"12517099",
          3062 => x"268938e0",
          3063 => x"127081ff",
          3064 => x"06535172",
          3065 => x"30709f2a",
          3066 => x"51517272",
          3067 => x"2e098106",
          3068 => x"853870ff",
          3069 => x"be387230",
          3070 => x"74773270",
          3071 => x"30707207",
          3072 => x"9f2a739f",
          3073 => x"2a075354",
          3074 => x"54517080",
          3075 => x"2e8f3881",
          3076 => x"15841959",
          3077 => x"55837525",
          3078 => x"ff94388b",
          3079 => x"39748324",
          3080 => x"86387476",
          3081 => x"7c0c5978",
          3082 => x"51863981",
          3083 => x"def03351",
          3084 => x"7081dec0",
          3085 => x"0c8c3d0d",
          3086 => x"04fa3d0d",
          3087 => x"7856800b",
          3088 => x"831734ff",
          3089 => x"0bb0170c",
          3090 => x"79527551",
          3091 => x"e2e03f84",
          3092 => x"5581dec0",
          3093 => x"08818038",
          3094 => x"84b21651",
          3095 => x"dfb43f81",
          3096 => x"dec00883",
          3097 => x"ffff0654",
          3098 => x"83557382",
          3099 => x"d4d52e09",
          3100 => x"810680e3",
          3101 => x"38800bb4",
          3102 => x"17335657",
          3103 => x"7481e92e",
          3104 => x"09810683",
          3105 => x"38815774",
          3106 => x"81eb3270",
          3107 => x"30708025",
          3108 => x"79075151",
          3109 => x"54738a38",
          3110 => x"7481e82e",
          3111 => x"098106b5",
          3112 => x"38835381",
          3113 => x"cce45280",
          3114 => x"ea1651e0",
          3115 => x"b13f81de",
          3116 => x"c0085581",
          3117 => x"dec00880",
          3118 => x"2e9d3885",
          3119 => x"5381cce8",
          3120 => x"52818616",
          3121 => x"51e0973f",
          3122 => x"81dec008",
          3123 => x"5581dec0",
          3124 => x"08802e83",
          3125 => x"38825574",
          3126 => x"81dec00c",
          3127 => x"883d0d04",
          3128 => x"f23d0d61",
          3129 => x"02840580",
          3130 => x"cb053358",
          3131 => x"5580750c",
          3132 => x"6051fce1",
          3133 => x"3f81dec0",
          3134 => x"08588b56",
          3135 => x"800b81de",
          3136 => x"c0082486",
          3137 => x"fc3881de",
          3138 => x"c0088429",
          3139 => x"81dedc05",
          3140 => x"70085553",
          3141 => x"8c567380",
          3142 => x"2e86e638",
          3143 => x"73750c76",
          3144 => x"81fe0674",
          3145 => x"33545772",
          3146 => x"802eae38",
          3147 => x"81143351",
          3148 => x"d7ca3f81",
          3149 => x"dec00881",
          3150 => x"ff067081",
          3151 => x"06545572",
          3152 => x"98387680",
          3153 => x"2e86b838",
          3154 => x"74822a70",
          3155 => x"81065153",
          3156 => x"8a567286",
          3157 => x"ac3886a7",
          3158 => x"39807434",
          3159 => x"77811534",
          3160 => x"81528114",
          3161 => x"3351d7b2",
          3162 => x"3f81dec0",
          3163 => x"0881ff06",
          3164 => x"70810654",
          3165 => x"55835672",
          3166 => x"86873876",
          3167 => x"802e8f38",
          3168 => x"74822a70",
          3169 => x"81065153",
          3170 => x"8a567285",
          3171 => x"f4388070",
          3172 => x"5374525b",
          3173 => x"fda33f81",
          3174 => x"dec00881",
          3175 => x"ff065776",
          3176 => x"822e0981",
          3177 => x"0680e238",
          3178 => x"8c3d7456",
          3179 => x"58835683",
          3180 => x"f6153370",
          3181 => x"58537280",
          3182 => x"2e8d3883",
          3183 => x"fa1551dc",
          3184 => x"e83f81de",
          3185 => x"c0085776",
          3186 => x"78708405",
          3187 => x"5a0cff16",
          3188 => x"90165656",
          3189 => x"758025d7",
          3190 => x"38800b8d",
          3191 => x"3d545672",
          3192 => x"70840554",
          3193 => x"085b8357",
          3194 => x"7a802e95",
          3195 => x"387a5273",
          3196 => x"51fcc63f",
          3197 => x"81dec008",
          3198 => x"81ff0657",
          3199 => x"81772789",
          3200 => x"38811656",
          3201 => x"837627d7",
          3202 => x"38815676",
          3203 => x"842e84f1",
          3204 => x"388d5676",
          3205 => x"812684e9",
          3206 => x"38bf1451",
          3207 => x"dbf43f81",
          3208 => x"dec00883",
          3209 => x"ffff0653",
          3210 => x"7284802e",
          3211 => x"09810684",
          3212 => x"d03880ca",
          3213 => x"1451dbda",
          3214 => x"3f81dec0",
          3215 => x"0883ffff",
          3216 => x"0658778d",
          3217 => x"3880d814",
          3218 => x"51dbde3f",
          3219 => x"81dec008",
          3220 => x"58779c15",
          3221 => x"0c80c414",
          3222 => x"33821534",
          3223 => x"80c41433",
          3224 => x"ff117081",
          3225 => x"ff065154",
          3226 => x"558d5672",
          3227 => x"81268491",
          3228 => x"387481ff",
          3229 => x"06787129",
          3230 => x"80c11633",
          3231 => x"52595372",
          3232 => x"8a152372",
          3233 => x"802e8b38",
          3234 => x"ff137306",
          3235 => x"5372802e",
          3236 => x"86388d56",
          3237 => x"83eb3980",
          3238 => x"c51451da",
          3239 => x"f53f81de",
          3240 => x"c0085381",
          3241 => x"dec00888",
          3242 => x"1523728f",
          3243 => x"06578d56",
          3244 => x"7683ce38",
          3245 => x"80c71451",
          3246 => x"dad83f81",
          3247 => x"dec00883",
          3248 => x"ffff0655",
          3249 => x"748d3880",
          3250 => x"d41451da",
          3251 => x"dc3f81de",
          3252 => x"c0085580",
          3253 => x"c21451da",
          3254 => x"b93f81de",
          3255 => x"c00883ff",
          3256 => x"ff06538d",
          3257 => x"5672802e",
          3258 => x"83973888",
          3259 => x"14227814",
          3260 => x"71842a05",
          3261 => x"5a5a7875",
          3262 => x"26838638",
          3263 => x"8a142252",
          3264 => x"74793151",
          3265 => x"ffacf03f",
          3266 => x"81dec008",
          3267 => x"5581dec0",
          3268 => x"08802e82",
          3269 => x"ec3881de",
          3270 => x"c00880ff",
          3271 => x"fffff526",
          3272 => x"83388357",
          3273 => x"7483fff5",
          3274 => x"26833882",
          3275 => x"57749ff5",
          3276 => x"26853881",
          3277 => x"5789398d",
          3278 => x"5676802e",
          3279 => x"82c33882",
          3280 => x"15709816",
          3281 => x"0c7ba016",
          3282 => x"0c731c70",
          3283 => x"a4170c7a",
          3284 => x"1dac170c",
          3285 => x"54557683",
          3286 => x"2e098106",
          3287 => x"af3880de",
          3288 => x"1451d9ae",
          3289 => x"3f81dec0",
          3290 => x"0883ffff",
          3291 => x"06538d56",
          3292 => x"72828e38",
          3293 => x"79828a38",
          3294 => x"80e01451",
          3295 => x"d9ab3f81",
          3296 => x"dec008a8",
          3297 => x"150c7482",
          3298 => x"2b53a239",
          3299 => x"8d567980",
          3300 => x"2e81ee38",
          3301 => x"7713a815",
          3302 => x"0c741553",
          3303 => x"76822e8d",
          3304 => x"38741015",
          3305 => x"70812a76",
          3306 => x"81060551",
          3307 => x"5383ff13",
          3308 => x"892a538d",
          3309 => x"56729c15",
          3310 => x"082681c5",
          3311 => x"38ff0b90",
          3312 => x"150cff0b",
          3313 => x"8c150cff",
          3314 => x"800b8415",
          3315 => x"3476832e",
          3316 => x"09810681",
          3317 => x"923880e4",
          3318 => x"1451d8b6",
          3319 => x"3f81dec0",
          3320 => x"0883ffff",
          3321 => x"06537281",
          3322 => x"2e098106",
          3323 => x"80f93881",
          3324 => x"1b527351",
          3325 => x"dbb83f81",
          3326 => x"dec00880",
          3327 => x"ea3881de",
          3328 => x"c0088415",
          3329 => x"3484b214",
          3330 => x"51d8873f",
          3331 => x"81dec008",
          3332 => x"83ffff06",
          3333 => x"537282d4",
          3334 => x"d52e0981",
          3335 => x"0680c838",
          3336 => x"b41451d8",
          3337 => x"843f81de",
          3338 => x"c008848b",
          3339 => x"85a4d22e",
          3340 => x"098106b3",
          3341 => x"38849814",
          3342 => x"51d7ee3f",
          3343 => x"81dec008",
          3344 => x"868a85e4",
          3345 => x"f22e0981",
          3346 => x"069d3884",
          3347 => x"9c1451d7",
          3348 => x"d83f81de",
          3349 => x"c0089015",
          3350 => x"0c84a014",
          3351 => x"51d7ca3f",
          3352 => x"81dec008",
          3353 => x"8c150c76",
          3354 => x"743481de",
          3355 => x"ec228105",
          3356 => x"537281de",
          3357 => x"ec237286",
          3358 => x"1523800b",
          3359 => x"94150c80",
          3360 => x"567581de",
          3361 => x"c00c903d",
          3362 => x"0d04fb3d",
          3363 => x"0d775489",
          3364 => x"5573802e",
          3365 => x"b9387308",
          3366 => x"5372802e",
          3367 => x"b1387233",
          3368 => x"5271802e",
          3369 => x"a9388613",
          3370 => x"22841522",
          3371 => x"57527176",
          3372 => x"2e098106",
          3373 => x"99388113",
          3374 => x"3351d0c0",
          3375 => x"3f81dec0",
          3376 => x"08810652",
          3377 => x"71883871",
          3378 => x"74085455",
          3379 => x"83398053",
          3380 => x"7873710c",
          3381 => x"527481de",
          3382 => x"c00c873d",
          3383 => x"0d04fa3d",
          3384 => x"0d02ab05",
          3385 => x"337a5889",
          3386 => x"3dfc0552",
          3387 => x"56f4e63f",
          3388 => x"8b54800b",
          3389 => x"81dec008",
          3390 => x"24bc3881",
          3391 => x"dec00884",
          3392 => x"2981dedc",
          3393 => x"05700855",
          3394 => x"5573802e",
          3395 => x"84388074",
          3396 => x"34785473",
          3397 => x"802e8438",
          3398 => x"80743478",
          3399 => x"750c7554",
          3400 => x"75802e92",
          3401 => x"38805389",
          3402 => x"3d705384",
          3403 => x"0551f7b0",
          3404 => x"3f81dec0",
          3405 => x"08547381",
          3406 => x"dec00c88",
          3407 => x"3d0d04eb",
          3408 => x"3d0d6702",
          3409 => x"840580e7",
          3410 => x"05335959",
          3411 => x"89547880",
          3412 => x"2e84c838",
          3413 => x"77bf0670",
          3414 => x"54983dd0",
          3415 => x"0553993d",
          3416 => x"84055258",
          3417 => x"f6fa3f81",
          3418 => x"dec00855",
          3419 => x"81dec008",
          3420 => x"84a4387a",
          3421 => x"5c68528c",
          3422 => x"3d705256",
          3423 => x"edc63f81",
          3424 => x"dec00855",
          3425 => x"81dec008",
          3426 => x"92380280",
          3427 => x"d7053370",
          3428 => x"982b5557",
          3429 => x"73802583",
          3430 => x"38865577",
          3431 => x"9c065473",
          3432 => x"802e81ab",
          3433 => x"3874802e",
          3434 => x"95387484",
          3435 => x"2e098106",
          3436 => x"aa387551",
          3437 => x"eaf83f81",
          3438 => x"dec00855",
          3439 => x"9e3902b2",
          3440 => x"05339106",
          3441 => x"547381b8",
          3442 => x"3877822a",
          3443 => x"70810651",
          3444 => x"5473802e",
          3445 => x"8e388855",
          3446 => x"83bc3977",
          3447 => x"88075874",
          3448 => x"83b43877",
          3449 => x"832a7081",
          3450 => x"06515473",
          3451 => x"802e81af",
          3452 => x"3862527a",
          3453 => x"51e8a53f",
          3454 => x"81dec008",
          3455 => x"568288b2",
          3456 => x"0a52628e",
          3457 => x"0551d4ea",
          3458 => x"3f6254a0",
          3459 => x"0b8b1534",
          3460 => x"80536252",
          3461 => x"7a51e8bd",
          3462 => x"3f805262",
          3463 => x"9c0551d4",
          3464 => x"d13f7a54",
          3465 => x"810b8315",
          3466 => x"3475802e",
          3467 => x"80f1387a",
          3468 => x"b0110851",
          3469 => x"54805375",
          3470 => x"52973dd4",
          3471 => x"0551ddbe",
          3472 => x"3f81dec0",
          3473 => x"085581de",
          3474 => x"c00882ca",
          3475 => x"38b73974",
          3476 => x"82c43802",
          3477 => x"b2053370",
          3478 => x"842a7081",
          3479 => x"06515556",
          3480 => x"73802e86",
          3481 => x"38845582",
          3482 => x"ad397781",
          3483 => x"2a708106",
          3484 => x"51547380",
          3485 => x"2ea93875",
          3486 => x"81065473",
          3487 => x"802ea038",
          3488 => x"87558292",
          3489 => x"3973527a",
          3490 => x"51d6a33f",
          3491 => x"81dec008",
          3492 => x"7bff188c",
          3493 => x"120c5555",
          3494 => x"81dec008",
          3495 => x"81f83877",
          3496 => x"832a7081",
          3497 => x"06515473",
          3498 => x"802e8638",
          3499 => x"7780c007",
          3500 => x"587ab011",
          3501 => x"08a01b0c",
          3502 => x"63a41b0c",
          3503 => x"63537052",
          3504 => x"57e6d93f",
          3505 => x"81dec008",
          3506 => x"81dec008",
          3507 => x"881b0c63",
          3508 => x"9c05525a",
          3509 => x"d2d33f81",
          3510 => x"dec00881",
          3511 => x"dec0088c",
          3512 => x"1b0c777a",
          3513 => x"0c568617",
          3514 => x"22841a23",
          3515 => x"77901a34",
          3516 => x"800b911a",
          3517 => x"34800b9c",
          3518 => x"1a0c800b",
          3519 => x"941a0c77",
          3520 => x"852a7081",
          3521 => x"06515473",
          3522 => x"802e818d",
          3523 => x"3881dec0",
          3524 => x"08802e81",
          3525 => x"843881de",
          3526 => x"c008941a",
          3527 => x"0c8a1722",
          3528 => x"70892b7b",
          3529 => x"525957a8",
          3530 => x"39765278",
          3531 => x"51d79f3f",
          3532 => x"81dec008",
          3533 => x"5781dec0",
          3534 => x"08812683",
          3535 => x"38825581",
          3536 => x"dec008ff",
          3537 => x"2e098106",
          3538 => x"83387955",
          3539 => x"75783156",
          3540 => x"74307076",
          3541 => x"07802551",
          3542 => x"54777627",
          3543 => x"8a388170",
          3544 => x"7506555a",
          3545 => x"73c33876",
          3546 => x"981a0c74",
          3547 => x"a9387583",
          3548 => x"ff065473",
          3549 => x"802ea238",
          3550 => x"76527a51",
          3551 => x"d6a63f81",
          3552 => x"dec00885",
          3553 => x"3882558e",
          3554 => x"3975892a",
          3555 => x"81dec008",
          3556 => x"059c1a0c",
          3557 => x"84398079",
          3558 => x"0c745473",
          3559 => x"81dec00c",
          3560 => x"973d0d04",
          3561 => x"f23d0d60",
          3562 => x"63656440",
          3563 => x"405d5980",
          3564 => x"7e0c903d",
          3565 => x"fc055278",
          3566 => x"51f9cf3f",
          3567 => x"81dec008",
          3568 => x"5581dec0",
          3569 => x"088a3891",
          3570 => x"19335574",
          3571 => x"802e8638",
          3572 => x"745682c4",
          3573 => x"39901933",
          3574 => x"81065587",
          3575 => x"5674802e",
          3576 => x"82b63895",
          3577 => x"39820b91",
          3578 => x"1a348256",
          3579 => x"82aa3981",
          3580 => x"0b911a34",
          3581 => x"815682a0",
          3582 => x"398c1908",
          3583 => x"941a0831",
          3584 => x"55747c27",
          3585 => x"8338745c",
          3586 => x"7b802e82",
          3587 => x"89389419",
          3588 => x"087083ff",
          3589 => x"06565674",
          3590 => x"81b2387e",
          3591 => x"8a1122ff",
          3592 => x"0577892a",
          3593 => x"065b5579",
          3594 => x"a8387587",
          3595 => x"38881908",
          3596 => x"558f3998",
          3597 => x"19085278",
          3598 => x"51d5933f",
          3599 => x"81dec008",
          3600 => x"55817527",
          3601 => x"ff9f3874",
          3602 => x"ff2effa3",
          3603 => x"3874981a",
          3604 => x"0c981908",
          3605 => x"527e51d4",
          3606 => x"cb3f81de",
          3607 => x"c008802e",
          3608 => x"ff833881",
          3609 => x"dec0081a",
          3610 => x"7c892a59",
          3611 => x"5777802e",
          3612 => x"80d63877",
          3613 => x"1a7f8a11",
          3614 => x"22585c55",
          3615 => x"75752785",
          3616 => x"38757a31",
          3617 => x"58775476",
          3618 => x"537c5281",
          3619 => x"1b3351ca",
          3620 => x"883f81de",
          3621 => x"c008fed7",
          3622 => x"387e8311",
          3623 => x"33565674",
          3624 => x"802e9f38",
          3625 => x"b0160877",
          3626 => x"31557478",
          3627 => x"27943884",
          3628 => x"8053b416",
          3629 => x"52b01608",
          3630 => x"7731892b",
          3631 => x"7d0551cf",
          3632 => x"e03f7789",
          3633 => x"2b56b939",
          3634 => x"769c1a0c",
          3635 => x"94190883",
          3636 => x"ff068480",
          3637 => x"71315755",
          3638 => x"7b762783",
          3639 => x"387b569c",
          3640 => x"1908527e",
          3641 => x"51d1c73f",
          3642 => x"81dec008",
          3643 => x"fe813875",
          3644 => x"53941908",
          3645 => x"83ff061f",
          3646 => x"b405527c",
          3647 => x"51cfa23f",
          3648 => x"7b76317e",
          3649 => x"08177f0c",
          3650 => x"761e941b",
          3651 => x"0818941c",
          3652 => x"0c5e5cfd",
          3653 => x"f3398056",
          3654 => x"7581dec0",
          3655 => x"0c903d0d",
          3656 => x"04f23d0d",
          3657 => x"60636564",
          3658 => x"40405d58",
          3659 => x"807e0c90",
          3660 => x"3dfc0552",
          3661 => x"7751f6d2",
          3662 => x"3f81dec0",
          3663 => x"085581de",
          3664 => x"c0088a38",
          3665 => x"91183355",
          3666 => x"74802e86",
          3667 => x"38745683",
          3668 => x"b8399018",
          3669 => x"3370812a",
          3670 => x"70810651",
          3671 => x"56568756",
          3672 => x"74802e83",
          3673 => x"a4389539",
          3674 => x"820b9119",
          3675 => x"34825683",
          3676 => x"9839810b",
          3677 => x"91193481",
          3678 => x"56838e39",
          3679 => x"9418087c",
          3680 => x"11565674",
          3681 => x"76278438",
          3682 => x"75095c7b",
          3683 => x"802e82ec",
          3684 => x"38941808",
          3685 => x"7083ff06",
          3686 => x"56567481",
          3687 => x"fd387e8a",
          3688 => x"1122ff05",
          3689 => x"77892a06",
          3690 => x"5c557abf",
          3691 => x"38758c38",
          3692 => x"88180855",
          3693 => x"749c387a",
          3694 => x"52853998",
          3695 => x"18085277",
          3696 => x"51d7e73f",
          3697 => x"81dec008",
          3698 => x"5581dec0",
          3699 => x"08802e82",
          3700 => x"ab387481",
          3701 => x"2eff9138",
          3702 => x"74ff2eff",
          3703 => x"95387498",
          3704 => x"190c8818",
          3705 => x"08853874",
          3706 => x"88190c7e",
          3707 => x"55b01508",
          3708 => x"9c19082e",
          3709 => x"0981068d",
          3710 => x"387451ce",
          3711 => x"c13f81de",
          3712 => x"c008feee",
          3713 => x"38981808",
          3714 => x"527e51d1",
          3715 => x"973f81de",
          3716 => x"c008802e",
          3717 => x"fed23881",
          3718 => x"dec0081b",
          3719 => x"7c892a5a",
          3720 => x"5778802e",
          3721 => x"80d53878",
          3722 => x"1b7f8a11",
          3723 => x"22585b55",
          3724 => x"75752785",
          3725 => x"38757b31",
          3726 => x"59785476",
          3727 => x"537c5281",
          3728 => x"1a3351c8",
          3729 => x"be3f81de",
          3730 => x"c008fea6",
          3731 => x"387eb011",
          3732 => x"08783156",
          3733 => x"56747927",
          3734 => x"9b388480",
          3735 => x"53b01608",
          3736 => x"7731892b",
          3737 => x"7d0552b4",
          3738 => x"1651ccb5",
          3739 => x"3f7e5580",
          3740 => x"0b831634",
          3741 => x"78892b56",
          3742 => x"80db398c",
          3743 => x"18089419",
          3744 => x"08269338",
          3745 => x"7e51cdb6",
          3746 => x"3f81dec0",
          3747 => x"08fde338",
          3748 => x"7e77b012",
          3749 => x"0c55769c",
          3750 => x"190c9418",
          3751 => x"0883ff06",
          3752 => x"84807131",
          3753 => x"57557b76",
          3754 => x"2783387b",
          3755 => x"569c1808",
          3756 => x"527e51cd",
          3757 => x"f93f81de",
          3758 => x"c008fdb6",
          3759 => x"3875537c",
          3760 => x"52941808",
          3761 => x"83ff061f",
          3762 => x"b40551cb",
          3763 => x"d43f7e55",
          3764 => x"810b8316",
          3765 => x"347b7631",
          3766 => x"7e08177f",
          3767 => x"0c761e94",
          3768 => x"1a081870",
          3769 => x"941c0c8c",
          3770 => x"1b085858",
          3771 => x"5e5c7476",
          3772 => x"27833875",
          3773 => x"55748c19",
          3774 => x"0cfd9039",
          3775 => x"90183380",
          3776 => x"c0075574",
          3777 => x"90193480",
          3778 => x"567581de",
          3779 => x"c00c903d",
          3780 => x"0d04f83d",
          3781 => x"0d7a8b3d",
          3782 => x"fc055370",
          3783 => x"5256f2ea",
          3784 => x"3f81dec0",
          3785 => x"085781de",
          3786 => x"c00880fb",
          3787 => x"38901633",
          3788 => x"70862a70",
          3789 => x"81065155",
          3790 => x"5573802e",
          3791 => x"80e938a0",
          3792 => x"16085278",
          3793 => x"51cce73f",
          3794 => x"81dec008",
          3795 => x"5781dec0",
          3796 => x"0880d438",
          3797 => x"a416088b",
          3798 => x"1133a007",
          3799 => x"5555738b",
          3800 => x"16348816",
          3801 => x"08537452",
          3802 => x"750851dd",
          3803 => x"e83f8c16",
          3804 => x"08529c15",
          3805 => x"51c9fb3f",
          3806 => x"8288b20a",
          3807 => x"52961551",
          3808 => x"c9f03f76",
          3809 => x"52921551",
          3810 => x"c9ca3f78",
          3811 => x"54810b83",
          3812 => x"15347851",
          3813 => x"ccdf3f81",
          3814 => x"dec00890",
          3815 => x"173381bf",
          3816 => x"06555773",
          3817 => x"90173476",
          3818 => x"81dec00c",
          3819 => x"8a3d0d04",
          3820 => x"fc3d0d76",
          3821 => x"705254fe",
          3822 => x"d93f81de",
          3823 => x"c0085381",
          3824 => x"dec0089c",
          3825 => x"38863dfc",
          3826 => x"05527351",
          3827 => x"f1bc3f81",
          3828 => x"dec00853",
          3829 => x"81dec008",
          3830 => x"873881de",
          3831 => x"c008740c",
          3832 => x"7281dec0",
          3833 => x"0c863d0d",
          3834 => x"04ff3d0d",
          3835 => x"843d51e6",
          3836 => x"e43f8b52",
          3837 => x"800b81de",
          3838 => x"c008248b",
          3839 => x"3881dec0",
          3840 => x"0881def0",
          3841 => x"34805271",
          3842 => x"81dec00c",
          3843 => x"833d0d04",
          3844 => x"ef3d0d80",
          3845 => x"53933dd0",
          3846 => x"0552943d",
          3847 => x"51e9c13f",
          3848 => x"81dec008",
          3849 => x"5581dec0",
          3850 => x"0880e038",
          3851 => x"76586352",
          3852 => x"933dd405",
          3853 => x"51e08d3f",
          3854 => x"81dec008",
          3855 => x"5581dec0",
          3856 => x"08bc3802",
          3857 => x"80c70533",
          3858 => x"70982b55",
          3859 => x"56738025",
          3860 => x"8938767a",
          3861 => x"94120c54",
          3862 => x"b23902a2",
          3863 => x"05337084",
          3864 => x"2a708106",
          3865 => x"51555673",
          3866 => x"802e9e38",
          3867 => x"767f5370",
          3868 => x"5254dba8",
          3869 => x"3f81dec0",
          3870 => x"0894150c",
          3871 => x"8e3981de",
          3872 => x"c008842e",
          3873 => x"09810683",
          3874 => x"38855574",
          3875 => x"81dec00c",
          3876 => x"933d0d04",
          3877 => x"e43d0d6f",
          3878 => x"6f5b5b80",
          3879 => x"7a348053",
          3880 => x"9e3dffb8",
          3881 => x"05529f3d",
          3882 => x"51e8b53f",
          3883 => x"81dec008",
          3884 => x"5781dec0",
          3885 => x"0882fc38",
          3886 => x"7b437a7c",
          3887 => x"94110847",
          3888 => x"55586454",
          3889 => x"73802e81",
          3890 => x"ed38a052",
          3891 => x"933d7052",
          3892 => x"55d5ea3f",
          3893 => x"81dec008",
          3894 => x"5781dec0",
          3895 => x"0882d438",
          3896 => x"68527b51",
          3897 => x"c9c83f81",
          3898 => x"dec00857",
          3899 => x"81dec008",
          3900 => x"82c13869",
          3901 => x"527b51da",
          3902 => x"a33f81de",
          3903 => x"c0084576",
          3904 => x"527451d5",
          3905 => x"b83f81de",
          3906 => x"c0085781",
          3907 => x"dec00882",
          3908 => x"a2388052",
          3909 => x"7451daeb",
          3910 => x"3f81dec0",
          3911 => x"085781de",
          3912 => x"c008a438",
          3913 => x"69527b51",
          3914 => x"d9f23f73",
          3915 => x"81dec008",
          3916 => x"2ea63876",
          3917 => x"527451d6",
          3918 => x"cf3f81de",
          3919 => x"c0085781",
          3920 => x"dec00880",
          3921 => x"2ecc3876",
          3922 => x"842e0981",
          3923 => x"06863882",
          3924 => x"5781e039",
          3925 => x"7681dc38",
          3926 => x"9e3dffbc",
          3927 => x"05527451",
          3928 => x"dcc93f76",
          3929 => x"903d7811",
          3930 => x"81113351",
          3931 => x"565a5673",
          3932 => x"802e9138",
          3933 => x"02b90555",
          3934 => x"81168116",
          3935 => x"70335656",
          3936 => x"5673f538",
          3937 => x"81165473",
          3938 => x"78268190",
          3939 => x"3875802e",
          3940 => x"99387816",
          3941 => x"810555ff",
          3942 => x"186f11ff",
          3943 => x"18ff1858",
          3944 => x"58555874",
          3945 => x"33743475",
          3946 => x"ee38ff18",
          3947 => x"6f115558",
          3948 => x"af7434fe",
          3949 => x"8d39777b",
          3950 => x"2e098106",
          3951 => x"8a38ff18",
          3952 => x"6f115558",
          3953 => x"af743480",
          3954 => x"0b81def0",
          3955 => x"33708429",
          3956 => x"81cda405",
          3957 => x"70087033",
          3958 => x"525c5656",
          3959 => x"5673762e",
          3960 => x"8d388116",
          3961 => x"701a7033",
          3962 => x"51555673",
          3963 => x"f5388216",
          3964 => x"54737826",
          3965 => x"a7388055",
          3966 => x"74762791",
          3967 => x"38741954",
          3968 => x"73337a70",
          3969 => x"81055c34",
          3970 => x"811555ec",
          3971 => x"39ba7a70",
          3972 => x"81055c34",
          3973 => x"74ff2e09",
          3974 => x"81068538",
          3975 => x"91579439",
          3976 => x"6e188119",
          3977 => x"59547333",
          3978 => x"7a708105",
          3979 => x"5c347a78",
          3980 => x"26ee3880",
          3981 => x"7a347681",
          3982 => x"dec00c9e",
          3983 => x"3d0d04f7",
          3984 => x"3d0d7b7d",
          3985 => x"8d3dfc05",
          3986 => x"54715357",
          3987 => x"55ecbb3f",
          3988 => x"81dec008",
          3989 => x"5381dec0",
          3990 => x"0882fa38",
          3991 => x"91153353",
          3992 => x"7282f238",
          3993 => x"8c150854",
          3994 => x"73762792",
          3995 => x"38901533",
          3996 => x"70812a70",
          3997 => x"81065154",
          3998 => x"57728338",
          3999 => x"73569415",
          4000 => x"08548070",
          4001 => x"94170c58",
          4002 => x"75782e82",
          4003 => x"9738798a",
          4004 => x"11227089",
          4005 => x"2b595153",
          4006 => x"73782eb7",
          4007 => x"387652ff",
          4008 => x"1651ff95",
          4009 => x"d23f81de",
          4010 => x"c008ff15",
          4011 => x"78547053",
          4012 => x"5553ff95",
          4013 => x"c23f81de",
          4014 => x"c0087326",
          4015 => x"96387630",
          4016 => x"70750670",
          4017 => x"94180c77",
          4018 => x"71319818",
          4019 => x"08575851",
          4020 => x"53b13988",
          4021 => x"15085473",
          4022 => x"a6387352",
          4023 => x"7451cdca",
          4024 => x"3f81dec0",
          4025 => x"085481de",
          4026 => x"c008812e",
          4027 => x"819a3881",
          4028 => x"dec008ff",
          4029 => x"2e819b38",
          4030 => x"81dec008",
          4031 => x"88160c73",
          4032 => x"98160c73",
          4033 => x"802e819c",
          4034 => x"38767627",
          4035 => x"80dc3875",
          4036 => x"77319416",
          4037 => x"08189417",
          4038 => x"0c901633",
          4039 => x"70812a70",
          4040 => x"81065155",
          4041 => x"5a567280",
          4042 => x"2e9a3873",
          4043 => x"527451cc",
          4044 => x"f93f81de",
          4045 => x"c0085481",
          4046 => x"dec00894",
          4047 => x"3881dec0",
          4048 => x"0856a739",
          4049 => x"73527451",
          4050 => x"c7843f81",
          4051 => x"dec00854",
          4052 => x"73ff2ebe",
          4053 => x"38817427",
          4054 => x"af387953",
          4055 => x"73981408",
          4056 => x"27a63873",
          4057 => x"98160cff",
          4058 => x"a0399415",
          4059 => x"08169416",
          4060 => x"0c7583ff",
          4061 => x"06537280",
          4062 => x"2eaa3873",
          4063 => x"527951c6",
          4064 => x"a33f81de",
          4065 => x"c0089438",
          4066 => x"820b9116",
          4067 => x"34825380",
          4068 => x"c439810b",
          4069 => x"91163481",
          4070 => x"53bb3975",
          4071 => x"892a81de",
          4072 => x"c0080558",
          4073 => x"94150854",
          4074 => x"8c150874",
          4075 => x"27903873",
          4076 => x"8c160c90",
          4077 => x"153380c0",
          4078 => x"07537290",
          4079 => x"16347383",
          4080 => x"ff065372",
          4081 => x"802e8c38",
          4082 => x"779c1608",
          4083 => x"2e853877",
          4084 => x"9c160c80",
          4085 => x"537281de",
          4086 => x"c00c8b3d",
          4087 => x"0d04f93d",
          4088 => x"0d795689",
          4089 => x"5475802e",
          4090 => x"818a3880",
          4091 => x"53893dfc",
          4092 => x"05528a3d",
          4093 => x"840551e1",
          4094 => x"e73f81de",
          4095 => x"c0085581",
          4096 => x"dec00880",
          4097 => x"ea387776",
          4098 => x"0c7a5275",
          4099 => x"51d8b53f",
          4100 => x"81dec008",
          4101 => x"5581dec0",
          4102 => x"0880c338",
          4103 => x"ab163370",
          4104 => x"982b5557",
          4105 => x"807424a2",
          4106 => x"38861633",
          4107 => x"70842a70",
          4108 => x"81065155",
          4109 => x"5773802e",
          4110 => x"ad389c16",
          4111 => x"08527751",
          4112 => x"d3da3f81",
          4113 => x"dec00888",
          4114 => x"170c7754",
          4115 => x"86142284",
          4116 => x"17237452",
          4117 => x"7551cee5",
          4118 => x"3f81dec0",
          4119 => x"08557484",
          4120 => x"2e098106",
          4121 => x"85388555",
          4122 => x"86397480",
          4123 => x"2e843880",
          4124 => x"760c7454",
          4125 => x"7381dec0",
          4126 => x"0c893d0d",
          4127 => x"04fc3d0d",
          4128 => x"76873dfc",
          4129 => x"05537052",
          4130 => x"53e7ff3f",
          4131 => x"81dec008",
          4132 => x"873881de",
          4133 => x"c008730c",
          4134 => x"863d0d04",
          4135 => x"fb3d0d77",
          4136 => x"79893dfc",
          4137 => x"05547153",
          4138 => x"5654e7de",
          4139 => x"3f81dec0",
          4140 => x"085381de",
          4141 => x"c00880df",
          4142 => x"38749338",
          4143 => x"81dec008",
          4144 => x"527351cd",
          4145 => x"f83f81de",
          4146 => x"c0085380",
          4147 => x"ca3981de",
          4148 => x"c0085273",
          4149 => x"51d3ac3f",
          4150 => x"81dec008",
          4151 => x"5381dec0",
          4152 => x"08842e09",
          4153 => x"81068538",
          4154 => x"80538739",
          4155 => x"81dec008",
          4156 => x"a6387452",
          4157 => x"7351d5b3",
          4158 => x"3f725273",
          4159 => x"51cf893f",
          4160 => x"81dec008",
          4161 => x"84327030",
          4162 => x"7072079f",
          4163 => x"2c7081de",
          4164 => x"c0080651",
          4165 => x"51545472",
          4166 => x"81dec00c",
          4167 => x"873d0d04",
          4168 => x"ee3d0d65",
          4169 => x"57805389",
          4170 => x"3d705396",
          4171 => x"3d5256df",
          4172 => x"af3f81de",
          4173 => x"c0085581",
          4174 => x"dec008b2",
          4175 => x"38645275",
          4176 => x"51d6813f",
          4177 => x"81dec008",
          4178 => x"5581dec0",
          4179 => x"08a03802",
          4180 => x"80cb0533",
          4181 => x"70982b55",
          4182 => x"58738025",
          4183 => x"85388655",
          4184 => x"8d397680",
          4185 => x"2e883876",
          4186 => x"527551d4",
          4187 => x"be3f7481",
          4188 => x"dec00c94",
          4189 => x"3d0d04f0",
          4190 => x"3d0d6365",
          4191 => x"555c8053",
          4192 => x"923dec05",
          4193 => x"52933d51",
          4194 => x"ded63f81",
          4195 => x"dec0085b",
          4196 => x"81dec008",
          4197 => x"8280387c",
          4198 => x"740c7308",
          4199 => x"981108fe",
          4200 => x"11901308",
          4201 => x"59565855",
          4202 => x"75742691",
          4203 => x"38757c0c",
          4204 => x"81e43981",
          4205 => x"5b81cc39",
          4206 => x"825b81c7",
          4207 => x"3981dec0",
          4208 => x"08753355",
          4209 => x"5973812e",
          4210 => x"098106bf",
          4211 => x"3882755f",
          4212 => x"57765292",
          4213 => x"3df00551",
          4214 => x"c1f43f81",
          4215 => x"dec008ff",
          4216 => x"2ed13881",
          4217 => x"dec00881",
          4218 => x"2ece3881",
          4219 => x"dec00830",
          4220 => x"7081dec0",
          4221 => x"08078025",
          4222 => x"7a058119",
          4223 => x"7f53595a",
          4224 => x"54981408",
          4225 => x"7726ca38",
          4226 => x"80f939a4",
          4227 => x"150881de",
          4228 => x"c0085758",
          4229 => x"75983877",
          4230 => x"5281187d",
          4231 => x"5258ffbf",
          4232 => x"8d3f81de",
          4233 => x"c0085b81",
          4234 => x"dec00880",
          4235 => x"d6387c70",
          4236 => x"337712ff",
          4237 => x"1a5d5256",
          4238 => x"5474822e",
          4239 => x"0981069e",
          4240 => x"38b41451",
          4241 => x"ffbbcb3f",
          4242 => x"81dec008",
          4243 => x"83ffff06",
          4244 => x"70307080",
          4245 => x"251b8219",
          4246 => x"595b5154",
          4247 => x"9b39b414",
          4248 => x"51ffbbc5",
          4249 => x"3f81dec0",
          4250 => x"08f00a06",
          4251 => x"70307080",
          4252 => x"251b8419",
          4253 => x"595b5154",
          4254 => x"7583ff06",
          4255 => x"7a585679",
          4256 => x"ff923878",
          4257 => x"7c0c7c79",
          4258 => x"90120c84",
          4259 => x"11338107",
          4260 => x"56547484",
          4261 => x"15347a81",
          4262 => x"dec00c92",
          4263 => x"3d0d04f9",
          4264 => x"3d0d798a",
          4265 => x"3dfc0553",
          4266 => x"705257e3",
          4267 => x"dd3f81de",
          4268 => x"c0085681",
          4269 => x"dec00881",
          4270 => x"a8389117",
          4271 => x"33567581",
          4272 => x"a0389017",
          4273 => x"3370812a",
          4274 => x"70810651",
          4275 => x"55558755",
          4276 => x"73802e81",
          4277 => x"8e389417",
          4278 => x"0854738c",
          4279 => x"18082781",
          4280 => x"8038739b",
          4281 => x"3881dec0",
          4282 => x"08538817",
          4283 => x"08527651",
          4284 => x"c48c3f81",
          4285 => x"dec00874",
          4286 => x"88190c56",
          4287 => x"80c93998",
          4288 => x"17085276",
          4289 => x"51ffbfc6",
          4290 => x"3f81dec0",
          4291 => x"08ff2e09",
          4292 => x"81068338",
          4293 => x"815681de",
          4294 => x"c008812e",
          4295 => x"09810685",
          4296 => x"388256a3",
          4297 => x"3975a038",
          4298 => x"775481de",
          4299 => x"c0089815",
          4300 => x"08279438",
          4301 => x"98170853",
          4302 => x"81dec008",
          4303 => x"527651c3",
          4304 => x"bd3f81de",
          4305 => x"c0085694",
          4306 => x"17088c18",
          4307 => x"0c901733",
          4308 => x"80c00754",
          4309 => x"73901834",
          4310 => x"75802e85",
          4311 => x"38759118",
          4312 => x"34755574",
          4313 => x"81dec00c",
          4314 => x"893d0d04",
          4315 => x"e23d0d82",
          4316 => x"53a03dff",
          4317 => x"a40552a1",
          4318 => x"3d51dae4",
          4319 => x"3f81dec0",
          4320 => x"085581de",
          4321 => x"c00881f5",
          4322 => x"387845a1",
          4323 => x"3d085295",
          4324 => x"3d705258",
          4325 => x"d1ae3f81",
          4326 => x"dec00855",
          4327 => x"81dec008",
          4328 => x"81db3802",
          4329 => x"80fb0533",
          4330 => x"70852a70",
          4331 => x"81065155",
          4332 => x"56865573",
          4333 => x"81c73875",
          4334 => x"982b5480",
          4335 => x"742481bd",
          4336 => x"380280d6",
          4337 => x"05337081",
          4338 => x"06585487",
          4339 => x"557681ad",
          4340 => x"386b5278",
          4341 => x"51ccc53f",
          4342 => x"81dec008",
          4343 => x"74842a70",
          4344 => x"81065155",
          4345 => x"5673802e",
          4346 => x"80d43878",
          4347 => x"5481dec0",
          4348 => x"08941508",
          4349 => x"2e818638",
          4350 => x"735a81de",
          4351 => x"c0085c76",
          4352 => x"528a3d70",
          4353 => x"5254c7b5",
          4354 => x"3f81dec0",
          4355 => x"085581de",
          4356 => x"c00880e9",
          4357 => x"3881dec0",
          4358 => x"08527351",
          4359 => x"cce53f81",
          4360 => x"dec00855",
          4361 => x"81dec008",
          4362 => x"86388755",
          4363 => x"80cf3981",
          4364 => x"dec00884",
          4365 => x"2e883881",
          4366 => x"dec00880",
          4367 => x"c0387751",
          4368 => x"cec23f81",
          4369 => x"dec00881",
          4370 => x"dec00830",
          4371 => x"7081dec0",
          4372 => x"08078025",
          4373 => x"51555575",
          4374 => x"802e9438",
          4375 => x"73802e8f",
          4376 => x"38805375",
          4377 => x"527751c1",
          4378 => x"953f81de",
          4379 => x"c0085574",
          4380 => x"8c387851",
          4381 => x"ffbafe3f",
          4382 => x"81dec008",
          4383 => x"557481de",
          4384 => x"c00ca03d",
          4385 => x"0d04e93d",
          4386 => x"0d825399",
          4387 => x"3dc00552",
          4388 => x"9a3d51d8",
          4389 => x"cb3f81de",
          4390 => x"c0085481",
          4391 => x"dec00882",
          4392 => x"b038785e",
          4393 => x"69528e3d",
          4394 => x"705258cf",
          4395 => x"973f81de",
          4396 => x"c0085481",
          4397 => x"dec00886",
          4398 => x"38885482",
          4399 => x"943981de",
          4400 => x"c008842e",
          4401 => x"09810682",
          4402 => x"88380280",
          4403 => x"df053370",
          4404 => x"852a8106",
          4405 => x"51558654",
          4406 => x"7481f638",
          4407 => x"785a7452",
          4408 => x"8a3d7052",
          4409 => x"57c1c33f",
          4410 => x"81dec008",
          4411 => x"75555681",
          4412 => x"dec00883",
          4413 => x"38875481",
          4414 => x"dec00881",
          4415 => x"2e098106",
          4416 => x"83388254",
          4417 => x"81dec008",
          4418 => x"ff2e0981",
          4419 => x"06863881",
          4420 => x"5481b439",
          4421 => x"7381b038",
          4422 => x"81dec008",
          4423 => x"527851c4",
          4424 => x"a43f81de",
          4425 => x"c0085481",
          4426 => x"dec00881",
          4427 => x"9a388b53",
          4428 => x"a052b419",
          4429 => x"51ffb78c",
          4430 => x"3f7854ae",
          4431 => x"0bb41534",
          4432 => x"7854900b",
          4433 => x"bf153482",
          4434 => x"88b20a52",
          4435 => x"80ca1951",
          4436 => x"ffb69f3f",
          4437 => x"755378b4",
          4438 => x"115351c9",
          4439 => x"f83fa053",
          4440 => x"78b41153",
          4441 => x"80d40551",
          4442 => x"ffb6b63f",
          4443 => x"7854ae0b",
          4444 => x"80d51534",
          4445 => x"7f537880",
          4446 => x"d4115351",
          4447 => x"c9d73f78",
          4448 => x"54810b83",
          4449 => x"15347751",
          4450 => x"cba43f81",
          4451 => x"dec00854",
          4452 => x"81dec008",
          4453 => x"b2388288",
          4454 => x"b20a5264",
          4455 => x"960551ff",
          4456 => x"b5d03f75",
          4457 => x"53645278",
          4458 => x"51c9aa3f",
          4459 => x"6454900b",
          4460 => x"8b153478",
          4461 => x"54810b83",
          4462 => x"15347851",
          4463 => x"ffb8b63f",
          4464 => x"81dec008",
          4465 => x"548b3980",
          4466 => x"53755276",
          4467 => x"51ffbeae",
          4468 => x"3f7381de",
          4469 => x"c00c993d",
          4470 => x"0d04da3d",
          4471 => x"0da93d84",
          4472 => x"0551d2f1",
          4473 => x"3f8253a8",
          4474 => x"3dff8405",
          4475 => x"52a93d51",
          4476 => x"d5ee3f81",
          4477 => x"dec00855",
          4478 => x"81dec008",
          4479 => x"82d33878",
          4480 => x"4da93d08",
          4481 => x"529d3d70",
          4482 => x"5258ccb8",
          4483 => x"3f81dec0",
          4484 => x"085581de",
          4485 => x"c00882b9",
          4486 => x"3802819b",
          4487 => x"053381a0",
          4488 => x"06548655",
          4489 => x"7382aa38",
          4490 => x"a053a43d",
          4491 => x"0852a83d",
          4492 => x"ff880551",
          4493 => x"ffb4ea3f",
          4494 => x"ac537752",
          4495 => x"923d7052",
          4496 => x"54ffb4dd",
          4497 => x"3faa3d08",
          4498 => x"527351cb",
          4499 => x"f73f81de",
          4500 => x"c0085581",
          4501 => x"dec00895",
          4502 => x"38636f2e",
          4503 => x"09810688",
          4504 => x"3865a23d",
          4505 => x"082e9238",
          4506 => x"885581e5",
          4507 => x"3981dec0",
          4508 => x"08842e09",
          4509 => x"810681b8",
          4510 => x"387351c9",
          4511 => x"b13f81de",
          4512 => x"c0085581",
          4513 => x"dec00881",
          4514 => x"c8386856",
          4515 => x"9353a83d",
          4516 => x"ff950552",
          4517 => x"8d1651ff",
          4518 => x"b4873f02",
          4519 => x"af05338b",
          4520 => x"17348b16",
          4521 => x"3370842a",
          4522 => x"70810651",
          4523 => x"55557389",
          4524 => x"3874a007",
          4525 => x"54738b17",
          4526 => x"34785481",
          4527 => x"0b831534",
          4528 => x"8b163370",
          4529 => x"842a7081",
          4530 => x"06515555",
          4531 => x"73802e80",
          4532 => x"e5386e64",
          4533 => x"2e80df38",
          4534 => x"75527851",
          4535 => x"c6be3f81",
          4536 => x"dec00852",
          4537 => x"7851ffb7",
          4538 => x"bb3f8255",
          4539 => x"81dec008",
          4540 => x"802e80dd",
          4541 => x"3881dec0",
          4542 => x"08527851",
          4543 => x"ffb5af3f",
          4544 => x"81dec008",
          4545 => x"7980d411",
          4546 => x"58585581",
          4547 => x"dec00880",
          4548 => x"c0388116",
          4549 => x"335473ae",
          4550 => x"2e098106",
          4551 => x"99386353",
          4552 => x"75527651",
          4553 => x"c6af3f78",
          4554 => x"54810b83",
          4555 => x"15348739",
          4556 => x"81dec008",
          4557 => x"9c387751",
          4558 => x"c8ca3f81",
          4559 => x"dec00855",
          4560 => x"81dec008",
          4561 => x"8c387851",
          4562 => x"ffb5aa3f",
          4563 => x"81dec008",
          4564 => x"557481de",
          4565 => x"c00ca83d",
          4566 => x"0d04ed3d",
          4567 => x"0d0280db",
          4568 => x"05330284",
          4569 => x"0580df05",
          4570 => x"33575782",
          4571 => x"53953dd0",
          4572 => x"0552963d",
          4573 => x"51d2e93f",
          4574 => x"81dec008",
          4575 => x"5581dec0",
          4576 => x"0880cf38",
          4577 => x"785a6552",
          4578 => x"953dd405",
          4579 => x"51c9b53f",
          4580 => x"81dec008",
          4581 => x"5581dec0",
          4582 => x"08b83802",
          4583 => x"80cf0533",
          4584 => x"81a00654",
          4585 => x"865573aa",
          4586 => x"3875a706",
          4587 => x"6171098b",
          4588 => x"12337106",
          4589 => x"7a740607",
          4590 => x"51575556",
          4591 => x"748b1534",
          4592 => x"7854810b",
          4593 => x"83153478",
          4594 => x"51ffb4a9",
          4595 => x"3f81dec0",
          4596 => x"08557481",
          4597 => x"dec00c95",
          4598 => x"3d0d04ef",
          4599 => x"3d0d6456",
          4600 => x"8253933d",
          4601 => x"d0055294",
          4602 => x"3d51d1f4",
          4603 => x"3f81dec0",
          4604 => x"085581de",
          4605 => x"c00880cb",
          4606 => x"38765863",
          4607 => x"52933dd4",
          4608 => x"0551c8c0",
          4609 => x"3f81dec0",
          4610 => x"085581de",
          4611 => x"c008b438",
          4612 => x"0280c705",
          4613 => x"3381a006",
          4614 => x"54865573",
          4615 => x"a6388416",
          4616 => x"22861722",
          4617 => x"71902b07",
          4618 => x"5354961f",
          4619 => x"51ffb0c2",
          4620 => x"3f765481",
          4621 => x"0b831534",
          4622 => x"7651ffb3",
          4623 => x"b83f81de",
          4624 => x"c0085574",
          4625 => x"81dec00c",
          4626 => x"933d0d04",
          4627 => x"ea3d0d69",
          4628 => x"6b5c5a80",
          4629 => x"53983dd0",
          4630 => x"0552993d",
          4631 => x"51d1813f",
          4632 => x"81dec008",
          4633 => x"81dec008",
          4634 => x"307081de",
          4635 => x"c0080780",
          4636 => x"25515557",
          4637 => x"79802e81",
          4638 => x"85388170",
          4639 => x"75065555",
          4640 => x"73802e80",
          4641 => x"f9387b5d",
          4642 => x"805f8052",
          4643 => x"8d3d7052",
          4644 => x"54ffbea9",
          4645 => x"3f81dec0",
          4646 => x"085781de",
          4647 => x"c00880d1",
          4648 => x"38745273",
          4649 => x"51c3dc3f",
          4650 => x"81dec008",
          4651 => x"5781dec0",
          4652 => x"08bf3881",
          4653 => x"dec00881",
          4654 => x"dec00865",
          4655 => x"5b595678",
          4656 => x"1881197b",
          4657 => x"18565955",
          4658 => x"74337434",
          4659 => x"8116568a",
          4660 => x"7827ec38",
          4661 => x"8b56751a",
          4662 => x"54807434",
          4663 => x"75802e9e",
          4664 => x"38ff1670",
          4665 => x"1b703351",
          4666 => x"555673a0",
          4667 => x"2ee8388e",
          4668 => x"3976842e",
          4669 => x"09810686",
          4670 => x"38807a34",
          4671 => x"80577630",
          4672 => x"70780780",
          4673 => x"2551547a",
          4674 => x"802e80c1",
          4675 => x"3873802e",
          4676 => x"bc387ba0",
          4677 => x"11085351",
          4678 => x"ffb1933f",
          4679 => x"81dec008",
          4680 => x"5781dec0",
          4681 => x"08a7387b",
          4682 => x"70335555",
          4683 => x"80c35673",
          4684 => x"832e8b38",
          4685 => x"80e45673",
          4686 => x"842e8338",
          4687 => x"a7567515",
          4688 => x"b40551ff",
          4689 => x"ade33f81",
          4690 => x"dec0087b",
          4691 => x"0c7681de",
          4692 => x"c00c983d",
          4693 => x"0d04e63d",
          4694 => x"0d82539c",
          4695 => x"3dffb805",
          4696 => x"529d3d51",
          4697 => x"cefa3f81",
          4698 => x"dec00881",
          4699 => x"dec00856",
          4700 => x"5481dec0",
          4701 => x"08839838",
          4702 => x"8b53a052",
          4703 => x"8b3d7052",
          4704 => x"59ffaec0",
          4705 => x"3f736d70",
          4706 => x"337081ff",
          4707 => x"06525755",
          4708 => x"579f7427",
          4709 => x"81bc3878",
          4710 => x"587481ff",
          4711 => x"066d8105",
          4712 => x"4e705255",
          4713 => x"ffaf893f",
          4714 => x"81dec008",
          4715 => x"802ea538",
          4716 => x"6c703370",
          4717 => x"535754ff",
          4718 => x"aefd3f81",
          4719 => x"dec00880",
          4720 => x"2e8d3874",
          4721 => x"882b7607",
          4722 => x"6d81054e",
          4723 => x"55863981",
          4724 => x"dec00855",
          4725 => x"ff9f1570",
          4726 => x"83ffff06",
          4727 => x"51547399",
          4728 => x"268a38e0",
          4729 => x"157083ff",
          4730 => x"ff065654",
          4731 => x"80ff7527",
          4732 => x"873881cc",
          4733 => x"b4153355",
          4734 => x"74802ea3",
          4735 => x"38745281",
          4736 => x"ceb451ff",
          4737 => x"ae893f81",
          4738 => x"dec00893",
          4739 => x"3881ff75",
          4740 => x"27883876",
          4741 => x"89268838",
          4742 => x"8b398a77",
          4743 => x"27863886",
          4744 => x"5581ec39",
          4745 => x"81ff7527",
          4746 => x"8f387488",
          4747 => x"2a547378",
          4748 => x"7081055a",
          4749 => x"34811757",
          4750 => x"74787081",
          4751 => x"055a3481",
          4752 => x"176d7033",
          4753 => x"7081ff06",
          4754 => x"52575557",
          4755 => x"739f26fe",
          4756 => x"c8388b3d",
          4757 => x"33548655",
          4758 => x"7381e52e",
          4759 => x"81b13876",
          4760 => x"802e9938",
          4761 => x"02a70555",
          4762 => x"76157033",
          4763 => x"515473a0",
          4764 => x"2e098106",
          4765 => x"8738ff17",
          4766 => x"5776ed38",
          4767 => x"79418043",
          4768 => x"8052913d",
          4769 => x"705255ff",
          4770 => x"bab33f81",
          4771 => x"dec00854",
          4772 => x"81dec008",
          4773 => x"80f73881",
          4774 => x"527451ff",
          4775 => x"bfe53f81",
          4776 => x"dec00854",
          4777 => x"81dec008",
          4778 => x"8d387680",
          4779 => x"c4386754",
          4780 => x"e5743480",
          4781 => x"c63981de",
          4782 => x"c008842e",
          4783 => x"09810680",
          4784 => x"cc388054",
          4785 => x"76742e80",
          4786 => x"c4388152",
          4787 => x"7451ffbd",
          4788 => x"b03f81de",
          4789 => x"c0085481",
          4790 => x"dec008b1",
          4791 => x"38a05381",
          4792 => x"dec00852",
          4793 => x"6751ffab",
          4794 => x"db3f6754",
          4795 => x"880b8b15",
          4796 => x"348b5378",
          4797 => x"526751ff",
          4798 => x"aba73f79",
          4799 => x"54810b83",
          4800 => x"15347951",
          4801 => x"ffadee3f",
          4802 => x"81dec008",
          4803 => x"54735574",
          4804 => x"81dec00c",
          4805 => x"9c3d0d04",
          4806 => x"f23d0d60",
          4807 => x"62028805",
          4808 => x"80cb0533",
          4809 => x"933dfc05",
          4810 => x"55725440",
          4811 => x"5e5ad2da",
          4812 => x"3f81dec0",
          4813 => x"085881de",
          4814 => x"c00882bd",
          4815 => x"38911a33",
          4816 => x"587782b5",
          4817 => x"387c802e",
          4818 => x"97388c1a",
          4819 => x"08597890",
          4820 => x"38901a33",
          4821 => x"70812a70",
          4822 => x"81065155",
          4823 => x"55739038",
          4824 => x"87548297",
          4825 => x"39825882",
          4826 => x"90398158",
          4827 => x"828b397e",
          4828 => x"8a112270",
          4829 => x"892b7055",
          4830 => x"7f545656",
          4831 => x"56fefbf7",
          4832 => x"3fff147d",
          4833 => x"06703070",
          4834 => x"72079f2a",
          4835 => x"81dec008",
          4836 => x"058c1908",
          4837 => x"7c405a5d",
          4838 => x"55558177",
          4839 => x"27883898",
          4840 => x"16087726",
          4841 => x"83388257",
          4842 => x"76775659",
          4843 => x"80567452",
          4844 => x"7951ffae",
          4845 => x"993f8115",
          4846 => x"7f555598",
          4847 => x"14087526",
          4848 => x"83388255",
          4849 => x"81dec008",
          4850 => x"812eff99",
          4851 => x"3881dec0",
          4852 => x"08ff2eff",
          4853 => x"953881de",
          4854 => x"c0088e38",
          4855 => x"81165675",
          4856 => x"7b2e0981",
          4857 => x"06873893",
          4858 => x"39745980",
          4859 => x"5674772e",
          4860 => x"098106ff",
          4861 => x"b9388758",
          4862 => x"80ff397d",
          4863 => x"802eba38",
          4864 => x"787b5555",
          4865 => x"7a802eb4",
          4866 => x"38811556",
          4867 => x"73812e09",
          4868 => x"81068338",
          4869 => x"ff567553",
          4870 => x"74527e51",
          4871 => x"ffafa83f",
          4872 => x"81dec008",
          4873 => x"5881dec0",
          4874 => x"0880ce38",
          4875 => x"748116ff",
          4876 => x"1656565c",
          4877 => x"73d33884",
          4878 => x"39ff195c",
          4879 => x"7e7c8c12",
          4880 => x"0c557d80",
          4881 => x"2eb33878",
          4882 => x"881b0c7c",
          4883 => x"8c1b0c90",
          4884 => x"1a3380c0",
          4885 => x"07547390",
          4886 => x"1b349815",
          4887 => x"08fe0590",
          4888 => x"16085754",
          4889 => x"75742691",
          4890 => x"38757b31",
          4891 => x"90160c84",
          4892 => x"15338107",
          4893 => x"54738416",
          4894 => x"34775473",
          4895 => x"81dec00c",
          4896 => x"903d0d04",
          4897 => x"e93d0d6b",
          4898 => x"6d028805",
          4899 => x"80eb0533",
          4900 => x"9d3d545a",
          4901 => x"5c59c5bd",
          4902 => x"3f8b5680",
          4903 => x"0b81dec0",
          4904 => x"08248bf8",
          4905 => x"3881dec0",
          4906 => x"08842981",
          4907 => x"dedc0570",
          4908 => x"08515574",
          4909 => x"802e8438",
          4910 => x"80753481",
          4911 => x"dec00881",
          4912 => x"ff065f81",
          4913 => x"527e51ff",
          4914 => x"a0d03f81",
          4915 => x"dec00881",
          4916 => x"ff067081",
          4917 => x"06565783",
          4918 => x"56748bc0",
          4919 => x"3876822a",
          4920 => x"70810651",
          4921 => x"558a5674",
          4922 => x"8bb23899",
          4923 => x"3dfc0553",
          4924 => x"83527e51",
          4925 => x"ffa4f03f",
          4926 => x"81dec008",
          4927 => x"99386755",
          4928 => x"74802e92",
          4929 => x"38748280",
          4930 => x"80268b38",
          4931 => x"ff157506",
          4932 => x"5574802e",
          4933 => x"83388148",
          4934 => x"78802e87",
          4935 => x"38848079",
          4936 => x"26923878",
          4937 => x"81800a26",
          4938 => x"8b38ff19",
          4939 => x"79065574",
          4940 => x"802e8638",
          4941 => x"93568ae4",
          4942 => x"3978892a",
          4943 => x"6e892a70",
          4944 => x"892b7759",
          4945 => x"4843597a",
          4946 => x"83388156",
          4947 => x"61307080",
          4948 => x"25770751",
          4949 => x"55915674",
          4950 => x"8ac23899",
          4951 => x"3df80553",
          4952 => x"81527e51",
          4953 => x"ffa4803f",
          4954 => x"815681de",
          4955 => x"c0088aac",
          4956 => x"3877832a",
          4957 => x"70770681",
          4958 => x"dec00843",
          4959 => x"56457483",
          4960 => x"38bf4166",
          4961 => x"558e5660",
          4962 => x"75268a90",
          4963 => x"38746131",
          4964 => x"70485580",
          4965 => x"ff75278a",
          4966 => x"83389356",
          4967 => x"78818026",
          4968 => x"89fa3877",
          4969 => x"812a7081",
          4970 => x"06564374",
          4971 => x"802e9538",
          4972 => x"77870655",
          4973 => x"74822e83",
          4974 => x"8d387781",
          4975 => x"06557480",
          4976 => x"2e838338",
          4977 => x"77810655",
          4978 => x"9356825e",
          4979 => x"74802e89",
          4980 => x"cb38785a",
          4981 => x"7d832e09",
          4982 => x"810680e1",
          4983 => x"3878ae38",
          4984 => x"66912a57",
          4985 => x"810b81ce",
          4986 => x"d822565a",
          4987 => x"74802e9d",
          4988 => x"38747726",
          4989 => x"983881ce",
          4990 => x"d8567910",
          4991 => x"82177022",
          4992 => x"57575a74",
          4993 => x"802e8638",
          4994 => x"767527ee",
          4995 => x"38795266",
          4996 => x"51fef6e3",
          4997 => x"3f81dec0",
          4998 => x"08842984",
          4999 => x"87057089",
          5000 => x"2a5e55a0",
          5001 => x"5c800b81",
          5002 => x"dec008fc",
          5003 => x"808a0556",
          5004 => x"44fdfff0",
          5005 => x"0a752780",
          5006 => x"ec3888d3",
          5007 => x"3978ae38",
          5008 => x"668c2a57",
          5009 => x"810b81ce",
          5010 => x"c822565a",
          5011 => x"74802e9d",
          5012 => x"38747726",
          5013 => x"983881ce",
          5014 => x"c8567910",
          5015 => x"82177022",
          5016 => x"57575a74",
          5017 => x"802e8638",
          5018 => x"767527ee",
          5019 => x"38795266",
          5020 => x"51fef683",
          5021 => x"3f81dec0",
          5022 => x"08108405",
          5023 => x"5781dec0",
          5024 => x"089ff526",
          5025 => x"9638810b",
          5026 => x"81dec008",
          5027 => x"1081dec0",
          5028 => x"08057111",
          5029 => x"722a8305",
          5030 => x"59565e83",
          5031 => x"ff17892a",
          5032 => x"5d815ca0",
          5033 => x"44601c7d",
          5034 => x"11650569",
          5035 => x"7012ff05",
          5036 => x"71307072",
          5037 => x"0674315c",
          5038 => x"52595759",
          5039 => x"407d832e",
          5040 => x"09810689",
          5041 => x"38761c60",
          5042 => x"18415c84",
          5043 => x"39761d5d",
          5044 => x"79902918",
          5045 => x"70623168",
          5046 => x"58515574",
          5047 => x"762687af",
          5048 => x"38757c31",
          5049 => x"7d317a53",
          5050 => x"70653152",
          5051 => x"55fef587",
          5052 => x"3f81dec0",
          5053 => x"08587d83",
          5054 => x"2e098106",
          5055 => x"9b3881de",
          5056 => x"c00883ff",
          5057 => x"f52680dd",
          5058 => x"38788783",
          5059 => x"3879812a",
          5060 => x"5978fdbe",
          5061 => x"3886f839",
          5062 => x"7d822e09",
          5063 => x"810680c5",
          5064 => x"3883fff5",
          5065 => x"0b81dec0",
          5066 => x"0827a038",
          5067 => x"788f3879",
          5068 => x"1a557480",
          5069 => x"c0268638",
          5070 => x"7459fd96",
          5071 => x"39628106",
          5072 => x"5574802e",
          5073 => x"8f38835e",
          5074 => x"fd883981",
          5075 => x"dec0089f",
          5076 => x"f5269238",
          5077 => x"7886b838",
          5078 => x"791a5981",
          5079 => x"807927fc",
          5080 => x"f13886ab",
          5081 => x"3980557d",
          5082 => x"812e0981",
          5083 => x"0683387d",
          5084 => x"559ff578",
          5085 => x"278b3874",
          5086 => x"8106558e",
          5087 => x"5674869c",
          5088 => x"38848053",
          5089 => x"80527a51",
          5090 => x"ffa2b93f",
          5091 => x"8b5381cc",
          5092 => x"f0527a51",
          5093 => x"ffa28a3f",
          5094 => x"8480528b",
          5095 => x"1b51ffa1",
          5096 => x"b33f798d",
          5097 => x"1c347b83",
          5098 => x"ffff0652",
          5099 => x"8e1b51ff",
          5100 => x"a1a23f81",
          5101 => x"0b901c34",
          5102 => x"7d833270",
          5103 => x"3070962a",
          5104 => x"84800654",
          5105 => x"5155911b",
          5106 => x"51ffa188",
          5107 => x"3f665574",
          5108 => x"83ffff26",
          5109 => x"90387483",
          5110 => x"ffff0652",
          5111 => x"931b51ff",
          5112 => x"a0f23f8a",
          5113 => x"397452a0",
          5114 => x"1b51ffa1",
          5115 => x"853ff80b",
          5116 => x"951c34bf",
          5117 => x"52981b51",
          5118 => x"ffa0d93f",
          5119 => x"81ff529a",
          5120 => x"1b51ffa0",
          5121 => x"cf3f6052",
          5122 => x"9c1b51ff",
          5123 => x"a0e43f7d",
          5124 => x"832e0981",
          5125 => x"0680cb38",
          5126 => x"8288b20a",
          5127 => x"5280c31b",
          5128 => x"51ffa0ce",
          5129 => x"3f7c52a4",
          5130 => x"1b51ffa0",
          5131 => x"c53f8252",
          5132 => x"ac1b51ff",
          5133 => x"a0bc3f81",
          5134 => x"52b01b51",
          5135 => x"ffa0953f",
          5136 => x"8652b21b",
          5137 => x"51ffa08c",
          5138 => x"3fff800b",
          5139 => x"80c01c34",
          5140 => x"a90b80c2",
          5141 => x"1c349353",
          5142 => x"81ccfc52",
          5143 => x"80c71b51",
          5144 => x"ae398288",
          5145 => x"b20a52a7",
          5146 => x"1b51ffa0",
          5147 => x"853f7c83",
          5148 => x"ffff0652",
          5149 => x"961b51ff",
          5150 => x"9fda3fff",
          5151 => x"800ba41c",
          5152 => x"34a90ba6",
          5153 => x"1c349353",
          5154 => x"81cd9052",
          5155 => x"ab1b51ff",
          5156 => x"a08f3f82",
          5157 => x"d4d55283",
          5158 => x"fe1b7052",
          5159 => x"59ff9fb4",
          5160 => x"3f815460",
          5161 => x"537a527e",
          5162 => x"51ff9bd7",
          5163 => x"3f815681",
          5164 => x"dec00883",
          5165 => x"e7387d83",
          5166 => x"2e098106",
          5167 => x"80ee3875",
          5168 => x"54608605",
          5169 => x"537a527e",
          5170 => x"51ff9bb7",
          5171 => x"3f848053",
          5172 => x"80527a51",
          5173 => x"ff9fed3f",
          5174 => x"848b85a4",
          5175 => x"d2527a51",
          5176 => x"ff9f8f3f",
          5177 => x"868a85e4",
          5178 => x"f25283e4",
          5179 => x"1b51ff9f",
          5180 => x"813fff18",
          5181 => x"5283e81b",
          5182 => x"51ff9ef6",
          5183 => x"3f825283",
          5184 => x"ec1b51ff",
          5185 => x"9eec3f82",
          5186 => x"d4d55278",
          5187 => x"51ff9ec4",
          5188 => x"3f755460",
          5189 => x"8705537a",
          5190 => x"527e51ff",
          5191 => x"9ae53f75",
          5192 => x"54601653",
          5193 => x"7a527e51",
          5194 => x"ff9ad83f",
          5195 => x"65538052",
          5196 => x"7a51ff9f",
          5197 => x"8f3f7f56",
          5198 => x"80587d83",
          5199 => x"2e098106",
          5200 => x"9a38f852",
          5201 => x"7a51ff9e",
          5202 => x"a93fff52",
          5203 => x"841b51ff",
          5204 => x"9ea03ff0",
          5205 => x"0a52881b",
          5206 => x"51913987",
          5207 => x"fffff855",
          5208 => x"7d812e83",
          5209 => x"38f85574",
          5210 => x"527a51ff",
          5211 => x"9e843f7c",
          5212 => x"55615774",
          5213 => x"62268338",
          5214 => x"74577654",
          5215 => x"75537a52",
          5216 => x"7e51ff99",
          5217 => x"fe3f81de",
          5218 => x"c0088287",
          5219 => x"38848053",
          5220 => x"81dec008",
          5221 => x"527a51ff",
          5222 => x"9eaa3f76",
          5223 => x"16757831",
          5224 => x"565674cd",
          5225 => x"38811858",
          5226 => x"77802eff",
          5227 => x"8d387955",
          5228 => x"7d832e83",
          5229 => x"38635561",
          5230 => x"57746226",
          5231 => x"83387457",
          5232 => x"76547553",
          5233 => x"7a527e51",
          5234 => x"ff99b83f",
          5235 => x"81dec008",
          5236 => x"81c13876",
          5237 => x"16757831",
          5238 => x"565674db",
          5239 => x"388c567d",
          5240 => x"832e9338",
          5241 => x"86566683",
          5242 => x"ffff268a",
          5243 => x"3884567d",
          5244 => x"822e8338",
          5245 => x"81566481",
          5246 => x"06587780",
          5247 => x"fe388480",
          5248 => x"5377527a",
          5249 => x"51ff9dbc",
          5250 => x"3f82d4d5",
          5251 => x"527851ff",
          5252 => x"9cc23f83",
          5253 => x"be1b5577",
          5254 => x"7534810b",
          5255 => x"81163481",
          5256 => x"0b821634",
          5257 => x"77831634",
          5258 => x"75841634",
          5259 => x"60670556",
          5260 => x"80fdc152",
          5261 => x"7551feee",
          5262 => x"be3ffe0b",
          5263 => x"85163481",
          5264 => x"dec00882",
          5265 => x"2abf0756",
          5266 => x"75861634",
          5267 => x"81dec008",
          5268 => x"87163460",
          5269 => x"5283c61b",
          5270 => x"51ff9c96",
          5271 => x"3f665283",
          5272 => x"ca1b51ff",
          5273 => x"9c8c3f81",
          5274 => x"5477537a",
          5275 => x"527e51ff",
          5276 => x"98913f81",
          5277 => x"5681dec0",
          5278 => x"08a23880",
          5279 => x"5380527e",
          5280 => x"51ff99e3",
          5281 => x"3f815681",
          5282 => x"dec00890",
          5283 => x"3889398e",
          5284 => x"568a3981",
          5285 => x"56863981",
          5286 => x"dec00856",
          5287 => x"7581dec0",
          5288 => x"0c993d0d",
          5289 => x"04f53d0d",
          5290 => x"7d605b59",
          5291 => x"807960ff",
          5292 => x"055a5757",
          5293 => x"767825b4",
          5294 => x"388d3df8",
          5295 => x"11555581",
          5296 => x"53fc1552",
          5297 => x"7951c9dc",
          5298 => x"3f7a812e",
          5299 => x"0981069c",
          5300 => x"388c3d33",
          5301 => x"55748d2e",
          5302 => x"db387476",
          5303 => x"70810558",
          5304 => x"34811757",
          5305 => x"748a2e09",
          5306 => x"8106c938",
          5307 => x"80763478",
          5308 => x"55768338",
          5309 => x"76557481",
          5310 => x"dec00c8d",
          5311 => x"3d0d04ff",
          5312 => x"3d0d7352",
          5313 => x"71932681",
          5314 => x"8e387184",
          5315 => x"2981c694",
          5316 => x"05527108",
          5317 => x"0481cff0",
          5318 => x"51818039",
          5319 => x"81cffc51",
          5320 => x"80f93981",
          5321 => x"d0905180",
          5322 => x"f23981d0",
          5323 => x"a45180eb",
          5324 => x"3981d0b4",
          5325 => x"5180e439",
          5326 => x"81d0c451",
          5327 => x"80dd3981",
          5328 => x"d0d85180",
          5329 => x"d63981d0",
          5330 => x"e85180cf",
          5331 => x"3981d180",
          5332 => x"5180c839",
          5333 => x"81d19851",
          5334 => x"80c13981",
          5335 => x"d1b051bb",
          5336 => x"3981d1cc",
          5337 => x"51b53981",
          5338 => x"d1e051af",
          5339 => x"3981d28c",
          5340 => x"51a93981",
          5341 => x"d2a051a3",
          5342 => x"3981d2c0",
          5343 => x"519d3981",
          5344 => x"d2d45197",
          5345 => x"3981d2ec",
          5346 => x"51913981",
          5347 => x"d384518b",
          5348 => x"3981d39c",
          5349 => x"51853981",
          5350 => x"d3a851ff",
          5351 => x"87a13f83",
          5352 => x"3d0d04fb",
          5353 => x"3d0d7779",
          5354 => x"56567487",
          5355 => x"e7268a38",
          5356 => x"74527587",
          5357 => x"e8295191",
          5358 => x"3987e852",
          5359 => x"7451feeb",
          5360 => x"b63f81de",
          5361 => x"c0085275",
          5362 => x"51feebab",
          5363 => x"3f81dec0",
          5364 => x"08547953",
          5365 => x"755281d3",
          5366 => x"b851ff8c",
          5367 => x"c63f873d",
          5368 => x"0d04f53d",
          5369 => x"0d7d7f61",
          5370 => x"028c0580",
          5371 => x"c7053373",
          5372 => x"7315665f",
          5373 => x"5d5a5a5c",
          5374 => x"5c5c7852",
          5375 => x"81d3dc51",
          5376 => x"ff8ca03f",
          5377 => x"81d3e451",
          5378 => x"ff86b43f",
          5379 => x"80557477",
          5380 => x"2780fc38",
          5381 => x"79902e89",
          5382 => x"3879a02e",
          5383 => x"a73880c6",
          5384 => x"39741653",
          5385 => x"7278278e",
          5386 => x"38722252",
          5387 => x"81d3e851",
          5388 => x"ff8bf03f",
          5389 => x"893981d3",
          5390 => x"f451ff86",
          5391 => x"823f8215",
          5392 => x"5580c339",
          5393 => x"74165372",
          5394 => x"78278e38",
          5395 => x"72085281",
          5396 => x"d3dc51ff",
          5397 => x"8bcd3f89",
          5398 => x"3981d3f0",
          5399 => x"51ff85df",
          5400 => x"3f841555",
          5401 => x"a1397416",
          5402 => x"53727827",
          5403 => x"8e387233",
          5404 => x"5281d3fc",
          5405 => x"51ff8bab",
          5406 => x"3f893981",
          5407 => x"d48451ff",
          5408 => x"85bd3f81",
          5409 => x"1555a051",
          5410 => x"fef6af3f",
          5411 => x"ff803981",
          5412 => x"d48851ff",
          5413 => x"85a93f80",
          5414 => x"55747727",
          5415 => x"aa387416",
          5416 => x"70337972",
          5417 => x"26525553",
          5418 => x"9f742790",
          5419 => x"3872802e",
          5420 => x"8b387380",
          5421 => x"fe268538",
          5422 => x"73518339",
          5423 => x"a051fef5",
          5424 => x"f93f8115",
          5425 => x"55d33981",
          5426 => x"d48c51ff",
          5427 => x"84f13f76",
          5428 => x"16771a5a",
          5429 => x"56fef9b4",
          5430 => x"3f81dec0",
          5431 => x"08982b70",
          5432 => x"982c5155",
          5433 => x"74a02e09",
          5434 => x"8106a538",
          5435 => x"fef99d3f",
          5436 => x"81dec008",
          5437 => x"982b7098",
          5438 => x"2c70a032",
          5439 => x"70307072",
          5440 => x"079f2a51",
          5441 => x"56565155",
          5442 => x"749b2e8c",
          5443 => x"3872dd38",
          5444 => x"749b2e09",
          5445 => x"81068538",
          5446 => x"80538c39",
          5447 => x"7a1c5372",
          5448 => x"7626fdd6",
          5449 => x"38ff5372",
          5450 => x"81dec00c",
          5451 => x"8d3d0d04",
          5452 => x"ec3d0d66",
          5453 => x"02840580",
          5454 => x"e3053369",
          5455 => x"72307074",
          5456 => x"07802570",
          5457 => x"87ff7427",
          5458 => x"07515158",
          5459 => x"5a5b5693",
          5460 => x"577480fc",
          5461 => x"38815375",
          5462 => x"528c3d70",
          5463 => x"5257ffbf",
          5464 => x"de3f81de",
          5465 => x"c0085681",
          5466 => x"dec008b8",
          5467 => x"3881dec0",
          5468 => x"0887c098",
          5469 => x"880c81de",
          5470 => x"c0085996",
          5471 => x"3dd40554",
          5472 => x"84805377",
          5473 => x"527651c4",
          5474 => x"9b3f81de",
          5475 => x"c0085681",
          5476 => x"dec00890",
          5477 => x"387a5574",
          5478 => x"802e8938",
          5479 => x"74197519",
          5480 => x"5959d839",
          5481 => x"963dd805",
          5482 => x"51cc853f",
          5483 => x"75307077",
          5484 => x"07802551",
          5485 => x"5579802e",
          5486 => x"95387480",
          5487 => x"2e903881",
          5488 => x"d4905387",
          5489 => x"c0988808",
          5490 => x"527851fb",
          5491 => x"d63f7557",
          5492 => x"7681dec0",
          5493 => x"0c963d0d",
          5494 => x"04f93d0d",
          5495 => x"7b028405",
          5496 => x"b3053357",
          5497 => x"58ff5780",
          5498 => x"537a5279",
          5499 => x"51fec13f",
          5500 => x"81dec008",
          5501 => x"a4387580",
          5502 => x"2e883875",
          5503 => x"812e9838",
          5504 => x"98396055",
          5505 => x"7f5481de",
          5506 => x"c0537e52",
          5507 => x"7d51772d",
          5508 => x"81dec008",
          5509 => x"57833977",
          5510 => x"047681de",
          5511 => x"c00c893d",
          5512 => x"0d04fc3d",
          5513 => x"0d029b05",
          5514 => x"3381d498",
          5515 => x"5381d4a0",
          5516 => x"5255ff87",
          5517 => x"ee3f81db",
          5518 => x"c02251ff",
          5519 => x"80893f81",
          5520 => x"d4ac5481",
          5521 => x"d4b85381",
          5522 => x"dbc13352",
          5523 => x"81d4c051",
          5524 => x"ff87d03f",
          5525 => x"74802e85",
          5526 => x"38fefbd4",
          5527 => x"3f863d0d",
          5528 => x"04fe3d0d",
          5529 => x"87c09680",
          5530 => x"0853ff80",
          5531 => x"a23f8151",
          5532 => x"fef2ad3f",
          5533 => x"81d4dc51",
          5534 => x"fef4a53f",
          5535 => x"8051fef2",
          5536 => x"9f3f7281",
          5537 => x"2a708106",
          5538 => x"51527180",
          5539 => x"2e953881",
          5540 => x"51fef28c",
          5541 => x"3f81d4f8",
          5542 => x"51fef484",
          5543 => x"3f8051fe",
          5544 => x"f1fe3f72",
          5545 => x"822a7081",
          5546 => x"06515271",
          5547 => x"802e9538",
          5548 => x"8151fef1",
          5549 => x"eb3f81d5",
          5550 => x"8c51fef3",
          5551 => x"e33f8051",
          5552 => x"fef1dd3f",
          5553 => x"72832a70",
          5554 => x"81065152",
          5555 => x"71802e95",
          5556 => x"388151fe",
          5557 => x"f1ca3f81",
          5558 => x"d59c51fe",
          5559 => x"f3c23f80",
          5560 => x"51fef1bc",
          5561 => x"3f72842a",
          5562 => x"70810651",
          5563 => x"5271802e",
          5564 => x"95388151",
          5565 => x"fef1a93f",
          5566 => x"81d5b051",
          5567 => x"fef3a13f",
          5568 => x"8051fef1",
          5569 => x"9b3f7285",
          5570 => x"2a708106",
          5571 => x"51527180",
          5572 => x"2e953881",
          5573 => x"51fef188",
          5574 => x"3f81d5c4",
          5575 => x"51fef380",
          5576 => x"3f8051fe",
          5577 => x"f0fa3f72",
          5578 => x"862a7081",
          5579 => x"06515271",
          5580 => x"802e9538",
          5581 => x"8151fef0",
          5582 => x"e73f81d5",
          5583 => x"d851fef2",
          5584 => x"df3f8051",
          5585 => x"fef0d93f",
          5586 => x"72872a70",
          5587 => x"81065152",
          5588 => x"71802e95",
          5589 => x"388151fe",
          5590 => x"f0c63f81",
          5591 => x"d5ec51fe",
          5592 => x"f2be3f80",
          5593 => x"51fef0b8",
          5594 => x"3f72882a",
          5595 => x"70810651",
          5596 => x"5271802e",
          5597 => x"95388151",
          5598 => x"fef0a53f",
          5599 => x"81d68051",
          5600 => x"fef29d3f",
          5601 => x"8051fef0",
          5602 => x"973ffefe",
          5603 => x"cb3f843d",
          5604 => x"0d04fa3d",
          5605 => x"0d787008",
          5606 => x"70555557",
          5607 => x"73802e80",
          5608 => x"f0388e39",
          5609 => x"73770c85",
          5610 => x"15335380",
          5611 => x"e4398114",
          5612 => x"54807433",
          5613 => x"7081ff06",
          5614 => x"57575374",
          5615 => x"a02e8338",
          5616 => x"81537480",
          5617 => x"2e843872",
          5618 => x"e5387581",
          5619 => x"ff065372",
          5620 => x"a02e0981",
          5621 => x"06883880",
          5622 => x"74708105",
          5623 => x"56348056",
          5624 => x"75902981",
          5625 => x"dbf00577",
          5626 => x"08537008",
          5627 => x"5255feea",
          5628 => x"9e3f81de",
          5629 => x"c0088b38",
          5630 => x"84153353",
          5631 => x"72812eff",
          5632 => x"a3388116",
          5633 => x"7081ff06",
          5634 => x"57539476",
          5635 => x"27d238ff",
          5636 => x"537281de",
          5637 => x"c00c883d",
          5638 => x"0d04fb3d",
          5639 => x"0d777970",
          5640 => x"55565680",
          5641 => x"527551fe",
          5642 => x"e8d43f81",
          5643 => x"dbec3354",
          5644 => x"73a73881",
          5645 => x"5381d6c0",
          5646 => x"5281f5c4",
          5647 => x"51ffb9ff",
          5648 => x"3f81dec0",
          5649 => x"08307081",
          5650 => x"dec00807",
          5651 => x"80258271",
          5652 => x"31515154",
          5653 => x"7381dbec",
          5654 => x"3481dbec",
          5655 => x"33547381",
          5656 => x"2e098106",
          5657 => x"ac3881f5",
          5658 => x"c4537452",
          5659 => x"7551f4b5",
          5660 => x"3f81dec0",
          5661 => x"08802e8c",
          5662 => x"3881dec0",
          5663 => x"0851fefd",
          5664 => x"be3f8e39",
          5665 => x"81f5c451",
          5666 => x"c6a63f82",
          5667 => x"0b81dbec",
          5668 => x"3481dbec",
          5669 => x"33547382",
          5670 => x"2e098106",
          5671 => x"89387452",
          5672 => x"7551ff83",
          5673 => x"d83f800b",
          5674 => x"81dec00c",
          5675 => x"873d0d04",
          5676 => x"cb3d0d80",
          5677 => x"707181f5",
          5678 => x"c00c405d",
          5679 => x"81527c51",
          5680 => x"ff88d73f",
          5681 => x"81dec008",
          5682 => x"81ff0659",
          5683 => x"787d2e09",
          5684 => x"8106a238",
          5685 => x"81d6d052",
          5686 => x"993d7052",
          5687 => x"59ff82d9",
          5688 => x"3f7c5378",
          5689 => x"5281dff0",
          5690 => x"51ffb7f2",
          5691 => x"3f81dec0",
          5692 => x"087d2e88",
          5693 => x"3881d6d4",
          5694 => x"5192bc39",
          5695 => x"8170405d",
          5696 => x"81d78c51",
          5697 => x"fefcb83f",
          5698 => x"993d7046",
          5699 => x"5a80f852",
          5700 => x"7951fe86",
          5701 => x"3fb73dfe",
          5702 => x"f80551fc",
          5703 => x"f53f81de",
          5704 => x"c008902b",
          5705 => x"70902c51",
          5706 => x"597880c3",
          5707 => x"2e8ace38",
          5708 => x"7880c324",
          5709 => x"80dc3878",
          5710 => x"ab2e83bc",
          5711 => x"3878ab24",
          5712 => x"a4387882",
          5713 => x"2e81af38",
          5714 => x"7882248a",
          5715 => x"3878802e",
          5716 => x"ffae388f",
          5717 => x"de397884",
          5718 => x"2e828238",
          5719 => x"78942e82",
          5720 => x"ad388fcf",
          5721 => x"397880c0",
          5722 => x"2e858738",
          5723 => x"7880c024",
          5724 => x"903878b0",
          5725 => x"2e83a938",
          5726 => x"78bc2e84",
          5727 => x"8b388fb3",
          5728 => x"397880c1",
          5729 => x"2e879e38",
          5730 => x"7880c22e",
          5731 => x"88bf388f",
          5732 => x"a2397880",
          5733 => x"d52e8df3",
          5734 => x"387880d5",
          5735 => x"24a93878",
          5736 => x"80d02e8d",
          5737 => x"a7387880",
          5738 => x"d0248b38",
          5739 => x"7880c52e",
          5740 => x"8aeb388e",
          5741 => x"fe397880",
          5742 => x"d12e8da1",
          5743 => x"387880d4",
          5744 => x"2e8dab38",
          5745 => x"8eed3978",
          5746 => x"81822e8e",
          5747 => x"c3387881",
          5748 => x"82249238",
          5749 => x"7880f82e",
          5750 => x"8dce3878",
          5751 => x"80f92e8d",
          5752 => x"ec388ecf",
          5753 => x"39788183",
          5754 => x"2e8eb438",
          5755 => x"7881852e",
          5756 => x"8eba388e",
          5757 => x"be39b73d",
          5758 => x"fef41153",
          5759 => x"fef80551",
          5760 => x"ff82953f",
          5761 => x"81dec008",
          5762 => x"883881d7",
          5763 => x"905190a7",
          5764 => x"39b73dfe",
          5765 => x"f01153fe",
          5766 => x"f80551ff",
          5767 => x"81fa3f81",
          5768 => x"dec00880",
          5769 => x"2e883881",
          5770 => x"63258338",
          5771 => x"80430280",
          5772 => x"cb053352",
          5773 => x"0280cf05",
          5774 => x"3351ff85",
          5775 => x"dd3f81de",
          5776 => x"c00881ff",
          5777 => x"0659788e",
          5778 => x"3881d7a0",
          5779 => x"51fef9ef",
          5780 => x"3f815ffd",
          5781 => x"ab3981d7",
          5782 => x"b0518ca8",
          5783 => x"39b73dfe",
          5784 => x"f41153fe",
          5785 => x"f80551ff",
          5786 => x"81ae3f81",
          5787 => x"dec00880",
          5788 => x"2efd8d38",
          5789 => x"80538052",
          5790 => x"0280cf05",
          5791 => x"3351ff89",
          5792 => x"e63f81de",
          5793 => x"c0085281",
          5794 => x"d7c8518c",
          5795 => x"fc39b73d",
          5796 => x"fef41153",
          5797 => x"fef80551",
          5798 => x"ff80fd3f",
          5799 => x"81dec008",
          5800 => x"802e8738",
          5801 => x"638926fc",
          5802 => x"d738b73d",
          5803 => x"fef01153",
          5804 => x"fef80551",
          5805 => x"ff80e13f",
          5806 => x"81dec008",
          5807 => x"863881de",
          5808 => x"c0084363",
          5809 => x"5381d7d0",
          5810 => x"527951fe",
          5811 => x"feeb3f02",
          5812 => x"80cb0533",
          5813 => x"53795263",
          5814 => x"84b42981",
          5815 => x"dff00551",
          5816 => x"ffb3fb3f",
          5817 => x"81dec008",
          5818 => x"81933881",
          5819 => x"d7a051fe",
          5820 => x"f8cd3f81",
          5821 => x"5dfc8939",
          5822 => x"b73dfef8",
          5823 => x"0551fee5",
          5824 => x"d03f81de",
          5825 => x"c008b83d",
          5826 => x"fef80552",
          5827 => x"5bfee6a3",
          5828 => x"3f815381",
          5829 => x"dec00852",
          5830 => x"7a51f494",
          5831 => x"3f80d539",
          5832 => x"b73dfef8",
          5833 => x"0551fee5",
          5834 => x"a83f81de",
          5835 => x"c008b83d",
          5836 => x"fef80552",
          5837 => x"5bfee5fb",
          5838 => x"3f81dec0",
          5839 => x"08b83dfe",
          5840 => x"f805525a",
          5841 => x"fee5ec3f",
          5842 => x"81dec008",
          5843 => x"b83dfef8",
          5844 => x"055259fe",
          5845 => x"e5dd3f81",
          5846 => x"db8c5881",
          5847 => x"def45780",
          5848 => x"56805581",
          5849 => x"dec00881",
          5850 => x"ff065478",
          5851 => x"5379527a",
          5852 => x"51f4e63f",
          5853 => x"81dec008",
          5854 => x"802efb84",
          5855 => x"3881dec0",
          5856 => x"0851eefb",
          5857 => x"3ffaf939",
          5858 => x"b73dfef4",
          5859 => x"1153fef8",
          5860 => x"0551feff",
          5861 => x"833f81de",
          5862 => x"c008802e",
          5863 => x"fae238b7",
          5864 => x"3dfef011",
          5865 => x"53fef805",
          5866 => x"51fefeec",
          5867 => x"3f81dec0",
          5868 => x"08802efa",
          5869 => x"cb38b73d",
          5870 => x"feec1153",
          5871 => x"fef80551",
          5872 => x"fefed53f",
          5873 => x"81dec008",
          5874 => x"863881de",
          5875 => x"c0084281",
          5876 => x"d7d451fe",
          5877 => x"f6e93f63",
          5878 => x"635c5a79",
          5879 => x"7b2788e6",
          5880 => x"38615978",
          5881 => x"7a708405",
          5882 => x"5c0c7a7a",
          5883 => x"26f53888",
          5884 => x"d539b73d",
          5885 => x"fef41153",
          5886 => x"fef80551",
          5887 => x"fefe993f",
          5888 => x"81dec008",
          5889 => x"80df3881",
          5890 => x"dbd43359",
          5891 => x"78802e89",
          5892 => x"3881db8c",
          5893 => x"084480cd",
          5894 => x"3981dbd5",
          5895 => x"33597880",
          5896 => x"2e883881",
          5897 => x"db940844",
          5898 => x"bc3981db",
          5899 => x"d6335978",
          5900 => x"802e8838",
          5901 => x"81db9c08",
          5902 => x"44ab3981",
          5903 => x"dbd73359",
          5904 => x"78802e88",
          5905 => x"3881dba4",
          5906 => x"08449a39",
          5907 => x"81dbd233",
          5908 => x"5978802e",
          5909 => x"883881db",
          5910 => x"ac084489",
          5911 => x"3981dbbc",
          5912 => x"08fc8005",
          5913 => x"44b73dfe",
          5914 => x"f01153fe",
          5915 => x"f80551fe",
          5916 => x"fda63f81",
          5917 => x"dec00880",
          5918 => x"de3881db",
          5919 => x"d4335978",
          5920 => x"802e8938",
          5921 => x"81db9008",
          5922 => x"4380cc39",
          5923 => x"81dbd533",
          5924 => x"5978802e",
          5925 => x"883881db",
          5926 => x"980843bb",
          5927 => x"3981dbd6",
          5928 => x"33597880",
          5929 => x"2e883881",
          5930 => x"dba00843",
          5931 => x"aa3981db",
          5932 => x"d7335978",
          5933 => x"802e8838",
          5934 => x"81dba808",
          5935 => x"43993981",
          5936 => x"dbd23359",
          5937 => x"78802e88",
          5938 => x"3881dbb0",
          5939 => x"08438839",
          5940 => x"81dbbc08",
          5941 => x"880543b7",
          5942 => x"3dfeec11",
          5943 => x"53fef805",
          5944 => x"51fefcb4",
          5945 => x"3f81dec0",
          5946 => x"08802e9b",
          5947 => x"3880625b",
          5948 => x"5979882e",
          5949 => x"83388159",
          5950 => x"79902e8d",
          5951 => x"3878802e",
          5952 => x"883879a0",
          5953 => x"2e833888",
          5954 => x"4281d7e4",
          5955 => x"51fef4af",
          5956 => x"3fa05563",
          5957 => x"54615362",
          5958 => x"526351ed",
          5959 => x"c53f81d7",
          5960 => x"f45186e0",
          5961 => x"39b73dfe",
          5962 => x"f41153fe",
          5963 => x"f80551fe",
          5964 => x"fbe63f81",
          5965 => x"dec00880",
          5966 => x"2ef7c538",
          5967 => x"b73dfef0",
          5968 => x"1153fef8",
          5969 => x"0551fefb",
          5970 => x"cf3f81de",
          5971 => x"c008802e",
          5972 => x"a5386359",
          5973 => x"0280cb05",
          5974 => x"33793463",
          5975 => x"810544b7",
          5976 => x"3dfef011",
          5977 => x"53fef805",
          5978 => x"51fefbac",
          5979 => x"3f81dec0",
          5980 => x"08e038f7",
          5981 => x"8b396370",
          5982 => x"33545281",
          5983 => x"d88051fe",
          5984 => x"f9a13f80",
          5985 => x"f8527951",
          5986 => x"fef9f23f",
          5987 => x"79457933",
          5988 => x"5978ae2e",
          5989 => x"f6ea389f",
          5990 => x"7927a038",
          5991 => x"b73dfef0",
          5992 => x"1153fef8",
          5993 => x"0551fefa",
          5994 => x"ef3f81de",
          5995 => x"c008802e",
          5996 => x"91386359",
          5997 => x"0280cb05",
          5998 => x"33793463",
          5999 => x"810544ff",
          6000 => x"b53981d8",
          6001 => x"8c51fef2",
          6002 => x"f63fffaa",
          6003 => x"39b73dfe",
          6004 => x"e81153fe",
          6005 => x"f80551fe",
          6006 => x"fcb03f81",
          6007 => x"dec00880",
          6008 => x"2ef69d38",
          6009 => x"b73dfee4",
          6010 => x"1153fef8",
          6011 => x"0551fefc",
          6012 => x"993f81de",
          6013 => x"c008802e",
          6014 => x"a6386059",
          6015 => x"02be0522",
          6016 => x"79708205",
          6017 => x"5b237841",
          6018 => x"b73dfee4",
          6019 => x"1153fef8",
          6020 => x"0551fefb",
          6021 => x"f53f81de",
          6022 => x"c008df38",
          6023 => x"f5e23960",
          6024 => x"70225452",
          6025 => x"81d89451",
          6026 => x"fef7f83f",
          6027 => x"80f85279",
          6028 => x"51fef8c9",
          6029 => x"3f794579",
          6030 => x"335978ae",
          6031 => x"2ef5c138",
          6032 => x"789f2687",
          6033 => x"38608205",
          6034 => x"41d539b7",
          6035 => x"3dfee411",
          6036 => x"53fef805",
          6037 => x"51fefbb2",
          6038 => x"3f81dec0",
          6039 => x"08802e92",
          6040 => x"38605902",
          6041 => x"be052279",
          6042 => x"7082055b",
          6043 => x"237841ff",
          6044 => x"ae3981d8",
          6045 => x"8c51fef1",
          6046 => x"c63fffa3",
          6047 => x"39b73dfe",
          6048 => x"e81153fe",
          6049 => x"f80551fe",
          6050 => x"fb803f81",
          6051 => x"dec00880",
          6052 => x"2ef4ed38",
          6053 => x"b73dfee4",
          6054 => x"1153fef8",
          6055 => x"0551fefa",
          6056 => x"e93f81de",
          6057 => x"c008802e",
          6058 => x"a1386060",
          6059 => x"710c5960",
          6060 => x"840541b7",
          6061 => x"3dfee411",
          6062 => x"53fef805",
          6063 => x"51fefaca",
          6064 => x"3f81dec0",
          6065 => x"08e438f4",
          6066 => x"b7396070",
          6067 => x"08545281",
          6068 => x"d8a051fe",
          6069 => x"f6cd3f80",
          6070 => x"f8527951",
          6071 => x"fef79e3f",
          6072 => x"79457933",
          6073 => x"5978ae2e",
          6074 => x"f496389f",
          6075 => x"79279c38",
          6076 => x"b73dfee4",
          6077 => x"1153fef8",
          6078 => x"0551fefa",
          6079 => x"8d3f81de",
          6080 => x"c008802e",
          6081 => x"8d386060",
          6082 => x"710c5960",
          6083 => x"840541ff",
          6084 => x"b93981d8",
          6085 => x"8c51fef0",
          6086 => x"a63fffae",
          6087 => x"39b73dfe",
          6088 => x"f41153fe",
          6089 => x"f80551fe",
          6090 => x"f7ee3f81",
          6091 => x"dec00880",
          6092 => x"df3881db",
          6093 => x"d4335978",
          6094 => x"802e8938",
          6095 => x"81db8c08",
          6096 => x"4480cd39",
          6097 => x"81dbd533",
          6098 => x"5978802e",
          6099 => x"883881db",
          6100 => x"940844bc",
          6101 => x"3981dbd6",
          6102 => x"33597880",
          6103 => x"2e883881",
          6104 => x"db9c0844",
          6105 => x"ab3981db",
          6106 => x"d7335978",
          6107 => x"802e8838",
          6108 => x"81dba408",
          6109 => x"449a3981",
          6110 => x"dbd23359",
          6111 => x"78802e88",
          6112 => x"3881dbac",
          6113 => x"08448939",
          6114 => x"81dbbc08",
          6115 => x"fc800544",
          6116 => x"b73dfef0",
          6117 => x"1153fef8",
          6118 => x"0551fef6",
          6119 => x"fb3f81de",
          6120 => x"c00880de",
          6121 => x"3881dbd4",
          6122 => x"33597880",
          6123 => x"2e893881",
          6124 => x"db900843",
          6125 => x"80cc3981",
          6126 => x"dbd53359",
          6127 => x"78802e88",
          6128 => x"3881db98",
          6129 => x"0843bb39",
          6130 => x"81dbd633",
          6131 => x"5978802e",
          6132 => x"883881db",
          6133 => x"a00843aa",
          6134 => x"3981dbd7",
          6135 => x"33597880",
          6136 => x"2e883881",
          6137 => x"dba80843",
          6138 => x"993981db",
          6139 => x"d2335978",
          6140 => x"802e8838",
          6141 => x"81dbb008",
          6142 => x"43883981",
          6143 => x"dbbc0888",
          6144 => x"0543b73d",
          6145 => x"feec1153",
          6146 => x"fef80551",
          6147 => x"fef6893f",
          6148 => x"81dec008",
          6149 => x"863881de",
          6150 => x"c0084281",
          6151 => x"d8ac51fe",
          6152 => x"ee9d3f63",
          6153 => x"5a796327",
          6154 => x"9d387908",
          6155 => x"5978622e",
          6156 => x"0981068d",
          6157 => x"38785379",
          6158 => x"5281d8bc",
          6159 => x"51fef3e3",
          6160 => x"3f841a5a",
          6161 => x"e03981d7",
          6162 => x"9c51b939",
          6163 => x"81d8cc51",
          6164 => x"feedec3f",
          6165 => x"8251feec",
          6166 => x"da3ff1a4",
          6167 => x"3981d8e4",
          6168 => x"51feeddb",
          6169 => x"3fa251fe",
          6170 => x"ecad3ff1",
          6171 => x"93398480",
          6172 => x"810b87c0",
          6173 => x"94840c84",
          6174 => x"80810b87",
          6175 => x"c094940c",
          6176 => x"81d8fc51",
          6177 => x"feedb83f",
          6178 => x"f0f63981",
          6179 => x"d99051fe",
          6180 => x"edad3f8c",
          6181 => x"80830b87",
          6182 => x"c094840c",
          6183 => x"8c80830b",
          6184 => x"87c09494",
          6185 => x"0cf0d939",
          6186 => x"b73dfef4",
          6187 => x"1153fef8",
          6188 => x"0551fef4",
          6189 => x"e33f81de",
          6190 => x"c008802e",
          6191 => x"f0c23863",
          6192 => x"5281d9a4",
          6193 => x"51fef2db",
          6194 => x"3f635978",
          6195 => x"04b73dfe",
          6196 => x"f41153fe",
          6197 => x"f80551fe",
          6198 => x"f4be3f81",
          6199 => x"dec00880",
          6200 => x"2ef09d38",
          6201 => x"635281d9",
          6202 => x"c051fef2",
          6203 => x"b63f6359",
          6204 => x"782d81de",
          6205 => x"c0085e81",
          6206 => x"dec00880",
          6207 => x"2ef08138",
          6208 => x"81dec008",
          6209 => x"5281d9dc",
          6210 => x"51fef297",
          6211 => x"3feff139",
          6212 => x"81d9f851",
          6213 => x"feeca83f",
          6214 => x"febde53f",
          6215 => x"efe23981",
          6216 => x"da9451fe",
          6217 => x"ec993f80",
          6218 => x"59ffa039",
          6219 => x"fee6813f",
          6220 => x"efce3964",
          6221 => x"70335159",
          6222 => x"78802eef",
          6223 => x"c3387c80",
          6224 => x"2e81dc38",
          6225 => x"81706006",
          6226 => x"5a5a7880",
          6227 => x"2e81d038",
          6228 => x"b73dfef8",
          6229 => x"0551fed8",
          6230 => x"f83f81de",
          6231 => x"c0087a5d",
          6232 => x"5b7b822e",
          6233 => x"b2387b82",
          6234 => x"2489387b",
          6235 => x"812e8c38",
          6236 => x"80cd397b",
          6237 => x"832eb038",
          6238 => x"80c53981",
          6239 => x"daa8567a",
          6240 => x"5581daac",
          6241 => x"54805381",
          6242 => x"dab052b7",
          6243 => x"3dffb005",
          6244 => x"51fef1a5",
          6245 => x"3fbb3981",
          6246 => x"dad052b7",
          6247 => x"3dffb005",
          6248 => x"51fef195",
          6249 => x"3fab397a",
          6250 => x"5581daac",
          6251 => x"54805381",
          6252 => x"dac052b7",
          6253 => x"3dffb005",
          6254 => x"51fef0fd",
          6255 => x"3f93397a",
          6256 => x"54805381",
          6257 => x"dacc52b7",
          6258 => x"3dffb005",
          6259 => x"51fef0e9",
          6260 => x"3f81db8c",
          6261 => x"5881def4",
          6262 => x"57805664",
          6263 => x"81114681",
          6264 => x"05558054",
          6265 => x"82808053",
          6266 => x"82808052",
          6267 => x"b73dffb0",
          6268 => x"0551e7e5",
          6269 => x"3f81dec0",
          6270 => x"0881dec0",
          6271 => x"08097030",
          6272 => x"70720780",
          6273 => x"25515b5b",
          6274 => x"5e7b8326",
          6275 => x"92387880",
          6276 => x"2e8d3881",
          6277 => x"1c7081ff",
          6278 => x"065d597b",
          6279 => x"fec3387e",
          6280 => x"81327d81",
          6281 => x"32075978",
          6282 => x"8a387dff",
          6283 => x"2e098106",
          6284 => x"edce3881",
          6285 => x"dad451fe",
          6286 => x"efe93fed",
          6287 => x"c339fc3d",
          6288 => x"0d800b81",
          6289 => x"def43487",
          6290 => x"c0948c70",
          6291 => x"08545587",
          6292 => x"84805272",
          6293 => x"51fece9f",
          6294 => x"3f81dec0",
          6295 => x"08902b75",
          6296 => x"08555387",
          6297 => x"84805273",
          6298 => x"51fece8b",
          6299 => x"3f7281de",
          6300 => x"c0080775",
          6301 => x"0c87c094",
          6302 => x"9c700854",
          6303 => x"55878480",
          6304 => x"527251fe",
          6305 => x"cdf13f81",
          6306 => x"dec00890",
          6307 => x"2b750855",
          6308 => x"53878480",
          6309 => x"527351fe",
          6310 => x"cddd3f72",
          6311 => x"81dec008",
          6312 => x"07750c8c",
          6313 => x"80830b87",
          6314 => x"c094840c",
          6315 => x"8c80830b",
          6316 => x"87c09494",
          6317 => x"0c9fba0b",
          6318 => x"81ded00c",
          6319 => x"a2bb0b81",
          6320 => x"ded40cfe",
          6321 => x"de9e3ffe",
          6322 => x"e7c53f81",
          6323 => x"dae451fe",
          6324 => x"dbce3f81",
          6325 => x"daf051fe",
          6326 => x"e8e53f81",
          6327 => x"ace151fe",
          6328 => x"e7a83f81",
          6329 => x"51e6bb3f",
          6330 => x"ebc63f80",
          6331 => x"04000000",
          6332 => x"00ffffff",
          6333 => x"ff00ffff",
          6334 => x"ffff00ff",
          6335 => x"ffffff00",
          6336 => x"00001661",
          6337 => x"00001667",
          6338 => x"0000166d",
          6339 => x"00001673",
          6340 => x"00001679",
          6341 => x"00005391",
          6342 => x"00005315",
          6343 => x"0000531c",
          6344 => x"00005323",
          6345 => x"0000532a",
          6346 => x"00005331",
          6347 => x"00005338",
          6348 => x"0000533f",
          6349 => x"00005346",
          6350 => x"0000534d",
          6351 => x"00005354",
          6352 => x"0000535b",
          6353 => x"00005361",
          6354 => x"00005367",
          6355 => x"0000536d",
          6356 => x"00005373",
          6357 => x"00005379",
          6358 => x"0000537f",
          6359 => x"00005385",
          6360 => x"0000538b",
          6361 => x"25642f25",
          6362 => x"642f2564",
          6363 => x"2025643a",
          6364 => x"25643a25",
          6365 => x"642e2564",
          6366 => x"25640a00",
          6367 => x"536f4320",
          6368 => x"436f6e66",
          6369 => x"69677572",
          6370 => x"6174696f",
          6371 => x"6e000000",
          6372 => x"20286672",
          6373 => x"6f6d2053",
          6374 => x"6f432063",
          6375 => x"6f6e6669",
          6376 => x"67290000",
          6377 => x"3a0a4465",
          6378 => x"76696365",
          6379 => x"7320696d",
          6380 => x"706c656d",
          6381 => x"656e7465",
          6382 => x"643a0a00",
          6383 => x"20202020",
          6384 => x"57422053",
          6385 => x"4452414d",
          6386 => x"20202825",
          6387 => x"3038583a",
          6388 => x"25303858",
          6389 => x"292e0a00",
          6390 => x"20202020",
          6391 => x"53445241",
          6392 => x"4d202020",
          6393 => x"20202825",
          6394 => x"3038583a",
          6395 => x"25303858",
          6396 => x"292e0a00",
          6397 => x"20202020",
          6398 => x"494e534e",
          6399 => x"20425241",
          6400 => x"4d202825",
          6401 => x"3038583a",
          6402 => x"25303858",
          6403 => x"292e0a00",
          6404 => x"20202020",
          6405 => x"4252414d",
          6406 => x"20202020",
          6407 => x"20202825",
          6408 => x"3038583a",
          6409 => x"25303858",
          6410 => x"292e0a00",
          6411 => x"20202020",
          6412 => x"52414d20",
          6413 => x"20202020",
          6414 => x"20202825",
          6415 => x"3038583a",
          6416 => x"25303858",
          6417 => x"292e0a00",
          6418 => x"20202020",
          6419 => x"53442043",
          6420 => x"41524420",
          6421 => x"20202844",
          6422 => x"65766963",
          6423 => x"6573203d",
          6424 => x"25303264",
          6425 => x"292e0a00",
          6426 => x"20202020",
          6427 => x"54494d45",
          6428 => x"52312020",
          6429 => x"20202854",
          6430 => x"696d6572",
          6431 => x"7320203d",
          6432 => x"25303264",
          6433 => x"292e0a00",
          6434 => x"20202020",
          6435 => x"494e5452",
          6436 => x"20435452",
          6437 => x"4c202843",
          6438 => x"68616e6e",
          6439 => x"656c733d",
          6440 => x"25303264",
          6441 => x"292e0a00",
          6442 => x"20202020",
          6443 => x"57495348",
          6444 => x"424f4e45",
          6445 => x"20425553",
          6446 => x"0a000000",
          6447 => x"20202020",
          6448 => x"57422049",
          6449 => x"32430a00",
          6450 => x"20202020",
          6451 => x"494f4354",
          6452 => x"4c0a0000",
          6453 => x"20202020",
          6454 => x"5053320a",
          6455 => x"00000000",
          6456 => x"20202020",
          6457 => x"5350490a",
          6458 => x"00000000",
          6459 => x"41646472",
          6460 => x"65737365",
          6461 => x"733a0a00",
          6462 => x"20202020",
          6463 => x"43505520",
          6464 => x"52657365",
          6465 => x"74205665",
          6466 => x"63746f72",
          6467 => x"20416464",
          6468 => x"72657373",
          6469 => x"203d2025",
          6470 => x"3038580a",
          6471 => x"00000000",
          6472 => x"20202020",
          6473 => x"43505520",
          6474 => x"4d656d6f",
          6475 => x"72792053",
          6476 => x"74617274",
          6477 => x"20416464",
          6478 => x"72657373",
          6479 => x"203d2025",
          6480 => x"3038580a",
          6481 => x"00000000",
          6482 => x"20202020",
          6483 => x"53746163",
          6484 => x"6b205374",
          6485 => x"61727420",
          6486 => x"41646472",
          6487 => x"65737320",
          6488 => x"20202020",
          6489 => x"203d2025",
          6490 => x"3038580a",
          6491 => x"00000000",
          6492 => x"4d697363",
          6493 => x"3a0a0000",
          6494 => x"20202020",
          6495 => x"5a505520",
          6496 => x"49642020",
          6497 => x"20202020",
          6498 => x"20202020",
          6499 => x"20202020",
          6500 => x"20202020",
          6501 => x"203d2025",
          6502 => x"3034580a",
          6503 => x"00000000",
          6504 => x"20202020",
          6505 => x"53797374",
          6506 => x"656d2043",
          6507 => x"6c6f636b",
          6508 => x"20467265",
          6509 => x"71202020",
          6510 => x"20202020",
          6511 => x"203d2025",
          6512 => x"642e2530",
          6513 => x"34644d48",
          6514 => x"7a0a0000",
          6515 => x"20202020",
          6516 => x"53445241",
          6517 => x"4d20436c",
          6518 => x"6f636b20",
          6519 => x"46726571",
          6520 => x"20202020",
          6521 => x"20202020",
          6522 => x"203d2025",
          6523 => x"642e2530",
          6524 => x"34644d48",
          6525 => x"7a0a0000",
          6526 => x"20202020",
          6527 => x"57697368",
          6528 => x"626f6e65",
          6529 => x"20534452",
          6530 => x"414d2043",
          6531 => x"6c6f636b",
          6532 => x"20467265",
          6533 => x"713d2025",
          6534 => x"642e2530",
          6535 => x"34644d48",
          6536 => x"7a0a0000",
          6537 => x"536d616c",
          6538 => x"6c000000",
          6539 => x"4d656469",
          6540 => x"756d0000",
          6541 => x"466c6578",
          6542 => x"00000000",
          6543 => x"45564f00",
          6544 => x"45564f6d",
          6545 => x"696e0000",
          6546 => x"556e6b6e",
          6547 => x"6f776e00",
          6548 => x"53440000",
          6549 => x"222a2b2c",
          6550 => x"3a3b3c3d",
          6551 => x"3e3f5b5d",
          6552 => x"7c7f0000",
          6553 => x"46415400",
          6554 => x"46415433",
          6555 => x"32000000",
          6556 => x"ebfe904d",
          6557 => x"53444f53",
          6558 => x"352e3000",
          6559 => x"4e4f204e",
          6560 => x"414d4520",
          6561 => x"20202046",
          6562 => x"41543332",
          6563 => x"20202000",
          6564 => x"4e4f204e",
          6565 => x"414d4520",
          6566 => x"20202046",
          6567 => x"41542020",
          6568 => x"20202000",
          6569 => x"00006650",
          6570 => x"00000000",
          6571 => x"00000000",
          6572 => x"00000000",
          6573 => x"809a4541",
          6574 => x"8e418f80",
          6575 => x"45454549",
          6576 => x"49498e8f",
          6577 => x"9092924f",
          6578 => x"994f5555",
          6579 => x"59999a9b",
          6580 => x"9c9d9e9f",
          6581 => x"41494f55",
          6582 => x"a5a5a6a7",
          6583 => x"a8a9aaab",
          6584 => x"acadaeaf",
          6585 => x"b0b1b2b3",
          6586 => x"b4b5b6b7",
          6587 => x"b8b9babb",
          6588 => x"bcbdbebf",
          6589 => x"c0c1c2c3",
          6590 => x"c4c5c6c7",
          6591 => x"c8c9cacb",
          6592 => x"cccdcecf",
          6593 => x"d0d1d2d3",
          6594 => x"d4d5d6d7",
          6595 => x"d8d9dadb",
          6596 => x"dcdddedf",
          6597 => x"e0e1e2e3",
          6598 => x"e4e5e6e7",
          6599 => x"e8e9eaeb",
          6600 => x"ecedeeef",
          6601 => x"f0f1f2f3",
          6602 => x"f4f5f6f7",
          6603 => x"f8f9fafb",
          6604 => x"fcfdfeff",
          6605 => x"2b2e2c3b",
          6606 => x"3d5b5d2f",
          6607 => x"5c222a3a",
          6608 => x"3c3e3f7c",
          6609 => x"7f000000",
          6610 => x"00010004",
          6611 => x"00100040",
          6612 => x"01000200",
          6613 => x"00000000",
          6614 => x"00010002",
          6615 => x"00040008",
          6616 => x"00100020",
          6617 => x"00000000",
          6618 => x"64696e69",
          6619 => x"74000000",
          6620 => x"64696f63",
          6621 => x"746c0000",
          6622 => x"66696e69",
          6623 => x"74000000",
          6624 => x"666c6f61",
          6625 => x"64000000",
          6626 => x"66657865",
          6627 => x"63000000",
          6628 => x"6d636c65",
          6629 => x"61720000",
          6630 => x"6d64756d",
          6631 => x"70000000",
          6632 => x"6d737263",
          6633 => x"68000000",
          6634 => x"6d656200",
          6635 => x"6d656800",
          6636 => x"6d657700",
          6637 => x"68696400",
          6638 => x"68696500",
          6639 => x"68666400",
          6640 => x"68666500",
          6641 => x"63616c6c",
          6642 => x"00000000",
          6643 => x"6a6d7000",
          6644 => x"72657374",
          6645 => x"61727400",
          6646 => x"72657365",
          6647 => x"74000000",
          6648 => x"696e666f",
          6649 => x"00000000",
          6650 => x"74657374",
          6651 => x"00000000",
          6652 => x"4469736b",
          6653 => x"20457272",
          6654 => x"6f720a00",
          6655 => x"496e7465",
          6656 => x"726e616c",
          6657 => x"20657272",
          6658 => x"6f722e0a",
          6659 => x"00000000",
          6660 => x"4469736b",
          6661 => x"206e6f74",
          6662 => x"20726561",
          6663 => x"64792e0a",
          6664 => x"00000000",
          6665 => x"4e6f2066",
          6666 => x"696c6520",
          6667 => x"666f756e",
          6668 => x"642e0a00",
          6669 => x"4e6f2070",
          6670 => x"61746820",
          6671 => x"666f756e",
          6672 => x"642e0a00",
          6673 => x"496e7661",
          6674 => x"6c696420",
          6675 => x"66696c65",
          6676 => x"6e616d65",
          6677 => x"2e0a0000",
          6678 => x"41636365",
          6679 => x"73732064",
          6680 => x"656e6965",
          6681 => x"642e0a00",
          6682 => x"46696c65",
          6683 => x"20616c72",
          6684 => x"65616479",
          6685 => x"20657869",
          6686 => x"7374732e",
          6687 => x"0a000000",
          6688 => x"46696c65",
          6689 => x"2068616e",
          6690 => x"646c6520",
          6691 => x"696e7661",
          6692 => x"6c69642e",
          6693 => x"0a000000",
          6694 => x"53442069",
          6695 => x"73207772",
          6696 => x"69746520",
          6697 => x"70726f74",
          6698 => x"65637465",
          6699 => x"642e0a00",
          6700 => x"44726976",
          6701 => x"65206e75",
          6702 => x"6d626572",
          6703 => x"20697320",
          6704 => x"696e7661",
          6705 => x"6c69642e",
          6706 => x"0a000000",
          6707 => x"4469736b",
          6708 => x"206e6f74",
          6709 => x"20656e61",
          6710 => x"626c6564",
          6711 => x"2e0a0000",
          6712 => x"4e6f2063",
          6713 => x"6f6d7061",
          6714 => x"7469626c",
          6715 => x"65206669",
          6716 => x"6c657379",
          6717 => x"7374656d",
          6718 => x"20666f75",
          6719 => x"6e64206f",
          6720 => x"6e206469",
          6721 => x"736b2e0a",
          6722 => x"00000000",
          6723 => x"466f726d",
          6724 => x"61742061",
          6725 => x"626f7274",
          6726 => x"65642e0a",
          6727 => x"00000000",
          6728 => x"54696d65",
          6729 => x"6f75742c",
          6730 => x"206f7065",
          6731 => x"72617469",
          6732 => x"6f6e2063",
          6733 => x"616e6365",
          6734 => x"6c6c6564",
          6735 => x"2e0a0000",
          6736 => x"46696c65",
          6737 => x"20697320",
          6738 => x"6c6f636b",
          6739 => x"65642e0a",
          6740 => x"00000000",
          6741 => x"496e7375",
          6742 => x"66666963",
          6743 => x"69656e74",
          6744 => x"206d656d",
          6745 => x"6f72792e",
          6746 => x"0a000000",
          6747 => x"546f6f20",
          6748 => x"6d616e79",
          6749 => x"206f7065",
          6750 => x"6e206669",
          6751 => x"6c65732e",
          6752 => x"0a000000",
          6753 => x"50617261",
          6754 => x"6d657465",
          6755 => x"72732069",
          6756 => x"6e636f72",
          6757 => x"72656374",
          6758 => x"2e0a0000",
          6759 => x"53756363",
          6760 => x"6573732e",
          6761 => x"0a000000",
          6762 => x"556e6b6e",
          6763 => x"6f776e20",
          6764 => x"6572726f",
          6765 => x"722e0a00",
          6766 => x"0a256c75",
          6767 => x"20627974",
          6768 => x"65732025",
          6769 => x"73206174",
          6770 => x"20256c75",
          6771 => x"20627974",
          6772 => x"65732f73",
          6773 => x"65632e0a",
          6774 => x"00000000",
          6775 => x"25303858",
          6776 => x"00000000",
          6777 => x"3a202000",
          6778 => x"25303458",
          6779 => x"00000000",
          6780 => x"20202020",
          6781 => x"20202020",
          6782 => x"00000000",
          6783 => x"25303258",
          6784 => x"00000000",
          6785 => x"20200000",
          6786 => x"207c0000",
          6787 => x"7c0d0a00",
          6788 => x"72656164",
          6789 => x"00000000",
          6790 => x"5a505554",
          6791 => x"41000000",
          6792 => x"0a2a2a20",
          6793 => x"25732028",
          6794 => x"00000000",
          6795 => x"32392f31",
          6796 => x"322f3230",
          6797 => x"31390000",
          6798 => x"76312e34",
          6799 => x"00000000",
          6800 => x"205a5055",
          6801 => x"2c207265",
          6802 => x"76202530",
          6803 => x"32782920",
          6804 => x"25732025",
          6805 => x"73202a2a",
          6806 => x"0a0a0000",
          6807 => x"5a505554",
          6808 => x"4120496e",
          6809 => x"74657272",
          6810 => x"75707420",
          6811 => x"48616e64",
          6812 => x"6c65720a",
          6813 => x"00000000",
          6814 => x"54696d65",
          6815 => x"7220696e",
          6816 => x"74657272",
          6817 => x"7570740a",
          6818 => x"00000000",
          6819 => x"50533220",
          6820 => x"696e7465",
          6821 => x"72727570",
          6822 => x"740a0000",
          6823 => x"494f4354",
          6824 => x"4c205244",
          6825 => x"20696e74",
          6826 => x"65727275",
          6827 => x"70740a00",
          6828 => x"494f4354",
          6829 => x"4c205752",
          6830 => x"20696e74",
          6831 => x"65727275",
          6832 => x"70740a00",
          6833 => x"55415254",
          6834 => x"30205258",
          6835 => x"20696e74",
          6836 => x"65727275",
          6837 => x"70740a00",
          6838 => x"55415254",
          6839 => x"30205458",
          6840 => x"20696e74",
          6841 => x"65727275",
          6842 => x"70740a00",
          6843 => x"55415254",
          6844 => x"31205258",
          6845 => x"20696e74",
          6846 => x"65727275",
          6847 => x"70740a00",
          6848 => x"55415254",
          6849 => x"31205458",
          6850 => x"20696e74",
          6851 => x"65727275",
          6852 => x"70740a00",
          6853 => x"53657474",
          6854 => x"696e6720",
          6855 => x"75702074",
          6856 => x"696d6572",
          6857 => x"2e2e2e0a",
          6858 => x"00000000",
          6859 => x"456e6162",
          6860 => x"6c696e67",
          6861 => x"2074696d",
          6862 => x"65722e2e",
          6863 => x"2e0a0000",
          6864 => x"6175746f",
          6865 => x"65786563",
          6866 => x"2e626174",
          6867 => x"00000000",
          6868 => x"303a0000",
          6869 => x"4661696c",
          6870 => x"65642074",
          6871 => x"6f20696e",
          6872 => x"69746961",
          6873 => x"6c697365",
          6874 => x"20736420",
          6875 => x"63617264",
          6876 => x"20302c20",
          6877 => x"706c6561",
          6878 => x"73652069",
          6879 => x"6e697420",
          6880 => x"6d616e75",
          6881 => x"616c6c79",
          6882 => x"2e0a0000",
          6883 => x"2a200000",
          6884 => x"42616420",
          6885 => x"6469736b",
          6886 => x"20696421",
          6887 => x"0a000000",
          6888 => x"496e6974",
          6889 => x"69616c69",
          6890 => x"7365642e",
          6891 => x"0a000000",
          6892 => x"4661696c",
          6893 => x"65642074",
          6894 => x"6f20696e",
          6895 => x"69746961",
          6896 => x"6c697365",
          6897 => x"2e0a0000",
          6898 => x"72633d25",
          6899 => x"640a0000",
          6900 => x"25753a00",
          6901 => x"436c6561",
          6902 => x"72696e67",
          6903 => x"2e2e2e2e",
          6904 => x"00000000",
          6905 => x"44756d70",
          6906 => x"204d656d",
          6907 => x"6f72790a",
          6908 => x"00000000",
          6909 => x"0a436f6d",
          6910 => x"706c6574",
          6911 => x"652e0a00",
          6912 => x"25303858",
          6913 => x"20253032",
          6914 => x"582d0000",
          6915 => x"3f3f3f0a",
          6916 => x"00000000",
          6917 => x"25303858",
          6918 => x"20253034",
          6919 => x"582d0000",
          6920 => x"25303858",
          6921 => x"20253038",
          6922 => x"582d0000",
          6923 => x"53656172",
          6924 => x"6368696e",
          6925 => x"672e2e0a",
          6926 => x"00000000",
          6927 => x"2530386c",
          6928 => x"782d3e25",
          6929 => x"30386c78",
          6930 => x"0a000000",
          6931 => x"44697361",
          6932 => x"626c696e",
          6933 => x"6720696e",
          6934 => x"74657272",
          6935 => x"75707473",
          6936 => x"0a000000",
          6937 => x"456e6162",
          6938 => x"6c696e67",
          6939 => x"20696e74",
          6940 => x"65727275",
          6941 => x"7074730a",
          6942 => x"00000000",
          6943 => x"44697361",
          6944 => x"626c6564",
          6945 => x"20756172",
          6946 => x"74206669",
          6947 => x"666f0a00",
          6948 => x"456e6162",
          6949 => x"6c696e67",
          6950 => x"20756172",
          6951 => x"74206669",
          6952 => x"666f0a00",
          6953 => x"45786563",
          6954 => x"7574696e",
          6955 => x"6720636f",
          6956 => x"64652040",
          6957 => x"20253038",
          6958 => x"78202e2e",
          6959 => x"2e0a0000",
          6960 => x"43616c6c",
          6961 => x"696e6720",
          6962 => x"636f6465",
          6963 => x"20402025",
          6964 => x"30387820",
          6965 => x"2e2e2e0a",
          6966 => x"00000000",
          6967 => x"43616c6c",
          6968 => x"20726574",
          6969 => x"75726e65",
          6970 => x"6420636f",
          6971 => x"64652028",
          6972 => x"2564292e",
          6973 => x"0a000000",
          6974 => x"52657374",
          6975 => x"61727469",
          6976 => x"6e672061",
          6977 => x"70706c69",
          6978 => x"63617469",
          6979 => x"6f6e2e2e",
          6980 => x"2e0a0000",
          6981 => x"436f6c64",
          6982 => x"20726562",
          6983 => x"6f6f7469",
          6984 => x"6e672e2e",
          6985 => x"2e0a0000",
          6986 => x"5a505500",
          6987 => x"62696e00",
          6988 => x"25643a5c",
          6989 => x"25735c25",
          6990 => x"732e2573",
          6991 => x"00000000",
          6992 => x"25643a5c",
          6993 => x"25735c25",
          6994 => x"73000000",
          6995 => x"25643a5c",
          6996 => x"25730000",
          6997 => x"42616420",
          6998 => x"636f6d6d",
          6999 => x"616e642e",
          7000 => x"0a000000",
          7001 => x"52756e6e",
          7002 => x"696e672e",
          7003 => x"2e2e0a00",
          7004 => x"456e6162",
          7005 => x"6c696e67",
          7006 => x"20696e74",
          7007 => x"65727275",
          7008 => x"7074732e",
          7009 => x"2e2e0a00",
          7010 => x"00000000",
          7011 => x"00000000",
          7012 => x"00007fff",
          7013 => x"00000000",
          7014 => x"00007fff",
          7015 => x"00010000",
          7016 => x"00007fff",
          7017 => x"00010000",
          7018 => x"00810000",
          7019 => x"01000000",
          7020 => x"017fffff",
          7021 => x"00000000",
          7022 => x"00000000",
          7023 => x"00007800",
          7024 => x"00000000",
          7025 => x"05f5e100",
          7026 => x"05f5e100",
          7027 => x"05f5e100",
          7028 => x"00000000",
          7029 => x"01010101",
          7030 => x"01010101",
          7031 => x"01011001",
          7032 => x"01000000",
          7033 => x"00000000",
          7034 => x"01000000",
          7035 => x"00000000",
          7036 => x"00006768",
          7037 => x"01020100",
          7038 => x"00000000",
          7039 => x"00000000",
          7040 => x"00006770",
          7041 => x"01040100",
          7042 => x"00000000",
          7043 => x"00000000",
          7044 => x"00006778",
          7045 => x"01140300",
          7046 => x"00000000",
          7047 => x"00000000",
          7048 => x"00006780",
          7049 => x"012b0300",
          7050 => x"00000000",
          7051 => x"00000000",
          7052 => x"00006788",
          7053 => x"01300300",
          7054 => x"00000000",
          7055 => x"00000000",
          7056 => x"00006790",
          7057 => x"013c0400",
          7058 => x"00000000",
          7059 => x"00000000",
          7060 => x"00006798",
          7061 => x"01400400",
          7062 => x"00000000",
          7063 => x"00000000",
          7064 => x"000067a0",
          7065 => x"01450400",
          7066 => x"00000000",
          7067 => x"00000000",
          7068 => x"000067a8",
          7069 => x"01410400",
          7070 => x"00000000",
          7071 => x"00000000",
          7072 => x"000067ac",
          7073 => x"01420400",
          7074 => x"00000000",
          7075 => x"00000000",
          7076 => x"000067b0",
          7077 => x"01430400",
          7078 => x"00000000",
          7079 => x"00000000",
          7080 => x"000067b4",
          7081 => x"01500500",
          7082 => x"00000000",
          7083 => x"00000000",
          7084 => x"000067b8",
          7085 => x"01510500",
          7086 => x"00000000",
          7087 => x"00000000",
          7088 => x"000067bc",
          7089 => x"01540500",
          7090 => x"00000000",
          7091 => x"00000000",
          7092 => x"000067c0",
          7093 => x"01550500",
          7094 => x"00000000",
          7095 => x"00000000",
          7096 => x"000067c4",
          7097 => x"01790700",
          7098 => x"00000000",
          7099 => x"00000000",
          7100 => x"000067cc",
          7101 => x"01780700",
          7102 => x"00000000",
          7103 => x"00000000",
          7104 => x"000067d0",
          7105 => x"01820800",
          7106 => x"00000000",
          7107 => x"00000000",
          7108 => x"000067d8",
          7109 => x"01830800",
          7110 => x"00000000",
          7111 => x"00000000",
          7112 => x"000067e0",
          7113 => x"01850800",
          7114 => x"00000000",
          7115 => x"00000000",
          7116 => x"000067e8",
          7117 => x"01870800",
          7118 => x"00000000",
          7119 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

