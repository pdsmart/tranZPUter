../../../../cpu/zpu_core_evo.vhd