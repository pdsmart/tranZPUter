-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"92",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"92",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"9f",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"c5",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"93",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"95",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"cc",
           386 => x"2d",
           387 => x"08",
           388 => x"04",
           389 => x"0c",
           390 => x"81",
           391 => x"82",
           392 => x"81",
           393 => x"ae",
           394 => x"de",
           395 => x"80",
           396 => x"de",
           397 => x"bf",
           398 => x"cc",
           399 => x"90",
           400 => x"cc",
           401 => x"2d",
           402 => x"08",
           403 => x"04",
           404 => x"0c",
           405 => x"81",
           406 => x"82",
           407 => x"81",
           408 => x"ae",
           409 => x"de",
           410 => x"80",
           411 => x"de",
           412 => x"98",
           413 => x"cc",
           414 => x"90",
           415 => x"cc",
           416 => x"2d",
           417 => x"08",
           418 => x"04",
           419 => x"0c",
           420 => x"81",
           421 => x"82",
           422 => x"81",
           423 => x"b4",
           424 => x"de",
           425 => x"80",
           426 => x"de",
           427 => x"dd",
           428 => x"cc",
           429 => x"90",
           430 => x"cc",
           431 => x"2d",
           432 => x"08",
           433 => x"04",
           434 => x"0c",
           435 => x"81",
           436 => x"82",
           437 => x"81",
           438 => x"9b",
           439 => x"de",
           440 => x"80",
           441 => x"de",
           442 => x"dd",
           443 => x"cc",
           444 => x"90",
           445 => x"cc",
           446 => x"2d",
           447 => x"08",
           448 => x"04",
           449 => x"0c",
           450 => x"2d",
           451 => x"08",
           452 => x"04",
           453 => x"0c",
           454 => x"2d",
           455 => x"08",
           456 => x"04",
           457 => x"0c",
           458 => x"2d",
           459 => x"08",
           460 => x"04",
           461 => x"0c",
           462 => x"2d",
           463 => x"08",
           464 => x"04",
           465 => x"0c",
           466 => x"2d",
           467 => x"08",
           468 => x"04",
           469 => x"0c",
           470 => x"2d",
           471 => x"08",
           472 => x"04",
           473 => x"0c",
           474 => x"2d",
           475 => x"08",
           476 => x"04",
           477 => x"0c",
           478 => x"2d",
           479 => x"08",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"04",
           485 => x"0c",
           486 => x"2d",
           487 => x"08",
           488 => x"04",
           489 => x"0c",
           490 => x"2d",
           491 => x"08",
           492 => x"04",
           493 => x"0c",
           494 => x"2d",
           495 => x"08",
           496 => x"04",
           497 => x"0c",
           498 => x"2d",
           499 => x"08",
           500 => x"04",
           501 => x"0c",
           502 => x"2d",
           503 => x"08",
           504 => x"04",
           505 => x"0c",
           506 => x"2d",
           507 => x"08",
           508 => x"04",
           509 => x"0c",
           510 => x"2d",
           511 => x"08",
           512 => x"04",
           513 => x"0c",
           514 => x"2d",
           515 => x"08",
           516 => x"04",
           517 => x"0c",
           518 => x"2d",
           519 => x"08",
           520 => x"04",
           521 => x"0c",
           522 => x"2d",
           523 => x"08",
           524 => x"04",
           525 => x"0c",
           526 => x"2d",
           527 => x"08",
           528 => x"04",
           529 => x"0c",
           530 => x"2d",
           531 => x"08",
           532 => x"04",
           533 => x"0c",
           534 => x"2d",
           535 => x"08",
           536 => x"04",
           537 => x"0c",
           538 => x"2d",
           539 => x"08",
           540 => x"04",
           541 => x"0c",
           542 => x"2d",
           543 => x"08",
           544 => x"04",
           545 => x"0c",
           546 => x"2d",
           547 => x"08",
           548 => x"04",
           549 => x"0c",
           550 => x"81",
           551 => x"82",
           552 => x"81",
           553 => x"bd",
           554 => x"de",
           555 => x"80",
           556 => x"de",
           557 => x"e7",
           558 => x"cc",
           559 => x"90",
           560 => x"cc",
           561 => x"2d",
           562 => x"08",
           563 => x"04",
           564 => x"0c",
           565 => x"81",
           566 => x"82",
           567 => x"81",
           568 => x"9f",
           569 => x"de",
           570 => x"80",
           571 => x"de",
           572 => x"a5",
           573 => x"de",
           574 => x"80",
           575 => x"04",
           576 => x"10",
           577 => x"10",
           578 => x"10",
           579 => x"10",
           580 => x"10",
           581 => x"10",
           582 => x"10",
           583 => x"53",
           584 => x"00",
           585 => x"06",
           586 => x"09",
           587 => x"05",
           588 => x"2b",
           589 => x"06",
           590 => x"04",
           591 => x"72",
           592 => x"05",
           593 => x"05",
           594 => x"72",
           595 => x"53",
           596 => x"51",
           597 => x"04",
           598 => x"70",
           599 => x"27",
           600 => x"71",
           601 => x"53",
           602 => x"0b",
           603 => x"8c",
           604 => x"c4",
           605 => x"81",
           606 => x"02",
           607 => x"0c",
           608 => x"80",
           609 => x"cc",
           610 => x"08",
           611 => x"cc",
           612 => x"08",
           613 => x"3f",
           614 => x"08",
           615 => x"c0",
           616 => x"3d",
           617 => x"cc",
           618 => x"de",
           619 => x"81",
           620 => x"fd",
           621 => x"53",
           622 => x"08",
           623 => x"52",
           624 => x"08",
           625 => x"51",
           626 => x"81",
           627 => x"70",
           628 => x"0c",
           629 => x"0d",
           630 => x"0c",
           631 => x"cc",
           632 => x"de",
           633 => x"3d",
           634 => x"81",
           635 => x"fc",
           636 => x"de",
           637 => x"05",
           638 => x"b9",
           639 => x"cc",
           640 => x"08",
           641 => x"cc",
           642 => x"0c",
           643 => x"de",
           644 => x"05",
           645 => x"cc",
           646 => x"08",
           647 => x"0b",
           648 => x"08",
           649 => x"81",
           650 => x"f4",
           651 => x"de",
           652 => x"05",
           653 => x"cc",
           654 => x"08",
           655 => x"38",
           656 => x"08",
           657 => x"30",
           658 => x"08",
           659 => x"80",
           660 => x"cc",
           661 => x"0c",
           662 => x"08",
           663 => x"8a",
           664 => x"81",
           665 => x"f0",
           666 => x"de",
           667 => x"05",
           668 => x"cc",
           669 => x"0c",
           670 => x"de",
           671 => x"05",
           672 => x"de",
           673 => x"05",
           674 => x"df",
           675 => x"c0",
           676 => x"de",
           677 => x"05",
           678 => x"de",
           679 => x"05",
           680 => x"90",
           681 => x"cc",
           682 => x"08",
           683 => x"cc",
           684 => x"0c",
           685 => x"08",
           686 => x"70",
           687 => x"0c",
           688 => x"0d",
           689 => x"0c",
           690 => x"cc",
           691 => x"de",
           692 => x"3d",
           693 => x"81",
           694 => x"fc",
           695 => x"de",
           696 => x"05",
           697 => x"99",
           698 => x"cc",
           699 => x"08",
           700 => x"cc",
           701 => x"0c",
           702 => x"de",
           703 => x"05",
           704 => x"cc",
           705 => x"08",
           706 => x"38",
           707 => x"08",
           708 => x"30",
           709 => x"08",
           710 => x"81",
           711 => x"cc",
           712 => x"08",
           713 => x"cc",
           714 => x"08",
           715 => x"81",
           716 => x"70",
           717 => x"08",
           718 => x"54",
           719 => x"08",
           720 => x"80",
           721 => x"81",
           722 => x"f8",
           723 => x"81",
           724 => x"f8",
           725 => x"de",
           726 => x"05",
           727 => x"de",
           728 => x"87",
           729 => x"de",
           730 => x"81",
           731 => x"02",
           732 => x"0c",
           733 => x"81",
           734 => x"cc",
           735 => x"0c",
           736 => x"de",
           737 => x"05",
           738 => x"cc",
           739 => x"08",
           740 => x"08",
           741 => x"27",
           742 => x"de",
           743 => x"05",
           744 => x"ae",
           745 => x"81",
           746 => x"8c",
           747 => x"a2",
           748 => x"cc",
           749 => x"08",
           750 => x"cc",
           751 => x"0c",
           752 => x"08",
           753 => x"10",
           754 => x"08",
           755 => x"ff",
           756 => x"de",
           757 => x"05",
           758 => x"80",
           759 => x"de",
           760 => x"05",
           761 => x"cc",
           762 => x"08",
           763 => x"81",
           764 => x"88",
           765 => x"de",
           766 => x"05",
           767 => x"de",
           768 => x"05",
           769 => x"cc",
           770 => x"08",
           771 => x"08",
           772 => x"07",
           773 => x"08",
           774 => x"81",
           775 => x"fc",
           776 => x"2a",
           777 => x"08",
           778 => x"81",
           779 => x"8c",
           780 => x"2a",
           781 => x"08",
           782 => x"ff",
           783 => x"de",
           784 => x"05",
           785 => x"93",
           786 => x"cc",
           787 => x"08",
           788 => x"cc",
           789 => x"0c",
           790 => x"81",
           791 => x"f8",
           792 => x"81",
           793 => x"f4",
           794 => x"81",
           795 => x"f4",
           796 => x"de",
           797 => x"3d",
           798 => x"cc",
           799 => x"3d",
           800 => x"71",
           801 => x"9f",
           802 => x"55",
           803 => x"72",
           804 => x"74",
           805 => x"70",
           806 => x"38",
           807 => x"71",
           808 => x"38",
           809 => x"81",
           810 => x"ff",
           811 => x"ff",
           812 => x"06",
           813 => x"81",
           814 => x"86",
           815 => x"74",
           816 => x"75",
           817 => x"90",
           818 => x"54",
           819 => x"27",
           820 => x"71",
           821 => x"53",
           822 => x"70",
           823 => x"0c",
           824 => x"84",
           825 => x"72",
           826 => x"05",
           827 => x"12",
           828 => x"26",
           829 => x"72",
           830 => x"72",
           831 => x"05",
           832 => x"12",
           833 => x"26",
           834 => x"53",
           835 => x"fb",
           836 => x"79",
           837 => x"83",
           838 => x"52",
           839 => x"71",
           840 => x"54",
           841 => x"73",
           842 => x"c6",
           843 => x"54",
           844 => x"70",
           845 => x"52",
           846 => x"2e",
           847 => x"33",
           848 => x"2e",
           849 => x"95",
           850 => x"81",
           851 => x"70",
           852 => x"54",
           853 => x"70",
           854 => x"33",
           855 => x"ff",
           856 => x"ff",
           857 => x"31",
           858 => x"0c",
           859 => x"3d",
           860 => x"09",
           861 => x"fd",
           862 => x"70",
           863 => x"81",
           864 => x"51",
           865 => x"38",
           866 => x"16",
           867 => x"56",
           868 => x"08",
           869 => x"73",
           870 => x"ff",
           871 => x"0b",
           872 => x"0c",
           873 => x"04",
           874 => x"80",
           875 => x"71",
           876 => x"87",
           877 => x"de",
           878 => x"ff",
           879 => x"ff",
           880 => x"72",
           881 => x"38",
           882 => x"c0",
           883 => x"0d",
           884 => x"0d",
           885 => x"70",
           886 => x"71",
           887 => x"ca",
           888 => x"51",
           889 => x"09",
           890 => x"38",
           891 => x"f1",
           892 => x"84",
           893 => x"53",
           894 => x"70",
           895 => x"53",
           896 => x"a0",
           897 => x"81",
           898 => x"2e",
           899 => x"e5",
           900 => x"ff",
           901 => x"a0",
           902 => x"06",
           903 => x"73",
           904 => x"55",
           905 => x"0c",
           906 => x"81",
           907 => x"87",
           908 => x"fc",
           909 => x"53",
           910 => x"2e",
           911 => x"3d",
           912 => x"72",
           913 => x"3f",
           914 => x"08",
           915 => x"53",
           916 => x"53",
           917 => x"c0",
           918 => x"0d",
           919 => x"0d",
           920 => x"33",
           921 => x"53",
           922 => x"8b",
           923 => x"38",
           924 => x"ff",
           925 => x"52",
           926 => x"81",
           927 => x"13",
           928 => x"52",
           929 => x"80",
           930 => x"13",
           931 => x"52",
           932 => x"80",
           933 => x"13",
           934 => x"52",
           935 => x"80",
           936 => x"13",
           937 => x"52",
           938 => x"26",
           939 => x"8a",
           940 => x"87",
           941 => x"e7",
           942 => x"38",
           943 => x"c0",
           944 => x"72",
           945 => x"98",
           946 => x"13",
           947 => x"98",
           948 => x"13",
           949 => x"98",
           950 => x"13",
           951 => x"98",
           952 => x"13",
           953 => x"98",
           954 => x"13",
           955 => x"98",
           956 => x"87",
           957 => x"0c",
           958 => x"98",
           959 => x"0b",
           960 => x"9c",
           961 => x"71",
           962 => x"0c",
           963 => x"04",
           964 => x"7f",
           965 => x"98",
           966 => x"7d",
           967 => x"98",
           968 => x"7d",
           969 => x"c0",
           970 => x"5a",
           971 => x"34",
           972 => x"b4",
           973 => x"83",
           974 => x"c0",
           975 => x"5a",
           976 => x"34",
           977 => x"ac",
           978 => x"85",
           979 => x"c0",
           980 => x"5a",
           981 => x"34",
           982 => x"a4",
           983 => x"88",
           984 => x"c0",
           985 => x"5a",
           986 => x"23",
           987 => x"79",
           988 => x"06",
           989 => x"ff",
           990 => x"86",
           991 => x"85",
           992 => x"84",
           993 => x"83",
           994 => x"82",
           995 => x"7d",
           996 => x"06",
           997 => x"e4",
           998 => x"3f",
           999 => x"04",
          1000 => x"02",
          1001 => x"70",
          1002 => x"2a",
          1003 => x"70",
          1004 => x"db",
          1005 => x"3d",
          1006 => x"3d",
          1007 => x"0b",
          1008 => x"33",
          1009 => x"06",
          1010 => x"87",
          1011 => x"51",
          1012 => x"86",
          1013 => x"94",
          1014 => x"08",
          1015 => x"70",
          1016 => x"54",
          1017 => x"2e",
          1018 => x"91",
          1019 => x"06",
          1020 => x"d7",
          1021 => x"32",
          1022 => x"51",
          1023 => x"2e",
          1024 => x"93",
          1025 => x"06",
          1026 => x"ff",
          1027 => x"81",
          1028 => x"87",
          1029 => x"52",
          1030 => x"86",
          1031 => x"94",
          1032 => x"72",
          1033 => x"de",
          1034 => x"3d",
          1035 => x"3d",
          1036 => x"05",
          1037 => x"81",
          1038 => x"70",
          1039 => x"57",
          1040 => x"c0",
          1041 => x"74",
          1042 => x"38",
          1043 => x"94",
          1044 => x"70",
          1045 => x"81",
          1046 => x"52",
          1047 => x"8c",
          1048 => x"2a",
          1049 => x"51",
          1050 => x"38",
          1051 => x"70",
          1052 => x"51",
          1053 => x"8d",
          1054 => x"2a",
          1055 => x"51",
          1056 => x"be",
          1057 => x"ff",
          1058 => x"c0",
          1059 => x"70",
          1060 => x"38",
          1061 => x"90",
          1062 => x"0c",
          1063 => x"04",
          1064 => x"79",
          1065 => x"33",
          1066 => x"06",
          1067 => x"70",
          1068 => x"fe",
          1069 => x"ff",
          1070 => x"0b",
          1071 => x"88",
          1072 => x"ff",
          1073 => x"55",
          1074 => x"94",
          1075 => x"80",
          1076 => x"87",
          1077 => x"51",
          1078 => x"96",
          1079 => x"06",
          1080 => x"70",
          1081 => x"38",
          1082 => x"70",
          1083 => x"51",
          1084 => x"72",
          1085 => x"81",
          1086 => x"70",
          1087 => x"38",
          1088 => x"70",
          1089 => x"51",
          1090 => x"38",
          1091 => x"06",
          1092 => x"94",
          1093 => x"80",
          1094 => x"87",
          1095 => x"52",
          1096 => x"81",
          1097 => x"70",
          1098 => x"53",
          1099 => x"ff",
          1100 => x"81",
          1101 => x"89",
          1102 => x"fe",
          1103 => x"0b",
          1104 => x"33",
          1105 => x"06",
          1106 => x"c0",
          1107 => x"72",
          1108 => x"38",
          1109 => x"94",
          1110 => x"70",
          1111 => x"81",
          1112 => x"51",
          1113 => x"e2",
          1114 => x"ff",
          1115 => x"c0",
          1116 => x"70",
          1117 => x"38",
          1118 => x"90",
          1119 => x"70",
          1120 => x"81",
          1121 => x"51",
          1122 => x"04",
          1123 => x"0b",
          1124 => x"88",
          1125 => x"ff",
          1126 => x"87",
          1127 => x"52",
          1128 => x"86",
          1129 => x"94",
          1130 => x"08",
          1131 => x"70",
          1132 => x"51",
          1133 => x"70",
          1134 => x"38",
          1135 => x"06",
          1136 => x"94",
          1137 => x"80",
          1138 => x"87",
          1139 => x"52",
          1140 => x"98",
          1141 => x"2c",
          1142 => x"71",
          1143 => x"0c",
          1144 => x"04",
          1145 => x"87",
          1146 => x"08",
          1147 => x"8a",
          1148 => x"70",
          1149 => x"b4",
          1150 => x"9e",
          1151 => x"db",
          1152 => x"c0",
          1153 => x"81",
          1154 => x"87",
          1155 => x"08",
          1156 => x"0c",
          1157 => x"98",
          1158 => x"98",
          1159 => x"9e",
          1160 => x"db",
          1161 => x"c0",
          1162 => x"81",
          1163 => x"87",
          1164 => x"08",
          1165 => x"0c",
          1166 => x"b0",
          1167 => x"a8",
          1168 => x"9e",
          1169 => x"db",
          1170 => x"c0",
          1171 => x"81",
          1172 => x"87",
          1173 => x"08",
          1174 => x"0c",
          1175 => x"c0",
          1176 => x"b8",
          1177 => x"9e",
          1178 => x"db",
          1179 => x"c0",
          1180 => x"51",
          1181 => x"c0",
          1182 => x"9e",
          1183 => x"db",
          1184 => x"c0",
          1185 => x"81",
          1186 => x"87",
          1187 => x"08",
          1188 => x"0c",
          1189 => x"db",
          1190 => x"0b",
          1191 => x"90",
          1192 => x"80",
          1193 => x"52",
          1194 => x"2e",
          1195 => x"52",
          1196 => x"d1",
          1197 => x"87",
          1198 => x"08",
          1199 => x"0a",
          1200 => x"52",
          1201 => x"83",
          1202 => x"71",
          1203 => x"34",
          1204 => x"c0",
          1205 => x"70",
          1206 => x"06",
          1207 => x"70",
          1208 => x"38",
          1209 => x"81",
          1210 => x"80",
          1211 => x"9e",
          1212 => x"88",
          1213 => x"51",
          1214 => x"80",
          1215 => x"81",
          1216 => x"db",
          1217 => x"0b",
          1218 => x"90",
          1219 => x"80",
          1220 => x"52",
          1221 => x"2e",
          1222 => x"52",
          1223 => x"d5",
          1224 => x"87",
          1225 => x"08",
          1226 => x"80",
          1227 => x"52",
          1228 => x"83",
          1229 => x"71",
          1230 => x"34",
          1231 => x"c0",
          1232 => x"70",
          1233 => x"06",
          1234 => x"70",
          1235 => x"38",
          1236 => x"81",
          1237 => x"80",
          1238 => x"9e",
          1239 => x"82",
          1240 => x"51",
          1241 => x"80",
          1242 => x"81",
          1243 => x"db",
          1244 => x"0b",
          1245 => x"90",
          1246 => x"80",
          1247 => x"52",
          1248 => x"2e",
          1249 => x"52",
          1250 => x"d9",
          1251 => x"87",
          1252 => x"08",
          1253 => x"80",
          1254 => x"52",
          1255 => x"83",
          1256 => x"71",
          1257 => x"34",
          1258 => x"c0",
          1259 => x"70",
          1260 => x"51",
          1261 => x"80",
          1262 => x"81",
          1263 => x"db",
          1264 => x"c0",
          1265 => x"70",
          1266 => x"70",
          1267 => x"51",
          1268 => x"db",
          1269 => x"0b",
          1270 => x"90",
          1271 => x"80",
          1272 => x"52",
          1273 => x"83",
          1274 => x"71",
          1275 => x"34",
          1276 => x"90",
          1277 => x"f0",
          1278 => x"2a",
          1279 => x"70",
          1280 => x"34",
          1281 => x"c0",
          1282 => x"70",
          1283 => x"52",
          1284 => x"2e",
          1285 => x"52",
          1286 => x"df",
          1287 => x"9e",
          1288 => x"87",
          1289 => x"70",
          1290 => x"34",
          1291 => x"04",
          1292 => x"81",
          1293 => x"86",
          1294 => x"db",
          1295 => x"73",
          1296 => x"38",
          1297 => x"51",
          1298 => x"81",
          1299 => x"85",
          1300 => x"db",
          1301 => x"73",
          1302 => x"38",
          1303 => x"08",
          1304 => x"08",
          1305 => x"81",
          1306 => x"8b",
          1307 => x"db",
          1308 => x"73",
          1309 => x"38",
          1310 => x"08",
          1311 => x"08",
          1312 => x"81",
          1313 => x"8b",
          1314 => x"db",
          1315 => x"73",
          1316 => x"38",
          1317 => x"08",
          1318 => x"08",
          1319 => x"81",
          1320 => x"8a",
          1321 => x"db",
          1322 => x"73",
          1323 => x"38",
          1324 => x"08",
          1325 => x"08",
          1326 => x"81",
          1327 => x"8a",
          1328 => x"db",
          1329 => x"73",
          1330 => x"38",
          1331 => x"08",
          1332 => x"08",
          1333 => x"81",
          1334 => x"8a",
          1335 => x"db",
          1336 => x"73",
          1337 => x"38",
          1338 => x"33",
          1339 => x"c8",
          1340 => x"3f",
          1341 => x"33",
          1342 => x"2e",
          1343 => x"db",
          1344 => x"81",
          1345 => x"8a",
          1346 => x"db",
          1347 => x"73",
          1348 => x"38",
          1349 => x"33",
          1350 => x"88",
          1351 => x"3f",
          1352 => x"33",
          1353 => x"2e",
          1354 => x"c9",
          1355 => x"8f",
          1356 => x"d3",
          1357 => x"80",
          1358 => x"81",
          1359 => x"83",
          1360 => x"db",
          1361 => x"73",
          1362 => x"38",
          1363 => x"51",
          1364 => x"81",
          1365 => x"54",
          1366 => x"88",
          1367 => x"d4",
          1368 => x"3f",
          1369 => x"33",
          1370 => x"2e",
          1371 => x"c9",
          1372 => x"cb",
          1373 => x"ec",
          1374 => x"3f",
          1375 => x"08",
          1376 => x"f8",
          1377 => x"3f",
          1378 => x"08",
          1379 => x"a0",
          1380 => x"3f",
          1381 => x"08",
          1382 => x"c8",
          1383 => x"3f",
          1384 => x"51",
          1385 => x"81",
          1386 => x"52",
          1387 => x"51",
          1388 => x"81",
          1389 => x"56",
          1390 => x"52",
          1391 => x"b7",
          1392 => x"c0",
          1393 => x"c0",
          1394 => x"31",
          1395 => x"de",
          1396 => x"81",
          1397 => x"88",
          1398 => x"db",
          1399 => x"73",
          1400 => x"38",
          1401 => x"08",
          1402 => x"c0",
          1403 => x"e7",
          1404 => x"de",
          1405 => x"84",
          1406 => x"71",
          1407 => x"81",
          1408 => x"52",
          1409 => x"51",
          1410 => x"81",
          1411 => x"54",
          1412 => x"a8",
          1413 => x"cc",
          1414 => x"84",
          1415 => x"51",
          1416 => x"81",
          1417 => x"bd",
          1418 => x"76",
          1419 => x"54",
          1420 => x"08",
          1421 => x"f8",
          1422 => x"3f",
          1423 => x"51",
          1424 => x"87",
          1425 => x"fe",
          1426 => x"92",
          1427 => x"05",
          1428 => x"26",
          1429 => x"84",
          1430 => x"80",
          1431 => x"08",
          1432 => x"a4",
          1433 => x"81",
          1434 => x"97",
          1435 => x"b4",
          1436 => x"81",
          1437 => x"8b",
          1438 => x"c0",
          1439 => x"81",
          1440 => x"f4",
          1441 => x"3d",
          1442 => x"88",
          1443 => x"80",
          1444 => x"96",
          1445 => x"ff",
          1446 => x"c0",
          1447 => x"08",
          1448 => x"72",
          1449 => x"07",
          1450 => x"e4",
          1451 => x"83",
          1452 => x"ff",
          1453 => x"c0",
          1454 => x"08",
          1455 => x"0c",
          1456 => x"0c",
          1457 => x"81",
          1458 => x"06",
          1459 => x"e4",
          1460 => x"51",
          1461 => x"04",
          1462 => x"08",
          1463 => x"84",
          1464 => x"3d",
          1465 => x"05",
          1466 => x"8a",
          1467 => x"06",
          1468 => x"51",
          1469 => x"de",
          1470 => x"71",
          1471 => x"38",
          1472 => x"81",
          1473 => x"81",
          1474 => x"d8",
          1475 => x"81",
          1476 => x"52",
          1477 => x"85",
          1478 => x"71",
          1479 => x"0d",
          1480 => x"0d",
          1481 => x"33",
          1482 => x"08",
          1483 => x"d0",
          1484 => x"ff",
          1485 => x"81",
          1486 => x"84",
          1487 => x"fd",
          1488 => x"54",
          1489 => x"81",
          1490 => x"53",
          1491 => x"8e",
          1492 => x"ff",
          1493 => x"14",
          1494 => x"3f",
          1495 => x"3d",
          1496 => x"3d",
          1497 => x"de",
          1498 => x"81",
          1499 => x"56",
          1500 => x"70",
          1501 => x"53",
          1502 => x"2e",
          1503 => x"81",
          1504 => x"81",
          1505 => x"da",
          1506 => x"74",
          1507 => x"0c",
          1508 => x"04",
          1509 => x"66",
          1510 => x"78",
          1511 => x"5a",
          1512 => x"80",
          1513 => x"38",
          1514 => x"09",
          1515 => x"de",
          1516 => x"7a",
          1517 => x"5c",
          1518 => x"5b",
          1519 => x"09",
          1520 => x"38",
          1521 => x"39",
          1522 => x"09",
          1523 => x"38",
          1524 => x"70",
          1525 => x"33",
          1526 => x"2e",
          1527 => x"92",
          1528 => x"19",
          1529 => x"70",
          1530 => x"33",
          1531 => x"53",
          1532 => x"16",
          1533 => x"26",
          1534 => x"88",
          1535 => x"05",
          1536 => x"05",
          1537 => x"05",
          1538 => x"5b",
          1539 => x"80",
          1540 => x"30",
          1541 => x"80",
          1542 => x"cc",
          1543 => x"70",
          1544 => x"25",
          1545 => x"54",
          1546 => x"53",
          1547 => x"8c",
          1548 => x"07",
          1549 => x"05",
          1550 => x"5a",
          1551 => x"83",
          1552 => x"54",
          1553 => x"27",
          1554 => x"16",
          1555 => x"06",
          1556 => x"80",
          1557 => x"aa",
          1558 => x"cf",
          1559 => x"73",
          1560 => x"81",
          1561 => x"80",
          1562 => x"38",
          1563 => x"2e",
          1564 => x"81",
          1565 => x"80",
          1566 => x"8a",
          1567 => x"39",
          1568 => x"2e",
          1569 => x"73",
          1570 => x"8a",
          1571 => x"d3",
          1572 => x"80",
          1573 => x"80",
          1574 => x"ee",
          1575 => x"39",
          1576 => x"71",
          1577 => x"53",
          1578 => x"54",
          1579 => x"2e",
          1580 => x"15",
          1581 => x"33",
          1582 => x"72",
          1583 => x"81",
          1584 => x"39",
          1585 => x"56",
          1586 => x"27",
          1587 => x"51",
          1588 => x"75",
          1589 => x"72",
          1590 => x"38",
          1591 => x"df",
          1592 => x"16",
          1593 => x"7b",
          1594 => x"38",
          1595 => x"f2",
          1596 => x"77",
          1597 => x"12",
          1598 => x"53",
          1599 => x"5c",
          1600 => x"5c",
          1601 => x"5c",
          1602 => x"5c",
          1603 => x"51",
          1604 => x"fd",
          1605 => x"82",
          1606 => x"06",
          1607 => x"80",
          1608 => x"77",
          1609 => x"53",
          1610 => x"18",
          1611 => x"72",
          1612 => x"c4",
          1613 => x"70",
          1614 => x"25",
          1615 => x"55",
          1616 => x"8d",
          1617 => x"2e",
          1618 => x"30",
          1619 => x"5b",
          1620 => x"8f",
          1621 => x"7b",
          1622 => x"e0",
          1623 => x"de",
          1624 => x"ff",
          1625 => x"75",
          1626 => x"8b",
          1627 => x"c0",
          1628 => x"74",
          1629 => x"a7",
          1630 => x"80",
          1631 => x"38",
          1632 => x"72",
          1633 => x"54",
          1634 => x"72",
          1635 => x"05",
          1636 => x"17",
          1637 => x"77",
          1638 => x"51",
          1639 => x"9f",
          1640 => x"72",
          1641 => x"79",
          1642 => x"81",
          1643 => x"72",
          1644 => x"38",
          1645 => x"05",
          1646 => x"ad",
          1647 => x"17",
          1648 => x"81",
          1649 => x"b0",
          1650 => x"38",
          1651 => x"81",
          1652 => x"06",
          1653 => x"9f",
          1654 => x"55",
          1655 => x"97",
          1656 => x"f9",
          1657 => x"81",
          1658 => x"8b",
          1659 => x"16",
          1660 => x"73",
          1661 => x"96",
          1662 => x"e0",
          1663 => x"17",
          1664 => x"33",
          1665 => x"f9",
          1666 => x"f2",
          1667 => x"16",
          1668 => x"7b",
          1669 => x"38",
          1670 => x"c6",
          1671 => x"96",
          1672 => x"fd",
          1673 => x"3d",
          1674 => x"05",
          1675 => x"52",
          1676 => x"e0",
          1677 => x"0d",
          1678 => x"0d",
          1679 => x"d8",
          1680 => x"88",
          1681 => x"51",
          1682 => x"81",
          1683 => x"53",
          1684 => x"80",
          1685 => x"d8",
          1686 => x"0d",
          1687 => x"0d",
          1688 => x"08",
          1689 => x"d0",
          1690 => x"88",
          1691 => x"52",
          1692 => x"3f",
          1693 => x"d0",
          1694 => x"0d",
          1695 => x"0d",
          1696 => x"de",
          1697 => x"56",
          1698 => x"80",
          1699 => x"2e",
          1700 => x"81",
          1701 => x"52",
          1702 => x"de",
          1703 => x"ff",
          1704 => x"80",
          1705 => x"38",
          1706 => x"b9",
          1707 => x"32",
          1708 => x"80",
          1709 => x"52",
          1710 => x"8b",
          1711 => x"2e",
          1712 => x"14",
          1713 => x"9f",
          1714 => x"38",
          1715 => x"73",
          1716 => x"38",
          1717 => x"72",
          1718 => x"14",
          1719 => x"f8",
          1720 => x"af",
          1721 => x"52",
          1722 => x"8a",
          1723 => x"3f",
          1724 => x"81",
          1725 => x"87",
          1726 => x"fe",
          1727 => x"de",
          1728 => x"81",
          1729 => x"77",
          1730 => x"53",
          1731 => x"72",
          1732 => x"0c",
          1733 => x"04",
          1734 => x"7a",
          1735 => x"80",
          1736 => x"58",
          1737 => x"33",
          1738 => x"a0",
          1739 => x"06",
          1740 => x"13",
          1741 => x"39",
          1742 => x"09",
          1743 => x"38",
          1744 => x"11",
          1745 => x"08",
          1746 => x"54",
          1747 => x"2e",
          1748 => x"80",
          1749 => x"08",
          1750 => x"0c",
          1751 => x"33",
          1752 => x"80",
          1753 => x"38",
          1754 => x"80",
          1755 => x"38",
          1756 => x"57",
          1757 => x"0c",
          1758 => x"33",
          1759 => x"39",
          1760 => x"74",
          1761 => x"38",
          1762 => x"80",
          1763 => x"89",
          1764 => x"38",
          1765 => x"d0",
          1766 => x"55",
          1767 => x"80",
          1768 => x"39",
          1769 => x"d9",
          1770 => x"80",
          1771 => x"27",
          1772 => x"80",
          1773 => x"89",
          1774 => x"70",
          1775 => x"55",
          1776 => x"70",
          1777 => x"55",
          1778 => x"27",
          1779 => x"14",
          1780 => x"06",
          1781 => x"74",
          1782 => x"73",
          1783 => x"38",
          1784 => x"14",
          1785 => x"05",
          1786 => x"08",
          1787 => x"54",
          1788 => x"39",
          1789 => x"84",
          1790 => x"55",
          1791 => x"81",
          1792 => x"de",
          1793 => x"3d",
          1794 => x"3d",
          1795 => x"5a",
          1796 => x"7a",
          1797 => x"08",
          1798 => x"53",
          1799 => x"09",
          1800 => x"38",
          1801 => x"0c",
          1802 => x"ad",
          1803 => x"06",
          1804 => x"76",
          1805 => x"0c",
          1806 => x"33",
          1807 => x"73",
          1808 => x"81",
          1809 => x"38",
          1810 => x"05",
          1811 => x"08",
          1812 => x"53",
          1813 => x"2e",
          1814 => x"57",
          1815 => x"2e",
          1816 => x"39",
          1817 => x"13",
          1818 => x"08",
          1819 => x"53",
          1820 => x"55",
          1821 => x"80",
          1822 => x"14",
          1823 => x"88",
          1824 => x"27",
          1825 => x"eb",
          1826 => x"53",
          1827 => x"89",
          1828 => x"38",
          1829 => x"55",
          1830 => x"8a",
          1831 => x"a0",
          1832 => x"c2",
          1833 => x"74",
          1834 => x"e0",
          1835 => x"ff",
          1836 => x"d0",
          1837 => x"ff",
          1838 => x"90",
          1839 => x"38",
          1840 => x"81",
          1841 => x"53",
          1842 => x"ca",
          1843 => x"27",
          1844 => x"77",
          1845 => x"08",
          1846 => x"0c",
          1847 => x"33",
          1848 => x"ff",
          1849 => x"80",
          1850 => x"74",
          1851 => x"79",
          1852 => x"74",
          1853 => x"0c",
          1854 => x"04",
          1855 => x"02",
          1856 => x"51",
          1857 => x"72",
          1858 => x"81",
          1859 => x"33",
          1860 => x"de",
          1861 => x"3d",
          1862 => x"3d",
          1863 => x"05",
          1864 => x"05",
          1865 => x"56",
          1866 => x"72",
          1867 => x"e0",
          1868 => x"2b",
          1869 => x"8c",
          1870 => x"88",
          1871 => x"2e",
          1872 => x"88",
          1873 => x"0c",
          1874 => x"8c",
          1875 => x"71",
          1876 => x"87",
          1877 => x"0c",
          1878 => x"08",
          1879 => x"51",
          1880 => x"2e",
          1881 => x"c0",
          1882 => x"51",
          1883 => x"71",
          1884 => x"80",
          1885 => x"92",
          1886 => x"98",
          1887 => x"70",
          1888 => x"38",
          1889 => x"e8",
          1890 => x"db",
          1891 => x"51",
          1892 => x"c0",
          1893 => x"0d",
          1894 => x"0d",
          1895 => x"02",
          1896 => x"05",
          1897 => x"58",
          1898 => x"52",
          1899 => x"3f",
          1900 => x"08",
          1901 => x"54",
          1902 => x"be",
          1903 => x"75",
          1904 => x"c0",
          1905 => x"87",
          1906 => x"12",
          1907 => x"84",
          1908 => x"40",
          1909 => x"85",
          1910 => x"98",
          1911 => x"7d",
          1912 => x"0c",
          1913 => x"85",
          1914 => x"06",
          1915 => x"71",
          1916 => x"38",
          1917 => x"71",
          1918 => x"05",
          1919 => x"19",
          1920 => x"a2",
          1921 => x"71",
          1922 => x"38",
          1923 => x"83",
          1924 => x"38",
          1925 => x"8a",
          1926 => x"98",
          1927 => x"71",
          1928 => x"c0",
          1929 => x"52",
          1930 => x"87",
          1931 => x"80",
          1932 => x"81",
          1933 => x"c0",
          1934 => x"53",
          1935 => x"82",
          1936 => x"71",
          1937 => x"1a",
          1938 => x"84",
          1939 => x"19",
          1940 => x"06",
          1941 => x"79",
          1942 => x"38",
          1943 => x"80",
          1944 => x"87",
          1945 => x"26",
          1946 => x"73",
          1947 => x"06",
          1948 => x"2e",
          1949 => x"52",
          1950 => x"81",
          1951 => x"8f",
          1952 => x"f3",
          1953 => x"62",
          1954 => x"05",
          1955 => x"57",
          1956 => x"83",
          1957 => x"52",
          1958 => x"3f",
          1959 => x"08",
          1960 => x"54",
          1961 => x"2e",
          1962 => x"81",
          1963 => x"74",
          1964 => x"c0",
          1965 => x"87",
          1966 => x"12",
          1967 => x"84",
          1968 => x"5f",
          1969 => x"0b",
          1970 => x"8c",
          1971 => x"0c",
          1972 => x"80",
          1973 => x"70",
          1974 => x"81",
          1975 => x"54",
          1976 => x"8c",
          1977 => x"81",
          1978 => x"7c",
          1979 => x"58",
          1980 => x"70",
          1981 => x"52",
          1982 => x"8a",
          1983 => x"98",
          1984 => x"71",
          1985 => x"c0",
          1986 => x"52",
          1987 => x"87",
          1988 => x"80",
          1989 => x"81",
          1990 => x"c0",
          1991 => x"53",
          1992 => x"82",
          1993 => x"71",
          1994 => x"19",
          1995 => x"81",
          1996 => x"ff",
          1997 => x"19",
          1998 => x"78",
          1999 => x"38",
          2000 => x"80",
          2001 => x"87",
          2002 => x"26",
          2003 => x"73",
          2004 => x"06",
          2005 => x"2e",
          2006 => x"52",
          2007 => x"81",
          2008 => x"8f",
          2009 => x"f6",
          2010 => x"02",
          2011 => x"05",
          2012 => x"05",
          2013 => x"71",
          2014 => x"57",
          2015 => x"81",
          2016 => x"81",
          2017 => x"54",
          2018 => x"38",
          2019 => x"c0",
          2020 => x"81",
          2021 => x"2e",
          2022 => x"71",
          2023 => x"38",
          2024 => x"87",
          2025 => x"11",
          2026 => x"80",
          2027 => x"80",
          2028 => x"83",
          2029 => x"38",
          2030 => x"72",
          2031 => x"2a",
          2032 => x"51",
          2033 => x"80",
          2034 => x"87",
          2035 => x"08",
          2036 => x"38",
          2037 => x"8c",
          2038 => x"96",
          2039 => x"0c",
          2040 => x"8c",
          2041 => x"08",
          2042 => x"51",
          2043 => x"38",
          2044 => x"56",
          2045 => x"80",
          2046 => x"85",
          2047 => x"77",
          2048 => x"83",
          2049 => x"75",
          2050 => x"de",
          2051 => x"3d",
          2052 => x"3d",
          2053 => x"11",
          2054 => x"71",
          2055 => x"81",
          2056 => x"53",
          2057 => x"0d",
          2058 => x"0d",
          2059 => x"33",
          2060 => x"71",
          2061 => x"88",
          2062 => x"14",
          2063 => x"07",
          2064 => x"33",
          2065 => x"de",
          2066 => x"53",
          2067 => x"52",
          2068 => x"04",
          2069 => x"73",
          2070 => x"92",
          2071 => x"52",
          2072 => x"81",
          2073 => x"70",
          2074 => x"70",
          2075 => x"3d",
          2076 => x"3d",
          2077 => x"52",
          2078 => x"70",
          2079 => x"34",
          2080 => x"51",
          2081 => x"81",
          2082 => x"70",
          2083 => x"70",
          2084 => x"05",
          2085 => x"88",
          2086 => x"72",
          2087 => x"0d",
          2088 => x"0d",
          2089 => x"54",
          2090 => x"80",
          2091 => x"71",
          2092 => x"53",
          2093 => x"81",
          2094 => x"ff",
          2095 => x"39",
          2096 => x"04",
          2097 => x"75",
          2098 => x"52",
          2099 => x"70",
          2100 => x"34",
          2101 => x"70",
          2102 => x"3d",
          2103 => x"3d",
          2104 => x"79",
          2105 => x"74",
          2106 => x"56",
          2107 => x"81",
          2108 => x"71",
          2109 => x"16",
          2110 => x"52",
          2111 => x"86",
          2112 => x"2e",
          2113 => x"81",
          2114 => x"86",
          2115 => x"fe",
          2116 => x"76",
          2117 => x"39",
          2118 => x"8a",
          2119 => x"51",
          2120 => x"71",
          2121 => x"33",
          2122 => x"0c",
          2123 => x"04",
          2124 => x"de",
          2125 => x"80",
          2126 => x"c0",
          2127 => x"3d",
          2128 => x"80",
          2129 => x"33",
          2130 => x"7a",
          2131 => x"38",
          2132 => x"16",
          2133 => x"16",
          2134 => x"17",
          2135 => x"fa",
          2136 => x"de",
          2137 => x"2e",
          2138 => x"b7",
          2139 => x"c0",
          2140 => x"34",
          2141 => x"70",
          2142 => x"31",
          2143 => x"59",
          2144 => x"77",
          2145 => x"82",
          2146 => x"74",
          2147 => x"81",
          2148 => x"81",
          2149 => x"53",
          2150 => x"16",
          2151 => x"e3",
          2152 => x"81",
          2153 => x"de",
          2154 => x"3d",
          2155 => x"3d",
          2156 => x"56",
          2157 => x"74",
          2158 => x"2e",
          2159 => x"51",
          2160 => x"81",
          2161 => x"57",
          2162 => x"08",
          2163 => x"54",
          2164 => x"16",
          2165 => x"33",
          2166 => x"3f",
          2167 => x"08",
          2168 => x"38",
          2169 => x"57",
          2170 => x"0c",
          2171 => x"c0",
          2172 => x"0d",
          2173 => x"0d",
          2174 => x"57",
          2175 => x"81",
          2176 => x"58",
          2177 => x"08",
          2178 => x"76",
          2179 => x"83",
          2180 => x"06",
          2181 => x"84",
          2182 => x"78",
          2183 => x"81",
          2184 => x"38",
          2185 => x"81",
          2186 => x"52",
          2187 => x"52",
          2188 => x"3f",
          2189 => x"52",
          2190 => x"51",
          2191 => x"84",
          2192 => x"d2",
          2193 => x"fc",
          2194 => x"8a",
          2195 => x"52",
          2196 => x"51",
          2197 => x"90",
          2198 => x"84",
          2199 => x"fc",
          2200 => x"17",
          2201 => x"a0",
          2202 => x"86",
          2203 => x"08",
          2204 => x"b0",
          2205 => x"55",
          2206 => x"81",
          2207 => x"f8",
          2208 => x"84",
          2209 => x"53",
          2210 => x"17",
          2211 => x"d7",
          2212 => x"c0",
          2213 => x"83",
          2214 => x"77",
          2215 => x"0c",
          2216 => x"04",
          2217 => x"77",
          2218 => x"12",
          2219 => x"55",
          2220 => x"56",
          2221 => x"8d",
          2222 => x"22",
          2223 => x"ac",
          2224 => x"57",
          2225 => x"de",
          2226 => x"3d",
          2227 => x"3d",
          2228 => x"70",
          2229 => x"57",
          2230 => x"81",
          2231 => x"98",
          2232 => x"81",
          2233 => x"74",
          2234 => x"72",
          2235 => x"f5",
          2236 => x"24",
          2237 => x"81",
          2238 => x"81",
          2239 => x"83",
          2240 => x"38",
          2241 => x"76",
          2242 => x"70",
          2243 => x"16",
          2244 => x"74",
          2245 => x"96",
          2246 => x"c0",
          2247 => x"38",
          2248 => x"06",
          2249 => x"33",
          2250 => x"89",
          2251 => x"08",
          2252 => x"54",
          2253 => x"fc",
          2254 => x"de",
          2255 => x"fe",
          2256 => x"ff",
          2257 => x"11",
          2258 => x"2b",
          2259 => x"81",
          2260 => x"2a",
          2261 => x"51",
          2262 => x"e2",
          2263 => x"ff",
          2264 => x"da",
          2265 => x"2a",
          2266 => x"05",
          2267 => x"fc",
          2268 => x"de",
          2269 => x"c6",
          2270 => x"83",
          2271 => x"05",
          2272 => x"f9",
          2273 => x"de",
          2274 => x"ff",
          2275 => x"ae",
          2276 => x"2a",
          2277 => x"05",
          2278 => x"fc",
          2279 => x"de",
          2280 => x"38",
          2281 => x"83",
          2282 => x"05",
          2283 => x"f8",
          2284 => x"de",
          2285 => x"0a",
          2286 => x"39",
          2287 => x"81",
          2288 => x"89",
          2289 => x"f8",
          2290 => x"7c",
          2291 => x"56",
          2292 => x"77",
          2293 => x"38",
          2294 => x"08",
          2295 => x"38",
          2296 => x"72",
          2297 => x"9d",
          2298 => x"24",
          2299 => x"81",
          2300 => x"82",
          2301 => x"83",
          2302 => x"38",
          2303 => x"76",
          2304 => x"70",
          2305 => x"18",
          2306 => x"76",
          2307 => x"9e",
          2308 => x"c0",
          2309 => x"de",
          2310 => x"d9",
          2311 => x"ff",
          2312 => x"05",
          2313 => x"81",
          2314 => x"54",
          2315 => x"80",
          2316 => x"77",
          2317 => x"f0",
          2318 => x"8f",
          2319 => x"51",
          2320 => x"34",
          2321 => x"17",
          2322 => x"2a",
          2323 => x"05",
          2324 => x"fa",
          2325 => x"de",
          2326 => x"81",
          2327 => x"81",
          2328 => x"83",
          2329 => x"b4",
          2330 => x"2a",
          2331 => x"8f",
          2332 => x"2a",
          2333 => x"f0",
          2334 => x"06",
          2335 => x"72",
          2336 => x"ec",
          2337 => x"2a",
          2338 => x"05",
          2339 => x"fa",
          2340 => x"de",
          2341 => x"81",
          2342 => x"80",
          2343 => x"83",
          2344 => x"52",
          2345 => x"fe",
          2346 => x"b4",
          2347 => x"a4",
          2348 => x"76",
          2349 => x"17",
          2350 => x"75",
          2351 => x"3f",
          2352 => x"08",
          2353 => x"c0",
          2354 => x"77",
          2355 => x"77",
          2356 => x"fc",
          2357 => x"b4",
          2358 => x"51",
          2359 => x"c9",
          2360 => x"c0",
          2361 => x"06",
          2362 => x"72",
          2363 => x"3f",
          2364 => x"17",
          2365 => x"de",
          2366 => x"3d",
          2367 => x"3d",
          2368 => x"7e",
          2369 => x"56",
          2370 => x"75",
          2371 => x"74",
          2372 => x"27",
          2373 => x"80",
          2374 => x"ff",
          2375 => x"75",
          2376 => x"3f",
          2377 => x"08",
          2378 => x"c0",
          2379 => x"38",
          2380 => x"54",
          2381 => x"81",
          2382 => x"39",
          2383 => x"08",
          2384 => x"39",
          2385 => x"51",
          2386 => x"81",
          2387 => x"58",
          2388 => x"08",
          2389 => x"c7",
          2390 => x"c0",
          2391 => x"d2",
          2392 => x"c0",
          2393 => x"cf",
          2394 => x"74",
          2395 => x"fc",
          2396 => x"de",
          2397 => x"38",
          2398 => x"fe",
          2399 => x"08",
          2400 => x"74",
          2401 => x"38",
          2402 => x"17",
          2403 => x"33",
          2404 => x"73",
          2405 => x"77",
          2406 => x"26",
          2407 => x"80",
          2408 => x"de",
          2409 => x"3d",
          2410 => x"3d",
          2411 => x"71",
          2412 => x"5b",
          2413 => x"8c",
          2414 => x"77",
          2415 => x"38",
          2416 => x"78",
          2417 => x"81",
          2418 => x"79",
          2419 => x"f9",
          2420 => x"55",
          2421 => x"c0",
          2422 => x"e0",
          2423 => x"c0",
          2424 => x"de",
          2425 => x"2e",
          2426 => x"98",
          2427 => x"de",
          2428 => x"82",
          2429 => x"58",
          2430 => x"70",
          2431 => x"80",
          2432 => x"38",
          2433 => x"09",
          2434 => x"e2",
          2435 => x"56",
          2436 => x"76",
          2437 => x"82",
          2438 => x"7a",
          2439 => x"3f",
          2440 => x"de",
          2441 => x"2e",
          2442 => x"86",
          2443 => x"c0",
          2444 => x"de",
          2445 => x"70",
          2446 => x"07",
          2447 => x"7c",
          2448 => x"c0",
          2449 => x"51",
          2450 => x"81",
          2451 => x"de",
          2452 => x"2e",
          2453 => x"17",
          2454 => x"74",
          2455 => x"73",
          2456 => x"27",
          2457 => x"58",
          2458 => x"80",
          2459 => x"56",
          2460 => x"98",
          2461 => x"26",
          2462 => x"56",
          2463 => x"81",
          2464 => x"52",
          2465 => x"c6",
          2466 => x"c0",
          2467 => x"b8",
          2468 => x"81",
          2469 => x"81",
          2470 => x"06",
          2471 => x"de",
          2472 => x"81",
          2473 => x"09",
          2474 => x"72",
          2475 => x"70",
          2476 => x"51",
          2477 => x"80",
          2478 => x"78",
          2479 => x"06",
          2480 => x"73",
          2481 => x"39",
          2482 => x"52",
          2483 => x"f7",
          2484 => x"c0",
          2485 => x"c0",
          2486 => x"81",
          2487 => x"07",
          2488 => x"55",
          2489 => x"2e",
          2490 => x"80",
          2491 => x"75",
          2492 => x"76",
          2493 => x"3f",
          2494 => x"08",
          2495 => x"38",
          2496 => x"0c",
          2497 => x"fe",
          2498 => x"08",
          2499 => x"74",
          2500 => x"ff",
          2501 => x"0c",
          2502 => x"81",
          2503 => x"84",
          2504 => x"39",
          2505 => x"81",
          2506 => x"8c",
          2507 => x"8c",
          2508 => x"c0",
          2509 => x"39",
          2510 => x"55",
          2511 => x"c0",
          2512 => x"0d",
          2513 => x"0d",
          2514 => x"55",
          2515 => x"81",
          2516 => x"58",
          2517 => x"de",
          2518 => x"d8",
          2519 => x"74",
          2520 => x"3f",
          2521 => x"08",
          2522 => x"08",
          2523 => x"59",
          2524 => x"77",
          2525 => x"70",
          2526 => x"c8",
          2527 => x"84",
          2528 => x"56",
          2529 => x"58",
          2530 => x"97",
          2531 => x"75",
          2532 => x"52",
          2533 => x"51",
          2534 => x"81",
          2535 => x"80",
          2536 => x"8a",
          2537 => x"32",
          2538 => x"72",
          2539 => x"2a",
          2540 => x"56",
          2541 => x"c0",
          2542 => x"0d",
          2543 => x"0d",
          2544 => x"08",
          2545 => x"74",
          2546 => x"26",
          2547 => x"74",
          2548 => x"72",
          2549 => x"74",
          2550 => x"88",
          2551 => x"73",
          2552 => x"33",
          2553 => x"27",
          2554 => x"16",
          2555 => x"9b",
          2556 => x"2a",
          2557 => x"88",
          2558 => x"58",
          2559 => x"80",
          2560 => x"16",
          2561 => x"0c",
          2562 => x"8a",
          2563 => x"89",
          2564 => x"72",
          2565 => x"38",
          2566 => x"51",
          2567 => x"81",
          2568 => x"54",
          2569 => x"08",
          2570 => x"38",
          2571 => x"de",
          2572 => x"8b",
          2573 => x"08",
          2574 => x"08",
          2575 => x"82",
          2576 => x"74",
          2577 => x"cb",
          2578 => x"75",
          2579 => x"3f",
          2580 => x"08",
          2581 => x"73",
          2582 => x"98",
          2583 => x"82",
          2584 => x"2e",
          2585 => x"39",
          2586 => x"39",
          2587 => x"13",
          2588 => x"74",
          2589 => x"16",
          2590 => x"18",
          2591 => x"77",
          2592 => x"0c",
          2593 => x"04",
          2594 => x"7a",
          2595 => x"12",
          2596 => x"59",
          2597 => x"80",
          2598 => x"86",
          2599 => x"98",
          2600 => x"14",
          2601 => x"55",
          2602 => x"81",
          2603 => x"83",
          2604 => x"77",
          2605 => x"81",
          2606 => x"0c",
          2607 => x"55",
          2608 => x"76",
          2609 => x"17",
          2610 => x"74",
          2611 => x"9b",
          2612 => x"39",
          2613 => x"ff",
          2614 => x"2a",
          2615 => x"81",
          2616 => x"52",
          2617 => x"e6",
          2618 => x"c0",
          2619 => x"55",
          2620 => x"de",
          2621 => x"80",
          2622 => x"55",
          2623 => x"08",
          2624 => x"f4",
          2625 => x"08",
          2626 => x"08",
          2627 => x"38",
          2628 => x"77",
          2629 => x"84",
          2630 => x"39",
          2631 => x"52",
          2632 => x"86",
          2633 => x"c0",
          2634 => x"55",
          2635 => x"08",
          2636 => x"c4",
          2637 => x"81",
          2638 => x"81",
          2639 => x"81",
          2640 => x"c0",
          2641 => x"b0",
          2642 => x"c0",
          2643 => x"51",
          2644 => x"81",
          2645 => x"a0",
          2646 => x"15",
          2647 => x"75",
          2648 => x"3f",
          2649 => x"08",
          2650 => x"76",
          2651 => x"77",
          2652 => x"9c",
          2653 => x"55",
          2654 => x"c0",
          2655 => x"0d",
          2656 => x"0d",
          2657 => x"08",
          2658 => x"80",
          2659 => x"fc",
          2660 => x"de",
          2661 => x"81",
          2662 => x"80",
          2663 => x"de",
          2664 => x"98",
          2665 => x"78",
          2666 => x"3f",
          2667 => x"08",
          2668 => x"c0",
          2669 => x"38",
          2670 => x"08",
          2671 => x"70",
          2672 => x"58",
          2673 => x"2e",
          2674 => x"83",
          2675 => x"81",
          2676 => x"55",
          2677 => x"81",
          2678 => x"07",
          2679 => x"2e",
          2680 => x"16",
          2681 => x"2e",
          2682 => x"88",
          2683 => x"81",
          2684 => x"56",
          2685 => x"51",
          2686 => x"81",
          2687 => x"54",
          2688 => x"08",
          2689 => x"9b",
          2690 => x"2e",
          2691 => x"83",
          2692 => x"73",
          2693 => x"0c",
          2694 => x"04",
          2695 => x"76",
          2696 => x"54",
          2697 => x"81",
          2698 => x"83",
          2699 => x"76",
          2700 => x"53",
          2701 => x"2e",
          2702 => x"90",
          2703 => x"51",
          2704 => x"81",
          2705 => x"90",
          2706 => x"53",
          2707 => x"c0",
          2708 => x"0d",
          2709 => x"0d",
          2710 => x"83",
          2711 => x"54",
          2712 => x"55",
          2713 => x"3f",
          2714 => x"51",
          2715 => x"2e",
          2716 => x"8b",
          2717 => x"2a",
          2718 => x"51",
          2719 => x"86",
          2720 => x"f7",
          2721 => x"7d",
          2722 => x"75",
          2723 => x"98",
          2724 => x"2e",
          2725 => x"98",
          2726 => x"78",
          2727 => x"3f",
          2728 => x"08",
          2729 => x"c0",
          2730 => x"38",
          2731 => x"70",
          2732 => x"73",
          2733 => x"58",
          2734 => x"8b",
          2735 => x"bf",
          2736 => x"ff",
          2737 => x"53",
          2738 => x"34",
          2739 => x"08",
          2740 => x"e5",
          2741 => x"81",
          2742 => x"2e",
          2743 => x"70",
          2744 => x"57",
          2745 => x"9e",
          2746 => x"2e",
          2747 => x"de",
          2748 => x"df",
          2749 => x"72",
          2750 => x"81",
          2751 => x"76",
          2752 => x"2e",
          2753 => x"52",
          2754 => x"fc",
          2755 => x"c0",
          2756 => x"de",
          2757 => x"38",
          2758 => x"fe",
          2759 => x"39",
          2760 => x"16",
          2761 => x"de",
          2762 => x"3d",
          2763 => x"3d",
          2764 => x"08",
          2765 => x"52",
          2766 => x"c5",
          2767 => x"c0",
          2768 => x"de",
          2769 => x"38",
          2770 => x"52",
          2771 => x"de",
          2772 => x"c0",
          2773 => x"de",
          2774 => x"38",
          2775 => x"de",
          2776 => x"9c",
          2777 => x"ea",
          2778 => x"53",
          2779 => x"9c",
          2780 => x"ea",
          2781 => x"0b",
          2782 => x"74",
          2783 => x"0c",
          2784 => x"04",
          2785 => x"75",
          2786 => x"12",
          2787 => x"53",
          2788 => x"9a",
          2789 => x"c0",
          2790 => x"9c",
          2791 => x"e5",
          2792 => x"0b",
          2793 => x"85",
          2794 => x"fa",
          2795 => x"7a",
          2796 => x"0b",
          2797 => x"98",
          2798 => x"2e",
          2799 => x"80",
          2800 => x"55",
          2801 => x"17",
          2802 => x"33",
          2803 => x"51",
          2804 => x"2e",
          2805 => x"85",
          2806 => x"06",
          2807 => x"e5",
          2808 => x"2e",
          2809 => x"8b",
          2810 => x"70",
          2811 => x"34",
          2812 => x"71",
          2813 => x"05",
          2814 => x"15",
          2815 => x"27",
          2816 => x"15",
          2817 => x"80",
          2818 => x"34",
          2819 => x"52",
          2820 => x"88",
          2821 => x"17",
          2822 => x"52",
          2823 => x"3f",
          2824 => x"08",
          2825 => x"12",
          2826 => x"3f",
          2827 => x"08",
          2828 => x"98",
          2829 => x"da",
          2830 => x"c0",
          2831 => x"23",
          2832 => x"04",
          2833 => x"7f",
          2834 => x"5b",
          2835 => x"33",
          2836 => x"73",
          2837 => x"38",
          2838 => x"80",
          2839 => x"38",
          2840 => x"8c",
          2841 => x"08",
          2842 => x"aa",
          2843 => x"41",
          2844 => x"33",
          2845 => x"73",
          2846 => x"81",
          2847 => x"81",
          2848 => x"dc",
          2849 => x"70",
          2850 => x"07",
          2851 => x"73",
          2852 => x"88",
          2853 => x"70",
          2854 => x"73",
          2855 => x"38",
          2856 => x"ab",
          2857 => x"52",
          2858 => x"91",
          2859 => x"c0",
          2860 => x"98",
          2861 => x"61",
          2862 => x"5a",
          2863 => x"a0",
          2864 => x"e7",
          2865 => x"70",
          2866 => x"79",
          2867 => x"73",
          2868 => x"81",
          2869 => x"38",
          2870 => x"33",
          2871 => x"ae",
          2872 => x"70",
          2873 => x"82",
          2874 => x"51",
          2875 => x"54",
          2876 => x"79",
          2877 => x"74",
          2878 => x"57",
          2879 => x"af",
          2880 => x"70",
          2881 => x"51",
          2882 => x"dc",
          2883 => x"73",
          2884 => x"38",
          2885 => x"82",
          2886 => x"19",
          2887 => x"54",
          2888 => x"82",
          2889 => x"54",
          2890 => x"78",
          2891 => x"81",
          2892 => x"54",
          2893 => x"81",
          2894 => x"af",
          2895 => x"77",
          2896 => x"70",
          2897 => x"25",
          2898 => x"07",
          2899 => x"51",
          2900 => x"2e",
          2901 => x"39",
          2902 => x"80",
          2903 => x"33",
          2904 => x"73",
          2905 => x"81",
          2906 => x"81",
          2907 => x"dc",
          2908 => x"70",
          2909 => x"07",
          2910 => x"73",
          2911 => x"b5",
          2912 => x"2e",
          2913 => x"83",
          2914 => x"76",
          2915 => x"07",
          2916 => x"2e",
          2917 => x"8b",
          2918 => x"77",
          2919 => x"30",
          2920 => x"71",
          2921 => x"53",
          2922 => x"55",
          2923 => x"38",
          2924 => x"5c",
          2925 => x"75",
          2926 => x"73",
          2927 => x"38",
          2928 => x"06",
          2929 => x"11",
          2930 => x"75",
          2931 => x"3f",
          2932 => x"08",
          2933 => x"38",
          2934 => x"33",
          2935 => x"54",
          2936 => x"e6",
          2937 => x"de",
          2938 => x"2e",
          2939 => x"ff",
          2940 => x"74",
          2941 => x"38",
          2942 => x"75",
          2943 => x"17",
          2944 => x"57",
          2945 => x"a7",
          2946 => x"81",
          2947 => x"e5",
          2948 => x"de",
          2949 => x"38",
          2950 => x"54",
          2951 => x"89",
          2952 => x"70",
          2953 => x"57",
          2954 => x"54",
          2955 => x"81",
          2956 => x"f7",
          2957 => x"7e",
          2958 => x"2e",
          2959 => x"33",
          2960 => x"e5",
          2961 => x"06",
          2962 => x"7a",
          2963 => x"a0",
          2964 => x"38",
          2965 => x"55",
          2966 => x"84",
          2967 => x"39",
          2968 => x"8b",
          2969 => x"7b",
          2970 => x"7a",
          2971 => x"3f",
          2972 => x"08",
          2973 => x"c0",
          2974 => x"38",
          2975 => x"52",
          2976 => x"aa",
          2977 => x"c0",
          2978 => x"de",
          2979 => x"c2",
          2980 => x"08",
          2981 => x"55",
          2982 => x"ff",
          2983 => x"15",
          2984 => x"54",
          2985 => x"34",
          2986 => x"70",
          2987 => x"81",
          2988 => x"58",
          2989 => x"8b",
          2990 => x"74",
          2991 => x"3f",
          2992 => x"08",
          2993 => x"38",
          2994 => x"51",
          2995 => x"ff",
          2996 => x"ab",
          2997 => x"55",
          2998 => x"bb",
          2999 => x"2e",
          3000 => x"80",
          3001 => x"85",
          3002 => x"06",
          3003 => x"58",
          3004 => x"80",
          3005 => x"75",
          3006 => x"73",
          3007 => x"b5",
          3008 => x"0b",
          3009 => x"80",
          3010 => x"39",
          3011 => x"54",
          3012 => x"85",
          3013 => x"75",
          3014 => x"81",
          3015 => x"73",
          3016 => x"1b",
          3017 => x"2a",
          3018 => x"51",
          3019 => x"80",
          3020 => x"90",
          3021 => x"ff",
          3022 => x"05",
          3023 => x"f5",
          3024 => x"de",
          3025 => x"1c",
          3026 => x"39",
          3027 => x"c0",
          3028 => x"0d",
          3029 => x"0d",
          3030 => x"7b",
          3031 => x"73",
          3032 => x"55",
          3033 => x"2e",
          3034 => x"75",
          3035 => x"57",
          3036 => x"26",
          3037 => x"ba",
          3038 => x"70",
          3039 => x"ba",
          3040 => x"06",
          3041 => x"73",
          3042 => x"70",
          3043 => x"51",
          3044 => x"89",
          3045 => x"82",
          3046 => x"ff",
          3047 => x"56",
          3048 => x"2e",
          3049 => x"80",
          3050 => x"a4",
          3051 => x"08",
          3052 => x"76",
          3053 => x"58",
          3054 => x"81",
          3055 => x"ff",
          3056 => x"53",
          3057 => x"26",
          3058 => x"13",
          3059 => x"06",
          3060 => x"9f",
          3061 => x"99",
          3062 => x"e0",
          3063 => x"ff",
          3064 => x"72",
          3065 => x"2a",
          3066 => x"72",
          3067 => x"06",
          3068 => x"ff",
          3069 => x"30",
          3070 => x"70",
          3071 => x"07",
          3072 => x"9f",
          3073 => x"54",
          3074 => x"80",
          3075 => x"81",
          3076 => x"59",
          3077 => x"25",
          3078 => x"8b",
          3079 => x"24",
          3080 => x"76",
          3081 => x"78",
          3082 => x"81",
          3083 => x"51",
          3084 => x"c0",
          3085 => x"0d",
          3086 => x"0d",
          3087 => x"0b",
          3088 => x"ff",
          3089 => x"0c",
          3090 => x"51",
          3091 => x"84",
          3092 => x"c0",
          3093 => x"38",
          3094 => x"51",
          3095 => x"81",
          3096 => x"83",
          3097 => x"54",
          3098 => x"82",
          3099 => x"09",
          3100 => x"e3",
          3101 => x"b4",
          3102 => x"57",
          3103 => x"2e",
          3104 => x"83",
          3105 => x"74",
          3106 => x"70",
          3107 => x"25",
          3108 => x"51",
          3109 => x"38",
          3110 => x"2e",
          3111 => x"b5",
          3112 => x"81",
          3113 => x"80",
          3114 => x"e0",
          3115 => x"de",
          3116 => x"81",
          3117 => x"80",
          3118 => x"85",
          3119 => x"e8",
          3120 => x"16",
          3121 => x"3f",
          3122 => x"08",
          3123 => x"c0",
          3124 => x"83",
          3125 => x"74",
          3126 => x"0c",
          3127 => x"04",
          3128 => x"61",
          3129 => x"80",
          3130 => x"58",
          3131 => x"0c",
          3132 => x"e1",
          3133 => x"c0",
          3134 => x"56",
          3135 => x"de",
          3136 => x"86",
          3137 => x"de",
          3138 => x"29",
          3139 => x"05",
          3140 => x"53",
          3141 => x"80",
          3142 => x"38",
          3143 => x"76",
          3144 => x"74",
          3145 => x"72",
          3146 => x"38",
          3147 => x"51",
          3148 => x"81",
          3149 => x"81",
          3150 => x"81",
          3151 => x"72",
          3152 => x"80",
          3153 => x"38",
          3154 => x"70",
          3155 => x"53",
          3156 => x"86",
          3157 => x"a7",
          3158 => x"34",
          3159 => x"34",
          3160 => x"14",
          3161 => x"b2",
          3162 => x"c0",
          3163 => x"06",
          3164 => x"54",
          3165 => x"72",
          3166 => x"76",
          3167 => x"38",
          3168 => x"70",
          3169 => x"53",
          3170 => x"85",
          3171 => x"70",
          3172 => x"5b",
          3173 => x"81",
          3174 => x"81",
          3175 => x"76",
          3176 => x"81",
          3177 => x"38",
          3178 => x"56",
          3179 => x"83",
          3180 => x"70",
          3181 => x"80",
          3182 => x"83",
          3183 => x"dc",
          3184 => x"de",
          3185 => x"76",
          3186 => x"05",
          3187 => x"16",
          3188 => x"56",
          3189 => x"d7",
          3190 => x"8d",
          3191 => x"72",
          3192 => x"54",
          3193 => x"57",
          3194 => x"95",
          3195 => x"73",
          3196 => x"3f",
          3197 => x"08",
          3198 => x"57",
          3199 => x"89",
          3200 => x"56",
          3201 => x"d7",
          3202 => x"76",
          3203 => x"f1",
          3204 => x"76",
          3205 => x"e9",
          3206 => x"51",
          3207 => x"81",
          3208 => x"83",
          3209 => x"53",
          3210 => x"2e",
          3211 => x"84",
          3212 => x"ca",
          3213 => x"da",
          3214 => x"c0",
          3215 => x"ff",
          3216 => x"8d",
          3217 => x"14",
          3218 => x"3f",
          3219 => x"08",
          3220 => x"15",
          3221 => x"14",
          3222 => x"34",
          3223 => x"33",
          3224 => x"81",
          3225 => x"54",
          3226 => x"72",
          3227 => x"91",
          3228 => x"ff",
          3229 => x"29",
          3230 => x"33",
          3231 => x"72",
          3232 => x"72",
          3233 => x"38",
          3234 => x"06",
          3235 => x"2e",
          3236 => x"56",
          3237 => x"80",
          3238 => x"da",
          3239 => x"de",
          3240 => x"81",
          3241 => x"88",
          3242 => x"8f",
          3243 => x"56",
          3244 => x"38",
          3245 => x"51",
          3246 => x"81",
          3247 => x"83",
          3248 => x"55",
          3249 => x"80",
          3250 => x"da",
          3251 => x"de",
          3252 => x"80",
          3253 => x"da",
          3254 => x"de",
          3255 => x"ff",
          3256 => x"8d",
          3257 => x"2e",
          3258 => x"88",
          3259 => x"14",
          3260 => x"05",
          3261 => x"75",
          3262 => x"38",
          3263 => x"52",
          3264 => x"51",
          3265 => x"3f",
          3266 => x"08",
          3267 => x"c0",
          3268 => x"82",
          3269 => x"de",
          3270 => x"ff",
          3271 => x"26",
          3272 => x"57",
          3273 => x"f5",
          3274 => x"82",
          3275 => x"f5",
          3276 => x"81",
          3277 => x"8d",
          3278 => x"2e",
          3279 => x"82",
          3280 => x"16",
          3281 => x"16",
          3282 => x"70",
          3283 => x"7a",
          3284 => x"0c",
          3285 => x"83",
          3286 => x"06",
          3287 => x"de",
          3288 => x"ae",
          3289 => x"c0",
          3290 => x"ff",
          3291 => x"56",
          3292 => x"38",
          3293 => x"38",
          3294 => x"51",
          3295 => x"81",
          3296 => x"a8",
          3297 => x"82",
          3298 => x"39",
          3299 => x"80",
          3300 => x"38",
          3301 => x"15",
          3302 => x"53",
          3303 => x"8d",
          3304 => x"15",
          3305 => x"76",
          3306 => x"51",
          3307 => x"13",
          3308 => x"8d",
          3309 => x"15",
          3310 => x"c5",
          3311 => x"90",
          3312 => x"0b",
          3313 => x"ff",
          3314 => x"15",
          3315 => x"2e",
          3316 => x"81",
          3317 => x"e4",
          3318 => x"b6",
          3319 => x"c0",
          3320 => x"ff",
          3321 => x"81",
          3322 => x"06",
          3323 => x"81",
          3324 => x"51",
          3325 => x"81",
          3326 => x"80",
          3327 => x"de",
          3328 => x"15",
          3329 => x"14",
          3330 => x"3f",
          3331 => x"08",
          3332 => x"06",
          3333 => x"d4",
          3334 => x"81",
          3335 => x"38",
          3336 => x"d8",
          3337 => x"de",
          3338 => x"8b",
          3339 => x"2e",
          3340 => x"b3",
          3341 => x"14",
          3342 => x"3f",
          3343 => x"08",
          3344 => x"e4",
          3345 => x"81",
          3346 => x"84",
          3347 => x"d7",
          3348 => x"de",
          3349 => x"15",
          3350 => x"14",
          3351 => x"3f",
          3352 => x"08",
          3353 => x"76",
          3354 => x"de",
          3355 => x"05",
          3356 => x"de",
          3357 => x"86",
          3358 => x"0b",
          3359 => x"80",
          3360 => x"de",
          3361 => x"3d",
          3362 => x"3d",
          3363 => x"89",
          3364 => x"2e",
          3365 => x"08",
          3366 => x"2e",
          3367 => x"33",
          3368 => x"2e",
          3369 => x"13",
          3370 => x"22",
          3371 => x"76",
          3372 => x"06",
          3373 => x"13",
          3374 => x"c0",
          3375 => x"c0",
          3376 => x"52",
          3377 => x"71",
          3378 => x"55",
          3379 => x"53",
          3380 => x"0c",
          3381 => x"de",
          3382 => x"3d",
          3383 => x"3d",
          3384 => x"05",
          3385 => x"89",
          3386 => x"52",
          3387 => x"3f",
          3388 => x"0b",
          3389 => x"08",
          3390 => x"81",
          3391 => x"84",
          3392 => x"dc",
          3393 => x"55",
          3394 => x"2e",
          3395 => x"74",
          3396 => x"73",
          3397 => x"38",
          3398 => x"78",
          3399 => x"54",
          3400 => x"92",
          3401 => x"89",
          3402 => x"84",
          3403 => x"b0",
          3404 => x"c0",
          3405 => x"81",
          3406 => x"88",
          3407 => x"eb",
          3408 => x"02",
          3409 => x"e7",
          3410 => x"59",
          3411 => x"80",
          3412 => x"38",
          3413 => x"70",
          3414 => x"d0",
          3415 => x"3d",
          3416 => x"58",
          3417 => x"81",
          3418 => x"55",
          3419 => x"08",
          3420 => x"7a",
          3421 => x"8c",
          3422 => x"56",
          3423 => x"81",
          3424 => x"55",
          3425 => x"08",
          3426 => x"80",
          3427 => x"70",
          3428 => x"57",
          3429 => x"83",
          3430 => x"77",
          3431 => x"73",
          3432 => x"ab",
          3433 => x"2e",
          3434 => x"84",
          3435 => x"06",
          3436 => x"51",
          3437 => x"81",
          3438 => x"55",
          3439 => x"b2",
          3440 => x"06",
          3441 => x"b8",
          3442 => x"2a",
          3443 => x"51",
          3444 => x"2e",
          3445 => x"55",
          3446 => x"77",
          3447 => x"74",
          3448 => x"77",
          3449 => x"81",
          3450 => x"73",
          3451 => x"af",
          3452 => x"7a",
          3453 => x"3f",
          3454 => x"08",
          3455 => x"b2",
          3456 => x"8e",
          3457 => x"ea",
          3458 => x"a0",
          3459 => x"34",
          3460 => x"52",
          3461 => x"bd",
          3462 => x"62",
          3463 => x"d4",
          3464 => x"54",
          3465 => x"15",
          3466 => x"2e",
          3467 => x"7a",
          3468 => x"51",
          3469 => x"75",
          3470 => x"d4",
          3471 => x"be",
          3472 => x"c0",
          3473 => x"de",
          3474 => x"ca",
          3475 => x"74",
          3476 => x"02",
          3477 => x"70",
          3478 => x"81",
          3479 => x"56",
          3480 => x"86",
          3481 => x"82",
          3482 => x"81",
          3483 => x"06",
          3484 => x"80",
          3485 => x"75",
          3486 => x"73",
          3487 => x"38",
          3488 => x"92",
          3489 => x"7a",
          3490 => x"3f",
          3491 => x"08",
          3492 => x"8c",
          3493 => x"55",
          3494 => x"08",
          3495 => x"77",
          3496 => x"81",
          3497 => x"73",
          3498 => x"38",
          3499 => x"07",
          3500 => x"11",
          3501 => x"0c",
          3502 => x"0c",
          3503 => x"52",
          3504 => x"3f",
          3505 => x"08",
          3506 => x"08",
          3507 => x"63",
          3508 => x"5a",
          3509 => x"81",
          3510 => x"81",
          3511 => x"8c",
          3512 => x"7a",
          3513 => x"17",
          3514 => x"23",
          3515 => x"34",
          3516 => x"1a",
          3517 => x"9c",
          3518 => x"0b",
          3519 => x"77",
          3520 => x"81",
          3521 => x"73",
          3522 => x"8d",
          3523 => x"c0",
          3524 => x"81",
          3525 => x"de",
          3526 => x"1a",
          3527 => x"22",
          3528 => x"7b",
          3529 => x"a8",
          3530 => x"78",
          3531 => x"3f",
          3532 => x"08",
          3533 => x"c0",
          3534 => x"83",
          3535 => x"81",
          3536 => x"ff",
          3537 => x"06",
          3538 => x"55",
          3539 => x"56",
          3540 => x"76",
          3541 => x"51",
          3542 => x"27",
          3543 => x"70",
          3544 => x"5a",
          3545 => x"76",
          3546 => x"74",
          3547 => x"83",
          3548 => x"73",
          3549 => x"38",
          3550 => x"51",
          3551 => x"81",
          3552 => x"85",
          3553 => x"8e",
          3554 => x"2a",
          3555 => x"08",
          3556 => x"0c",
          3557 => x"79",
          3558 => x"73",
          3559 => x"0c",
          3560 => x"04",
          3561 => x"60",
          3562 => x"40",
          3563 => x"80",
          3564 => x"3d",
          3565 => x"78",
          3566 => x"3f",
          3567 => x"08",
          3568 => x"c0",
          3569 => x"91",
          3570 => x"74",
          3571 => x"38",
          3572 => x"c4",
          3573 => x"33",
          3574 => x"87",
          3575 => x"2e",
          3576 => x"95",
          3577 => x"91",
          3578 => x"56",
          3579 => x"81",
          3580 => x"34",
          3581 => x"a0",
          3582 => x"08",
          3583 => x"31",
          3584 => x"27",
          3585 => x"5c",
          3586 => x"82",
          3587 => x"19",
          3588 => x"ff",
          3589 => x"74",
          3590 => x"7e",
          3591 => x"ff",
          3592 => x"2a",
          3593 => x"79",
          3594 => x"87",
          3595 => x"08",
          3596 => x"98",
          3597 => x"78",
          3598 => x"3f",
          3599 => x"08",
          3600 => x"27",
          3601 => x"74",
          3602 => x"a3",
          3603 => x"1a",
          3604 => x"08",
          3605 => x"d4",
          3606 => x"de",
          3607 => x"2e",
          3608 => x"81",
          3609 => x"1a",
          3610 => x"59",
          3611 => x"2e",
          3612 => x"77",
          3613 => x"11",
          3614 => x"55",
          3615 => x"85",
          3616 => x"31",
          3617 => x"76",
          3618 => x"81",
          3619 => x"ca",
          3620 => x"de",
          3621 => x"d7",
          3622 => x"11",
          3623 => x"74",
          3624 => x"38",
          3625 => x"77",
          3626 => x"78",
          3627 => x"84",
          3628 => x"16",
          3629 => x"08",
          3630 => x"2b",
          3631 => x"cf",
          3632 => x"89",
          3633 => x"39",
          3634 => x"0c",
          3635 => x"83",
          3636 => x"80",
          3637 => x"55",
          3638 => x"83",
          3639 => x"9c",
          3640 => x"7e",
          3641 => x"3f",
          3642 => x"08",
          3643 => x"75",
          3644 => x"08",
          3645 => x"1f",
          3646 => x"7c",
          3647 => x"3f",
          3648 => x"7e",
          3649 => x"0c",
          3650 => x"1b",
          3651 => x"1c",
          3652 => x"fd",
          3653 => x"56",
          3654 => x"c0",
          3655 => x"0d",
          3656 => x"0d",
          3657 => x"64",
          3658 => x"58",
          3659 => x"90",
          3660 => x"52",
          3661 => x"d2",
          3662 => x"c0",
          3663 => x"de",
          3664 => x"38",
          3665 => x"55",
          3666 => x"86",
          3667 => x"83",
          3668 => x"18",
          3669 => x"2a",
          3670 => x"51",
          3671 => x"56",
          3672 => x"83",
          3673 => x"39",
          3674 => x"19",
          3675 => x"83",
          3676 => x"0b",
          3677 => x"81",
          3678 => x"39",
          3679 => x"7c",
          3680 => x"74",
          3681 => x"38",
          3682 => x"7b",
          3683 => x"ec",
          3684 => x"08",
          3685 => x"06",
          3686 => x"81",
          3687 => x"8a",
          3688 => x"05",
          3689 => x"06",
          3690 => x"bf",
          3691 => x"38",
          3692 => x"55",
          3693 => x"7a",
          3694 => x"98",
          3695 => x"77",
          3696 => x"3f",
          3697 => x"08",
          3698 => x"c0",
          3699 => x"82",
          3700 => x"81",
          3701 => x"38",
          3702 => x"ff",
          3703 => x"98",
          3704 => x"18",
          3705 => x"74",
          3706 => x"7e",
          3707 => x"08",
          3708 => x"2e",
          3709 => x"8d",
          3710 => x"ce",
          3711 => x"de",
          3712 => x"ee",
          3713 => x"08",
          3714 => x"d1",
          3715 => x"de",
          3716 => x"2e",
          3717 => x"81",
          3718 => x"1b",
          3719 => x"5a",
          3720 => x"2e",
          3721 => x"78",
          3722 => x"11",
          3723 => x"55",
          3724 => x"85",
          3725 => x"31",
          3726 => x"76",
          3727 => x"81",
          3728 => x"c8",
          3729 => x"de",
          3730 => x"a6",
          3731 => x"11",
          3732 => x"56",
          3733 => x"27",
          3734 => x"80",
          3735 => x"08",
          3736 => x"2b",
          3737 => x"b4",
          3738 => x"b5",
          3739 => x"80",
          3740 => x"34",
          3741 => x"56",
          3742 => x"8c",
          3743 => x"19",
          3744 => x"38",
          3745 => x"b6",
          3746 => x"c0",
          3747 => x"38",
          3748 => x"12",
          3749 => x"9c",
          3750 => x"18",
          3751 => x"06",
          3752 => x"31",
          3753 => x"76",
          3754 => x"7b",
          3755 => x"08",
          3756 => x"cd",
          3757 => x"de",
          3758 => x"b6",
          3759 => x"7c",
          3760 => x"08",
          3761 => x"1f",
          3762 => x"cb",
          3763 => x"55",
          3764 => x"16",
          3765 => x"31",
          3766 => x"7f",
          3767 => x"94",
          3768 => x"70",
          3769 => x"8c",
          3770 => x"58",
          3771 => x"76",
          3772 => x"75",
          3773 => x"19",
          3774 => x"39",
          3775 => x"80",
          3776 => x"74",
          3777 => x"80",
          3778 => x"de",
          3779 => x"3d",
          3780 => x"3d",
          3781 => x"3d",
          3782 => x"70",
          3783 => x"ea",
          3784 => x"c0",
          3785 => x"de",
          3786 => x"fb",
          3787 => x"33",
          3788 => x"70",
          3789 => x"55",
          3790 => x"2e",
          3791 => x"a0",
          3792 => x"78",
          3793 => x"3f",
          3794 => x"08",
          3795 => x"c0",
          3796 => x"38",
          3797 => x"8b",
          3798 => x"07",
          3799 => x"8b",
          3800 => x"16",
          3801 => x"52",
          3802 => x"dd",
          3803 => x"16",
          3804 => x"15",
          3805 => x"3f",
          3806 => x"0a",
          3807 => x"51",
          3808 => x"76",
          3809 => x"51",
          3810 => x"78",
          3811 => x"83",
          3812 => x"51",
          3813 => x"81",
          3814 => x"90",
          3815 => x"bf",
          3816 => x"73",
          3817 => x"76",
          3818 => x"0c",
          3819 => x"04",
          3820 => x"76",
          3821 => x"fe",
          3822 => x"de",
          3823 => x"81",
          3824 => x"9c",
          3825 => x"fc",
          3826 => x"51",
          3827 => x"81",
          3828 => x"53",
          3829 => x"08",
          3830 => x"de",
          3831 => x"0c",
          3832 => x"c0",
          3833 => x"0d",
          3834 => x"0d",
          3835 => x"e6",
          3836 => x"52",
          3837 => x"de",
          3838 => x"8b",
          3839 => x"c0",
          3840 => x"f0",
          3841 => x"71",
          3842 => x"0c",
          3843 => x"04",
          3844 => x"80",
          3845 => x"d0",
          3846 => x"3d",
          3847 => x"3f",
          3848 => x"08",
          3849 => x"c0",
          3850 => x"38",
          3851 => x"52",
          3852 => x"05",
          3853 => x"3f",
          3854 => x"08",
          3855 => x"c0",
          3856 => x"02",
          3857 => x"33",
          3858 => x"55",
          3859 => x"25",
          3860 => x"7a",
          3861 => x"54",
          3862 => x"a2",
          3863 => x"84",
          3864 => x"06",
          3865 => x"73",
          3866 => x"38",
          3867 => x"70",
          3868 => x"a8",
          3869 => x"c0",
          3870 => x"0c",
          3871 => x"de",
          3872 => x"2e",
          3873 => x"83",
          3874 => x"74",
          3875 => x"0c",
          3876 => x"04",
          3877 => x"6f",
          3878 => x"80",
          3879 => x"53",
          3880 => x"b8",
          3881 => x"3d",
          3882 => x"3f",
          3883 => x"08",
          3884 => x"c0",
          3885 => x"38",
          3886 => x"7c",
          3887 => x"47",
          3888 => x"54",
          3889 => x"81",
          3890 => x"52",
          3891 => x"52",
          3892 => x"3f",
          3893 => x"08",
          3894 => x"c0",
          3895 => x"38",
          3896 => x"51",
          3897 => x"81",
          3898 => x"57",
          3899 => x"08",
          3900 => x"69",
          3901 => x"da",
          3902 => x"de",
          3903 => x"76",
          3904 => x"d5",
          3905 => x"de",
          3906 => x"81",
          3907 => x"82",
          3908 => x"52",
          3909 => x"eb",
          3910 => x"c0",
          3911 => x"de",
          3912 => x"38",
          3913 => x"51",
          3914 => x"73",
          3915 => x"08",
          3916 => x"76",
          3917 => x"d6",
          3918 => x"de",
          3919 => x"81",
          3920 => x"80",
          3921 => x"76",
          3922 => x"81",
          3923 => x"82",
          3924 => x"39",
          3925 => x"38",
          3926 => x"bc",
          3927 => x"51",
          3928 => x"76",
          3929 => x"11",
          3930 => x"51",
          3931 => x"73",
          3932 => x"38",
          3933 => x"55",
          3934 => x"16",
          3935 => x"56",
          3936 => x"38",
          3937 => x"73",
          3938 => x"90",
          3939 => x"2e",
          3940 => x"16",
          3941 => x"ff",
          3942 => x"ff",
          3943 => x"58",
          3944 => x"74",
          3945 => x"75",
          3946 => x"18",
          3947 => x"58",
          3948 => x"fe",
          3949 => x"7b",
          3950 => x"06",
          3951 => x"18",
          3952 => x"58",
          3953 => x"80",
          3954 => x"f0",
          3955 => x"29",
          3956 => x"05",
          3957 => x"33",
          3958 => x"56",
          3959 => x"2e",
          3960 => x"16",
          3961 => x"33",
          3962 => x"73",
          3963 => x"16",
          3964 => x"26",
          3965 => x"55",
          3966 => x"91",
          3967 => x"54",
          3968 => x"70",
          3969 => x"34",
          3970 => x"ec",
          3971 => x"70",
          3972 => x"34",
          3973 => x"09",
          3974 => x"38",
          3975 => x"39",
          3976 => x"19",
          3977 => x"33",
          3978 => x"05",
          3979 => x"78",
          3980 => x"80",
          3981 => x"81",
          3982 => x"9e",
          3983 => x"f7",
          3984 => x"7d",
          3985 => x"05",
          3986 => x"57",
          3987 => x"3f",
          3988 => x"08",
          3989 => x"c0",
          3990 => x"38",
          3991 => x"53",
          3992 => x"38",
          3993 => x"54",
          3994 => x"92",
          3995 => x"33",
          3996 => x"70",
          3997 => x"54",
          3998 => x"38",
          3999 => x"15",
          4000 => x"70",
          4001 => x"58",
          4002 => x"82",
          4003 => x"8a",
          4004 => x"89",
          4005 => x"53",
          4006 => x"b7",
          4007 => x"ff",
          4008 => x"95",
          4009 => x"de",
          4010 => x"15",
          4011 => x"53",
          4012 => x"95",
          4013 => x"de",
          4014 => x"26",
          4015 => x"30",
          4016 => x"70",
          4017 => x"77",
          4018 => x"18",
          4019 => x"51",
          4020 => x"88",
          4021 => x"73",
          4022 => x"52",
          4023 => x"ca",
          4024 => x"c0",
          4025 => x"de",
          4026 => x"2e",
          4027 => x"81",
          4028 => x"ff",
          4029 => x"38",
          4030 => x"08",
          4031 => x"73",
          4032 => x"73",
          4033 => x"9c",
          4034 => x"27",
          4035 => x"75",
          4036 => x"16",
          4037 => x"17",
          4038 => x"33",
          4039 => x"70",
          4040 => x"55",
          4041 => x"80",
          4042 => x"73",
          4043 => x"cc",
          4044 => x"de",
          4045 => x"81",
          4046 => x"94",
          4047 => x"c0",
          4048 => x"39",
          4049 => x"51",
          4050 => x"81",
          4051 => x"54",
          4052 => x"be",
          4053 => x"27",
          4054 => x"53",
          4055 => x"08",
          4056 => x"73",
          4057 => x"ff",
          4058 => x"15",
          4059 => x"16",
          4060 => x"ff",
          4061 => x"80",
          4062 => x"73",
          4063 => x"c6",
          4064 => x"de",
          4065 => x"38",
          4066 => x"16",
          4067 => x"80",
          4068 => x"0b",
          4069 => x"81",
          4070 => x"75",
          4071 => x"de",
          4072 => x"58",
          4073 => x"54",
          4074 => x"74",
          4075 => x"73",
          4076 => x"90",
          4077 => x"c0",
          4078 => x"90",
          4079 => x"83",
          4080 => x"72",
          4081 => x"38",
          4082 => x"08",
          4083 => x"77",
          4084 => x"80",
          4085 => x"de",
          4086 => x"3d",
          4087 => x"3d",
          4088 => x"89",
          4089 => x"2e",
          4090 => x"80",
          4091 => x"fc",
          4092 => x"3d",
          4093 => x"e1",
          4094 => x"de",
          4095 => x"81",
          4096 => x"80",
          4097 => x"76",
          4098 => x"75",
          4099 => x"3f",
          4100 => x"08",
          4101 => x"c0",
          4102 => x"38",
          4103 => x"70",
          4104 => x"57",
          4105 => x"a2",
          4106 => x"33",
          4107 => x"70",
          4108 => x"55",
          4109 => x"2e",
          4110 => x"16",
          4111 => x"51",
          4112 => x"81",
          4113 => x"88",
          4114 => x"54",
          4115 => x"84",
          4116 => x"52",
          4117 => x"e5",
          4118 => x"c0",
          4119 => x"84",
          4120 => x"06",
          4121 => x"55",
          4122 => x"80",
          4123 => x"80",
          4124 => x"54",
          4125 => x"c0",
          4126 => x"0d",
          4127 => x"0d",
          4128 => x"fc",
          4129 => x"52",
          4130 => x"3f",
          4131 => x"08",
          4132 => x"de",
          4133 => x"0c",
          4134 => x"04",
          4135 => x"77",
          4136 => x"fc",
          4137 => x"53",
          4138 => x"de",
          4139 => x"c0",
          4140 => x"de",
          4141 => x"df",
          4142 => x"38",
          4143 => x"08",
          4144 => x"cd",
          4145 => x"de",
          4146 => x"80",
          4147 => x"de",
          4148 => x"73",
          4149 => x"3f",
          4150 => x"08",
          4151 => x"c0",
          4152 => x"09",
          4153 => x"38",
          4154 => x"39",
          4155 => x"08",
          4156 => x"52",
          4157 => x"b3",
          4158 => x"73",
          4159 => x"3f",
          4160 => x"08",
          4161 => x"30",
          4162 => x"9f",
          4163 => x"de",
          4164 => x"51",
          4165 => x"72",
          4166 => x"0c",
          4167 => x"04",
          4168 => x"65",
          4169 => x"89",
          4170 => x"96",
          4171 => x"df",
          4172 => x"de",
          4173 => x"81",
          4174 => x"b2",
          4175 => x"75",
          4176 => x"3f",
          4177 => x"08",
          4178 => x"c0",
          4179 => x"02",
          4180 => x"33",
          4181 => x"55",
          4182 => x"25",
          4183 => x"55",
          4184 => x"80",
          4185 => x"76",
          4186 => x"d4",
          4187 => x"81",
          4188 => x"94",
          4189 => x"f0",
          4190 => x"65",
          4191 => x"53",
          4192 => x"05",
          4193 => x"51",
          4194 => x"81",
          4195 => x"5b",
          4196 => x"08",
          4197 => x"7c",
          4198 => x"08",
          4199 => x"fe",
          4200 => x"08",
          4201 => x"55",
          4202 => x"91",
          4203 => x"0c",
          4204 => x"81",
          4205 => x"39",
          4206 => x"c7",
          4207 => x"c0",
          4208 => x"55",
          4209 => x"2e",
          4210 => x"bf",
          4211 => x"5f",
          4212 => x"92",
          4213 => x"51",
          4214 => x"81",
          4215 => x"ff",
          4216 => x"81",
          4217 => x"81",
          4218 => x"81",
          4219 => x"30",
          4220 => x"c0",
          4221 => x"25",
          4222 => x"19",
          4223 => x"5a",
          4224 => x"08",
          4225 => x"38",
          4226 => x"a4",
          4227 => x"de",
          4228 => x"58",
          4229 => x"77",
          4230 => x"7d",
          4231 => x"bf",
          4232 => x"de",
          4233 => x"81",
          4234 => x"80",
          4235 => x"70",
          4236 => x"ff",
          4237 => x"56",
          4238 => x"2e",
          4239 => x"9e",
          4240 => x"51",
          4241 => x"3f",
          4242 => x"08",
          4243 => x"06",
          4244 => x"80",
          4245 => x"19",
          4246 => x"54",
          4247 => x"14",
          4248 => x"c5",
          4249 => x"c0",
          4250 => x"06",
          4251 => x"80",
          4252 => x"19",
          4253 => x"54",
          4254 => x"06",
          4255 => x"79",
          4256 => x"78",
          4257 => x"79",
          4258 => x"84",
          4259 => x"07",
          4260 => x"84",
          4261 => x"81",
          4262 => x"92",
          4263 => x"f9",
          4264 => x"8a",
          4265 => x"53",
          4266 => x"e3",
          4267 => x"de",
          4268 => x"81",
          4269 => x"81",
          4270 => x"17",
          4271 => x"81",
          4272 => x"17",
          4273 => x"2a",
          4274 => x"51",
          4275 => x"55",
          4276 => x"81",
          4277 => x"17",
          4278 => x"8c",
          4279 => x"81",
          4280 => x"9b",
          4281 => x"c0",
          4282 => x"17",
          4283 => x"51",
          4284 => x"81",
          4285 => x"74",
          4286 => x"56",
          4287 => x"98",
          4288 => x"76",
          4289 => x"c6",
          4290 => x"c0",
          4291 => x"09",
          4292 => x"38",
          4293 => x"de",
          4294 => x"2e",
          4295 => x"85",
          4296 => x"a3",
          4297 => x"38",
          4298 => x"de",
          4299 => x"15",
          4300 => x"38",
          4301 => x"53",
          4302 => x"08",
          4303 => x"c3",
          4304 => x"de",
          4305 => x"94",
          4306 => x"18",
          4307 => x"33",
          4308 => x"54",
          4309 => x"34",
          4310 => x"85",
          4311 => x"18",
          4312 => x"74",
          4313 => x"0c",
          4314 => x"04",
          4315 => x"82",
          4316 => x"ff",
          4317 => x"a1",
          4318 => x"e4",
          4319 => x"c0",
          4320 => x"de",
          4321 => x"f5",
          4322 => x"a1",
          4323 => x"95",
          4324 => x"58",
          4325 => x"81",
          4326 => x"55",
          4327 => x"08",
          4328 => x"02",
          4329 => x"33",
          4330 => x"70",
          4331 => x"55",
          4332 => x"73",
          4333 => x"75",
          4334 => x"80",
          4335 => x"bd",
          4336 => x"d6",
          4337 => x"81",
          4338 => x"87",
          4339 => x"ad",
          4340 => x"78",
          4341 => x"3f",
          4342 => x"08",
          4343 => x"70",
          4344 => x"55",
          4345 => x"2e",
          4346 => x"78",
          4347 => x"c0",
          4348 => x"08",
          4349 => x"38",
          4350 => x"de",
          4351 => x"76",
          4352 => x"70",
          4353 => x"b5",
          4354 => x"c0",
          4355 => x"de",
          4356 => x"e9",
          4357 => x"c0",
          4358 => x"51",
          4359 => x"81",
          4360 => x"55",
          4361 => x"08",
          4362 => x"55",
          4363 => x"81",
          4364 => x"84",
          4365 => x"81",
          4366 => x"80",
          4367 => x"51",
          4368 => x"81",
          4369 => x"81",
          4370 => x"30",
          4371 => x"c0",
          4372 => x"25",
          4373 => x"75",
          4374 => x"38",
          4375 => x"8f",
          4376 => x"75",
          4377 => x"c1",
          4378 => x"de",
          4379 => x"74",
          4380 => x"51",
          4381 => x"3f",
          4382 => x"08",
          4383 => x"de",
          4384 => x"3d",
          4385 => x"3d",
          4386 => x"99",
          4387 => x"52",
          4388 => x"d8",
          4389 => x"de",
          4390 => x"81",
          4391 => x"82",
          4392 => x"5e",
          4393 => x"3d",
          4394 => x"cf",
          4395 => x"de",
          4396 => x"81",
          4397 => x"86",
          4398 => x"82",
          4399 => x"de",
          4400 => x"2e",
          4401 => x"82",
          4402 => x"80",
          4403 => x"70",
          4404 => x"06",
          4405 => x"54",
          4406 => x"38",
          4407 => x"52",
          4408 => x"52",
          4409 => x"3f",
          4410 => x"08",
          4411 => x"81",
          4412 => x"83",
          4413 => x"81",
          4414 => x"81",
          4415 => x"06",
          4416 => x"54",
          4417 => x"08",
          4418 => x"81",
          4419 => x"81",
          4420 => x"39",
          4421 => x"38",
          4422 => x"08",
          4423 => x"c4",
          4424 => x"de",
          4425 => x"81",
          4426 => x"81",
          4427 => x"53",
          4428 => x"19",
          4429 => x"8c",
          4430 => x"ae",
          4431 => x"34",
          4432 => x"0b",
          4433 => x"82",
          4434 => x"52",
          4435 => x"51",
          4436 => x"3f",
          4437 => x"b4",
          4438 => x"c9",
          4439 => x"53",
          4440 => x"53",
          4441 => x"51",
          4442 => x"3f",
          4443 => x"0b",
          4444 => x"34",
          4445 => x"80",
          4446 => x"51",
          4447 => x"78",
          4448 => x"83",
          4449 => x"51",
          4450 => x"81",
          4451 => x"54",
          4452 => x"08",
          4453 => x"88",
          4454 => x"64",
          4455 => x"ff",
          4456 => x"75",
          4457 => x"78",
          4458 => x"3f",
          4459 => x"0b",
          4460 => x"78",
          4461 => x"83",
          4462 => x"51",
          4463 => x"3f",
          4464 => x"08",
          4465 => x"80",
          4466 => x"76",
          4467 => x"ae",
          4468 => x"de",
          4469 => x"3d",
          4470 => x"3d",
          4471 => x"84",
          4472 => x"f1",
          4473 => x"a8",
          4474 => x"05",
          4475 => x"51",
          4476 => x"81",
          4477 => x"55",
          4478 => x"08",
          4479 => x"78",
          4480 => x"08",
          4481 => x"70",
          4482 => x"b8",
          4483 => x"c0",
          4484 => x"de",
          4485 => x"b9",
          4486 => x"9b",
          4487 => x"a0",
          4488 => x"55",
          4489 => x"38",
          4490 => x"3d",
          4491 => x"3d",
          4492 => x"51",
          4493 => x"3f",
          4494 => x"52",
          4495 => x"52",
          4496 => x"dd",
          4497 => x"08",
          4498 => x"cb",
          4499 => x"de",
          4500 => x"81",
          4501 => x"95",
          4502 => x"2e",
          4503 => x"88",
          4504 => x"3d",
          4505 => x"38",
          4506 => x"e5",
          4507 => x"c0",
          4508 => x"09",
          4509 => x"b8",
          4510 => x"c9",
          4511 => x"de",
          4512 => x"81",
          4513 => x"81",
          4514 => x"56",
          4515 => x"3d",
          4516 => x"52",
          4517 => x"ff",
          4518 => x"02",
          4519 => x"8b",
          4520 => x"16",
          4521 => x"2a",
          4522 => x"51",
          4523 => x"89",
          4524 => x"07",
          4525 => x"17",
          4526 => x"81",
          4527 => x"34",
          4528 => x"70",
          4529 => x"81",
          4530 => x"55",
          4531 => x"80",
          4532 => x"64",
          4533 => x"38",
          4534 => x"51",
          4535 => x"81",
          4536 => x"52",
          4537 => x"b7",
          4538 => x"55",
          4539 => x"08",
          4540 => x"dd",
          4541 => x"c0",
          4542 => x"51",
          4543 => x"3f",
          4544 => x"08",
          4545 => x"11",
          4546 => x"81",
          4547 => x"80",
          4548 => x"16",
          4549 => x"ae",
          4550 => x"06",
          4551 => x"53",
          4552 => x"51",
          4553 => x"78",
          4554 => x"83",
          4555 => x"39",
          4556 => x"08",
          4557 => x"51",
          4558 => x"81",
          4559 => x"55",
          4560 => x"08",
          4561 => x"51",
          4562 => x"3f",
          4563 => x"08",
          4564 => x"de",
          4565 => x"3d",
          4566 => x"3d",
          4567 => x"db",
          4568 => x"84",
          4569 => x"05",
          4570 => x"82",
          4571 => x"d0",
          4572 => x"3d",
          4573 => x"3f",
          4574 => x"08",
          4575 => x"c0",
          4576 => x"38",
          4577 => x"52",
          4578 => x"05",
          4579 => x"3f",
          4580 => x"08",
          4581 => x"c0",
          4582 => x"02",
          4583 => x"33",
          4584 => x"54",
          4585 => x"aa",
          4586 => x"06",
          4587 => x"8b",
          4588 => x"06",
          4589 => x"07",
          4590 => x"56",
          4591 => x"34",
          4592 => x"0b",
          4593 => x"78",
          4594 => x"a9",
          4595 => x"c0",
          4596 => x"81",
          4597 => x"95",
          4598 => x"ef",
          4599 => x"56",
          4600 => x"3d",
          4601 => x"94",
          4602 => x"f4",
          4603 => x"c0",
          4604 => x"de",
          4605 => x"cb",
          4606 => x"63",
          4607 => x"d4",
          4608 => x"c0",
          4609 => x"c0",
          4610 => x"de",
          4611 => x"38",
          4612 => x"05",
          4613 => x"06",
          4614 => x"73",
          4615 => x"16",
          4616 => x"22",
          4617 => x"07",
          4618 => x"1f",
          4619 => x"c2",
          4620 => x"81",
          4621 => x"34",
          4622 => x"b3",
          4623 => x"de",
          4624 => x"74",
          4625 => x"0c",
          4626 => x"04",
          4627 => x"69",
          4628 => x"80",
          4629 => x"d0",
          4630 => x"3d",
          4631 => x"3f",
          4632 => x"08",
          4633 => x"08",
          4634 => x"de",
          4635 => x"80",
          4636 => x"57",
          4637 => x"81",
          4638 => x"70",
          4639 => x"55",
          4640 => x"80",
          4641 => x"5d",
          4642 => x"52",
          4643 => x"52",
          4644 => x"a9",
          4645 => x"c0",
          4646 => x"de",
          4647 => x"d1",
          4648 => x"73",
          4649 => x"3f",
          4650 => x"08",
          4651 => x"c0",
          4652 => x"81",
          4653 => x"81",
          4654 => x"65",
          4655 => x"78",
          4656 => x"7b",
          4657 => x"55",
          4658 => x"34",
          4659 => x"8a",
          4660 => x"38",
          4661 => x"1a",
          4662 => x"34",
          4663 => x"9e",
          4664 => x"70",
          4665 => x"51",
          4666 => x"a0",
          4667 => x"8e",
          4668 => x"2e",
          4669 => x"86",
          4670 => x"34",
          4671 => x"30",
          4672 => x"80",
          4673 => x"7a",
          4674 => x"c1",
          4675 => x"2e",
          4676 => x"a0",
          4677 => x"51",
          4678 => x"3f",
          4679 => x"08",
          4680 => x"c0",
          4681 => x"7b",
          4682 => x"55",
          4683 => x"73",
          4684 => x"38",
          4685 => x"73",
          4686 => x"38",
          4687 => x"15",
          4688 => x"ff",
          4689 => x"81",
          4690 => x"7b",
          4691 => x"de",
          4692 => x"3d",
          4693 => x"3d",
          4694 => x"9c",
          4695 => x"05",
          4696 => x"51",
          4697 => x"81",
          4698 => x"81",
          4699 => x"56",
          4700 => x"c0",
          4701 => x"38",
          4702 => x"52",
          4703 => x"52",
          4704 => x"c0",
          4705 => x"70",
          4706 => x"ff",
          4707 => x"55",
          4708 => x"27",
          4709 => x"78",
          4710 => x"ff",
          4711 => x"05",
          4712 => x"55",
          4713 => x"3f",
          4714 => x"08",
          4715 => x"38",
          4716 => x"70",
          4717 => x"ff",
          4718 => x"81",
          4719 => x"80",
          4720 => x"74",
          4721 => x"07",
          4722 => x"4e",
          4723 => x"81",
          4724 => x"55",
          4725 => x"70",
          4726 => x"06",
          4727 => x"99",
          4728 => x"e0",
          4729 => x"ff",
          4730 => x"54",
          4731 => x"27",
          4732 => x"cc",
          4733 => x"55",
          4734 => x"a3",
          4735 => x"81",
          4736 => x"ff",
          4737 => x"81",
          4738 => x"93",
          4739 => x"75",
          4740 => x"76",
          4741 => x"38",
          4742 => x"77",
          4743 => x"86",
          4744 => x"39",
          4745 => x"27",
          4746 => x"88",
          4747 => x"78",
          4748 => x"5a",
          4749 => x"57",
          4750 => x"81",
          4751 => x"81",
          4752 => x"33",
          4753 => x"06",
          4754 => x"57",
          4755 => x"fe",
          4756 => x"3d",
          4757 => x"55",
          4758 => x"2e",
          4759 => x"76",
          4760 => x"38",
          4761 => x"55",
          4762 => x"33",
          4763 => x"a0",
          4764 => x"06",
          4765 => x"17",
          4766 => x"38",
          4767 => x"43",
          4768 => x"3d",
          4769 => x"ff",
          4770 => x"81",
          4771 => x"54",
          4772 => x"08",
          4773 => x"81",
          4774 => x"ff",
          4775 => x"81",
          4776 => x"54",
          4777 => x"08",
          4778 => x"80",
          4779 => x"54",
          4780 => x"80",
          4781 => x"de",
          4782 => x"2e",
          4783 => x"80",
          4784 => x"54",
          4785 => x"80",
          4786 => x"52",
          4787 => x"bd",
          4788 => x"de",
          4789 => x"81",
          4790 => x"b1",
          4791 => x"81",
          4792 => x"52",
          4793 => x"ab",
          4794 => x"54",
          4795 => x"15",
          4796 => x"78",
          4797 => x"ff",
          4798 => x"79",
          4799 => x"83",
          4800 => x"51",
          4801 => x"3f",
          4802 => x"08",
          4803 => x"74",
          4804 => x"0c",
          4805 => x"04",
          4806 => x"60",
          4807 => x"05",
          4808 => x"33",
          4809 => x"05",
          4810 => x"40",
          4811 => x"da",
          4812 => x"c0",
          4813 => x"de",
          4814 => x"bd",
          4815 => x"33",
          4816 => x"b5",
          4817 => x"2e",
          4818 => x"1a",
          4819 => x"90",
          4820 => x"33",
          4821 => x"70",
          4822 => x"55",
          4823 => x"38",
          4824 => x"97",
          4825 => x"82",
          4826 => x"58",
          4827 => x"7e",
          4828 => x"70",
          4829 => x"55",
          4830 => x"56",
          4831 => x"f7",
          4832 => x"7d",
          4833 => x"70",
          4834 => x"2a",
          4835 => x"08",
          4836 => x"08",
          4837 => x"5d",
          4838 => x"77",
          4839 => x"98",
          4840 => x"26",
          4841 => x"57",
          4842 => x"59",
          4843 => x"52",
          4844 => x"ae",
          4845 => x"15",
          4846 => x"98",
          4847 => x"26",
          4848 => x"55",
          4849 => x"08",
          4850 => x"99",
          4851 => x"c0",
          4852 => x"ff",
          4853 => x"de",
          4854 => x"38",
          4855 => x"75",
          4856 => x"81",
          4857 => x"93",
          4858 => x"80",
          4859 => x"2e",
          4860 => x"ff",
          4861 => x"58",
          4862 => x"7d",
          4863 => x"38",
          4864 => x"55",
          4865 => x"b4",
          4866 => x"56",
          4867 => x"09",
          4868 => x"38",
          4869 => x"53",
          4870 => x"51",
          4871 => x"3f",
          4872 => x"08",
          4873 => x"c0",
          4874 => x"38",
          4875 => x"ff",
          4876 => x"5c",
          4877 => x"84",
          4878 => x"5c",
          4879 => x"12",
          4880 => x"80",
          4881 => x"78",
          4882 => x"7c",
          4883 => x"90",
          4884 => x"c0",
          4885 => x"90",
          4886 => x"15",
          4887 => x"90",
          4888 => x"54",
          4889 => x"91",
          4890 => x"31",
          4891 => x"84",
          4892 => x"07",
          4893 => x"16",
          4894 => x"73",
          4895 => x"0c",
          4896 => x"04",
          4897 => x"6b",
          4898 => x"05",
          4899 => x"33",
          4900 => x"5a",
          4901 => x"bd",
          4902 => x"80",
          4903 => x"c0",
          4904 => x"f8",
          4905 => x"c0",
          4906 => x"81",
          4907 => x"70",
          4908 => x"74",
          4909 => x"38",
          4910 => x"81",
          4911 => x"81",
          4912 => x"81",
          4913 => x"ff",
          4914 => x"81",
          4915 => x"81",
          4916 => x"81",
          4917 => x"83",
          4918 => x"c0",
          4919 => x"2a",
          4920 => x"51",
          4921 => x"74",
          4922 => x"99",
          4923 => x"53",
          4924 => x"51",
          4925 => x"3f",
          4926 => x"08",
          4927 => x"55",
          4928 => x"92",
          4929 => x"80",
          4930 => x"38",
          4931 => x"06",
          4932 => x"2e",
          4933 => x"48",
          4934 => x"87",
          4935 => x"79",
          4936 => x"78",
          4937 => x"26",
          4938 => x"19",
          4939 => x"74",
          4940 => x"38",
          4941 => x"e4",
          4942 => x"2a",
          4943 => x"70",
          4944 => x"59",
          4945 => x"7a",
          4946 => x"56",
          4947 => x"80",
          4948 => x"51",
          4949 => x"74",
          4950 => x"99",
          4951 => x"53",
          4952 => x"51",
          4953 => x"3f",
          4954 => x"de",
          4955 => x"ac",
          4956 => x"2a",
          4957 => x"81",
          4958 => x"43",
          4959 => x"83",
          4960 => x"66",
          4961 => x"60",
          4962 => x"90",
          4963 => x"31",
          4964 => x"80",
          4965 => x"8a",
          4966 => x"56",
          4967 => x"26",
          4968 => x"77",
          4969 => x"81",
          4970 => x"74",
          4971 => x"38",
          4972 => x"55",
          4973 => x"83",
          4974 => x"81",
          4975 => x"80",
          4976 => x"38",
          4977 => x"55",
          4978 => x"5e",
          4979 => x"89",
          4980 => x"5a",
          4981 => x"09",
          4982 => x"e1",
          4983 => x"38",
          4984 => x"57",
          4985 => x"ce",
          4986 => x"5a",
          4987 => x"9d",
          4988 => x"26",
          4989 => x"ce",
          4990 => x"10",
          4991 => x"22",
          4992 => x"74",
          4993 => x"38",
          4994 => x"ee",
          4995 => x"66",
          4996 => x"e3",
          4997 => x"c0",
          4998 => x"84",
          4999 => x"89",
          5000 => x"a0",
          5001 => x"81",
          5002 => x"fc",
          5003 => x"56",
          5004 => x"f0",
          5005 => x"80",
          5006 => x"d3",
          5007 => x"38",
          5008 => x"57",
          5009 => x"ce",
          5010 => x"5a",
          5011 => x"9d",
          5012 => x"26",
          5013 => x"ce",
          5014 => x"10",
          5015 => x"22",
          5016 => x"74",
          5017 => x"38",
          5018 => x"ee",
          5019 => x"66",
          5020 => x"83",
          5021 => x"c0",
          5022 => x"05",
          5023 => x"c0",
          5024 => x"26",
          5025 => x"0b",
          5026 => x"08",
          5027 => x"c0",
          5028 => x"11",
          5029 => x"05",
          5030 => x"83",
          5031 => x"2a",
          5032 => x"a0",
          5033 => x"7d",
          5034 => x"69",
          5035 => x"05",
          5036 => x"72",
          5037 => x"5c",
          5038 => x"59",
          5039 => x"2e",
          5040 => x"89",
          5041 => x"60",
          5042 => x"84",
          5043 => x"5d",
          5044 => x"18",
          5045 => x"68",
          5046 => x"74",
          5047 => x"af",
          5048 => x"31",
          5049 => x"53",
          5050 => x"52",
          5051 => x"87",
          5052 => x"c0",
          5053 => x"83",
          5054 => x"06",
          5055 => x"de",
          5056 => x"ff",
          5057 => x"dd",
          5058 => x"83",
          5059 => x"2a",
          5060 => x"be",
          5061 => x"39",
          5062 => x"09",
          5063 => x"c5",
          5064 => x"f5",
          5065 => x"c0",
          5066 => x"38",
          5067 => x"79",
          5068 => x"80",
          5069 => x"38",
          5070 => x"96",
          5071 => x"06",
          5072 => x"2e",
          5073 => x"5e",
          5074 => x"81",
          5075 => x"9f",
          5076 => x"38",
          5077 => x"38",
          5078 => x"81",
          5079 => x"fc",
          5080 => x"ab",
          5081 => x"7d",
          5082 => x"81",
          5083 => x"7d",
          5084 => x"78",
          5085 => x"74",
          5086 => x"8e",
          5087 => x"9c",
          5088 => x"53",
          5089 => x"51",
          5090 => x"3f",
          5091 => x"cc",
          5092 => x"51",
          5093 => x"3f",
          5094 => x"8b",
          5095 => x"a1",
          5096 => x"8d",
          5097 => x"83",
          5098 => x"52",
          5099 => x"ff",
          5100 => x"81",
          5101 => x"34",
          5102 => x"70",
          5103 => x"2a",
          5104 => x"54",
          5105 => x"1b",
          5106 => x"88",
          5107 => x"74",
          5108 => x"26",
          5109 => x"83",
          5110 => x"52",
          5111 => x"ff",
          5112 => x"8a",
          5113 => x"a0",
          5114 => x"a1",
          5115 => x"0b",
          5116 => x"bf",
          5117 => x"51",
          5118 => x"3f",
          5119 => x"9a",
          5120 => x"a0",
          5121 => x"52",
          5122 => x"ff",
          5123 => x"7d",
          5124 => x"81",
          5125 => x"38",
          5126 => x"0a",
          5127 => x"1b",
          5128 => x"ce",
          5129 => x"a4",
          5130 => x"a0",
          5131 => x"52",
          5132 => x"ff",
          5133 => x"81",
          5134 => x"51",
          5135 => x"3f",
          5136 => x"1b",
          5137 => x"8c",
          5138 => x"0b",
          5139 => x"34",
          5140 => x"c2",
          5141 => x"53",
          5142 => x"52",
          5143 => x"51",
          5144 => x"88",
          5145 => x"a7",
          5146 => x"a0",
          5147 => x"83",
          5148 => x"52",
          5149 => x"ff",
          5150 => x"ff",
          5151 => x"1c",
          5152 => x"a6",
          5153 => x"53",
          5154 => x"52",
          5155 => x"ff",
          5156 => x"82",
          5157 => x"83",
          5158 => x"52",
          5159 => x"b4",
          5160 => x"60",
          5161 => x"7e",
          5162 => x"d7",
          5163 => x"81",
          5164 => x"83",
          5165 => x"83",
          5166 => x"06",
          5167 => x"75",
          5168 => x"05",
          5169 => x"7e",
          5170 => x"b7",
          5171 => x"53",
          5172 => x"51",
          5173 => x"3f",
          5174 => x"a4",
          5175 => x"51",
          5176 => x"3f",
          5177 => x"e4",
          5178 => x"e4",
          5179 => x"9f",
          5180 => x"18",
          5181 => x"1b",
          5182 => x"f6",
          5183 => x"83",
          5184 => x"ff",
          5185 => x"82",
          5186 => x"78",
          5187 => x"c4",
          5188 => x"60",
          5189 => x"7a",
          5190 => x"ff",
          5191 => x"75",
          5192 => x"53",
          5193 => x"51",
          5194 => x"3f",
          5195 => x"52",
          5196 => x"9f",
          5197 => x"56",
          5198 => x"83",
          5199 => x"06",
          5200 => x"52",
          5201 => x"9e",
          5202 => x"52",
          5203 => x"ff",
          5204 => x"f0",
          5205 => x"1b",
          5206 => x"87",
          5207 => x"55",
          5208 => x"83",
          5209 => x"74",
          5210 => x"ff",
          5211 => x"7c",
          5212 => x"74",
          5213 => x"38",
          5214 => x"54",
          5215 => x"52",
          5216 => x"99",
          5217 => x"de",
          5218 => x"87",
          5219 => x"53",
          5220 => x"08",
          5221 => x"ff",
          5222 => x"76",
          5223 => x"31",
          5224 => x"cd",
          5225 => x"58",
          5226 => x"ff",
          5227 => x"55",
          5228 => x"83",
          5229 => x"61",
          5230 => x"26",
          5231 => x"57",
          5232 => x"53",
          5233 => x"51",
          5234 => x"3f",
          5235 => x"08",
          5236 => x"76",
          5237 => x"31",
          5238 => x"db",
          5239 => x"7d",
          5240 => x"38",
          5241 => x"83",
          5242 => x"8a",
          5243 => x"7d",
          5244 => x"38",
          5245 => x"81",
          5246 => x"80",
          5247 => x"80",
          5248 => x"7a",
          5249 => x"bc",
          5250 => x"d5",
          5251 => x"ff",
          5252 => x"83",
          5253 => x"77",
          5254 => x"0b",
          5255 => x"81",
          5256 => x"34",
          5257 => x"34",
          5258 => x"34",
          5259 => x"56",
          5260 => x"52",
          5261 => x"ee",
          5262 => x"0b",
          5263 => x"81",
          5264 => x"82",
          5265 => x"56",
          5266 => x"34",
          5267 => x"08",
          5268 => x"60",
          5269 => x"1b",
          5270 => x"96",
          5271 => x"83",
          5272 => x"ff",
          5273 => x"81",
          5274 => x"7a",
          5275 => x"ff",
          5276 => x"81",
          5277 => x"c0",
          5278 => x"80",
          5279 => x"7e",
          5280 => x"e3",
          5281 => x"81",
          5282 => x"90",
          5283 => x"8e",
          5284 => x"81",
          5285 => x"81",
          5286 => x"56",
          5287 => x"c0",
          5288 => x"0d",
          5289 => x"0d",
          5290 => x"59",
          5291 => x"ff",
          5292 => x"57",
          5293 => x"b4",
          5294 => x"f8",
          5295 => x"81",
          5296 => x"52",
          5297 => x"dc",
          5298 => x"2e",
          5299 => x"9c",
          5300 => x"33",
          5301 => x"2e",
          5302 => x"76",
          5303 => x"58",
          5304 => x"57",
          5305 => x"09",
          5306 => x"38",
          5307 => x"78",
          5308 => x"38",
          5309 => x"81",
          5310 => x"8d",
          5311 => x"ff",
          5312 => x"52",
          5313 => x"81",
          5314 => x"84",
          5315 => x"94",
          5316 => x"08",
          5317 => x"f0",
          5318 => x"39",
          5319 => x"51",
          5320 => x"81",
          5321 => x"80",
          5322 => x"d0",
          5323 => x"eb",
          5324 => x"b4",
          5325 => x"39",
          5326 => x"51",
          5327 => x"81",
          5328 => x"80",
          5329 => x"d0",
          5330 => x"cf",
          5331 => x"80",
          5332 => x"39",
          5333 => x"51",
          5334 => x"81",
          5335 => x"bb",
          5336 => x"cc",
          5337 => x"81",
          5338 => x"af",
          5339 => x"8c",
          5340 => x"81",
          5341 => x"a3",
          5342 => x"c0",
          5343 => x"81",
          5344 => x"97",
          5345 => x"ec",
          5346 => x"81",
          5347 => x"8b",
          5348 => x"9c",
          5349 => x"81",
          5350 => x"ff",
          5351 => x"83",
          5352 => x"fb",
          5353 => x"79",
          5354 => x"87",
          5355 => x"38",
          5356 => x"87",
          5357 => x"91",
          5358 => x"52",
          5359 => x"eb",
          5360 => x"de",
          5361 => x"75",
          5362 => x"ab",
          5363 => x"c0",
          5364 => x"53",
          5365 => x"d3",
          5366 => x"8c",
          5367 => x"3d",
          5368 => x"3d",
          5369 => x"61",
          5370 => x"80",
          5371 => x"73",
          5372 => x"5f",
          5373 => x"5c",
          5374 => x"52",
          5375 => x"51",
          5376 => x"3f",
          5377 => x"51",
          5378 => x"3f",
          5379 => x"77",
          5380 => x"38",
          5381 => x"89",
          5382 => x"2e",
          5383 => x"c6",
          5384 => x"53",
          5385 => x"8e",
          5386 => x"52",
          5387 => x"51",
          5388 => x"3f",
          5389 => x"d3",
          5390 => x"86",
          5391 => x"15",
          5392 => x"39",
          5393 => x"72",
          5394 => x"38",
          5395 => x"81",
          5396 => x"ff",
          5397 => x"89",
          5398 => x"f0",
          5399 => x"df",
          5400 => x"55",
          5401 => x"16",
          5402 => x"27",
          5403 => x"33",
          5404 => x"fc",
          5405 => x"ab",
          5406 => x"81",
          5407 => x"ff",
          5408 => x"81",
          5409 => x"51",
          5410 => x"3f",
          5411 => x"81",
          5412 => x"ff",
          5413 => x"80",
          5414 => x"27",
          5415 => x"16",
          5416 => x"72",
          5417 => x"53",
          5418 => x"90",
          5419 => x"2e",
          5420 => x"80",
          5421 => x"38",
          5422 => x"39",
          5423 => x"f5",
          5424 => x"15",
          5425 => x"81",
          5426 => x"ff",
          5427 => x"76",
          5428 => x"5a",
          5429 => x"b4",
          5430 => x"c0",
          5431 => x"70",
          5432 => x"55",
          5433 => x"09",
          5434 => x"38",
          5435 => x"3f",
          5436 => x"08",
          5437 => x"98",
          5438 => x"32",
          5439 => x"72",
          5440 => x"51",
          5441 => x"55",
          5442 => x"8c",
          5443 => x"38",
          5444 => x"09",
          5445 => x"38",
          5446 => x"39",
          5447 => x"72",
          5448 => x"d6",
          5449 => x"72",
          5450 => x"0c",
          5451 => x"04",
          5452 => x"66",
          5453 => x"80",
          5454 => x"69",
          5455 => x"74",
          5456 => x"70",
          5457 => x"27",
          5458 => x"58",
          5459 => x"93",
          5460 => x"fc",
          5461 => x"75",
          5462 => x"70",
          5463 => x"bf",
          5464 => x"de",
          5465 => x"81",
          5466 => x"b8",
          5467 => x"c0",
          5468 => x"98",
          5469 => x"de",
          5470 => x"96",
          5471 => x"54",
          5472 => x"77",
          5473 => x"c4",
          5474 => x"de",
          5475 => x"81",
          5476 => x"90",
          5477 => x"74",
          5478 => x"38",
          5479 => x"19",
          5480 => x"39",
          5481 => x"05",
          5482 => x"3f",
          5483 => x"77",
          5484 => x"51",
          5485 => x"2e",
          5486 => x"80",
          5487 => x"81",
          5488 => x"87",
          5489 => x"08",
          5490 => x"fb",
          5491 => x"57",
          5492 => x"c0",
          5493 => x"0d",
          5494 => x"0d",
          5495 => x"05",
          5496 => x"57",
          5497 => x"80",
          5498 => x"79",
          5499 => x"3f",
          5500 => x"08",
          5501 => x"80",
          5502 => x"75",
          5503 => x"38",
          5504 => x"55",
          5505 => x"de",
          5506 => x"52",
          5507 => x"2d",
          5508 => x"08",
          5509 => x"77",
          5510 => x"de",
          5511 => x"3d",
          5512 => x"3d",
          5513 => x"05",
          5514 => x"98",
          5515 => x"a0",
          5516 => x"87",
          5517 => x"db",
          5518 => x"ff",
          5519 => x"81",
          5520 => x"81",
          5521 => x"81",
          5522 => x"52",
          5523 => x"51",
          5524 => x"3f",
          5525 => x"85",
          5526 => x"d4",
          5527 => x"0d",
          5528 => x"0d",
          5529 => x"80",
          5530 => x"80",
          5531 => x"51",
          5532 => x"3f",
          5533 => x"51",
          5534 => x"3f",
          5535 => x"f2",
          5536 => x"81",
          5537 => x"06",
          5538 => x"80",
          5539 => x"81",
          5540 => x"8c",
          5541 => x"f8",
          5542 => x"84",
          5543 => x"fe",
          5544 => x"72",
          5545 => x"81",
          5546 => x"71",
          5547 => x"38",
          5548 => x"f1",
          5549 => x"d5",
          5550 => x"f3",
          5551 => x"51",
          5552 => x"3f",
          5553 => x"70",
          5554 => x"52",
          5555 => x"95",
          5556 => x"fe",
          5557 => x"81",
          5558 => x"fe",
          5559 => x"80",
          5560 => x"bc",
          5561 => x"2a",
          5562 => x"51",
          5563 => x"2e",
          5564 => x"51",
          5565 => x"3f",
          5566 => x"51",
          5567 => x"3f",
          5568 => x"f1",
          5569 => x"85",
          5570 => x"06",
          5571 => x"80",
          5572 => x"81",
          5573 => x"88",
          5574 => x"c4",
          5575 => x"80",
          5576 => x"fe",
          5577 => x"72",
          5578 => x"81",
          5579 => x"71",
          5580 => x"38",
          5581 => x"f0",
          5582 => x"d5",
          5583 => x"f2",
          5584 => x"51",
          5585 => x"3f",
          5586 => x"70",
          5587 => x"52",
          5588 => x"95",
          5589 => x"fe",
          5590 => x"81",
          5591 => x"fe",
          5592 => x"80",
          5593 => x"b8",
          5594 => x"2a",
          5595 => x"51",
          5596 => x"2e",
          5597 => x"51",
          5598 => x"3f",
          5599 => x"51",
          5600 => x"3f",
          5601 => x"f0",
          5602 => x"fe",
          5603 => x"3d",
          5604 => x"3d",
          5605 => x"08",
          5606 => x"57",
          5607 => x"80",
          5608 => x"39",
          5609 => x"85",
          5610 => x"80",
          5611 => x"14",
          5612 => x"33",
          5613 => x"06",
          5614 => x"74",
          5615 => x"38",
          5616 => x"80",
          5617 => x"72",
          5618 => x"81",
          5619 => x"72",
          5620 => x"81",
          5621 => x"80",
          5622 => x"05",
          5623 => x"56",
          5624 => x"81",
          5625 => x"77",
          5626 => x"08",
          5627 => x"ea",
          5628 => x"de",
          5629 => x"38",
          5630 => x"53",
          5631 => x"ff",
          5632 => x"16",
          5633 => x"06",
          5634 => x"76",
          5635 => x"ff",
          5636 => x"de",
          5637 => x"3d",
          5638 => x"3d",
          5639 => x"70",
          5640 => x"80",
          5641 => x"fe",
          5642 => x"81",
          5643 => x"54",
          5644 => x"81",
          5645 => x"c0",
          5646 => x"c4",
          5647 => x"ff",
          5648 => x"c0",
          5649 => x"81",
          5650 => x"07",
          5651 => x"71",
          5652 => x"54",
          5653 => x"ec",
          5654 => x"ec",
          5655 => x"81",
          5656 => x"06",
          5657 => x"f5",
          5658 => x"52",
          5659 => x"b5",
          5660 => x"c0",
          5661 => x"8c",
          5662 => x"c0",
          5663 => x"fd",
          5664 => x"39",
          5665 => x"51",
          5666 => x"82",
          5667 => x"ec",
          5668 => x"ec",
          5669 => x"82",
          5670 => x"06",
          5671 => x"52",
          5672 => x"83",
          5673 => x"0b",
          5674 => x"0c",
          5675 => x"04",
          5676 => x"80",
          5677 => x"f5",
          5678 => x"5d",
          5679 => x"51",
          5680 => x"3f",
          5681 => x"08",
          5682 => x"59",
          5683 => x"09",
          5684 => x"38",
          5685 => x"52",
          5686 => x"52",
          5687 => x"d9",
          5688 => x"78",
          5689 => x"f0",
          5690 => x"f2",
          5691 => x"c0",
          5692 => x"88",
          5693 => x"d4",
          5694 => x"39",
          5695 => x"5d",
          5696 => x"51",
          5697 => x"3f",
          5698 => x"46",
          5699 => x"52",
          5700 => x"86",
          5701 => x"fe",
          5702 => x"fc",
          5703 => x"de",
          5704 => x"2b",
          5705 => x"51",
          5706 => x"c3",
          5707 => x"38",
          5708 => x"24",
          5709 => x"78",
          5710 => x"bc",
          5711 => x"24",
          5712 => x"82",
          5713 => x"38",
          5714 => x"8a",
          5715 => x"2e",
          5716 => x"8f",
          5717 => x"84",
          5718 => x"38",
          5719 => x"82",
          5720 => x"cf",
          5721 => x"c0",
          5722 => x"38",
          5723 => x"24",
          5724 => x"b0",
          5725 => x"38",
          5726 => x"84",
          5727 => x"b3",
          5728 => x"c1",
          5729 => x"38",
          5730 => x"2e",
          5731 => x"8f",
          5732 => x"80",
          5733 => x"f3",
          5734 => x"d5",
          5735 => x"78",
          5736 => x"8d",
          5737 => x"80",
          5738 => x"38",
          5739 => x"2e",
          5740 => x"8e",
          5741 => x"80",
          5742 => x"a1",
          5743 => x"d4",
          5744 => x"38",
          5745 => x"78",
          5746 => x"8e",
          5747 => x"81",
          5748 => x"38",
          5749 => x"2e",
          5750 => x"78",
          5751 => x"8d",
          5752 => x"cf",
          5753 => x"83",
          5754 => x"38",
          5755 => x"2e",
          5756 => x"8e",
          5757 => x"3d",
          5758 => x"53",
          5759 => x"51",
          5760 => x"3f",
          5761 => x"08",
          5762 => x"d7",
          5763 => x"a7",
          5764 => x"fe",
          5765 => x"fe",
          5766 => x"ff",
          5767 => x"81",
          5768 => x"80",
          5769 => x"81",
          5770 => x"38",
          5771 => x"80",
          5772 => x"52",
          5773 => x"05",
          5774 => x"85",
          5775 => x"de",
          5776 => x"ff",
          5777 => x"8e",
          5778 => x"a0",
          5779 => x"ef",
          5780 => x"fd",
          5781 => x"d7",
          5782 => x"a8",
          5783 => x"fe",
          5784 => x"fe",
          5785 => x"ff",
          5786 => x"81",
          5787 => x"80",
          5788 => x"38",
          5789 => x"52",
          5790 => x"05",
          5791 => x"89",
          5792 => x"de",
          5793 => x"81",
          5794 => x"8c",
          5795 => x"3d",
          5796 => x"53",
          5797 => x"51",
          5798 => x"3f",
          5799 => x"08",
          5800 => x"38",
          5801 => x"fc",
          5802 => x"3d",
          5803 => x"53",
          5804 => x"51",
          5805 => x"3f",
          5806 => x"08",
          5807 => x"de",
          5808 => x"63",
          5809 => x"d0",
          5810 => x"fe",
          5811 => x"02",
          5812 => x"33",
          5813 => x"63",
          5814 => x"81",
          5815 => x"51",
          5816 => x"3f",
          5817 => x"08",
          5818 => x"81",
          5819 => x"fe",
          5820 => x"81",
          5821 => x"39",
          5822 => x"f8",
          5823 => x"e5",
          5824 => x"de",
          5825 => x"3d",
          5826 => x"52",
          5827 => x"a3",
          5828 => x"81",
          5829 => x"52",
          5830 => x"94",
          5831 => x"39",
          5832 => x"f8",
          5833 => x"e5",
          5834 => x"de",
          5835 => x"3d",
          5836 => x"52",
          5837 => x"fb",
          5838 => x"c0",
          5839 => x"fe",
          5840 => x"5a",
          5841 => x"3f",
          5842 => x"08",
          5843 => x"f8",
          5844 => x"fe",
          5845 => x"81",
          5846 => x"81",
          5847 => x"80",
          5848 => x"81",
          5849 => x"81",
          5850 => x"78",
          5851 => x"7a",
          5852 => x"3f",
          5853 => x"08",
          5854 => x"84",
          5855 => x"c0",
          5856 => x"fb",
          5857 => x"39",
          5858 => x"f4",
          5859 => x"f8",
          5860 => x"ff",
          5861 => x"de",
          5862 => x"2e",
          5863 => x"b7",
          5864 => x"11",
          5865 => x"05",
          5866 => x"ec",
          5867 => x"c0",
          5868 => x"fa",
          5869 => x"3d",
          5870 => x"53",
          5871 => x"51",
          5872 => x"3f",
          5873 => x"08",
          5874 => x"de",
          5875 => x"81",
          5876 => x"fe",
          5877 => x"63",
          5878 => x"79",
          5879 => x"e6",
          5880 => x"78",
          5881 => x"05",
          5882 => x"7a",
          5883 => x"88",
          5884 => x"3d",
          5885 => x"53",
          5886 => x"51",
          5887 => x"3f",
          5888 => x"08",
          5889 => x"81",
          5890 => x"59",
          5891 => x"89",
          5892 => x"8c",
          5893 => x"cd",
          5894 => x"d5",
          5895 => x"80",
          5896 => x"81",
          5897 => x"44",
          5898 => x"db",
          5899 => x"78",
          5900 => x"38",
          5901 => x"08",
          5902 => x"81",
          5903 => x"59",
          5904 => x"88",
          5905 => x"a4",
          5906 => x"39",
          5907 => x"33",
          5908 => x"2e",
          5909 => x"db",
          5910 => x"89",
          5911 => x"bc",
          5912 => x"05",
          5913 => x"fe",
          5914 => x"fe",
          5915 => x"fe",
          5916 => x"81",
          5917 => x"80",
          5918 => x"db",
          5919 => x"78",
          5920 => x"38",
          5921 => x"08",
          5922 => x"39",
          5923 => x"33",
          5924 => x"2e",
          5925 => x"db",
          5926 => x"bb",
          5927 => x"d6",
          5928 => x"80",
          5929 => x"81",
          5930 => x"43",
          5931 => x"db",
          5932 => x"78",
          5933 => x"38",
          5934 => x"08",
          5935 => x"81",
          5936 => x"59",
          5937 => x"88",
          5938 => x"b0",
          5939 => x"39",
          5940 => x"08",
          5941 => x"b7",
          5942 => x"11",
          5943 => x"05",
          5944 => x"b4",
          5945 => x"c0",
          5946 => x"9b",
          5947 => x"5b",
          5948 => x"2e",
          5949 => x"59",
          5950 => x"8d",
          5951 => x"2e",
          5952 => x"a0",
          5953 => x"88",
          5954 => x"e4",
          5955 => x"af",
          5956 => x"63",
          5957 => x"62",
          5958 => x"ed",
          5959 => x"d7",
          5960 => x"e0",
          5961 => x"fe",
          5962 => x"fe",
          5963 => x"fe",
          5964 => x"81",
          5965 => x"80",
          5966 => x"38",
          5967 => x"f0",
          5968 => x"f8",
          5969 => x"fb",
          5970 => x"de",
          5971 => x"2e",
          5972 => x"59",
          5973 => x"05",
          5974 => x"63",
          5975 => x"b7",
          5976 => x"11",
          5977 => x"05",
          5978 => x"ac",
          5979 => x"c0",
          5980 => x"f7",
          5981 => x"70",
          5982 => x"81",
          5983 => x"fe",
          5984 => x"80",
          5985 => x"51",
          5986 => x"3f",
          5987 => x"33",
          5988 => x"2e",
          5989 => x"9f",
          5990 => x"38",
          5991 => x"f0",
          5992 => x"f8",
          5993 => x"fa",
          5994 => x"de",
          5995 => x"2e",
          5996 => x"59",
          5997 => x"05",
          5998 => x"63",
          5999 => x"ff",
          6000 => x"d8",
          6001 => x"f2",
          6002 => x"aa",
          6003 => x"fe",
          6004 => x"fe",
          6005 => x"fe",
          6006 => x"81",
          6007 => x"80",
          6008 => x"38",
          6009 => x"e4",
          6010 => x"f8",
          6011 => x"fc",
          6012 => x"de",
          6013 => x"2e",
          6014 => x"59",
          6015 => x"22",
          6016 => x"05",
          6017 => x"41",
          6018 => x"e4",
          6019 => x"f8",
          6020 => x"fb",
          6021 => x"de",
          6022 => x"38",
          6023 => x"60",
          6024 => x"52",
          6025 => x"51",
          6026 => x"3f",
          6027 => x"79",
          6028 => x"c9",
          6029 => x"79",
          6030 => x"ae",
          6031 => x"38",
          6032 => x"87",
          6033 => x"05",
          6034 => x"b7",
          6035 => x"11",
          6036 => x"05",
          6037 => x"b2",
          6038 => x"c0",
          6039 => x"92",
          6040 => x"02",
          6041 => x"79",
          6042 => x"5b",
          6043 => x"ff",
          6044 => x"d8",
          6045 => x"f1",
          6046 => x"a3",
          6047 => x"fe",
          6048 => x"fe",
          6049 => x"fe",
          6050 => x"81",
          6051 => x"80",
          6052 => x"38",
          6053 => x"e4",
          6054 => x"f8",
          6055 => x"fa",
          6056 => x"de",
          6057 => x"2e",
          6058 => x"60",
          6059 => x"60",
          6060 => x"b7",
          6061 => x"11",
          6062 => x"05",
          6063 => x"ca",
          6064 => x"c0",
          6065 => x"f4",
          6066 => x"70",
          6067 => x"81",
          6068 => x"fe",
          6069 => x"80",
          6070 => x"51",
          6071 => x"3f",
          6072 => x"33",
          6073 => x"2e",
          6074 => x"9f",
          6075 => x"38",
          6076 => x"e4",
          6077 => x"f8",
          6078 => x"fa",
          6079 => x"de",
          6080 => x"2e",
          6081 => x"60",
          6082 => x"60",
          6083 => x"ff",
          6084 => x"d8",
          6085 => x"f0",
          6086 => x"ae",
          6087 => x"fe",
          6088 => x"fe",
          6089 => x"fe",
          6090 => x"81",
          6091 => x"80",
          6092 => x"db",
          6093 => x"78",
          6094 => x"38",
          6095 => x"08",
          6096 => x"39",
          6097 => x"33",
          6098 => x"2e",
          6099 => x"db",
          6100 => x"bc",
          6101 => x"d6",
          6102 => x"80",
          6103 => x"81",
          6104 => x"44",
          6105 => x"db",
          6106 => x"78",
          6107 => x"38",
          6108 => x"08",
          6109 => x"81",
          6110 => x"59",
          6111 => x"88",
          6112 => x"ac",
          6113 => x"39",
          6114 => x"08",
          6115 => x"44",
          6116 => x"f0",
          6117 => x"f8",
          6118 => x"f6",
          6119 => x"de",
          6120 => x"de",
          6121 => x"d4",
          6122 => x"80",
          6123 => x"81",
          6124 => x"43",
          6125 => x"81",
          6126 => x"59",
          6127 => x"88",
          6128 => x"98",
          6129 => x"39",
          6130 => x"33",
          6131 => x"2e",
          6132 => x"db",
          6133 => x"aa",
          6134 => x"d7",
          6135 => x"80",
          6136 => x"81",
          6137 => x"43",
          6138 => x"db",
          6139 => x"78",
          6140 => x"38",
          6141 => x"08",
          6142 => x"81",
          6143 => x"88",
          6144 => x"3d",
          6145 => x"53",
          6146 => x"51",
          6147 => x"3f",
          6148 => x"08",
          6149 => x"de",
          6150 => x"81",
          6151 => x"fe",
          6152 => x"63",
          6153 => x"27",
          6154 => x"08",
          6155 => x"2e",
          6156 => x"8d",
          6157 => x"79",
          6158 => x"bc",
          6159 => x"e3",
          6160 => x"5a",
          6161 => x"d7",
          6162 => x"39",
          6163 => x"51",
          6164 => x"3f",
          6165 => x"ec",
          6166 => x"a4",
          6167 => x"e4",
          6168 => x"db",
          6169 => x"fe",
          6170 => x"f1",
          6171 => x"80",
          6172 => x"c0",
          6173 => x"84",
          6174 => x"87",
          6175 => x"0c",
          6176 => x"51",
          6177 => x"3f",
          6178 => x"81",
          6179 => x"fe",
          6180 => x"8c",
          6181 => x"87",
          6182 => x"0c",
          6183 => x"0b",
          6184 => x"94",
          6185 => x"39",
          6186 => x"f4",
          6187 => x"f8",
          6188 => x"f4",
          6189 => x"de",
          6190 => x"2e",
          6191 => x"63",
          6192 => x"a4",
          6193 => x"db",
          6194 => x"78",
          6195 => x"fe",
          6196 => x"fe",
          6197 => x"fe",
          6198 => x"81",
          6199 => x"80",
          6200 => x"38",
          6201 => x"d9",
          6202 => x"f2",
          6203 => x"59",
          6204 => x"de",
          6205 => x"81",
          6206 => x"80",
          6207 => x"38",
          6208 => x"08",
          6209 => x"dc",
          6210 => x"97",
          6211 => x"39",
          6212 => x"51",
          6213 => x"3f",
          6214 => x"3f",
          6215 => x"81",
          6216 => x"fe",
          6217 => x"80",
          6218 => x"39",
          6219 => x"3f",
          6220 => x"64",
          6221 => x"59",
          6222 => x"ef",
          6223 => x"80",
          6224 => x"38",
          6225 => x"06",
          6226 => x"80",
          6227 => x"38",
          6228 => x"f8",
          6229 => x"d8",
          6230 => x"de",
          6231 => x"5d",
          6232 => x"2e",
          6233 => x"82",
          6234 => x"7b",
          6235 => x"38",
          6236 => x"7b",
          6237 => x"38",
          6238 => x"81",
          6239 => x"7a",
          6240 => x"ac",
          6241 => x"81",
          6242 => x"b7",
          6243 => x"05",
          6244 => x"a5",
          6245 => x"81",
          6246 => x"b7",
          6247 => x"05",
          6248 => x"95",
          6249 => x"7a",
          6250 => x"ac",
          6251 => x"81",
          6252 => x"b7",
          6253 => x"05",
          6254 => x"fd",
          6255 => x"7a",
          6256 => x"81",
          6257 => x"b7",
          6258 => x"05",
          6259 => x"e9",
          6260 => x"8c",
          6261 => x"f4",
          6262 => x"64",
          6263 => x"81",
          6264 => x"54",
          6265 => x"53",
          6266 => x"52",
          6267 => x"b0",
          6268 => x"e5",
          6269 => x"c0",
          6270 => x"c0",
          6271 => x"30",
          6272 => x"80",
          6273 => x"5b",
          6274 => x"26",
          6275 => x"80",
          6276 => x"81",
          6277 => x"ff",
          6278 => x"7b",
          6279 => x"7e",
          6280 => x"81",
          6281 => x"78",
          6282 => x"ff",
          6283 => x"06",
          6284 => x"81",
          6285 => x"fe",
          6286 => x"ed",
          6287 => x"3d",
          6288 => x"81",
          6289 => x"87",
          6290 => x"70",
          6291 => x"87",
          6292 => x"72",
          6293 => x"9f",
          6294 => x"c0",
          6295 => x"75",
          6296 => x"87",
          6297 => x"73",
          6298 => x"8b",
          6299 => x"de",
          6300 => x"75",
          6301 => x"94",
          6302 => x"54",
          6303 => x"80",
          6304 => x"fe",
          6305 => x"81",
          6306 => x"90",
          6307 => x"55",
          6308 => x"80",
          6309 => x"fe",
          6310 => x"72",
          6311 => x"08",
          6312 => x"8c",
          6313 => x"87",
          6314 => x"0c",
          6315 => x"0b",
          6316 => x"94",
          6317 => x"0b",
          6318 => x"0c",
          6319 => x"81",
          6320 => x"fe",
          6321 => x"fe",
          6322 => x"81",
          6323 => x"fe",
          6324 => x"81",
          6325 => x"fe",
          6326 => x"81",
          6327 => x"fe",
          6328 => x"81",
          6329 => x"3f",
          6330 => x"80",
          6331 => x"00",
          6332 => x"ff",
          6333 => x"ff",
          6334 => x"ff",
          6335 => x"00",
          6336 => x"61",
          6337 => x"67",
          6338 => x"6d",
          6339 => x"73",
          6340 => x"79",
          6341 => x"91",
          6342 => x"15",
          6343 => x"1c",
          6344 => x"23",
          6345 => x"2a",
          6346 => x"31",
          6347 => x"38",
          6348 => x"3f",
          6349 => x"46",
          6350 => x"4d",
          6351 => x"54",
          6352 => x"5b",
          6353 => x"61",
          6354 => x"67",
          6355 => x"6d",
          6356 => x"73",
          6357 => x"79",
          6358 => x"7f",
          6359 => x"85",
          6360 => x"8b",
          6361 => x"25",
          6362 => x"64",
          6363 => x"3a",
          6364 => x"25",
          6365 => x"64",
          6366 => x"00",
          6367 => x"20",
          6368 => x"66",
          6369 => x"72",
          6370 => x"6f",
          6371 => x"00",
          6372 => x"72",
          6373 => x"53",
          6374 => x"63",
          6375 => x"69",
          6376 => x"00",
          6377 => x"65",
          6378 => x"65",
          6379 => x"6d",
          6380 => x"6d",
          6381 => x"65",
          6382 => x"00",
          6383 => x"20",
          6384 => x"53",
          6385 => x"4d",
          6386 => x"25",
          6387 => x"3a",
          6388 => x"58",
          6389 => x"00",
          6390 => x"20",
          6391 => x"41",
          6392 => x"20",
          6393 => x"25",
          6394 => x"3a",
          6395 => x"58",
          6396 => x"00",
          6397 => x"20",
          6398 => x"4e",
          6399 => x"41",
          6400 => x"25",
          6401 => x"3a",
          6402 => x"58",
          6403 => x"00",
          6404 => x"20",
          6405 => x"4d",
          6406 => x"20",
          6407 => x"25",
          6408 => x"3a",
          6409 => x"58",
          6410 => x"00",
          6411 => x"20",
          6412 => x"20",
          6413 => x"20",
          6414 => x"25",
          6415 => x"3a",
          6416 => x"58",
          6417 => x"00",
          6418 => x"20",
          6419 => x"43",
          6420 => x"20",
          6421 => x"44",
          6422 => x"63",
          6423 => x"3d",
          6424 => x"64",
          6425 => x"00",
          6426 => x"20",
          6427 => x"45",
          6428 => x"20",
          6429 => x"54",
          6430 => x"72",
          6431 => x"3d",
          6432 => x"64",
          6433 => x"00",
          6434 => x"20",
          6435 => x"52",
          6436 => x"52",
          6437 => x"43",
          6438 => x"6e",
          6439 => x"3d",
          6440 => x"64",
          6441 => x"00",
          6442 => x"20",
          6443 => x"48",
          6444 => x"45",
          6445 => x"53",
          6446 => x"00",
          6447 => x"20",
          6448 => x"49",
          6449 => x"00",
          6450 => x"20",
          6451 => x"54",
          6452 => x"00",
          6453 => x"20",
          6454 => x"0a",
          6455 => x"00",
          6456 => x"20",
          6457 => x"0a",
          6458 => x"00",
          6459 => x"72",
          6460 => x"65",
          6461 => x"00",
          6462 => x"20",
          6463 => x"20",
          6464 => x"65",
          6465 => x"65",
          6466 => x"72",
          6467 => x"64",
          6468 => x"73",
          6469 => x"25",
          6470 => x"0a",
          6471 => x"00",
          6472 => x"20",
          6473 => x"20",
          6474 => x"6f",
          6475 => x"53",
          6476 => x"74",
          6477 => x"64",
          6478 => x"73",
          6479 => x"25",
          6480 => x"0a",
          6481 => x"00",
          6482 => x"20",
          6483 => x"63",
          6484 => x"74",
          6485 => x"20",
          6486 => x"72",
          6487 => x"20",
          6488 => x"20",
          6489 => x"25",
          6490 => x"0a",
          6491 => x"00",
          6492 => x"63",
          6493 => x"00",
          6494 => x"20",
          6495 => x"20",
          6496 => x"20",
          6497 => x"20",
          6498 => x"20",
          6499 => x"20",
          6500 => x"20",
          6501 => x"25",
          6502 => x"0a",
          6503 => x"00",
          6504 => x"20",
          6505 => x"74",
          6506 => x"43",
          6507 => x"6b",
          6508 => x"65",
          6509 => x"20",
          6510 => x"20",
          6511 => x"25",
          6512 => x"30",
          6513 => x"48",
          6514 => x"00",
          6515 => x"20",
          6516 => x"41",
          6517 => x"6c",
          6518 => x"20",
          6519 => x"71",
          6520 => x"20",
          6521 => x"20",
          6522 => x"25",
          6523 => x"30",
          6524 => x"48",
          6525 => x"00",
          6526 => x"20",
          6527 => x"68",
          6528 => x"65",
          6529 => x"52",
          6530 => x"43",
          6531 => x"6b",
          6532 => x"65",
          6533 => x"25",
          6534 => x"30",
          6535 => x"48",
          6536 => x"00",
          6537 => x"6c",
          6538 => x"00",
          6539 => x"69",
          6540 => x"00",
          6541 => x"78",
          6542 => x"00",
          6543 => x"00",
          6544 => x"6d",
          6545 => x"00",
          6546 => x"6e",
          6547 => x"00",
          6548 => x"00",
          6549 => x"2c",
          6550 => x"3d",
          6551 => x"5d",
          6552 => x"00",
          6553 => x"00",
          6554 => x"33",
          6555 => x"00",
          6556 => x"4d",
          6557 => x"53",
          6558 => x"00",
          6559 => x"4e",
          6560 => x"20",
          6561 => x"46",
          6562 => x"32",
          6563 => x"00",
          6564 => x"4e",
          6565 => x"20",
          6566 => x"46",
          6567 => x"20",
          6568 => x"00",
          6569 => x"50",
          6570 => x"00",
          6571 => x"00",
          6572 => x"00",
          6573 => x"41",
          6574 => x"80",
          6575 => x"49",
          6576 => x"8f",
          6577 => x"4f",
          6578 => x"55",
          6579 => x"9b",
          6580 => x"9f",
          6581 => x"55",
          6582 => x"a7",
          6583 => x"ab",
          6584 => x"af",
          6585 => x"b3",
          6586 => x"b7",
          6587 => x"bb",
          6588 => x"bf",
          6589 => x"c3",
          6590 => x"c7",
          6591 => x"cb",
          6592 => x"cf",
          6593 => x"d3",
          6594 => x"d7",
          6595 => x"db",
          6596 => x"df",
          6597 => x"e3",
          6598 => x"e7",
          6599 => x"eb",
          6600 => x"ef",
          6601 => x"f3",
          6602 => x"f7",
          6603 => x"fb",
          6604 => x"ff",
          6605 => x"3b",
          6606 => x"2f",
          6607 => x"3a",
          6608 => x"7c",
          6609 => x"00",
          6610 => x"04",
          6611 => x"40",
          6612 => x"00",
          6613 => x"00",
          6614 => x"02",
          6615 => x"08",
          6616 => x"20",
          6617 => x"00",
          6618 => x"69",
          6619 => x"00",
          6620 => x"63",
          6621 => x"00",
          6622 => x"69",
          6623 => x"00",
          6624 => x"61",
          6625 => x"00",
          6626 => x"65",
          6627 => x"00",
          6628 => x"65",
          6629 => x"00",
          6630 => x"6d",
          6631 => x"00",
          6632 => x"63",
          6633 => x"00",
          6634 => x"00",
          6635 => x"00",
          6636 => x"00",
          6637 => x"00",
          6638 => x"00",
          6639 => x"00",
          6640 => x"00",
          6641 => x"6c",
          6642 => x"00",
          6643 => x"00",
          6644 => x"74",
          6645 => x"00",
          6646 => x"65",
          6647 => x"00",
          6648 => x"6f",
          6649 => x"00",
          6650 => x"74",
          6651 => x"00",
          6652 => x"6b",
          6653 => x"72",
          6654 => x"00",
          6655 => x"65",
          6656 => x"6c",
          6657 => x"72",
          6658 => x"0a",
          6659 => x"00",
          6660 => x"6b",
          6661 => x"74",
          6662 => x"61",
          6663 => x"0a",
          6664 => x"00",
          6665 => x"66",
          6666 => x"20",
          6667 => x"6e",
          6668 => x"00",
          6669 => x"70",
          6670 => x"20",
          6671 => x"6e",
          6672 => x"00",
          6673 => x"61",
          6674 => x"20",
          6675 => x"65",
          6676 => x"65",
          6677 => x"00",
          6678 => x"65",
          6679 => x"64",
          6680 => x"65",
          6681 => x"00",
          6682 => x"65",
          6683 => x"72",
          6684 => x"79",
          6685 => x"69",
          6686 => x"2e",
          6687 => x"00",
          6688 => x"65",
          6689 => x"6e",
          6690 => x"20",
          6691 => x"61",
          6692 => x"2e",
          6693 => x"00",
          6694 => x"69",
          6695 => x"72",
          6696 => x"20",
          6697 => x"74",
          6698 => x"65",
          6699 => x"00",
          6700 => x"76",
          6701 => x"75",
          6702 => x"72",
          6703 => x"20",
          6704 => x"61",
          6705 => x"2e",
          6706 => x"00",
          6707 => x"6b",
          6708 => x"74",
          6709 => x"61",
          6710 => x"64",
          6711 => x"00",
          6712 => x"63",
          6713 => x"61",
          6714 => x"6c",
          6715 => x"69",
          6716 => x"79",
          6717 => x"6d",
          6718 => x"75",
          6719 => x"6f",
          6720 => x"69",
          6721 => x"0a",
          6722 => x"00",
          6723 => x"6d",
          6724 => x"61",
          6725 => x"74",
          6726 => x"0a",
          6727 => x"00",
          6728 => x"65",
          6729 => x"2c",
          6730 => x"65",
          6731 => x"69",
          6732 => x"63",
          6733 => x"65",
          6734 => x"64",
          6735 => x"00",
          6736 => x"65",
          6737 => x"20",
          6738 => x"6b",
          6739 => x"0a",
          6740 => x"00",
          6741 => x"75",
          6742 => x"63",
          6743 => x"74",
          6744 => x"6d",
          6745 => x"2e",
          6746 => x"00",
          6747 => x"20",
          6748 => x"79",
          6749 => x"65",
          6750 => x"69",
          6751 => x"2e",
          6752 => x"00",
          6753 => x"61",
          6754 => x"65",
          6755 => x"69",
          6756 => x"72",
          6757 => x"74",
          6758 => x"00",
          6759 => x"63",
          6760 => x"2e",
          6761 => x"00",
          6762 => x"6e",
          6763 => x"20",
          6764 => x"6f",
          6765 => x"00",
          6766 => x"75",
          6767 => x"74",
          6768 => x"25",
          6769 => x"74",
          6770 => x"75",
          6771 => x"74",
          6772 => x"73",
          6773 => x"0a",
          6774 => x"00",
          6775 => x"58",
          6776 => x"00",
          6777 => x"00",
          6778 => x"58",
          6779 => x"00",
          6780 => x"20",
          6781 => x"20",
          6782 => x"00",
          6783 => x"58",
          6784 => x"00",
          6785 => x"00",
          6786 => x"00",
          6787 => x"00",
          6788 => x"64",
          6789 => x"00",
          6790 => x"54",
          6791 => x"00",
          6792 => x"20",
          6793 => x"28",
          6794 => x"00",
          6795 => x"31",
          6796 => x"30",
          6797 => x"00",
          6798 => x"34",
          6799 => x"00",
          6800 => x"55",
          6801 => x"65",
          6802 => x"30",
          6803 => x"20",
          6804 => x"25",
          6805 => x"2a",
          6806 => x"00",
          6807 => x"54",
          6808 => x"6e",
          6809 => x"72",
          6810 => x"20",
          6811 => x"64",
          6812 => x"0a",
          6813 => x"00",
          6814 => x"65",
          6815 => x"6e",
          6816 => x"72",
          6817 => x"0a",
          6818 => x"00",
          6819 => x"20",
          6820 => x"65",
          6821 => x"70",
          6822 => x"00",
          6823 => x"54",
          6824 => x"44",
          6825 => x"74",
          6826 => x"75",
          6827 => x"00",
          6828 => x"54",
          6829 => x"52",
          6830 => x"74",
          6831 => x"75",
          6832 => x"00",
          6833 => x"54",
          6834 => x"58",
          6835 => x"74",
          6836 => x"75",
          6837 => x"00",
          6838 => x"54",
          6839 => x"58",
          6840 => x"74",
          6841 => x"75",
          6842 => x"00",
          6843 => x"54",
          6844 => x"58",
          6845 => x"74",
          6846 => x"75",
          6847 => x"00",
          6848 => x"54",
          6849 => x"58",
          6850 => x"74",
          6851 => x"75",
          6852 => x"00",
          6853 => x"74",
          6854 => x"20",
          6855 => x"74",
          6856 => x"72",
          6857 => x"0a",
          6858 => x"00",
          6859 => x"62",
          6860 => x"67",
          6861 => x"6d",
          6862 => x"2e",
          6863 => x"00",
          6864 => x"6f",
          6865 => x"63",
          6866 => x"74",
          6867 => x"00",
          6868 => x"00",
          6869 => x"6c",
          6870 => x"74",
          6871 => x"6e",
          6872 => x"61",
          6873 => x"65",
          6874 => x"20",
          6875 => x"64",
          6876 => x"20",
          6877 => x"61",
          6878 => x"69",
          6879 => x"20",
          6880 => x"75",
          6881 => x"79",
          6882 => x"00",
          6883 => x"00",
          6884 => x"20",
          6885 => x"6b",
          6886 => x"21",
          6887 => x"00",
          6888 => x"74",
          6889 => x"69",
          6890 => x"2e",
          6891 => x"00",
          6892 => x"6c",
          6893 => x"74",
          6894 => x"6e",
          6895 => x"61",
          6896 => x"65",
          6897 => x"00",
          6898 => x"25",
          6899 => x"00",
          6900 => x"00",
          6901 => x"61",
          6902 => x"67",
          6903 => x"2e",
          6904 => x"00",
          6905 => x"70",
          6906 => x"6d",
          6907 => x"0a",
          6908 => x"00",
          6909 => x"6d",
          6910 => x"74",
          6911 => x"00",
          6912 => x"58",
          6913 => x"32",
          6914 => x"00",
          6915 => x"0a",
          6916 => x"00",
          6917 => x"58",
          6918 => x"34",
          6919 => x"00",
          6920 => x"58",
          6921 => x"38",
          6922 => x"00",
          6923 => x"72",
          6924 => x"6e",
          6925 => x"0a",
          6926 => x"00",
          6927 => x"6c",
          6928 => x"25",
          6929 => x"78",
          6930 => x"00",
          6931 => x"61",
          6932 => x"6e",
          6933 => x"6e",
          6934 => x"72",
          6935 => x"73",
          6936 => x"00",
          6937 => x"62",
          6938 => x"67",
          6939 => x"74",
          6940 => x"75",
          6941 => x"0a",
          6942 => x"00",
          6943 => x"61",
          6944 => x"64",
          6945 => x"72",
          6946 => x"69",
          6947 => x"00",
          6948 => x"62",
          6949 => x"67",
          6950 => x"72",
          6951 => x"69",
          6952 => x"00",
          6953 => x"63",
          6954 => x"6e",
          6955 => x"6f",
          6956 => x"40",
          6957 => x"38",
          6958 => x"2e",
          6959 => x"00",
          6960 => x"6c",
          6961 => x"20",
          6962 => x"65",
          6963 => x"25",
          6964 => x"20",
          6965 => x"0a",
          6966 => x"00",
          6967 => x"6c",
          6968 => x"74",
          6969 => x"65",
          6970 => x"6f",
          6971 => x"28",
          6972 => x"2e",
          6973 => x"00",
          6974 => x"74",
          6975 => x"69",
          6976 => x"61",
          6977 => x"69",
          6978 => x"69",
          6979 => x"2e",
          6980 => x"00",
          6981 => x"64",
          6982 => x"62",
          6983 => x"69",
          6984 => x"2e",
          6985 => x"00",
          6986 => x"00",
          6987 => x"00",
          6988 => x"5c",
          6989 => x"25",
          6990 => x"73",
          6991 => x"00",
          6992 => x"5c",
          6993 => x"25",
          6994 => x"00",
          6995 => x"5c",
          6996 => x"00",
          6997 => x"20",
          6998 => x"6d",
          6999 => x"2e",
          7000 => x"00",
          7001 => x"6e",
          7002 => x"2e",
          7003 => x"00",
          7004 => x"62",
          7005 => x"67",
          7006 => x"74",
          7007 => x"75",
          7008 => x"2e",
          7009 => x"00",
          7010 => x"00",
          7011 => x"00",
          7012 => x"ff",
          7013 => x"00",
          7014 => x"ff",
          7015 => x"00",
          7016 => x"ff",
          7017 => x"00",
          7018 => x"00",
          7019 => x"00",
          7020 => x"ff",
          7021 => x"00",
          7022 => x"00",
          7023 => x"00",
          7024 => x"00",
          7025 => x"00",
          7026 => x"00",
          7027 => x"00",
          7028 => x"00",
          7029 => x"01",
          7030 => x"01",
          7031 => x"01",
          7032 => x"00",
          7033 => x"00",
          7034 => x"00",
          7035 => x"00",
          7036 => x"68",
          7037 => x"00",
          7038 => x"00",
          7039 => x"00",
          7040 => x"70",
          7041 => x"00",
          7042 => x"00",
          7043 => x"00",
          7044 => x"78",
          7045 => x"00",
          7046 => x"00",
          7047 => x"00",
          7048 => x"80",
          7049 => x"00",
          7050 => x"00",
          7051 => x"00",
          7052 => x"88",
          7053 => x"00",
          7054 => x"00",
          7055 => x"00",
          7056 => x"90",
          7057 => x"00",
          7058 => x"00",
          7059 => x"00",
          7060 => x"98",
          7061 => x"00",
          7062 => x"00",
          7063 => x"00",
          7064 => x"a0",
          7065 => x"00",
          7066 => x"00",
          7067 => x"00",
          7068 => x"a8",
          7069 => x"00",
          7070 => x"00",
          7071 => x"00",
          7072 => x"ac",
          7073 => x"00",
          7074 => x"00",
          7075 => x"00",
          7076 => x"b0",
          7077 => x"00",
          7078 => x"00",
          7079 => x"00",
          7080 => x"b4",
          7081 => x"00",
          7082 => x"00",
          7083 => x"00",
          7084 => x"b8",
          7085 => x"00",
          7086 => x"00",
          7087 => x"00",
          7088 => x"bc",
          7089 => x"00",
          7090 => x"00",
          7091 => x"00",
          7092 => x"c0",
          7093 => x"00",
          7094 => x"00",
          7095 => x"00",
          7096 => x"c4",
          7097 => x"00",
          7098 => x"00",
          7099 => x"00",
          7100 => x"cc",
          7101 => x"00",
          7102 => x"00",
          7103 => x"00",
          7104 => x"d0",
          7105 => x"00",
          7106 => x"00",
          7107 => x"00",
          7108 => x"d8",
          7109 => x"00",
          7110 => x"00",
          7111 => x"00",
          7112 => x"e0",
          7113 => x"00",
          7114 => x"00",
          7115 => x"00",
          7116 => x"e8",
          7117 => x"00",
          7118 => x"00",
          7119 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"92",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"81",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a3",
           270 => x"0b",
           271 => x"0b",
           272 => x"c1",
           273 => x"0b",
           274 => x"0b",
           275 => x"df",
           276 => x"0b",
           277 => x"0b",
           278 => x"fd",
           279 => x"0b",
           280 => x"0b",
           281 => x"9b",
           282 => x"0b",
           283 => x"0b",
           284 => x"b9",
           285 => x"0b",
           286 => x"0b",
           287 => x"d7",
           288 => x"0b",
           289 => x"0b",
           290 => x"f5",
           291 => x"0b",
           292 => x"0b",
           293 => x"94",
           294 => x"0b",
           295 => x"0b",
           296 => x"b4",
           297 => x"0b",
           298 => x"0b",
           299 => x"d4",
           300 => x"0b",
           301 => x"0b",
           302 => x"f4",
           303 => x"0b",
           304 => x"0b",
           305 => x"94",
           306 => x"0b",
           307 => x"0b",
           308 => x"b4",
           309 => x"0b",
           310 => x"0b",
           311 => x"d4",
           312 => x"0b",
           313 => x"0b",
           314 => x"f4",
           315 => x"0b",
           316 => x"0b",
           317 => x"94",
           318 => x"0b",
           319 => x"0b",
           320 => x"b4",
           321 => x"0b",
           322 => x"0b",
           323 => x"d4",
           324 => x"0b",
           325 => x"0b",
           326 => x"f4",
           327 => x"0b",
           328 => x"0b",
           329 => x"94",
           330 => x"0b",
           331 => x"0b",
           332 => x"b2",
           333 => x"0b",
           334 => x"0b",
           335 => x"d0",
           336 => x"0b",
           337 => x"0b",
           338 => x"ee",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"de",
           386 => x"ae",
           387 => x"cc",
           388 => x"90",
           389 => x"cc",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"81",
           395 => x"82",
           396 => x"81",
           397 => x"ae",
           398 => x"de",
           399 => x"80",
           400 => x"de",
           401 => x"fd",
           402 => x"cc",
           403 => x"90",
           404 => x"cc",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"81",
           410 => x"82",
           411 => x"81",
           412 => x"b6",
           413 => x"de",
           414 => x"80",
           415 => x"de",
           416 => x"8a",
           417 => x"cc",
           418 => x"90",
           419 => x"cc",
           420 => x"2d",
           421 => x"08",
           422 => x"04",
           423 => x"0c",
           424 => x"81",
           425 => x"82",
           426 => x"81",
           427 => x"b4",
           428 => x"de",
           429 => x"80",
           430 => x"de",
           431 => x"bb",
           432 => x"cc",
           433 => x"90",
           434 => x"cc",
           435 => x"2d",
           436 => x"08",
           437 => x"04",
           438 => x"0c",
           439 => x"81",
           440 => x"82",
           441 => x"81",
           442 => x"9c",
           443 => x"de",
           444 => x"80",
           445 => x"de",
           446 => x"90",
           447 => x"cc",
           448 => x"90",
           449 => x"cc",
           450 => x"bf",
           451 => x"cc",
           452 => x"90",
           453 => x"cc",
           454 => x"b0",
           455 => x"cc",
           456 => x"90",
           457 => x"cc",
           458 => x"a4",
           459 => x"cc",
           460 => x"90",
           461 => x"cc",
           462 => x"a1",
           463 => x"cc",
           464 => x"90",
           465 => x"cc",
           466 => x"bf",
           467 => x"cc",
           468 => x"90",
           469 => x"cc",
           470 => x"9f",
           471 => x"cc",
           472 => x"90",
           473 => x"cc",
           474 => x"92",
           475 => x"cc",
           476 => x"90",
           477 => x"cc",
           478 => x"de",
           479 => x"cc",
           480 => x"90",
           481 => x"cc",
           482 => x"fd",
           483 => x"cc",
           484 => x"90",
           485 => x"cc",
           486 => x"9c",
           487 => x"cc",
           488 => x"90",
           489 => x"cc",
           490 => x"86",
           491 => x"cc",
           492 => x"90",
           493 => x"cc",
           494 => x"ec",
           495 => x"cc",
           496 => x"90",
           497 => x"cc",
           498 => x"da",
           499 => x"cc",
           500 => x"90",
           501 => x"cc",
           502 => x"a0",
           503 => x"cc",
           504 => x"90",
           505 => x"cc",
           506 => x"da",
           507 => x"cc",
           508 => x"90",
           509 => x"cc",
           510 => x"db",
           511 => x"cc",
           512 => x"90",
           513 => x"cc",
           514 => x"90",
           515 => x"cc",
           516 => x"90",
           517 => x"cc",
           518 => x"e9",
           519 => x"cc",
           520 => x"90",
           521 => x"cc",
           522 => x"94",
           523 => x"cc",
           524 => x"90",
           525 => x"cc",
           526 => x"f7",
           527 => x"cc",
           528 => x"90",
           529 => x"cc",
           530 => x"cc",
           531 => x"cc",
           532 => x"90",
           533 => x"cc",
           534 => x"d6",
           535 => x"cc",
           536 => x"90",
           537 => x"cc",
           538 => x"98",
           539 => x"cc",
           540 => x"90",
           541 => x"cc",
           542 => x"de",
           543 => x"cc",
           544 => x"90",
           545 => x"cc",
           546 => x"84",
           547 => x"cc",
           548 => x"90",
           549 => x"cc",
           550 => x"2d",
           551 => x"08",
           552 => x"04",
           553 => x"0c",
           554 => x"81",
           555 => x"82",
           556 => x"81",
           557 => x"be",
           558 => x"de",
           559 => x"80",
           560 => x"de",
           561 => x"d1",
           562 => x"cc",
           563 => x"90",
           564 => x"cc",
           565 => x"2d",
           566 => x"08",
           567 => x"04",
           568 => x"0c",
           569 => x"81",
           570 => x"82",
           571 => x"81",
           572 => x"81",
           573 => x"81",
           574 => x"82",
           575 => x"3c",
           576 => x"10",
           577 => x"10",
           578 => x"10",
           579 => x"10",
           580 => x"10",
           581 => x"10",
           582 => x"10",
           583 => x"10",
           584 => x"00",
           585 => x"ff",
           586 => x"06",
           587 => x"83",
           588 => x"10",
           589 => x"fc",
           590 => x"51",
           591 => x"80",
           592 => x"ff",
           593 => x"06",
           594 => x"52",
           595 => x"0a",
           596 => x"38",
           597 => x"51",
           598 => x"c0",
           599 => x"ec",
           600 => x"80",
           601 => x"05",
           602 => x"0b",
           603 => x"04",
           604 => x"81",
           605 => x"00",
           606 => x"08",
           607 => x"cc",
           608 => x"0d",
           609 => x"de",
           610 => x"05",
           611 => x"de",
           612 => x"05",
           613 => x"d4",
           614 => x"c0",
           615 => x"de",
           616 => x"85",
           617 => x"de",
           618 => x"81",
           619 => x"02",
           620 => x"0c",
           621 => x"81",
           622 => x"cc",
           623 => x"08",
           624 => x"cc",
           625 => x"08",
           626 => x"3f",
           627 => x"08",
           628 => x"c0",
           629 => x"3d",
           630 => x"cc",
           631 => x"de",
           632 => x"81",
           633 => x"f9",
           634 => x"0b",
           635 => x"08",
           636 => x"81",
           637 => x"88",
           638 => x"25",
           639 => x"de",
           640 => x"05",
           641 => x"de",
           642 => x"05",
           643 => x"81",
           644 => x"f4",
           645 => x"de",
           646 => x"05",
           647 => x"81",
           648 => x"cc",
           649 => x"0c",
           650 => x"08",
           651 => x"81",
           652 => x"fc",
           653 => x"de",
           654 => x"05",
           655 => x"b9",
           656 => x"cc",
           657 => x"08",
           658 => x"cc",
           659 => x"0c",
           660 => x"de",
           661 => x"05",
           662 => x"cc",
           663 => x"08",
           664 => x"0b",
           665 => x"08",
           666 => x"81",
           667 => x"f0",
           668 => x"de",
           669 => x"05",
           670 => x"81",
           671 => x"8c",
           672 => x"81",
           673 => x"88",
           674 => x"81",
           675 => x"de",
           676 => x"81",
           677 => x"f8",
           678 => x"81",
           679 => x"fc",
           680 => x"2e",
           681 => x"de",
           682 => x"05",
           683 => x"de",
           684 => x"05",
           685 => x"cc",
           686 => x"08",
           687 => x"c0",
           688 => x"3d",
           689 => x"cc",
           690 => x"de",
           691 => x"81",
           692 => x"fb",
           693 => x"0b",
           694 => x"08",
           695 => x"81",
           696 => x"88",
           697 => x"25",
           698 => x"de",
           699 => x"05",
           700 => x"de",
           701 => x"05",
           702 => x"81",
           703 => x"fc",
           704 => x"de",
           705 => x"05",
           706 => x"90",
           707 => x"cc",
           708 => x"08",
           709 => x"cc",
           710 => x"0c",
           711 => x"de",
           712 => x"05",
           713 => x"de",
           714 => x"05",
           715 => x"3f",
           716 => x"08",
           717 => x"cc",
           718 => x"0c",
           719 => x"cc",
           720 => x"08",
           721 => x"38",
           722 => x"08",
           723 => x"30",
           724 => x"08",
           725 => x"81",
           726 => x"f8",
           727 => x"81",
           728 => x"54",
           729 => x"81",
           730 => x"04",
           731 => x"08",
           732 => x"cc",
           733 => x"0d",
           734 => x"de",
           735 => x"05",
           736 => x"81",
           737 => x"f8",
           738 => x"de",
           739 => x"05",
           740 => x"cc",
           741 => x"08",
           742 => x"81",
           743 => x"fc",
           744 => x"2e",
           745 => x"0b",
           746 => x"08",
           747 => x"24",
           748 => x"de",
           749 => x"05",
           750 => x"de",
           751 => x"05",
           752 => x"cc",
           753 => x"08",
           754 => x"cc",
           755 => x"0c",
           756 => x"81",
           757 => x"fc",
           758 => x"2e",
           759 => x"81",
           760 => x"8c",
           761 => x"de",
           762 => x"05",
           763 => x"38",
           764 => x"08",
           765 => x"81",
           766 => x"8c",
           767 => x"81",
           768 => x"88",
           769 => x"de",
           770 => x"05",
           771 => x"cc",
           772 => x"08",
           773 => x"cc",
           774 => x"0c",
           775 => x"08",
           776 => x"81",
           777 => x"cc",
           778 => x"0c",
           779 => x"08",
           780 => x"81",
           781 => x"cc",
           782 => x"0c",
           783 => x"81",
           784 => x"90",
           785 => x"2e",
           786 => x"de",
           787 => x"05",
           788 => x"de",
           789 => x"05",
           790 => x"39",
           791 => x"08",
           792 => x"70",
           793 => x"08",
           794 => x"51",
           795 => x"08",
           796 => x"81",
           797 => x"85",
           798 => x"de",
           799 => x"fc",
           800 => x"79",
           801 => x"05",
           802 => x"57",
           803 => x"83",
           804 => x"38",
           805 => x"51",
           806 => x"a4",
           807 => x"52",
           808 => x"93",
           809 => x"70",
           810 => x"34",
           811 => x"71",
           812 => x"81",
           813 => x"74",
           814 => x"0c",
           815 => x"04",
           816 => x"2b",
           817 => x"71",
           818 => x"51",
           819 => x"72",
           820 => x"72",
           821 => x"05",
           822 => x"71",
           823 => x"53",
           824 => x"70",
           825 => x"0c",
           826 => x"84",
           827 => x"f0",
           828 => x"8f",
           829 => x"83",
           830 => x"38",
           831 => x"84",
           832 => x"fc",
           833 => x"83",
           834 => x"70",
           835 => x"39",
           836 => x"77",
           837 => x"07",
           838 => x"54",
           839 => x"38",
           840 => x"08",
           841 => x"71",
           842 => x"80",
           843 => x"75",
           844 => x"33",
           845 => x"06",
           846 => x"80",
           847 => x"72",
           848 => x"75",
           849 => x"06",
           850 => x"12",
           851 => x"33",
           852 => x"06",
           853 => x"52",
           854 => x"72",
           855 => x"81",
           856 => x"81",
           857 => x"71",
           858 => x"c0",
           859 => x"87",
           860 => x"71",
           861 => x"fb",
           862 => x"06",
           863 => x"82",
           864 => x"51",
           865 => x"97",
           866 => x"84",
           867 => x"54",
           868 => x"75",
           869 => x"38",
           870 => x"52",
           871 => x"80",
           872 => x"c0",
           873 => x"0d",
           874 => x"0d",
           875 => x"53",
           876 => x"52",
           877 => x"81",
           878 => x"81",
           879 => x"07",
           880 => x"52",
           881 => x"e8",
           882 => x"de",
           883 => x"3d",
           884 => x"3d",
           885 => x"08",
           886 => x"56",
           887 => x"80",
           888 => x"33",
           889 => x"2e",
           890 => x"86",
           891 => x"52",
           892 => x"53",
           893 => x"13",
           894 => x"33",
           895 => x"06",
           896 => x"70",
           897 => x"38",
           898 => x"80",
           899 => x"74",
           900 => x"81",
           901 => x"70",
           902 => x"81",
           903 => x"80",
           904 => x"05",
           905 => x"76",
           906 => x"70",
           907 => x"0c",
           908 => x"04",
           909 => x"76",
           910 => x"80",
           911 => x"86",
           912 => x"52",
           913 => x"c3",
           914 => x"c0",
           915 => x"80",
           916 => x"74",
           917 => x"de",
           918 => x"3d",
           919 => x"3d",
           920 => x"11",
           921 => x"52",
           922 => x"70",
           923 => x"98",
           924 => x"33",
           925 => x"82",
           926 => x"26",
           927 => x"84",
           928 => x"83",
           929 => x"26",
           930 => x"85",
           931 => x"84",
           932 => x"26",
           933 => x"86",
           934 => x"85",
           935 => x"26",
           936 => x"88",
           937 => x"86",
           938 => x"e7",
           939 => x"38",
           940 => x"54",
           941 => x"87",
           942 => x"cc",
           943 => x"87",
           944 => x"0c",
           945 => x"c0",
           946 => x"82",
           947 => x"c0",
           948 => x"83",
           949 => x"c0",
           950 => x"84",
           951 => x"c0",
           952 => x"85",
           953 => x"c0",
           954 => x"86",
           955 => x"c0",
           956 => x"74",
           957 => x"a4",
           958 => x"c0",
           959 => x"80",
           960 => x"98",
           961 => x"52",
           962 => x"c0",
           963 => x"0d",
           964 => x"0d",
           965 => x"c0",
           966 => x"81",
           967 => x"c0",
           968 => x"5e",
           969 => x"87",
           970 => x"08",
           971 => x"1c",
           972 => x"98",
           973 => x"79",
           974 => x"87",
           975 => x"08",
           976 => x"1c",
           977 => x"98",
           978 => x"79",
           979 => x"87",
           980 => x"08",
           981 => x"1c",
           982 => x"98",
           983 => x"7b",
           984 => x"87",
           985 => x"08",
           986 => x"1c",
           987 => x"0c",
           988 => x"ff",
           989 => x"83",
           990 => x"58",
           991 => x"57",
           992 => x"56",
           993 => x"55",
           994 => x"54",
           995 => x"53",
           996 => x"ff",
           997 => x"c6",
           998 => x"88",
           999 => x"0d",
          1000 => x"0d",
          1001 => x"33",
          1002 => x"9f",
          1003 => x"52",
          1004 => x"81",
          1005 => x"83",
          1006 => x"fb",
          1007 => x"0b",
          1008 => x"88",
          1009 => x"ff",
          1010 => x"56",
          1011 => x"84",
          1012 => x"2e",
          1013 => x"c0",
          1014 => x"70",
          1015 => x"2a",
          1016 => x"53",
          1017 => x"80",
          1018 => x"71",
          1019 => x"81",
          1020 => x"70",
          1021 => x"81",
          1022 => x"06",
          1023 => x"80",
          1024 => x"71",
          1025 => x"81",
          1026 => x"70",
          1027 => x"73",
          1028 => x"51",
          1029 => x"80",
          1030 => x"2e",
          1031 => x"c0",
          1032 => x"75",
          1033 => x"81",
          1034 => x"87",
          1035 => x"fb",
          1036 => x"9f",
          1037 => x"0b",
          1038 => x"33",
          1039 => x"06",
          1040 => x"87",
          1041 => x"51",
          1042 => x"86",
          1043 => x"94",
          1044 => x"08",
          1045 => x"70",
          1046 => x"54",
          1047 => x"2e",
          1048 => x"91",
          1049 => x"06",
          1050 => x"d7",
          1051 => x"32",
          1052 => x"51",
          1053 => x"2e",
          1054 => x"93",
          1055 => x"06",
          1056 => x"ff",
          1057 => x"81",
          1058 => x"87",
          1059 => x"52",
          1060 => x"86",
          1061 => x"94",
          1062 => x"72",
          1063 => x"0d",
          1064 => x"0d",
          1065 => x"74",
          1066 => x"ff",
          1067 => x"57",
          1068 => x"80",
          1069 => x"81",
          1070 => x"15",
          1071 => x"db",
          1072 => x"81",
          1073 => x"57",
          1074 => x"c0",
          1075 => x"75",
          1076 => x"38",
          1077 => x"94",
          1078 => x"70",
          1079 => x"81",
          1080 => x"52",
          1081 => x"8c",
          1082 => x"2a",
          1083 => x"51",
          1084 => x"38",
          1085 => x"70",
          1086 => x"51",
          1087 => x"8d",
          1088 => x"2a",
          1089 => x"51",
          1090 => x"be",
          1091 => x"ff",
          1092 => x"c0",
          1093 => x"70",
          1094 => x"38",
          1095 => x"90",
          1096 => x"0c",
          1097 => x"33",
          1098 => x"06",
          1099 => x"70",
          1100 => x"76",
          1101 => x"0c",
          1102 => x"04",
          1103 => x"0b",
          1104 => x"88",
          1105 => x"ff",
          1106 => x"87",
          1107 => x"51",
          1108 => x"86",
          1109 => x"94",
          1110 => x"08",
          1111 => x"70",
          1112 => x"51",
          1113 => x"2e",
          1114 => x"81",
          1115 => x"87",
          1116 => x"52",
          1117 => x"86",
          1118 => x"94",
          1119 => x"08",
          1120 => x"06",
          1121 => x"0c",
          1122 => x"0d",
          1123 => x"0d",
          1124 => x"db",
          1125 => x"81",
          1126 => x"53",
          1127 => x"84",
          1128 => x"2e",
          1129 => x"c0",
          1130 => x"71",
          1131 => x"2a",
          1132 => x"51",
          1133 => x"52",
          1134 => x"a0",
          1135 => x"ff",
          1136 => x"c0",
          1137 => x"70",
          1138 => x"38",
          1139 => x"90",
          1140 => x"70",
          1141 => x"98",
          1142 => x"51",
          1143 => x"c0",
          1144 => x"0d",
          1145 => x"0d",
          1146 => x"80",
          1147 => x"2a",
          1148 => x"51",
          1149 => x"84",
          1150 => x"c0",
          1151 => x"81",
          1152 => x"87",
          1153 => x"08",
          1154 => x"0c",
          1155 => x"94",
          1156 => x"94",
          1157 => x"9e",
          1158 => x"db",
          1159 => x"c0",
          1160 => x"81",
          1161 => x"87",
          1162 => x"08",
          1163 => x"0c",
          1164 => x"ac",
          1165 => x"a4",
          1166 => x"9e",
          1167 => x"db",
          1168 => x"c0",
          1169 => x"81",
          1170 => x"87",
          1171 => x"08",
          1172 => x"0c",
          1173 => x"bc",
          1174 => x"b4",
          1175 => x"9e",
          1176 => x"db",
          1177 => x"c0",
          1178 => x"81",
          1179 => x"87",
          1180 => x"08",
          1181 => x"db",
          1182 => x"c0",
          1183 => x"81",
          1184 => x"87",
          1185 => x"08",
          1186 => x"0c",
          1187 => x"8c",
          1188 => x"cc",
          1189 => x"81",
          1190 => x"80",
          1191 => x"9e",
          1192 => x"84",
          1193 => x"51",
          1194 => x"80",
          1195 => x"81",
          1196 => x"db",
          1197 => x"0b",
          1198 => x"90",
          1199 => x"80",
          1200 => x"52",
          1201 => x"2e",
          1202 => x"52",
          1203 => x"d2",
          1204 => x"87",
          1205 => x"08",
          1206 => x"0a",
          1207 => x"52",
          1208 => x"83",
          1209 => x"71",
          1210 => x"34",
          1211 => x"c0",
          1212 => x"70",
          1213 => x"06",
          1214 => x"70",
          1215 => x"38",
          1216 => x"81",
          1217 => x"80",
          1218 => x"9e",
          1219 => x"a0",
          1220 => x"51",
          1221 => x"80",
          1222 => x"81",
          1223 => x"db",
          1224 => x"0b",
          1225 => x"90",
          1226 => x"80",
          1227 => x"52",
          1228 => x"2e",
          1229 => x"52",
          1230 => x"d6",
          1231 => x"87",
          1232 => x"08",
          1233 => x"80",
          1234 => x"52",
          1235 => x"83",
          1236 => x"71",
          1237 => x"34",
          1238 => x"c0",
          1239 => x"70",
          1240 => x"06",
          1241 => x"70",
          1242 => x"38",
          1243 => x"81",
          1244 => x"80",
          1245 => x"9e",
          1246 => x"81",
          1247 => x"51",
          1248 => x"80",
          1249 => x"81",
          1250 => x"db",
          1251 => x"0b",
          1252 => x"90",
          1253 => x"c0",
          1254 => x"52",
          1255 => x"2e",
          1256 => x"52",
          1257 => x"da",
          1258 => x"87",
          1259 => x"08",
          1260 => x"06",
          1261 => x"70",
          1262 => x"38",
          1263 => x"81",
          1264 => x"87",
          1265 => x"08",
          1266 => x"06",
          1267 => x"51",
          1268 => x"81",
          1269 => x"80",
          1270 => x"9e",
          1271 => x"84",
          1272 => x"52",
          1273 => x"2e",
          1274 => x"52",
          1275 => x"dd",
          1276 => x"9e",
          1277 => x"83",
          1278 => x"84",
          1279 => x"51",
          1280 => x"de",
          1281 => x"87",
          1282 => x"08",
          1283 => x"51",
          1284 => x"80",
          1285 => x"81",
          1286 => x"db",
          1287 => x"c0",
          1288 => x"70",
          1289 => x"51",
          1290 => x"e0",
          1291 => x"0d",
          1292 => x"0d",
          1293 => x"51",
          1294 => x"81",
          1295 => x"54",
          1296 => x"88",
          1297 => x"90",
          1298 => x"3f",
          1299 => x"51",
          1300 => x"81",
          1301 => x"54",
          1302 => x"93",
          1303 => x"ac",
          1304 => x"b0",
          1305 => x"52",
          1306 => x"51",
          1307 => x"81",
          1308 => x"54",
          1309 => x"93",
          1310 => x"a4",
          1311 => x"a8",
          1312 => x"52",
          1313 => x"51",
          1314 => x"81",
          1315 => x"54",
          1316 => x"93",
          1317 => x"8c",
          1318 => x"90",
          1319 => x"52",
          1320 => x"51",
          1321 => x"81",
          1322 => x"54",
          1323 => x"93",
          1324 => x"94",
          1325 => x"98",
          1326 => x"52",
          1327 => x"51",
          1328 => x"81",
          1329 => x"54",
          1330 => x"93",
          1331 => x"9c",
          1332 => x"a0",
          1333 => x"52",
          1334 => x"51",
          1335 => x"81",
          1336 => x"54",
          1337 => x"8d",
          1338 => x"dc",
          1339 => x"c8",
          1340 => x"b0",
          1341 => x"df",
          1342 => x"80",
          1343 => x"81",
          1344 => x"52",
          1345 => x"51",
          1346 => x"81",
          1347 => x"54",
          1348 => x"8d",
          1349 => x"de",
          1350 => x"c9",
          1351 => x"84",
          1352 => x"d1",
          1353 => x"80",
          1354 => x"81",
          1355 => x"84",
          1356 => x"db",
          1357 => x"73",
          1358 => x"38",
          1359 => x"51",
          1360 => x"81",
          1361 => x"54",
          1362 => x"88",
          1363 => x"c8",
          1364 => x"3f",
          1365 => x"33",
          1366 => x"2e",
          1367 => x"c9",
          1368 => x"dc",
          1369 => x"da",
          1370 => x"80",
          1371 => x"81",
          1372 => x"83",
          1373 => x"c9",
          1374 => x"c4",
          1375 => x"b4",
          1376 => x"c9",
          1377 => x"9c",
          1378 => x"b8",
          1379 => x"ca",
          1380 => x"90",
          1381 => x"bc",
          1382 => x"ca",
          1383 => x"84",
          1384 => x"f0",
          1385 => x"3f",
          1386 => x"22",
          1387 => x"f8",
          1388 => x"3f",
          1389 => x"08",
          1390 => x"c0",
          1391 => x"e7",
          1392 => x"de",
          1393 => x"84",
          1394 => x"71",
          1395 => x"81",
          1396 => x"52",
          1397 => x"51",
          1398 => x"81",
          1399 => x"54",
          1400 => x"a8",
          1401 => x"c8",
          1402 => x"84",
          1403 => x"51",
          1404 => x"81",
          1405 => x"bd",
          1406 => x"76",
          1407 => x"54",
          1408 => x"08",
          1409 => x"cc",
          1410 => x"3f",
          1411 => x"33",
          1412 => x"2e",
          1413 => x"db",
          1414 => x"bd",
          1415 => x"75",
          1416 => x"3f",
          1417 => x"08",
          1418 => x"29",
          1419 => x"54",
          1420 => x"c0",
          1421 => x"cb",
          1422 => x"e8",
          1423 => x"9c",
          1424 => x"3f",
          1425 => x"04",
          1426 => x"02",
          1427 => x"ff",
          1428 => x"84",
          1429 => x"71",
          1430 => x"c6",
          1431 => x"71",
          1432 => x"cc",
          1433 => x"39",
          1434 => x"51",
          1435 => x"cc",
          1436 => x"39",
          1437 => x"51",
          1438 => x"cc",
          1439 => x"39",
          1440 => x"51",
          1441 => x"84",
          1442 => x"71",
          1443 => x"04",
          1444 => x"c0",
          1445 => x"04",
          1446 => x"87",
          1447 => x"70",
          1448 => x"80",
          1449 => x"74",
          1450 => x"db",
          1451 => x"0c",
          1452 => x"04",
          1453 => x"87",
          1454 => x"70",
          1455 => x"e4",
          1456 => x"72",
          1457 => x"70",
          1458 => x"08",
          1459 => x"db",
          1460 => x"0c",
          1461 => x"0d",
          1462 => x"e4",
          1463 => x"96",
          1464 => x"fe",
          1465 => x"93",
          1466 => x"72",
          1467 => x"81",
          1468 => x"8d",
          1469 => x"81",
          1470 => x"52",
          1471 => x"90",
          1472 => x"34",
          1473 => x"08",
          1474 => x"de",
          1475 => x"39",
          1476 => x"08",
          1477 => x"2e",
          1478 => x"51",
          1479 => x"3d",
          1480 => x"3d",
          1481 => x"05",
          1482 => x"d0",
          1483 => x"de",
          1484 => x"51",
          1485 => x"72",
          1486 => x"0c",
          1487 => x"04",
          1488 => x"75",
          1489 => x"70",
          1490 => x"53",
          1491 => x"2e",
          1492 => x"81",
          1493 => x"81",
          1494 => x"87",
          1495 => x"85",
          1496 => x"fc",
          1497 => x"81",
          1498 => x"78",
          1499 => x"0c",
          1500 => x"33",
          1501 => x"06",
          1502 => x"80",
          1503 => x"72",
          1504 => x"51",
          1505 => x"fe",
          1506 => x"39",
          1507 => x"d0",
          1508 => x"0d",
          1509 => x"0d",
          1510 => x"59",
          1511 => x"05",
          1512 => x"75",
          1513 => x"f8",
          1514 => x"2e",
          1515 => x"82",
          1516 => x"70",
          1517 => x"05",
          1518 => x"5b",
          1519 => x"2e",
          1520 => x"85",
          1521 => x"8b",
          1522 => x"2e",
          1523 => x"8a",
          1524 => x"78",
          1525 => x"5a",
          1526 => x"aa",
          1527 => x"06",
          1528 => x"84",
          1529 => x"7b",
          1530 => x"5d",
          1531 => x"59",
          1532 => x"d0",
          1533 => x"89",
          1534 => x"7a",
          1535 => x"10",
          1536 => x"d0",
          1537 => x"81",
          1538 => x"57",
          1539 => x"75",
          1540 => x"70",
          1541 => x"07",
          1542 => x"80",
          1543 => x"30",
          1544 => x"80",
          1545 => x"53",
          1546 => x"55",
          1547 => x"2e",
          1548 => x"84",
          1549 => x"81",
          1550 => x"57",
          1551 => x"2e",
          1552 => x"75",
          1553 => x"76",
          1554 => x"e0",
          1555 => x"ff",
          1556 => x"73",
          1557 => x"81",
          1558 => x"80",
          1559 => x"38",
          1560 => x"2e",
          1561 => x"73",
          1562 => x"8b",
          1563 => x"c2",
          1564 => x"38",
          1565 => x"73",
          1566 => x"81",
          1567 => x"8f",
          1568 => x"d5",
          1569 => x"38",
          1570 => x"24",
          1571 => x"80",
          1572 => x"38",
          1573 => x"73",
          1574 => x"80",
          1575 => x"ef",
          1576 => x"19",
          1577 => x"59",
          1578 => x"33",
          1579 => x"75",
          1580 => x"81",
          1581 => x"70",
          1582 => x"55",
          1583 => x"79",
          1584 => x"90",
          1585 => x"16",
          1586 => x"7b",
          1587 => x"a0",
          1588 => x"3f",
          1589 => x"53",
          1590 => x"e9",
          1591 => x"fc",
          1592 => x"81",
          1593 => x"72",
          1594 => x"b0",
          1595 => x"fb",
          1596 => x"39",
          1597 => x"83",
          1598 => x"59",
          1599 => x"82",
          1600 => x"88",
          1601 => x"8a",
          1602 => x"90",
          1603 => x"75",
          1604 => x"3f",
          1605 => x"79",
          1606 => x"81",
          1607 => x"72",
          1608 => x"38",
          1609 => x"59",
          1610 => x"84",
          1611 => x"58",
          1612 => x"80",
          1613 => x"30",
          1614 => x"80",
          1615 => x"55",
          1616 => x"25",
          1617 => x"80",
          1618 => x"74",
          1619 => x"07",
          1620 => x"0b",
          1621 => x"57",
          1622 => x"51",
          1623 => x"81",
          1624 => x"81",
          1625 => x"53",
          1626 => x"e0",
          1627 => x"de",
          1628 => x"89",
          1629 => x"38",
          1630 => x"75",
          1631 => x"84",
          1632 => x"53",
          1633 => x"06",
          1634 => x"53",
          1635 => x"81",
          1636 => x"81",
          1637 => x"70",
          1638 => x"2a",
          1639 => x"76",
          1640 => x"38",
          1641 => x"38",
          1642 => x"70",
          1643 => x"53",
          1644 => x"8e",
          1645 => x"77",
          1646 => x"53",
          1647 => x"81",
          1648 => x"7a",
          1649 => x"55",
          1650 => x"83",
          1651 => x"79",
          1652 => x"81",
          1653 => x"72",
          1654 => x"17",
          1655 => x"27",
          1656 => x"51",
          1657 => x"75",
          1658 => x"72",
          1659 => x"81",
          1660 => x"7a",
          1661 => x"38",
          1662 => x"05",
          1663 => x"ff",
          1664 => x"70",
          1665 => x"57",
          1666 => x"76",
          1667 => x"81",
          1668 => x"72",
          1669 => x"84",
          1670 => x"f9",
          1671 => x"39",
          1672 => x"04",
          1673 => x"86",
          1674 => x"84",
          1675 => x"55",
          1676 => x"fa",
          1677 => x"3d",
          1678 => x"3d",
          1679 => x"de",
          1680 => x"3d",
          1681 => x"75",
          1682 => x"3f",
          1683 => x"08",
          1684 => x"34",
          1685 => x"de",
          1686 => x"3d",
          1687 => x"3d",
          1688 => x"d0",
          1689 => x"de",
          1690 => x"3d",
          1691 => x"77",
          1692 => x"a1",
          1693 => x"de",
          1694 => x"3d",
          1695 => x"3d",
          1696 => x"81",
          1697 => x"70",
          1698 => x"55",
          1699 => x"80",
          1700 => x"38",
          1701 => x"08",
          1702 => x"81",
          1703 => x"81",
          1704 => x"72",
          1705 => x"cb",
          1706 => x"2e",
          1707 => x"88",
          1708 => x"70",
          1709 => x"51",
          1710 => x"2e",
          1711 => x"80",
          1712 => x"ff",
          1713 => x"39",
          1714 => x"c8",
          1715 => x"52",
          1716 => x"c0",
          1717 => x"52",
          1718 => x"81",
          1719 => x"51",
          1720 => x"ff",
          1721 => x"15",
          1722 => x"34",
          1723 => x"f3",
          1724 => x"72",
          1725 => x"0c",
          1726 => x"04",
          1727 => x"81",
          1728 => x"75",
          1729 => x"0c",
          1730 => x"52",
          1731 => x"3f",
          1732 => x"d4",
          1733 => x"0d",
          1734 => x"0d",
          1735 => x"56",
          1736 => x"0c",
          1737 => x"70",
          1738 => x"73",
          1739 => x"81",
          1740 => x"81",
          1741 => x"ed",
          1742 => x"2e",
          1743 => x"8e",
          1744 => x"08",
          1745 => x"76",
          1746 => x"56",
          1747 => x"b0",
          1748 => x"06",
          1749 => x"75",
          1750 => x"76",
          1751 => x"70",
          1752 => x"73",
          1753 => x"8b",
          1754 => x"73",
          1755 => x"85",
          1756 => x"82",
          1757 => x"76",
          1758 => x"70",
          1759 => x"ac",
          1760 => x"a0",
          1761 => x"fa",
          1762 => x"53",
          1763 => x"57",
          1764 => x"98",
          1765 => x"39",
          1766 => x"80",
          1767 => x"26",
          1768 => x"86",
          1769 => x"80",
          1770 => x"57",
          1771 => x"74",
          1772 => x"38",
          1773 => x"27",
          1774 => x"14",
          1775 => x"06",
          1776 => x"14",
          1777 => x"06",
          1778 => x"74",
          1779 => x"f9",
          1780 => x"ff",
          1781 => x"89",
          1782 => x"38",
          1783 => x"c5",
          1784 => x"29",
          1785 => x"81",
          1786 => x"76",
          1787 => x"56",
          1788 => x"ba",
          1789 => x"2e",
          1790 => x"30",
          1791 => x"0c",
          1792 => x"81",
          1793 => x"8a",
          1794 => x"f8",
          1795 => x"7c",
          1796 => x"70",
          1797 => x"75",
          1798 => x"55",
          1799 => x"2e",
          1800 => x"87",
          1801 => x"76",
          1802 => x"73",
          1803 => x"81",
          1804 => x"81",
          1805 => x"77",
          1806 => x"70",
          1807 => x"58",
          1808 => x"09",
          1809 => x"c2",
          1810 => x"81",
          1811 => x"75",
          1812 => x"55",
          1813 => x"e2",
          1814 => x"90",
          1815 => x"f8",
          1816 => x"8f",
          1817 => x"81",
          1818 => x"75",
          1819 => x"55",
          1820 => x"81",
          1821 => x"27",
          1822 => x"d0",
          1823 => x"55",
          1824 => x"73",
          1825 => x"80",
          1826 => x"14",
          1827 => x"72",
          1828 => x"e0",
          1829 => x"80",
          1830 => x"39",
          1831 => x"55",
          1832 => x"80",
          1833 => x"e0",
          1834 => x"38",
          1835 => x"81",
          1836 => x"53",
          1837 => x"81",
          1838 => x"53",
          1839 => x"8e",
          1840 => x"70",
          1841 => x"55",
          1842 => x"27",
          1843 => x"77",
          1844 => x"74",
          1845 => x"76",
          1846 => x"77",
          1847 => x"70",
          1848 => x"55",
          1849 => x"77",
          1850 => x"38",
          1851 => x"74",
          1852 => x"55",
          1853 => x"c0",
          1854 => x"0d",
          1855 => x"0d",
          1856 => x"33",
          1857 => x"70",
          1858 => x"38",
          1859 => x"11",
          1860 => x"81",
          1861 => x"83",
          1862 => x"fc",
          1863 => x"9b",
          1864 => x"84",
          1865 => x"33",
          1866 => x"51",
          1867 => x"80",
          1868 => x"84",
          1869 => x"92",
          1870 => x"51",
          1871 => x"80",
          1872 => x"81",
          1873 => x"72",
          1874 => x"92",
          1875 => x"81",
          1876 => x"0b",
          1877 => x"8c",
          1878 => x"71",
          1879 => x"06",
          1880 => x"80",
          1881 => x"87",
          1882 => x"08",
          1883 => x"38",
          1884 => x"80",
          1885 => x"71",
          1886 => x"c0",
          1887 => x"51",
          1888 => x"87",
          1889 => x"db",
          1890 => x"81",
          1891 => x"33",
          1892 => x"de",
          1893 => x"3d",
          1894 => x"3d",
          1895 => x"64",
          1896 => x"bf",
          1897 => x"40",
          1898 => x"74",
          1899 => x"cd",
          1900 => x"c0",
          1901 => x"7a",
          1902 => x"81",
          1903 => x"72",
          1904 => x"87",
          1905 => x"11",
          1906 => x"8c",
          1907 => x"92",
          1908 => x"5a",
          1909 => x"58",
          1910 => x"c0",
          1911 => x"76",
          1912 => x"76",
          1913 => x"70",
          1914 => x"81",
          1915 => x"54",
          1916 => x"8e",
          1917 => x"52",
          1918 => x"81",
          1919 => x"81",
          1920 => x"74",
          1921 => x"53",
          1922 => x"83",
          1923 => x"78",
          1924 => x"8f",
          1925 => x"2e",
          1926 => x"c0",
          1927 => x"52",
          1928 => x"87",
          1929 => x"08",
          1930 => x"2e",
          1931 => x"84",
          1932 => x"38",
          1933 => x"87",
          1934 => x"15",
          1935 => x"70",
          1936 => x"52",
          1937 => x"ff",
          1938 => x"39",
          1939 => x"81",
          1940 => x"ff",
          1941 => x"57",
          1942 => x"90",
          1943 => x"80",
          1944 => x"71",
          1945 => x"78",
          1946 => x"38",
          1947 => x"80",
          1948 => x"80",
          1949 => x"81",
          1950 => x"72",
          1951 => x"0c",
          1952 => x"04",
          1953 => x"60",
          1954 => x"8c",
          1955 => x"33",
          1956 => x"5b",
          1957 => x"74",
          1958 => x"e1",
          1959 => x"c0",
          1960 => x"79",
          1961 => x"78",
          1962 => x"06",
          1963 => x"77",
          1964 => x"87",
          1965 => x"11",
          1966 => x"8c",
          1967 => x"92",
          1968 => x"59",
          1969 => x"85",
          1970 => x"98",
          1971 => x"7d",
          1972 => x"0c",
          1973 => x"08",
          1974 => x"70",
          1975 => x"53",
          1976 => x"2e",
          1977 => x"70",
          1978 => x"33",
          1979 => x"18",
          1980 => x"2a",
          1981 => x"51",
          1982 => x"2e",
          1983 => x"c0",
          1984 => x"52",
          1985 => x"87",
          1986 => x"08",
          1987 => x"2e",
          1988 => x"84",
          1989 => x"38",
          1990 => x"87",
          1991 => x"15",
          1992 => x"70",
          1993 => x"52",
          1994 => x"ff",
          1995 => x"39",
          1996 => x"81",
          1997 => x"80",
          1998 => x"52",
          1999 => x"90",
          2000 => x"80",
          2001 => x"71",
          2002 => x"7a",
          2003 => x"38",
          2004 => x"80",
          2005 => x"80",
          2006 => x"81",
          2007 => x"72",
          2008 => x"0c",
          2009 => x"04",
          2010 => x"7e",
          2011 => x"b3",
          2012 => x"88",
          2013 => x"33",
          2014 => x"56",
          2015 => x"3f",
          2016 => x"08",
          2017 => x"83",
          2018 => x"fe",
          2019 => x"87",
          2020 => x"0c",
          2021 => x"76",
          2022 => x"38",
          2023 => x"93",
          2024 => x"2b",
          2025 => x"8c",
          2026 => x"71",
          2027 => x"38",
          2028 => x"71",
          2029 => x"c6",
          2030 => x"39",
          2031 => x"81",
          2032 => x"06",
          2033 => x"71",
          2034 => x"38",
          2035 => x"8c",
          2036 => x"e8",
          2037 => x"98",
          2038 => x"71",
          2039 => x"73",
          2040 => x"92",
          2041 => x"72",
          2042 => x"06",
          2043 => x"f7",
          2044 => x"80",
          2045 => x"88",
          2046 => x"0c",
          2047 => x"80",
          2048 => x"56",
          2049 => x"56",
          2050 => x"81",
          2051 => x"8c",
          2052 => x"fe",
          2053 => x"81",
          2054 => x"33",
          2055 => x"07",
          2056 => x"0c",
          2057 => x"3d",
          2058 => x"3d",
          2059 => x"11",
          2060 => x"33",
          2061 => x"71",
          2062 => x"81",
          2063 => x"72",
          2064 => x"75",
          2065 => x"81",
          2066 => x"52",
          2067 => x"54",
          2068 => x"0d",
          2069 => x"0d",
          2070 => x"05",
          2071 => x"52",
          2072 => x"70",
          2073 => x"34",
          2074 => x"51",
          2075 => x"83",
          2076 => x"ff",
          2077 => x"75",
          2078 => x"72",
          2079 => x"54",
          2080 => x"2a",
          2081 => x"70",
          2082 => x"34",
          2083 => x"51",
          2084 => x"81",
          2085 => x"70",
          2086 => x"70",
          2087 => x"3d",
          2088 => x"3d",
          2089 => x"77",
          2090 => x"70",
          2091 => x"38",
          2092 => x"05",
          2093 => x"70",
          2094 => x"34",
          2095 => x"eb",
          2096 => x"0d",
          2097 => x"0d",
          2098 => x"54",
          2099 => x"72",
          2100 => x"54",
          2101 => x"51",
          2102 => x"84",
          2103 => x"fc",
          2104 => x"77",
          2105 => x"53",
          2106 => x"05",
          2107 => x"70",
          2108 => x"33",
          2109 => x"ff",
          2110 => x"52",
          2111 => x"2e",
          2112 => x"80",
          2113 => x"71",
          2114 => x"0c",
          2115 => x"04",
          2116 => x"74",
          2117 => x"89",
          2118 => x"2e",
          2119 => x"11",
          2120 => x"52",
          2121 => x"70",
          2122 => x"c0",
          2123 => x"0d",
          2124 => x"81",
          2125 => x"04",
          2126 => x"de",
          2127 => x"f7",
          2128 => x"56",
          2129 => x"17",
          2130 => x"74",
          2131 => x"d6",
          2132 => x"b0",
          2133 => x"b4",
          2134 => x"81",
          2135 => x"59",
          2136 => x"81",
          2137 => x"7a",
          2138 => x"06",
          2139 => x"de",
          2140 => x"17",
          2141 => x"08",
          2142 => x"08",
          2143 => x"08",
          2144 => x"74",
          2145 => x"38",
          2146 => x"55",
          2147 => x"09",
          2148 => x"38",
          2149 => x"18",
          2150 => x"81",
          2151 => x"f9",
          2152 => x"39",
          2153 => x"81",
          2154 => x"8b",
          2155 => x"fa",
          2156 => x"7a",
          2157 => x"57",
          2158 => x"08",
          2159 => x"75",
          2160 => x"3f",
          2161 => x"08",
          2162 => x"c0",
          2163 => x"81",
          2164 => x"b4",
          2165 => x"16",
          2166 => x"be",
          2167 => x"c0",
          2168 => x"85",
          2169 => x"81",
          2170 => x"17",
          2171 => x"de",
          2172 => x"3d",
          2173 => x"3d",
          2174 => x"52",
          2175 => x"3f",
          2176 => x"08",
          2177 => x"c0",
          2178 => x"38",
          2179 => x"74",
          2180 => x"81",
          2181 => x"38",
          2182 => x"59",
          2183 => x"09",
          2184 => x"e3",
          2185 => x"53",
          2186 => x"08",
          2187 => x"70",
          2188 => x"91",
          2189 => x"d5",
          2190 => x"17",
          2191 => x"3f",
          2192 => x"a4",
          2193 => x"51",
          2194 => x"86",
          2195 => x"f2",
          2196 => x"17",
          2197 => x"3f",
          2198 => x"52",
          2199 => x"51",
          2200 => x"8c",
          2201 => x"84",
          2202 => x"fc",
          2203 => x"17",
          2204 => x"70",
          2205 => x"79",
          2206 => x"52",
          2207 => x"51",
          2208 => x"77",
          2209 => x"80",
          2210 => x"81",
          2211 => x"f9",
          2212 => x"de",
          2213 => x"2e",
          2214 => x"58",
          2215 => x"c0",
          2216 => x"0d",
          2217 => x"0d",
          2218 => x"98",
          2219 => x"05",
          2220 => x"80",
          2221 => x"27",
          2222 => x"14",
          2223 => x"29",
          2224 => x"05",
          2225 => x"81",
          2226 => x"87",
          2227 => x"f9",
          2228 => x"7a",
          2229 => x"54",
          2230 => x"27",
          2231 => x"76",
          2232 => x"27",
          2233 => x"ff",
          2234 => x"58",
          2235 => x"80",
          2236 => x"82",
          2237 => x"72",
          2238 => x"38",
          2239 => x"72",
          2240 => x"8e",
          2241 => x"39",
          2242 => x"17",
          2243 => x"a4",
          2244 => x"53",
          2245 => x"fd",
          2246 => x"de",
          2247 => x"9f",
          2248 => x"ff",
          2249 => x"11",
          2250 => x"70",
          2251 => x"18",
          2252 => x"76",
          2253 => x"53",
          2254 => x"81",
          2255 => x"80",
          2256 => x"83",
          2257 => x"b4",
          2258 => x"88",
          2259 => x"79",
          2260 => x"84",
          2261 => x"58",
          2262 => x"80",
          2263 => x"9f",
          2264 => x"80",
          2265 => x"88",
          2266 => x"08",
          2267 => x"51",
          2268 => x"81",
          2269 => x"80",
          2270 => x"10",
          2271 => x"74",
          2272 => x"51",
          2273 => x"81",
          2274 => x"83",
          2275 => x"58",
          2276 => x"87",
          2277 => x"08",
          2278 => x"51",
          2279 => x"81",
          2280 => x"9b",
          2281 => x"2b",
          2282 => x"74",
          2283 => x"51",
          2284 => x"81",
          2285 => x"f0",
          2286 => x"83",
          2287 => x"77",
          2288 => x"0c",
          2289 => x"04",
          2290 => x"7a",
          2291 => x"58",
          2292 => x"81",
          2293 => x"9e",
          2294 => x"17",
          2295 => x"96",
          2296 => x"53",
          2297 => x"81",
          2298 => x"79",
          2299 => x"72",
          2300 => x"38",
          2301 => x"72",
          2302 => x"b8",
          2303 => x"39",
          2304 => x"17",
          2305 => x"a4",
          2306 => x"53",
          2307 => x"fb",
          2308 => x"de",
          2309 => x"81",
          2310 => x"81",
          2311 => x"83",
          2312 => x"b4",
          2313 => x"78",
          2314 => x"56",
          2315 => x"76",
          2316 => x"38",
          2317 => x"9f",
          2318 => x"33",
          2319 => x"07",
          2320 => x"74",
          2321 => x"83",
          2322 => x"89",
          2323 => x"08",
          2324 => x"51",
          2325 => x"81",
          2326 => x"59",
          2327 => x"08",
          2328 => x"74",
          2329 => x"16",
          2330 => x"84",
          2331 => x"76",
          2332 => x"88",
          2333 => x"81",
          2334 => x"8f",
          2335 => x"53",
          2336 => x"80",
          2337 => x"88",
          2338 => x"08",
          2339 => x"51",
          2340 => x"81",
          2341 => x"59",
          2342 => x"08",
          2343 => x"77",
          2344 => x"06",
          2345 => x"83",
          2346 => x"05",
          2347 => x"f7",
          2348 => x"39",
          2349 => x"a4",
          2350 => x"52",
          2351 => x"ef",
          2352 => x"c0",
          2353 => x"de",
          2354 => x"38",
          2355 => x"06",
          2356 => x"83",
          2357 => x"18",
          2358 => x"54",
          2359 => x"f6",
          2360 => x"de",
          2361 => x"0a",
          2362 => x"52",
          2363 => x"83",
          2364 => x"83",
          2365 => x"81",
          2366 => x"8a",
          2367 => x"f8",
          2368 => x"7c",
          2369 => x"59",
          2370 => x"81",
          2371 => x"38",
          2372 => x"08",
          2373 => x"73",
          2374 => x"38",
          2375 => x"52",
          2376 => x"a4",
          2377 => x"c0",
          2378 => x"de",
          2379 => x"f2",
          2380 => x"82",
          2381 => x"39",
          2382 => x"e6",
          2383 => x"c0",
          2384 => x"de",
          2385 => x"78",
          2386 => x"3f",
          2387 => x"08",
          2388 => x"c0",
          2389 => x"80",
          2390 => x"de",
          2391 => x"2e",
          2392 => x"de",
          2393 => x"2e",
          2394 => x"53",
          2395 => x"51",
          2396 => x"81",
          2397 => x"c5",
          2398 => x"08",
          2399 => x"18",
          2400 => x"57",
          2401 => x"90",
          2402 => x"90",
          2403 => x"16",
          2404 => x"54",
          2405 => x"34",
          2406 => x"78",
          2407 => x"38",
          2408 => x"81",
          2409 => x"8a",
          2410 => x"f6",
          2411 => x"7e",
          2412 => x"5b",
          2413 => x"38",
          2414 => x"58",
          2415 => x"88",
          2416 => x"08",
          2417 => x"38",
          2418 => x"39",
          2419 => x"51",
          2420 => x"81",
          2421 => x"de",
          2422 => x"82",
          2423 => x"de",
          2424 => x"81",
          2425 => x"ff",
          2426 => x"38",
          2427 => x"81",
          2428 => x"26",
          2429 => x"79",
          2430 => x"08",
          2431 => x"73",
          2432 => x"b9",
          2433 => x"2e",
          2434 => x"80",
          2435 => x"1a",
          2436 => x"08",
          2437 => x"38",
          2438 => x"52",
          2439 => x"af",
          2440 => x"81",
          2441 => x"81",
          2442 => x"06",
          2443 => x"de",
          2444 => x"81",
          2445 => x"09",
          2446 => x"72",
          2447 => x"70",
          2448 => x"de",
          2449 => x"51",
          2450 => x"73",
          2451 => x"81",
          2452 => x"80",
          2453 => x"8c",
          2454 => x"81",
          2455 => x"38",
          2456 => x"08",
          2457 => x"73",
          2458 => x"75",
          2459 => x"77",
          2460 => x"56",
          2461 => x"76",
          2462 => x"82",
          2463 => x"26",
          2464 => x"75",
          2465 => x"f8",
          2466 => x"de",
          2467 => x"2e",
          2468 => x"59",
          2469 => x"08",
          2470 => x"81",
          2471 => x"81",
          2472 => x"59",
          2473 => x"08",
          2474 => x"70",
          2475 => x"25",
          2476 => x"51",
          2477 => x"73",
          2478 => x"75",
          2479 => x"81",
          2480 => x"38",
          2481 => x"f5",
          2482 => x"75",
          2483 => x"f9",
          2484 => x"de",
          2485 => x"de",
          2486 => x"70",
          2487 => x"08",
          2488 => x"51",
          2489 => x"80",
          2490 => x"73",
          2491 => x"38",
          2492 => x"52",
          2493 => x"d0",
          2494 => x"c0",
          2495 => x"a5",
          2496 => x"18",
          2497 => x"08",
          2498 => x"18",
          2499 => x"74",
          2500 => x"38",
          2501 => x"18",
          2502 => x"33",
          2503 => x"73",
          2504 => x"97",
          2505 => x"74",
          2506 => x"38",
          2507 => x"55",
          2508 => x"de",
          2509 => x"85",
          2510 => x"75",
          2511 => x"de",
          2512 => x"3d",
          2513 => x"3d",
          2514 => x"52",
          2515 => x"3f",
          2516 => x"08",
          2517 => x"81",
          2518 => x"80",
          2519 => x"52",
          2520 => x"c1",
          2521 => x"c0",
          2522 => x"c0",
          2523 => x"0c",
          2524 => x"53",
          2525 => x"15",
          2526 => x"f2",
          2527 => x"56",
          2528 => x"16",
          2529 => x"22",
          2530 => x"27",
          2531 => x"54",
          2532 => x"76",
          2533 => x"33",
          2534 => x"3f",
          2535 => x"08",
          2536 => x"38",
          2537 => x"76",
          2538 => x"70",
          2539 => x"9f",
          2540 => x"56",
          2541 => x"de",
          2542 => x"3d",
          2543 => x"3d",
          2544 => x"71",
          2545 => x"57",
          2546 => x"0a",
          2547 => x"38",
          2548 => x"53",
          2549 => x"38",
          2550 => x"0c",
          2551 => x"54",
          2552 => x"75",
          2553 => x"73",
          2554 => x"a8",
          2555 => x"73",
          2556 => x"85",
          2557 => x"0b",
          2558 => x"5a",
          2559 => x"27",
          2560 => x"a8",
          2561 => x"18",
          2562 => x"39",
          2563 => x"70",
          2564 => x"58",
          2565 => x"b2",
          2566 => x"76",
          2567 => x"3f",
          2568 => x"08",
          2569 => x"c0",
          2570 => x"bd",
          2571 => x"81",
          2572 => x"27",
          2573 => x"16",
          2574 => x"c0",
          2575 => x"38",
          2576 => x"39",
          2577 => x"55",
          2578 => x"52",
          2579 => x"d5",
          2580 => x"c0",
          2581 => x"0c",
          2582 => x"0c",
          2583 => x"53",
          2584 => x"80",
          2585 => x"85",
          2586 => x"94",
          2587 => x"2a",
          2588 => x"0c",
          2589 => x"06",
          2590 => x"9c",
          2591 => x"58",
          2592 => x"c0",
          2593 => x"0d",
          2594 => x"0d",
          2595 => x"90",
          2596 => x"05",
          2597 => x"f0",
          2598 => x"27",
          2599 => x"0b",
          2600 => x"98",
          2601 => x"84",
          2602 => x"2e",
          2603 => x"76",
          2604 => x"58",
          2605 => x"38",
          2606 => x"15",
          2607 => x"08",
          2608 => x"38",
          2609 => x"88",
          2610 => x"53",
          2611 => x"81",
          2612 => x"c0",
          2613 => x"22",
          2614 => x"89",
          2615 => x"72",
          2616 => x"74",
          2617 => x"f3",
          2618 => x"de",
          2619 => x"82",
          2620 => x"81",
          2621 => x"27",
          2622 => x"81",
          2623 => x"c0",
          2624 => x"80",
          2625 => x"16",
          2626 => x"c0",
          2627 => x"ca",
          2628 => x"38",
          2629 => x"0c",
          2630 => x"dd",
          2631 => x"08",
          2632 => x"f9",
          2633 => x"de",
          2634 => x"87",
          2635 => x"c0",
          2636 => x"80",
          2637 => x"55",
          2638 => x"08",
          2639 => x"38",
          2640 => x"de",
          2641 => x"2e",
          2642 => x"de",
          2643 => x"75",
          2644 => x"3f",
          2645 => x"08",
          2646 => x"94",
          2647 => x"52",
          2648 => x"c1",
          2649 => x"c0",
          2650 => x"0c",
          2651 => x"0c",
          2652 => x"05",
          2653 => x"80",
          2654 => x"de",
          2655 => x"3d",
          2656 => x"3d",
          2657 => x"71",
          2658 => x"57",
          2659 => x"51",
          2660 => x"81",
          2661 => x"54",
          2662 => x"08",
          2663 => x"81",
          2664 => x"56",
          2665 => x"52",
          2666 => x"83",
          2667 => x"c0",
          2668 => x"de",
          2669 => x"d2",
          2670 => x"c0",
          2671 => x"08",
          2672 => x"54",
          2673 => x"e5",
          2674 => x"06",
          2675 => x"58",
          2676 => x"08",
          2677 => x"38",
          2678 => x"75",
          2679 => x"80",
          2680 => x"81",
          2681 => x"7a",
          2682 => x"06",
          2683 => x"39",
          2684 => x"08",
          2685 => x"76",
          2686 => x"3f",
          2687 => x"08",
          2688 => x"c0",
          2689 => x"ff",
          2690 => x"84",
          2691 => x"06",
          2692 => x"54",
          2693 => x"c0",
          2694 => x"0d",
          2695 => x"0d",
          2696 => x"52",
          2697 => x"3f",
          2698 => x"08",
          2699 => x"06",
          2700 => x"51",
          2701 => x"83",
          2702 => x"06",
          2703 => x"14",
          2704 => x"3f",
          2705 => x"08",
          2706 => x"07",
          2707 => x"de",
          2708 => x"3d",
          2709 => x"3d",
          2710 => x"70",
          2711 => x"06",
          2712 => x"53",
          2713 => x"ed",
          2714 => x"33",
          2715 => x"83",
          2716 => x"06",
          2717 => x"90",
          2718 => x"15",
          2719 => x"3f",
          2720 => x"04",
          2721 => x"7b",
          2722 => x"84",
          2723 => x"58",
          2724 => x"80",
          2725 => x"38",
          2726 => x"52",
          2727 => x"8f",
          2728 => x"c0",
          2729 => x"de",
          2730 => x"f5",
          2731 => x"08",
          2732 => x"53",
          2733 => x"84",
          2734 => x"39",
          2735 => x"70",
          2736 => x"81",
          2737 => x"51",
          2738 => x"16",
          2739 => x"c0",
          2740 => x"81",
          2741 => x"38",
          2742 => x"ae",
          2743 => x"81",
          2744 => x"54",
          2745 => x"2e",
          2746 => x"8f",
          2747 => x"81",
          2748 => x"76",
          2749 => x"54",
          2750 => x"09",
          2751 => x"38",
          2752 => x"7a",
          2753 => x"80",
          2754 => x"fa",
          2755 => x"de",
          2756 => x"81",
          2757 => x"89",
          2758 => x"08",
          2759 => x"86",
          2760 => x"98",
          2761 => x"81",
          2762 => x"8b",
          2763 => x"fb",
          2764 => x"70",
          2765 => x"81",
          2766 => x"fc",
          2767 => x"de",
          2768 => x"81",
          2769 => x"b4",
          2770 => x"08",
          2771 => x"ec",
          2772 => x"de",
          2773 => x"81",
          2774 => x"a0",
          2775 => x"81",
          2776 => x"52",
          2777 => x"51",
          2778 => x"8b",
          2779 => x"52",
          2780 => x"51",
          2781 => x"81",
          2782 => x"34",
          2783 => x"c0",
          2784 => x"0d",
          2785 => x"0d",
          2786 => x"98",
          2787 => x"70",
          2788 => x"ec",
          2789 => x"de",
          2790 => x"38",
          2791 => x"53",
          2792 => x"81",
          2793 => x"34",
          2794 => x"04",
          2795 => x"78",
          2796 => x"80",
          2797 => x"34",
          2798 => x"80",
          2799 => x"38",
          2800 => x"18",
          2801 => x"9c",
          2802 => x"70",
          2803 => x"56",
          2804 => x"a0",
          2805 => x"71",
          2806 => x"81",
          2807 => x"81",
          2808 => x"89",
          2809 => x"06",
          2810 => x"73",
          2811 => x"55",
          2812 => x"55",
          2813 => x"81",
          2814 => x"81",
          2815 => x"74",
          2816 => x"75",
          2817 => x"52",
          2818 => x"13",
          2819 => x"08",
          2820 => x"33",
          2821 => x"9c",
          2822 => x"11",
          2823 => x"8a",
          2824 => x"c0",
          2825 => x"96",
          2826 => x"e7",
          2827 => x"c0",
          2828 => x"23",
          2829 => x"e7",
          2830 => x"de",
          2831 => x"17",
          2832 => x"0d",
          2833 => x"0d",
          2834 => x"5e",
          2835 => x"70",
          2836 => x"55",
          2837 => x"83",
          2838 => x"73",
          2839 => x"91",
          2840 => x"2e",
          2841 => x"1d",
          2842 => x"0c",
          2843 => x"15",
          2844 => x"70",
          2845 => x"56",
          2846 => x"09",
          2847 => x"38",
          2848 => x"80",
          2849 => x"30",
          2850 => x"78",
          2851 => x"54",
          2852 => x"73",
          2853 => x"60",
          2854 => x"54",
          2855 => x"96",
          2856 => x"0b",
          2857 => x"80",
          2858 => x"f6",
          2859 => x"de",
          2860 => x"85",
          2861 => x"3d",
          2862 => x"5c",
          2863 => x"53",
          2864 => x"51",
          2865 => x"80",
          2866 => x"88",
          2867 => x"5c",
          2868 => x"09",
          2869 => x"d4",
          2870 => x"70",
          2871 => x"71",
          2872 => x"30",
          2873 => x"73",
          2874 => x"51",
          2875 => x"57",
          2876 => x"38",
          2877 => x"75",
          2878 => x"17",
          2879 => x"75",
          2880 => x"30",
          2881 => x"51",
          2882 => x"80",
          2883 => x"38",
          2884 => x"87",
          2885 => x"26",
          2886 => x"77",
          2887 => x"a4",
          2888 => x"27",
          2889 => x"a0",
          2890 => x"39",
          2891 => x"33",
          2892 => x"57",
          2893 => x"27",
          2894 => x"75",
          2895 => x"30",
          2896 => x"32",
          2897 => x"80",
          2898 => x"25",
          2899 => x"56",
          2900 => x"80",
          2901 => x"84",
          2902 => x"58",
          2903 => x"70",
          2904 => x"55",
          2905 => x"09",
          2906 => x"38",
          2907 => x"80",
          2908 => x"30",
          2909 => x"77",
          2910 => x"54",
          2911 => x"81",
          2912 => x"ae",
          2913 => x"06",
          2914 => x"54",
          2915 => x"74",
          2916 => x"80",
          2917 => x"7b",
          2918 => x"30",
          2919 => x"70",
          2920 => x"25",
          2921 => x"07",
          2922 => x"51",
          2923 => x"a7",
          2924 => x"8b",
          2925 => x"39",
          2926 => x"54",
          2927 => x"8c",
          2928 => x"ff",
          2929 => x"b4",
          2930 => x"54",
          2931 => x"e1",
          2932 => x"c0",
          2933 => x"b2",
          2934 => x"70",
          2935 => x"71",
          2936 => x"54",
          2937 => x"81",
          2938 => x"80",
          2939 => x"38",
          2940 => x"76",
          2941 => x"df",
          2942 => x"54",
          2943 => x"81",
          2944 => x"55",
          2945 => x"34",
          2946 => x"52",
          2947 => x"51",
          2948 => x"81",
          2949 => x"bf",
          2950 => x"16",
          2951 => x"26",
          2952 => x"16",
          2953 => x"06",
          2954 => x"17",
          2955 => x"34",
          2956 => x"fd",
          2957 => x"19",
          2958 => x"80",
          2959 => x"79",
          2960 => x"81",
          2961 => x"81",
          2962 => x"85",
          2963 => x"54",
          2964 => x"8f",
          2965 => x"86",
          2966 => x"39",
          2967 => x"f3",
          2968 => x"73",
          2969 => x"80",
          2970 => x"52",
          2971 => x"ce",
          2972 => x"c0",
          2973 => x"de",
          2974 => x"d7",
          2975 => x"08",
          2976 => x"e6",
          2977 => x"de",
          2978 => x"81",
          2979 => x"80",
          2980 => x"1b",
          2981 => x"55",
          2982 => x"2e",
          2983 => x"8b",
          2984 => x"06",
          2985 => x"1c",
          2986 => x"33",
          2987 => x"70",
          2988 => x"55",
          2989 => x"38",
          2990 => x"52",
          2991 => x"9f",
          2992 => x"c0",
          2993 => x"8b",
          2994 => x"7a",
          2995 => x"3f",
          2996 => x"75",
          2997 => x"57",
          2998 => x"2e",
          2999 => x"84",
          3000 => x"06",
          3001 => x"75",
          3002 => x"81",
          3003 => x"2a",
          3004 => x"73",
          3005 => x"38",
          3006 => x"54",
          3007 => x"fb",
          3008 => x"80",
          3009 => x"34",
          3010 => x"c1",
          3011 => x"06",
          3012 => x"38",
          3013 => x"39",
          3014 => x"70",
          3015 => x"54",
          3016 => x"86",
          3017 => x"84",
          3018 => x"06",
          3019 => x"73",
          3020 => x"38",
          3021 => x"83",
          3022 => x"b4",
          3023 => x"51",
          3024 => x"81",
          3025 => x"88",
          3026 => x"ea",
          3027 => x"de",
          3028 => x"3d",
          3029 => x"3d",
          3030 => x"ff",
          3031 => x"71",
          3032 => x"5c",
          3033 => x"80",
          3034 => x"38",
          3035 => x"05",
          3036 => x"a0",
          3037 => x"71",
          3038 => x"38",
          3039 => x"71",
          3040 => x"81",
          3041 => x"38",
          3042 => x"11",
          3043 => x"06",
          3044 => x"70",
          3045 => x"38",
          3046 => x"81",
          3047 => x"05",
          3048 => x"76",
          3049 => x"38",
          3050 => x"cd",
          3051 => x"77",
          3052 => x"57",
          3053 => x"05",
          3054 => x"70",
          3055 => x"33",
          3056 => x"53",
          3057 => x"99",
          3058 => x"e0",
          3059 => x"ff",
          3060 => x"ff",
          3061 => x"70",
          3062 => x"38",
          3063 => x"81",
          3064 => x"51",
          3065 => x"9f",
          3066 => x"72",
          3067 => x"81",
          3068 => x"70",
          3069 => x"72",
          3070 => x"32",
          3071 => x"72",
          3072 => x"73",
          3073 => x"53",
          3074 => x"70",
          3075 => x"38",
          3076 => x"19",
          3077 => x"75",
          3078 => x"38",
          3079 => x"83",
          3080 => x"74",
          3081 => x"59",
          3082 => x"39",
          3083 => x"33",
          3084 => x"de",
          3085 => x"3d",
          3086 => x"3d",
          3087 => x"80",
          3088 => x"34",
          3089 => x"17",
          3090 => x"75",
          3091 => x"3f",
          3092 => x"de",
          3093 => x"80",
          3094 => x"16",
          3095 => x"3f",
          3096 => x"08",
          3097 => x"06",
          3098 => x"73",
          3099 => x"2e",
          3100 => x"80",
          3101 => x"0b",
          3102 => x"56",
          3103 => x"e9",
          3104 => x"06",
          3105 => x"57",
          3106 => x"32",
          3107 => x"80",
          3108 => x"51",
          3109 => x"8a",
          3110 => x"e8",
          3111 => x"06",
          3112 => x"53",
          3113 => x"52",
          3114 => x"51",
          3115 => x"81",
          3116 => x"55",
          3117 => x"08",
          3118 => x"38",
          3119 => x"cc",
          3120 => x"86",
          3121 => x"97",
          3122 => x"c0",
          3123 => x"de",
          3124 => x"2e",
          3125 => x"55",
          3126 => x"c0",
          3127 => x"0d",
          3128 => x"0d",
          3129 => x"05",
          3130 => x"33",
          3131 => x"75",
          3132 => x"fc",
          3133 => x"de",
          3134 => x"8b",
          3135 => x"81",
          3136 => x"24",
          3137 => x"81",
          3138 => x"84",
          3139 => x"dc",
          3140 => x"55",
          3141 => x"73",
          3142 => x"e6",
          3143 => x"0c",
          3144 => x"06",
          3145 => x"57",
          3146 => x"ae",
          3147 => x"33",
          3148 => x"3f",
          3149 => x"08",
          3150 => x"70",
          3151 => x"55",
          3152 => x"76",
          3153 => x"b8",
          3154 => x"2a",
          3155 => x"51",
          3156 => x"72",
          3157 => x"86",
          3158 => x"74",
          3159 => x"15",
          3160 => x"81",
          3161 => x"d7",
          3162 => x"de",
          3163 => x"ff",
          3164 => x"06",
          3165 => x"56",
          3166 => x"38",
          3167 => x"8f",
          3168 => x"2a",
          3169 => x"51",
          3170 => x"72",
          3171 => x"80",
          3172 => x"52",
          3173 => x"3f",
          3174 => x"08",
          3175 => x"57",
          3176 => x"09",
          3177 => x"e2",
          3178 => x"74",
          3179 => x"56",
          3180 => x"33",
          3181 => x"72",
          3182 => x"38",
          3183 => x"51",
          3184 => x"81",
          3185 => x"57",
          3186 => x"84",
          3187 => x"ff",
          3188 => x"56",
          3189 => x"25",
          3190 => x"0b",
          3191 => x"56",
          3192 => x"05",
          3193 => x"83",
          3194 => x"2e",
          3195 => x"52",
          3196 => x"c6",
          3197 => x"c0",
          3198 => x"06",
          3199 => x"27",
          3200 => x"16",
          3201 => x"27",
          3202 => x"56",
          3203 => x"84",
          3204 => x"56",
          3205 => x"84",
          3206 => x"14",
          3207 => x"3f",
          3208 => x"08",
          3209 => x"06",
          3210 => x"80",
          3211 => x"06",
          3212 => x"80",
          3213 => x"db",
          3214 => x"de",
          3215 => x"ff",
          3216 => x"77",
          3217 => x"d8",
          3218 => x"de",
          3219 => x"c0",
          3220 => x"9c",
          3221 => x"c4",
          3222 => x"15",
          3223 => x"14",
          3224 => x"70",
          3225 => x"51",
          3226 => x"56",
          3227 => x"84",
          3228 => x"81",
          3229 => x"71",
          3230 => x"16",
          3231 => x"53",
          3232 => x"23",
          3233 => x"8b",
          3234 => x"73",
          3235 => x"80",
          3236 => x"8d",
          3237 => x"39",
          3238 => x"51",
          3239 => x"81",
          3240 => x"53",
          3241 => x"08",
          3242 => x"72",
          3243 => x"8d",
          3244 => x"ce",
          3245 => x"14",
          3246 => x"3f",
          3247 => x"08",
          3248 => x"06",
          3249 => x"38",
          3250 => x"51",
          3251 => x"81",
          3252 => x"55",
          3253 => x"51",
          3254 => x"81",
          3255 => x"83",
          3256 => x"53",
          3257 => x"80",
          3258 => x"38",
          3259 => x"78",
          3260 => x"2a",
          3261 => x"78",
          3262 => x"86",
          3263 => x"22",
          3264 => x"31",
          3265 => x"f0",
          3266 => x"c0",
          3267 => x"de",
          3268 => x"2e",
          3269 => x"81",
          3270 => x"80",
          3271 => x"f5",
          3272 => x"83",
          3273 => x"ff",
          3274 => x"38",
          3275 => x"9f",
          3276 => x"38",
          3277 => x"39",
          3278 => x"80",
          3279 => x"38",
          3280 => x"98",
          3281 => x"a0",
          3282 => x"1c",
          3283 => x"0c",
          3284 => x"17",
          3285 => x"76",
          3286 => x"81",
          3287 => x"80",
          3288 => x"d9",
          3289 => x"de",
          3290 => x"ff",
          3291 => x"8d",
          3292 => x"8e",
          3293 => x"8a",
          3294 => x"14",
          3295 => x"3f",
          3296 => x"08",
          3297 => x"74",
          3298 => x"a2",
          3299 => x"79",
          3300 => x"ee",
          3301 => x"a8",
          3302 => x"15",
          3303 => x"2e",
          3304 => x"10",
          3305 => x"2a",
          3306 => x"05",
          3307 => x"ff",
          3308 => x"53",
          3309 => x"9c",
          3310 => x"81",
          3311 => x"0b",
          3312 => x"ff",
          3313 => x"0c",
          3314 => x"84",
          3315 => x"83",
          3316 => x"06",
          3317 => x"80",
          3318 => x"d8",
          3319 => x"de",
          3320 => x"ff",
          3321 => x"72",
          3322 => x"81",
          3323 => x"38",
          3324 => x"73",
          3325 => x"3f",
          3326 => x"08",
          3327 => x"81",
          3328 => x"84",
          3329 => x"b2",
          3330 => x"87",
          3331 => x"c0",
          3332 => x"ff",
          3333 => x"82",
          3334 => x"09",
          3335 => x"c8",
          3336 => x"51",
          3337 => x"81",
          3338 => x"84",
          3339 => x"d2",
          3340 => x"06",
          3341 => x"98",
          3342 => x"ee",
          3343 => x"c0",
          3344 => x"85",
          3345 => x"09",
          3346 => x"38",
          3347 => x"51",
          3348 => x"81",
          3349 => x"90",
          3350 => x"a0",
          3351 => x"ca",
          3352 => x"c0",
          3353 => x"0c",
          3354 => x"81",
          3355 => x"81",
          3356 => x"81",
          3357 => x"72",
          3358 => x"80",
          3359 => x"0c",
          3360 => x"81",
          3361 => x"90",
          3362 => x"fb",
          3363 => x"54",
          3364 => x"80",
          3365 => x"73",
          3366 => x"80",
          3367 => x"72",
          3368 => x"80",
          3369 => x"86",
          3370 => x"15",
          3371 => x"71",
          3372 => x"81",
          3373 => x"81",
          3374 => x"d0",
          3375 => x"de",
          3376 => x"06",
          3377 => x"38",
          3378 => x"54",
          3379 => x"80",
          3380 => x"71",
          3381 => x"81",
          3382 => x"87",
          3383 => x"fa",
          3384 => x"ab",
          3385 => x"58",
          3386 => x"05",
          3387 => x"e6",
          3388 => x"80",
          3389 => x"c0",
          3390 => x"38",
          3391 => x"08",
          3392 => x"de",
          3393 => x"08",
          3394 => x"80",
          3395 => x"80",
          3396 => x"54",
          3397 => x"84",
          3398 => x"34",
          3399 => x"75",
          3400 => x"2e",
          3401 => x"53",
          3402 => x"53",
          3403 => x"f7",
          3404 => x"de",
          3405 => x"73",
          3406 => x"0c",
          3407 => x"04",
          3408 => x"67",
          3409 => x"80",
          3410 => x"59",
          3411 => x"78",
          3412 => x"c8",
          3413 => x"06",
          3414 => x"3d",
          3415 => x"99",
          3416 => x"52",
          3417 => x"3f",
          3418 => x"08",
          3419 => x"c0",
          3420 => x"38",
          3421 => x"52",
          3422 => x"52",
          3423 => x"3f",
          3424 => x"08",
          3425 => x"c0",
          3426 => x"02",
          3427 => x"33",
          3428 => x"55",
          3429 => x"25",
          3430 => x"55",
          3431 => x"54",
          3432 => x"81",
          3433 => x"80",
          3434 => x"74",
          3435 => x"81",
          3436 => x"75",
          3437 => x"3f",
          3438 => x"08",
          3439 => x"02",
          3440 => x"91",
          3441 => x"81",
          3442 => x"82",
          3443 => x"06",
          3444 => x"80",
          3445 => x"88",
          3446 => x"39",
          3447 => x"58",
          3448 => x"38",
          3449 => x"70",
          3450 => x"54",
          3451 => x"81",
          3452 => x"52",
          3453 => x"a5",
          3454 => x"c0",
          3455 => x"88",
          3456 => x"62",
          3457 => x"d4",
          3458 => x"54",
          3459 => x"15",
          3460 => x"62",
          3461 => x"e8",
          3462 => x"52",
          3463 => x"51",
          3464 => x"7a",
          3465 => x"83",
          3466 => x"80",
          3467 => x"38",
          3468 => x"08",
          3469 => x"53",
          3470 => x"3d",
          3471 => x"dd",
          3472 => x"de",
          3473 => x"81",
          3474 => x"82",
          3475 => x"39",
          3476 => x"38",
          3477 => x"33",
          3478 => x"70",
          3479 => x"55",
          3480 => x"2e",
          3481 => x"55",
          3482 => x"77",
          3483 => x"81",
          3484 => x"73",
          3485 => x"38",
          3486 => x"54",
          3487 => x"a0",
          3488 => x"82",
          3489 => x"52",
          3490 => x"a3",
          3491 => x"c0",
          3492 => x"18",
          3493 => x"55",
          3494 => x"c0",
          3495 => x"38",
          3496 => x"70",
          3497 => x"54",
          3498 => x"86",
          3499 => x"c0",
          3500 => x"b0",
          3501 => x"1b",
          3502 => x"1b",
          3503 => x"70",
          3504 => x"d9",
          3505 => x"c0",
          3506 => x"c0",
          3507 => x"0c",
          3508 => x"52",
          3509 => x"3f",
          3510 => x"08",
          3511 => x"08",
          3512 => x"77",
          3513 => x"86",
          3514 => x"1a",
          3515 => x"1a",
          3516 => x"91",
          3517 => x"0b",
          3518 => x"80",
          3519 => x"0c",
          3520 => x"70",
          3521 => x"54",
          3522 => x"81",
          3523 => x"de",
          3524 => x"2e",
          3525 => x"81",
          3526 => x"94",
          3527 => x"17",
          3528 => x"2b",
          3529 => x"57",
          3530 => x"52",
          3531 => x"9f",
          3532 => x"c0",
          3533 => x"de",
          3534 => x"26",
          3535 => x"55",
          3536 => x"08",
          3537 => x"81",
          3538 => x"79",
          3539 => x"31",
          3540 => x"70",
          3541 => x"25",
          3542 => x"76",
          3543 => x"81",
          3544 => x"55",
          3545 => x"38",
          3546 => x"0c",
          3547 => x"75",
          3548 => x"54",
          3549 => x"a2",
          3550 => x"7a",
          3551 => x"3f",
          3552 => x"08",
          3553 => x"55",
          3554 => x"89",
          3555 => x"c0",
          3556 => x"1a",
          3557 => x"80",
          3558 => x"54",
          3559 => x"c0",
          3560 => x"0d",
          3561 => x"0d",
          3562 => x"64",
          3563 => x"59",
          3564 => x"90",
          3565 => x"52",
          3566 => x"cf",
          3567 => x"c0",
          3568 => x"de",
          3569 => x"38",
          3570 => x"55",
          3571 => x"86",
          3572 => x"82",
          3573 => x"19",
          3574 => x"55",
          3575 => x"80",
          3576 => x"38",
          3577 => x"0b",
          3578 => x"82",
          3579 => x"39",
          3580 => x"1a",
          3581 => x"82",
          3582 => x"19",
          3583 => x"08",
          3584 => x"7c",
          3585 => x"74",
          3586 => x"2e",
          3587 => x"94",
          3588 => x"83",
          3589 => x"56",
          3590 => x"38",
          3591 => x"22",
          3592 => x"89",
          3593 => x"55",
          3594 => x"75",
          3595 => x"19",
          3596 => x"39",
          3597 => x"52",
          3598 => x"93",
          3599 => x"c0",
          3600 => x"75",
          3601 => x"38",
          3602 => x"ff",
          3603 => x"98",
          3604 => x"19",
          3605 => x"51",
          3606 => x"81",
          3607 => x"80",
          3608 => x"38",
          3609 => x"08",
          3610 => x"2a",
          3611 => x"80",
          3612 => x"38",
          3613 => x"8a",
          3614 => x"5c",
          3615 => x"27",
          3616 => x"7a",
          3617 => x"54",
          3618 => x"52",
          3619 => x"51",
          3620 => x"81",
          3621 => x"fe",
          3622 => x"83",
          3623 => x"56",
          3624 => x"9f",
          3625 => x"08",
          3626 => x"74",
          3627 => x"38",
          3628 => x"b4",
          3629 => x"16",
          3630 => x"89",
          3631 => x"51",
          3632 => x"77",
          3633 => x"b9",
          3634 => x"1a",
          3635 => x"08",
          3636 => x"84",
          3637 => x"57",
          3638 => x"27",
          3639 => x"56",
          3640 => x"52",
          3641 => x"c7",
          3642 => x"c0",
          3643 => x"38",
          3644 => x"19",
          3645 => x"06",
          3646 => x"52",
          3647 => x"a2",
          3648 => x"31",
          3649 => x"7f",
          3650 => x"94",
          3651 => x"94",
          3652 => x"5c",
          3653 => x"80",
          3654 => x"de",
          3655 => x"3d",
          3656 => x"3d",
          3657 => x"65",
          3658 => x"5d",
          3659 => x"0c",
          3660 => x"05",
          3661 => x"f6",
          3662 => x"de",
          3663 => x"81",
          3664 => x"8a",
          3665 => x"33",
          3666 => x"2e",
          3667 => x"56",
          3668 => x"90",
          3669 => x"81",
          3670 => x"06",
          3671 => x"87",
          3672 => x"2e",
          3673 => x"95",
          3674 => x"91",
          3675 => x"56",
          3676 => x"81",
          3677 => x"34",
          3678 => x"8e",
          3679 => x"08",
          3680 => x"56",
          3681 => x"84",
          3682 => x"5c",
          3683 => x"82",
          3684 => x"18",
          3685 => x"ff",
          3686 => x"74",
          3687 => x"7e",
          3688 => x"ff",
          3689 => x"2a",
          3690 => x"7a",
          3691 => x"8c",
          3692 => x"08",
          3693 => x"38",
          3694 => x"39",
          3695 => x"52",
          3696 => x"e7",
          3697 => x"c0",
          3698 => x"de",
          3699 => x"2e",
          3700 => x"74",
          3701 => x"91",
          3702 => x"2e",
          3703 => x"74",
          3704 => x"88",
          3705 => x"38",
          3706 => x"0c",
          3707 => x"15",
          3708 => x"08",
          3709 => x"06",
          3710 => x"51",
          3711 => x"81",
          3712 => x"fe",
          3713 => x"18",
          3714 => x"51",
          3715 => x"81",
          3716 => x"80",
          3717 => x"38",
          3718 => x"08",
          3719 => x"2a",
          3720 => x"80",
          3721 => x"38",
          3722 => x"8a",
          3723 => x"5b",
          3724 => x"27",
          3725 => x"7b",
          3726 => x"54",
          3727 => x"52",
          3728 => x"51",
          3729 => x"81",
          3730 => x"fe",
          3731 => x"b0",
          3732 => x"31",
          3733 => x"79",
          3734 => x"84",
          3735 => x"16",
          3736 => x"89",
          3737 => x"52",
          3738 => x"cc",
          3739 => x"55",
          3740 => x"16",
          3741 => x"2b",
          3742 => x"39",
          3743 => x"94",
          3744 => x"93",
          3745 => x"cd",
          3746 => x"de",
          3747 => x"e3",
          3748 => x"b0",
          3749 => x"76",
          3750 => x"94",
          3751 => x"ff",
          3752 => x"71",
          3753 => x"7b",
          3754 => x"38",
          3755 => x"18",
          3756 => x"51",
          3757 => x"81",
          3758 => x"fd",
          3759 => x"53",
          3760 => x"18",
          3761 => x"06",
          3762 => x"51",
          3763 => x"7e",
          3764 => x"83",
          3765 => x"76",
          3766 => x"17",
          3767 => x"1e",
          3768 => x"18",
          3769 => x"0c",
          3770 => x"58",
          3771 => x"74",
          3772 => x"38",
          3773 => x"8c",
          3774 => x"90",
          3775 => x"33",
          3776 => x"55",
          3777 => x"34",
          3778 => x"81",
          3779 => x"90",
          3780 => x"f8",
          3781 => x"8b",
          3782 => x"53",
          3783 => x"f2",
          3784 => x"de",
          3785 => x"81",
          3786 => x"80",
          3787 => x"16",
          3788 => x"2a",
          3789 => x"51",
          3790 => x"80",
          3791 => x"38",
          3792 => x"52",
          3793 => x"e7",
          3794 => x"c0",
          3795 => x"de",
          3796 => x"d4",
          3797 => x"08",
          3798 => x"a0",
          3799 => x"73",
          3800 => x"88",
          3801 => x"74",
          3802 => x"51",
          3803 => x"8c",
          3804 => x"9c",
          3805 => x"fb",
          3806 => x"b2",
          3807 => x"15",
          3808 => x"3f",
          3809 => x"15",
          3810 => x"3f",
          3811 => x"0b",
          3812 => x"78",
          3813 => x"3f",
          3814 => x"08",
          3815 => x"81",
          3816 => x"57",
          3817 => x"34",
          3818 => x"c0",
          3819 => x"0d",
          3820 => x"0d",
          3821 => x"54",
          3822 => x"81",
          3823 => x"53",
          3824 => x"08",
          3825 => x"3d",
          3826 => x"73",
          3827 => x"3f",
          3828 => x"08",
          3829 => x"c0",
          3830 => x"81",
          3831 => x"74",
          3832 => x"de",
          3833 => x"3d",
          3834 => x"3d",
          3835 => x"51",
          3836 => x"8b",
          3837 => x"81",
          3838 => x"24",
          3839 => x"de",
          3840 => x"de",
          3841 => x"52",
          3842 => x"c0",
          3843 => x"0d",
          3844 => x"0d",
          3845 => x"3d",
          3846 => x"94",
          3847 => x"c1",
          3848 => x"c0",
          3849 => x"de",
          3850 => x"e0",
          3851 => x"63",
          3852 => x"d4",
          3853 => x"8d",
          3854 => x"c0",
          3855 => x"de",
          3856 => x"38",
          3857 => x"05",
          3858 => x"2b",
          3859 => x"80",
          3860 => x"76",
          3861 => x"0c",
          3862 => x"02",
          3863 => x"70",
          3864 => x"81",
          3865 => x"56",
          3866 => x"9e",
          3867 => x"53",
          3868 => x"db",
          3869 => x"de",
          3870 => x"15",
          3871 => x"81",
          3872 => x"84",
          3873 => x"06",
          3874 => x"55",
          3875 => x"c0",
          3876 => x"0d",
          3877 => x"0d",
          3878 => x"5b",
          3879 => x"80",
          3880 => x"ff",
          3881 => x"9f",
          3882 => x"b5",
          3883 => x"c0",
          3884 => x"de",
          3885 => x"fc",
          3886 => x"7a",
          3887 => x"08",
          3888 => x"64",
          3889 => x"2e",
          3890 => x"a0",
          3891 => x"70",
          3892 => x"ea",
          3893 => x"c0",
          3894 => x"de",
          3895 => x"d4",
          3896 => x"7b",
          3897 => x"3f",
          3898 => x"08",
          3899 => x"c0",
          3900 => x"38",
          3901 => x"51",
          3902 => x"81",
          3903 => x"45",
          3904 => x"51",
          3905 => x"81",
          3906 => x"57",
          3907 => x"08",
          3908 => x"80",
          3909 => x"da",
          3910 => x"de",
          3911 => x"81",
          3912 => x"a4",
          3913 => x"7b",
          3914 => x"3f",
          3915 => x"c0",
          3916 => x"38",
          3917 => x"51",
          3918 => x"81",
          3919 => x"57",
          3920 => x"08",
          3921 => x"38",
          3922 => x"09",
          3923 => x"38",
          3924 => x"e0",
          3925 => x"dc",
          3926 => x"ff",
          3927 => x"74",
          3928 => x"3f",
          3929 => x"78",
          3930 => x"33",
          3931 => x"56",
          3932 => x"91",
          3933 => x"05",
          3934 => x"81",
          3935 => x"56",
          3936 => x"f5",
          3937 => x"54",
          3938 => x"81",
          3939 => x"80",
          3940 => x"78",
          3941 => x"55",
          3942 => x"11",
          3943 => x"18",
          3944 => x"58",
          3945 => x"34",
          3946 => x"ff",
          3947 => x"55",
          3948 => x"34",
          3949 => x"77",
          3950 => x"81",
          3951 => x"ff",
          3952 => x"55",
          3953 => x"34",
          3954 => x"de",
          3955 => x"84",
          3956 => x"a4",
          3957 => x"70",
          3958 => x"56",
          3959 => x"76",
          3960 => x"81",
          3961 => x"70",
          3962 => x"56",
          3963 => x"82",
          3964 => x"78",
          3965 => x"80",
          3966 => x"27",
          3967 => x"19",
          3968 => x"7a",
          3969 => x"5c",
          3970 => x"55",
          3971 => x"7a",
          3972 => x"5c",
          3973 => x"2e",
          3974 => x"85",
          3975 => x"94",
          3976 => x"81",
          3977 => x"73",
          3978 => x"81",
          3979 => x"7a",
          3980 => x"38",
          3981 => x"76",
          3982 => x"0c",
          3983 => x"04",
          3984 => x"7b",
          3985 => x"fc",
          3986 => x"53",
          3987 => x"bb",
          3988 => x"c0",
          3989 => x"de",
          3990 => x"fa",
          3991 => x"33",
          3992 => x"f2",
          3993 => x"08",
          3994 => x"27",
          3995 => x"15",
          3996 => x"2a",
          3997 => x"51",
          3998 => x"83",
          3999 => x"94",
          4000 => x"80",
          4001 => x"0c",
          4002 => x"2e",
          4003 => x"79",
          4004 => x"70",
          4005 => x"51",
          4006 => x"2e",
          4007 => x"52",
          4008 => x"ff",
          4009 => x"81",
          4010 => x"ff",
          4011 => x"70",
          4012 => x"ff",
          4013 => x"81",
          4014 => x"73",
          4015 => x"76",
          4016 => x"06",
          4017 => x"0c",
          4018 => x"98",
          4019 => x"58",
          4020 => x"39",
          4021 => x"54",
          4022 => x"73",
          4023 => x"cd",
          4024 => x"de",
          4025 => x"81",
          4026 => x"81",
          4027 => x"38",
          4028 => x"08",
          4029 => x"9b",
          4030 => x"c0",
          4031 => x"0c",
          4032 => x"0c",
          4033 => x"81",
          4034 => x"76",
          4035 => x"38",
          4036 => x"94",
          4037 => x"94",
          4038 => x"16",
          4039 => x"2a",
          4040 => x"51",
          4041 => x"72",
          4042 => x"38",
          4043 => x"51",
          4044 => x"81",
          4045 => x"54",
          4046 => x"08",
          4047 => x"de",
          4048 => x"a7",
          4049 => x"74",
          4050 => x"3f",
          4051 => x"08",
          4052 => x"2e",
          4053 => x"74",
          4054 => x"79",
          4055 => x"14",
          4056 => x"38",
          4057 => x"0c",
          4058 => x"94",
          4059 => x"94",
          4060 => x"83",
          4061 => x"72",
          4062 => x"38",
          4063 => x"51",
          4064 => x"81",
          4065 => x"94",
          4066 => x"91",
          4067 => x"53",
          4068 => x"81",
          4069 => x"34",
          4070 => x"39",
          4071 => x"81",
          4072 => x"05",
          4073 => x"08",
          4074 => x"08",
          4075 => x"38",
          4076 => x"0c",
          4077 => x"80",
          4078 => x"72",
          4079 => x"73",
          4080 => x"53",
          4081 => x"8c",
          4082 => x"16",
          4083 => x"38",
          4084 => x"0c",
          4085 => x"81",
          4086 => x"8b",
          4087 => x"f9",
          4088 => x"56",
          4089 => x"80",
          4090 => x"38",
          4091 => x"3d",
          4092 => x"8a",
          4093 => x"51",
          4094 => x"81",
          4095 => x"55",
          4096 => x"08",
          4097 => x"77",
          4098 => x"52",
          4099 => x"b5",
          4100 => x"c0",
          4101 => x"de",
          4102 => x"c3",
          4103 => x"33",
          4104 => x"55",
          4105 => x"24",
          4106 => x"16",
          4107 => x"2a",
          4108 => x"51",
          4109 => x"80",
          4110 => x"9c",
          4111 => x"77",
          4112 => x"3f",
          4113 => x"08",
          4114 => x"77",
          4115 => x"22",
          4116 => x"74",
          4117 => x"ce",
          4118 => x"de",
          4119 => x"74",
          4120 => x"81",
          4121 => x"85",
          4122 => x"74",
          4123 => x"38",
          4124 => x"74",
          4125 => x"de",
          4126 => x"3d",
          4127 => x"3d",
          4128 => x"3d",
          4129 => x"70",
          4130 => x"ff",
          4131 => x"c0",
          4132 => x"81",
          4133 => x"73",
          4134 => x"0d",
          4135 => x"0d",
          4136 => x"3d",
          4137 => x"71",
          4138 => x"e7",
          4139 => x"de",
          4140 => x"81",
          4141 => x"80",
          4142 => x"93",
          4143 => x"c0",
          4144 => x"51",
          4145 => x"81",
          4146 => x"53",
          4147 => x"81",
          4148 => x"52",
          4149 => x"ac",
          4150 => x"c0",
          4151 => x"de",
          4152 => x"2e",
          4153 => x"85",
          4154 => x"87",
          4155 => x"c0",
          4156 => x"74",
          4157 => x"d5",
          4158 => x"52",
          4159 => x"89",
          4160 => x"c0",
          4161 => x"70",
          4162 => x"07",
          4163 => x"81",
          4164 => x"06",
          4165 => x"54",
          4166 => x"c0",
          4167 => x"0d",
          4168 => x"0d",
          4169 => x"53",
          4170 => x"53",
          4171 => x"56",
          4172 => x"81",
          4173 => x"55",
          4174 => x"08",
          4175 => x"52",
          4176 => x"81",
          4177 => x"c0",
          4178 => x"de",
          4179 => x"38",
          4180 => x"05",
          4181 => x"2b",
          4182 => x"80",
          4183 => x"86",
          4184 => x"76",
          4185 => x"38",
          4186 => x"51",
          4187 => x"74",
          4188 => x"0c",
          4189 => x"04",
          4190 => x"63",
          4191 => x"80",
          4192 => x"ec",
          4193 => x"3d",
          4194 => x"3f",
          4195 => x"08",
          4196 => x"c0",
          4197 => x"38",
          4198 => x"73",
          4199 => x"08",
          4200 => x"13",
          4201 => x"58",
          4202 => x"26",
          4203 => x"7c",
          4204 => x"39",
          4205 => x"cc",
          4206 => x"81",
          4207 => x"de",
          4208 => x"33",
          4209 => x"81",
          4210 => x"06",
          4211 => x"75",
          4212 => x"52",
          4213 => x"05",
          4214 => x"3f",
          4215 => x"08",
          4216 => x"38",
          4217 => x"08",
          4218 => x"38",
          4219 => x"08",
          4220 => x"de",
          4221 => x"80",
          4222 => x"81",
          4223 => x"59",
          4224 => x"14",
          4225 => x"ca",
          4226 => x"39",
          4227 => x"81",
          4228 => x"57",
          4229 => x"38",
          4230 => x"18",
          4231 => x"ff",
          4232 => x"81",
          4233 => x"5b",
          4234 => x"08",
          4235 => x"7c",
          4236 => x"12",
          4237 => x"52",
          4238 => x"82",
          4239 => x"06",
          4240 => x"14",
          4241 => x"cb",
          4242 => x"c0",
          4243 => x"ff",
          4244 => x"70",
          4245 => x"82",
          4246 => x"51",
          4247 => x"b4",
          4248 => x"bb",
          4249 => x"de",
          4250 => x"0a",
          4251 => x"70",
          4252 => x"84",
          4253 => x"51",
          4254 => x"ff",
          4255 => x"56",
          4256 => x"38",
          4257 => x"7c",
          4258 => x"0c",
          4259 => x"81",
          4260 => x"74",
          4261 => x"7a",
          4262 => x"0c",
          4263 => x"04",
          4264 => x"79",
          4265 => x"05",
          4266 => x"57",
          4267 => x"81",
          4268 => x"56",
          4269 => x"08",
          4270 => x"91",
          4271 => x"75",
          4272 => x"90",
          4273 => x"81",
          4274 => x"06",
          4275 => x"87",
          4276 => x"2e",
          4277 => x"94",
          4278 => x"73",
          4279 => x"27",
          4280 => x"73",
          4281 => x"de",
          4282 => x"88",
          4283 => x"76",
          4284 => x"3f",
          4285 => x"08",
          4286 => x"0c",
          4287 => x"39",
          4288 => x"52",
          4289 => x"bf",
          4290 => x"de",
          4291 => x"2e",
          4292 => x"83",
          4293 => x"81",
          4294 => x"81",
          4295 => x"06",
          4296 => x"56",
          4297 => x"a0",
          4298 => x"81",
          4299 => x"98",
          4300 => x"94",
          4301 => x"08",
          4302 => x"c0",
          4303 => x"51",
          4304 => x"81",
          4305 => x"56",
          4306 => x"8c",
          4307 => x"17",
          4308 => x"07",
          4309 => x"18",
          4310 => x"2e",
          4311 => x"91",
          4312 => x"55",
          4313 => x"c0",
          4314 => x"0d",
          4315 => x"0d",
          4316 => x"3d",
          4317 => x"52",
          4318 => x"da",
          4319 => x"de",
          4320 => x"81",
          4321 => x"81",
          4322 => x"45",
          4323 => x"52",
          4324 => x"52",
          4325 => x"3f",
          4326 => x"08",
          4327 => x"c0",
          4328 => x"38",
          4329 => x"05",
          4330 => x"2a",
          4331 => x"51",
          4332 => x"55",
          4333 => x"38",
          4334 => x"54",
          4335 => x"81",
          4336 => x"80",
          4337 => x"70",
          4338 => x"54",
          4339 => x"81",
          4340 => x"52",
          4341 => x"c5",
          4342 => x"c0",
          4343 => x"2a",
          4344 => x"51",
          4345 => x"80",
          4346 => x"38",
          4347 => x"de",
          4348 => x"15",
          4349 => x"86",
          4350 => x"81",
          4351 => x"5c",
          4352 => x"3d",
          4353 => x"c7",
          4354 => x"de",
          4355 => x"81",
          4356 => x"80",
          4357 => x"de",
          4358 => x"73",
          4359 => x"3f",
          4360 => x"08",
          4361 => x"c0",
          4362 => x"87",
          4363 => x"39",
          4364 => x"08",
          4365 => x"38",
          4366 => x"08",
          4367 => x"77",
          4368 => x"3f",
          4369 => x"08",
          4370 => x"08",
          4371 => x"de",
          4372 => x"80",
          4373 => x"55",
          4374 => x"94",
          4375 => x"2e",
          4376 => x"53",
          4377 => x"51",
          4378 => x"81",
          4379 => x"55",
          4380 => x"78",
          4381 => x"fe",
          4382 => x"c0",
          4383 => x"81",
          4384 => x"a0",
          4385 => x"e9",
          4386 => x"53",
          4387 => x"05",
          4388 => x"51",
          4389 => x"81",
          4390 => x"54",
          4391 => x"08",
          4392 => x"78",
          4393 => x"8e",
          4394 => x"58",
          4395 => x"81",
          4396 => x"54",
          4397 => x"08",
          4398 => x"54",
          4399 => x"81",
          4400 => x"84",
          4401 => x"06",
          4402 => x"02",
          4403 => x"33",
          4404 => x"81",
          4405 => x"86",
          4406 => x"f6",
          4407 => x"74",
          4408 => x"70",
          4409 => x"c3",
          4410 => x"c0",
          4411 => x"56",
          4412 => x"08",
          4413 => x"54",
          4414 => x"08",
          4415 => x"81",
          4416 => x"82",
          4417 => x"c0",
          4418 => x"09",
          4419 => x"38",
          4420 => x"b4",
          4421 => x"b0",
          4422 => x"c0",
          4423 => x"51",
          4424 => x"81",
          4425 => x"54",
          4426 => x"08",
          4427 => x"8b",
          4428 => x"b4",
          4429 => x"b7",
          4430 => x"54",
          4431 => x"15",
          4432 => x"90",
          4433 => x"34",
          4434 => x"0a",
          4435 => x"19",
          4436 => x"9f",
          4437 => x"78",
          4438 => x"51",
          4439 => x"a0",
          4440 => x"11",
          4441 => x"05",
          4442 => x"b6",
          4443 => x"ae",
          4444 => x"15",
          4445 => x"78",
          4446 => x"53",
          4447 => x"3f",
          4448 => x"0b",
          4449 => x"77",
          4450 => x"3f",
          4451 => x"08",
          4452 => x"c0",
          4453 => x"82",
          4454 => x"52",
          4455 => x"51",
          4456 => x"3f",
          4457 => x"52",
          4458 => x"aa",
          4459 => x"90",
          4460 => x"34",
          4461 => x"0b",
          4462 => x"78",
          4463 => x"b6",
          4464 => x"c0",
          4465 => x"39",
          4466 => x"52",
          4467 => x"be",
          4468 => x"81",
          4469 => x"99",
          4470 => x"da",
          4471 => x"3d",
          4472 => x"d2",
          4473 => x"53",
          4474 => x"84",
          4475 => x"3d",
          4476 => x"3f",
          4477 => x"08",
          4478 => x"c0",
          4479 => x"38",
          4480 => x"3d",
          4481 => x"3d",
          4482 => x"cc",
          4483 => x"de",
          4484 => x"81",
          4485 => x"82",
          4486 => x"81",
          4487 => x"81",
          4488 => x"86",
          4489 => x"aa",
          4490 => x"a4",
          4491 => x"a8",
          4492 => x"05",
          4493 => x"ea",
          4494 => x"77",
          4495 => x"70",
          4496 => x"b4",
          4497 => x"3d",
          4498 => x"51",
          4499 => x"81",
          4500 => x"55",
          4501 => x"08",
          4502 => x"6f",
          4503 => x"06",
          4504 => x"a2",
          4505 => x"92",
          4506 => x"81",
          4507 => x"de",
          4508 => x"2e",
          4509 => x"81",
          4510 => x"51",
          4511 => x"81",
          4512 => x"55",
          4513 => x"08",
          4514 => x"68",
          4515 => x"a8",
          4516 => x"05",
          4517 => x"51",
          4518 => x"3f",
          4519 => x"33",
          4520 => x"8b",
          4521 => x"84",
          4522 => x"06",
          4523 => x"73",
          4524 => x"a0",
          4525 => x"8b",
          4526 => x"54",
          4527 => x"15",
          4528 => x"33",
          4529 => x"70",
          4530 => x"55",
          4531 => x"2e",
          4532 => x"6e",
          4533 => x"df",
          4534 => x"78",
          4535 => x"3f",
          4536 => x"08",
          4537 => x"ff",
          4538 => x"82",
          4539 => x"c0",
          4540 => x"80",
          4541 => x"de",
          4542 => x"78",
          4543 => x"af",
          4544 => x"c0",
          4545 => x"d4",
          4546 => x"55",
          4547 => x"08",
          4548 => x"81",
          4549 => x"73",
          4550 => x"81",
          4551 => x"63",
          4552 => x"76",
          4553 => x"3f",
          4554 => x"0b",
          4555 => x"87",
          4556 => x"c0",
          4557 => x"77",
          4558 => x"3f",
          4559 => x"08",
          4560 => x"c0",
          4561 => x"78",
          4562 => x"aa",
          4563 => x"c0",
          4564 => x"81",
          4565 => x"a8",
          4566 => x"ed",
          4567 => x"80",
          4568 => x"02",
          4569 => x"df",
          4570 => x"57",
          4571 => x"3d",
          4572 => x"96",
          4573 => x"e9",
          4574 => x"c0",
          4575 => x"de",
          4576 => x"cf",
          4577 => x"65",
          4578 => x"d4",
          4579 => x"b5",
          4580 => x"c0",
          4581 => x"de",
          4582 => x"38",
          4583 => x"05",
          4584 => x"06",
          4585 => x"73",
          4586 => x"a7",
          4587 => x"09",
          4588 => x"71",
          4589 => x"06",
          4590 => x"55",
          4591 => x"15",
          4592 => x"81",
          4593 => x"34",
          4594 => x"b4",
          4595 => x"de",
          4596 => x"74",
          4597 => x"0c",
          4598 => x"04",
          4599 => x"64",
          4600 => x"93",
          4601 => x"52",
          4602 => x"d1",
          4603 => x"de",
          4604 => x"81",
          4605 => x"80",
          4606 => x"58",
          4607 => x"3d",
          4608 => x"c8",
          4609 => x"de",
          4610 => x"81",
          4611 => x"b4",
          4612 => x"c7",
          4613 => x"a0",
          4614 => x"55",
          4615 => x"84",
          4616 => x"17",
          4617 => x"2b",
          4618 => x"96",
          4619 => x"b0",
          4620 => x"54",
          4621 => x"15",
          4622 => x"ff",
          4623 => x"81",
          4624 => x"55",
          4625 => x"c0",
          4626 => x"0d",
          4627 => x"0d",
          4628 => x"5a",
          4629 => x"3d",
          4630 => x"99",
          4631 => x"81",
          4632 => x"c0",
          4633 => x"c0",
          4634 => x"81",
          4635 => x"07",
          4636 => x"55",
          4637 => x"2e",
          4638 => x"81",
          4639 => x"55",
          4640 => x"2e",
          4641 => x"7b",
          4642 => x"80",
          4643 => x"70",
          4644 => x"be",
          4645 => x"de",
          4646 => x"81",
          4647 => x"80",
          4648 => x"52",
          4649 => x"dc",
          4650 => x"c0",
          4651 => x"de",
          4652 => x"38",
          4653 => x"08",
          4654 => x"08",
          4655 => x"56",
          4656 => x"19",
          4657 => x"59",
          4658 => x"74",
          4659 => x"56",
          4660 => x"ec",
          4661 => x"75",
          4662 => x"74",
          4663 => x"2e",
          4664 => x"16",
          4665 => x"33",
          4666 => x"73",
          4667 => x"38",
          4668 => x"84",
          4669 => x"06",
          4670 => x"7a",
          4671 => x"76",
          4672 => x"07",
          4673 => x"54",
          4674 => x"80",
          4675 => x"80",
          4676 => x"7b",
          4677 => x"53",
          4678 => x"93",
          4679 => x"c0",
          4680 => x"de",
          4681 => x"38",
          4682 => x"55",
          4683 => x"56",
          4684 => x"8b",
          4685 => x"56",
          4686 => x"83",
          4687 => x"75",
          4688 => x"51",
          4689 => x"3f",
          4690 => x"08",
          4691 => x"81",
          4692 => x"98",
          4693 => x"e6",
          4694 => x"53",
          4695 => x"b8",
          4696 => x"3d",
          4697 => x"3f",
          4698 => x"08",
          4699 => x"08",
          4700 => x"de",
          4701 => x"98",
          4702 => x"a0",
          4703 => x"70",
          4704 => x"ae",
          4705 => x"6d",
          4706 => x"81",
          4707 => x"57",
          4708 => x"74",
          4709 => x"38",
          4710 => x"81",
          4711 => x"81",
          4712 => x"52",
          4713 => x"89",
          4714 => x"c0",
          4715 => x"a5",
          4716 => x"33",
          4717 => x"54",
          4718 => x"3f",
          4719 => x"08",
          4720 => x"38",
          4721 => x"76",
          4722 => x"05",
          4723 => x"39",
          4724 => x"08",
          4725 => x"15",
          4726 => x"ff",
          4727 => x"73",
          4728 => x"38",
          4729 => x"83",
          4730 => x"56",
          4731 => x"75",
          4732 => x"81",
          4733 => x"33",
          4734 => x"2e",
          4735 => x"52",
          4736 => x"51",
          4737 => x"3f",
          4738 => x"08",
          4739 => x"ff",
          4740 => x"38",
          4741 => x"88",
          4742 => x"8a",
          4743 => x"38",
          4744 => x"ec",
          4745 => x"75",
          4746 => x"74",
          4747 => x"73",
          4748 => x"05",
          4749 => x"17",
          4750 => x"70",
          4751 => x"34",
          4752 => x"70",
          4753 => x"ff",
          4754 => x"55",
          4755 => x"26",
          4756 => x"8b",
          4757 => x"86",
          4758 => x"e5",
          4759 => x"38",
          4760 => x"99",
          4761 => x"05",
          4762 => x"70",
          4763 => x"73",
          4764 => x"81",
          4765 => x"ff",
          4766 => x"ed",
          4767 => x"80",
          4768 => x"91",
          4769 => x"55",
          4770 => x"3f",
          4771 => x"08",
          4772 => x"c0",
          4773 => x"38",
          4774 => x"51",
          4775 => x"3f",
          4776 => x"08",
          4777 => x"c0",
          4778 => x"76",
          4779 => x"67",
          4780 => x"34",
          4781 => x"81",
          4782 => x"84",
          4783 => x"06",
          4784 => x"80",
          4785 => x"2e",
          4786 => x"81",
          4787 => x"ff",
          4788 => x"81",
          4789 => x"54",
          4790 => x"08",
          4791 => x"53",
          4792 => x"08",
          4793 => x"ff",
          4794 => x"67",
          4795 => x"8b",
          4796 => x"53",
          4797 => x"51",
          4798 => x"3f",
          4799 => x"0b",
          4800 => x"79",
          4801 => x"ee",
          4802 => x"c0",
          4803 => x"55",
          4804 => x"c0",
          4805 => x"0d",
          4806 => x"0d",
          4807 => x"88",
          4808 => x"05",
          4809 => x"fc",
          4810 => x"54",
          4811 => x"d2",
          4812 => x"de",
          4813 => x"81",
          4814 => x"82",
          4815 => x"1a",
          4816 => x"82",
          4817 => x"80",
          4818 => x"8c",
          4819 => x"78",
          4820 => x"1a",
          4821 => x"2a",
          4822 => x"51",
          4823 => x"90",
          4824 => x"82",
          4825 => x"58",
          4826 => x"81",
          4827 => x"39",
          4828 => x"22",
          4829 => x"70",
          4830 => x"56",
          4831 => x"fb",
          4832 => x"14",
          4833 => x"30",
          4834 => x"9f",
          4835 => x"c0",
          4836 => x"19",
          4837 => x"5a",
          4838 => x"81",
          4839 => x"38",
          4840 => x"77",
          4841 => x"82",
          4842 => x"56",
          4843 => x"74",
          4844 => x"ff",
          4845 => x"81",
          4846 => x"55",
          4847 => x"75",
          4848 => x"82",
          4849 => x"c0",
          4850 => x"ff",
          4851 => x"de",
          4852 => x"2e",
          4853 => x"81",
          4854 => x"8e",
          4855 => x"56",
          4856 => x"09",
          4857 => x"38",
          4858 => x"59",
          4859 => x"77",
          4860 => x"06",
          4861 => x"87",
          4862 => x"39",
          4863 => x"ba",
          4864 => x"55",
          4865 => x"2e",
          4866 => x"15",
          4867 => x"2e",
          4868 => x"83",
          4869 => x"75",
          4870 => x"7e",
          4871 => x"a8",
          4872 => x"c0",
          4873 => x"de",
          4874 => x"ce",
          4875 => x"16",
          4876 => x"56",
          4877 => x"38",
          4878 => x"19",
          4879 => x"8c",
          4880 => x"7d",
          4881 => x"38",
          4882 => x"0c",
          4883 => x"0c",
          4884 => x"80",
          4885 => x"73",
          4886 => x"98",
          4887 => x"05",
          4888 => x"57",
          4889 => x"26",
          4890 => x"7b",
          4891 => x"0c",
          4892 => x"81",
          4893 => x"84",
          4894 => x"54",
          4895 => x"c0",
          4896 => x"0d",
          4897 => x"0d",
          4898 => x"88",
          4899 => x"05",
          4900 => x"54",
          4901 => x"c5",
          4902 => x"56",
          4903 => x"de",
          4904 => x"8b",
          4905 => x"de",
          4906 => x"29",
          4907 => x"05",
          4908 => x"55",
          4909 => x"84",
          4910 => x"34",
          4911 => x"08",
          4912 => x"5f",
          4913 => x"51",
          4914 => x"3f",
          4915 => x"08",
          4916 => x"70",
          4917 => x"57",
          4918 => x"8b",
          4919 => x"82",
          4920 => x"06",
          4921 => x"56",
          4922 => x"38",
          4923 => x"05",
          4924 => x"7e",
          4925 => x"f0",
          4926 => x"c0",
          4927 => x"67",
          4928 => x"2e",
          4929 => x"82",
          4930 => x"8b",
          4931 => x"75",
          4932 => x"80",
          4933 => x"81",
          4934 => x"2e",
          4935 => x"80",
          4936 => x"38",
          4937 => x"0a",
          4938 => x"ff",
          4939 => x"55",
          4940 => x"86",
          4941 => x"8a",
          4942 => x"89",
          4943 => x"2a",
          4944 => x"77",
          4945 => x"59",
          4946 => x"81",
          4947 => x"70",
          4948 => x"07",
          4949 => x"56",
          4950 => x"38",
          4951 => x"05",
          4952 => x"7e",
          4953 => x"80",
          4954 => x"81",
          4955 => x"8a",
          4956 => x"83",
          4957 => x"06",
          4958 => x"08",
          4959 => x"74",
          4960 => x"41",
          4961 => x"56",
          4962 => x"8a",
          4963 => x"61",
          4964 => x"55",
          4965 => x"27",
          4966 => x"93",
          4967 => x"80",
          4968 => x"38",
          4969 => x"70",
          4970 => x"43",
          4971 => x"95",
          4972 => x"06",
          4973 => x"2e",
          4974 => x"77",
          4975 => x"74",
          4976 => x"83",
          4977 => x"06",
          4978 => x"82",
          4979 => x"2e",
          4980 => x"78",
          4981 => x"2e",
          4982 => x"80",
          4983 => x"ae",
          4984 => x"2a",
          4985 => x"81",
          4986 => x"56",
          4987 => x"2e",
          4988 => x"77",
          4989 => x"81",
          4990 => x"79",
          4991 => x"70",
          4992 => x"5a",
          4993 => x"86",
          4994 => x"27",
          4995 => x"52",
          4996 => x"f6",
          4997 => x"de",
          4998 => x"29",
          4999 => x"70",
          5000 => x"55",
          5001 => x"0b",
          5002 => x"08",
          5003 => x"05",
          5004 => x"ff",
          5005 => x"27",
          5006 => x"88",
          5007 => x"ae",
          5008 => x"2a",
          5009 => x"81",
          5010 => x"56",
          5011 => x"2e",
          5012 => x"77",
          5013 => x"81",
          5014 => x"79",
          5015 => x"70",
          5016 => x"5a",
          5017 => x"86",
          5018 => x"27",
          5019 => x"52",
          5020 => x"f6",
          5021 => x"de",
          5022 => x"84",
          5023 => x"de",
          5024 => x"f5",
          5025 => x"81",
          5026 => x"c0",
          5027 => x"de",
          5028 => x"71",
          5029 => x"83",
          5030 => x"5e",
          5031 => x"89",
          5032 => x"5c",
          5033 => x"1c",
          5034 => x"05",
          5035 => x"ff",
          5036 => x"70",
          5037 => x"31",
          5038 => x"57",
          5039 => x"83",
          5040 => x"06",
          5041 => x"1c",
          5042 => x"5c",
          5043 => x"1d",
          5044 => x"29",
          5045 => x"31",
          5046 => x"55",
          5047 => x"87",
          5048 => x"7c",
          5049 => x"7a",
          5050 => x"31",
          5051 => x"f5",
          5052 => x"de",
          5053 => x"7d",
          5054 => x"81",
          5055 => x"81",
          5056 => x"83",
          5057 => x"80",
          5058 => x"87",
          5059 => x"81",
          5060 => x"fd",
          5061 => x"f8",
          5062 => x"2e",
          5063 => x"80",
          5064 => x"ff",
          5065 => x"de",
          5066 => x"a0",
          5067 => x"38",
          5068 => x"74",
          5069 => x"86",
          5070 => x"fd",
          5071 => x"81",
          5072 => x"80",
          5073 => x"83",
          5074 => x"39",
          5075 => x"08",
          5076 => x"92",
          5077 => x"b8",
          5078 => x"59",
          5079 => x"27",
          5080 => x"86",
          5081 => x"55",
          5082 => x"09",
          5083 => x"38",
          5084 => x"f5",
          5085 => x"38",
          5086 => x"55",
          5087 => x"86",
          5088 => x"80",
          5089 => x"7a",
          5090 => x"b9",
          5091 => x"81",
          5092 => x"7a",
          5093 => x"8a",
          5094 => x"52",
          5095 => x"ff",
          5096 => x"79",
          5097 => x"7b",
          5098 => x"06",
          5099 => x"51",
          5100 => x"3f",
          5101 => x"1c",
          5102 => x"32",
          5103 => x"96",
          5104 => x"06",
          5105 => x"91",
          5106 => x"a1",
          5107 => x"55",
          5108 => x"ff",
          5109 => x"74",
          5110 => x"06",
          5111 => x"51",
          5112 => x"3f",
          5113 => x"52",
          5114 => x"ff",
          5115 => x"f8",
          5116 => x"34",
          5117 => x"1b",
          5118 => x"d9",
          5119 => x"52",
          5120 => x"ff",
          5121 => x"60",
          5122 => x"51",
          5123 => x"3f",
          5124 => x"09",
          5125 => x"cb",
          5126 => x"b2",
          5127 => x"c3",
          5128 => x"a0",
          5129 => x"52",
          5130 => x"ff",
          5131 => x"82",
          5132 => x"51",
          5133 => x"3f",
          5134 => x"1b",
          5135 => x"95",
          5136 => x"b2",
          5137 => x"a0",
          5138 => x"80",
          5139 => x"1c",
          5140 => x"80",
          5141 => x"93",
          5142 => x"fc",
          5143 => x"1b",
          5144 => x"82",
          5145 => x"52",
          5146 => x"ff",
          5147 => x"7c",
          5148 => x"06",
          5149 => x"51",
          5150 => x"3f",
          5151 => x"a4",
          5152 => x"0b",
          5153 => x"93",
          5154 => x"90",
          5155 => x"51",
          5156 => x"3f",
          5157 => x"52",
          5158 => x"70",
          5159 => x"9f",
          5160 => x"54",
          5161 => x"52",
          5162 => x"9b",
          5163 => x"56",
          5164 => x"08",
          5165 => x"7d",
          5166 => x"81",
          5167 => x"38",
          5168 => x"86",
          5169 => x"52",
          5170 => x"9b",
          5171 => x"80",
          5172 => x"7a",
          5173 => x"ed",
          5174 => x"85",
          5175 => x"7a",
          5176 => x"8f",
          5177 => x"85",
          5178 => x"83",
          5179 => x"ff",
          5180 => x"ff",
          5181 => x"e8",
          5182 => x"9e",
          5183 => x"52",
          5184 => x"51",
          5185 => x"3f",
          5186 => x"52",
          5187 => x"9e",
          5188 => x"54",
          5189 => x"53",
          5190 => x"51",
          5191 => x"3f",
          5192 => x"16",
          5193 => x"7e",
          5194 => x"d8",
          5195 => x"80",
          5196 => x"ff",
          5197 => x"7f",
          5198 => x"7d",
          5199 => x"81",
          5200 => x"f8",
          5201 => x"ff",
          5202 => x"ff",
          5203 => x"51",
          5204 => x"3f",
          5205 => x"88",
          5206 => x"39",
          5207 => x"f8",
          5208 => x"2e",
          5209 => x"55",
          5210 => x"51",
          5211 => x"3f",
          5212 => x"57",
          5213 => x"83",
          5214 => x"76",
          5215 => x"7a",
          5216 => x"ff",
          5217 => x"81",
          5218 => x"82",
          5219 => x"80",
          5220 => x"c0",
          5221 => x"51",
          5222 => x"3f",
          5223 => x"78",
          5224 => x"74",
          5225 => x"18",
          5226 => x"2e",
          5227 => x"79",
          5228 => x"2e",
          5229 => x"55",
          5230 => x"62",
          5231 => x"74",
          5232 => x"75",
          5233 => x"7e",
          5234 => x"b8",
          5235 => x"c0",
          5236 => x"38",
          5237 => x"78",
          5238 => x"74",
          5239 => x"56",
          5240 => x"93",
          5241 => x"66",
          5242 => x"26",
          5243 => x"56",
          5244 => x"83",
          5245 => x"64",
          5246 => x"77",
          5247 => x"84",
          5248 => x"52",
          5249 => x"9d",
          5250 => x"d4",
          5251 => x"51",
          5252 => x"3f",
          5253 => x"55",
          5254 => x"81",
          5255 => x"34",
          5256 => x"16",
          5257 => x"16",
          5258 => x"16",
          5259 => x"05",
          5260 => x"c1",
          5261 => x"fe",
          5262 => x"fe",
          5263 => x"34",
          5264 => x"08",
          5265 => x"07",
          5266 => x"16",
          5267 => x"c0",
          5268 => x"34",
          5269 => x"c6",
          5270 => x"9c",
          5271 => x"52",
          5272 => x"51",
          5273 => x"3f",
          5274 => x"53",
          5275 => x"51",
          5276 => x"3f",
          5277 => x"de",
          5278 => x"38",
          5279 => x"52",
          5280 => x"99",
          5281 => x"56",
          5282 => x"08",
          5283 => x"39",
          5284 => x"39",
          5285 => x"39",
          5286 => x"08",
          5287 => x"de",
          5288 => x"3d",
          5289 => x"3d",
          5290 => x"5b",
          5291 => x"60",
          5292 => x"57",
          5293 => x"25",
          5294 => x"3d",
          5295 => x"55",
          5296 => x"15",
          5297 => x"c9",
          5298 => x"81",
          5299 => x"06",
          5300 => x"3d",
          5301 => x"8d",
          5302 => x"74",
          5303 => x"05",
          5304 => x"17",
          5305 => x"2e",
          5306 => x"c9",
          5307 => x"34",
          5308 => x"83",
          5309 => x"74",
          5310 => x"0c",
          5311 => x"04",
          5312 => x"73",
          5313 => x"26",
          5314 => x"71",
          5315 => x"c6",
          5316 => x"71",
          5317 => x"cf",
          5318 => x"80",
          5319 => x"fc",
          5320 => x"39",
          5321 => x"51",
          5322 => x"81",
          5323 => x"80",
          5324 => x"d0",
          5325 => x"e4",
          5326 => x"c4",
          5327 => x"39",
          5328 => x"51",
          5329 => x"81",
          5330 => x"80",
          5331 => x"d1",
          5332 => x"c8",
          5333 => x"98",
          5334 => x"39",
          5335 => x"51",
          5336 => x"d1",
          5337 => x"39",
          5338 => x"51",
          5339 => x"d2",
          5340 => x"39",
          5341 => x"51",
          5342 => x"d2",
          5343 => x"39",
          5344 => x"51",
          5345 => x"d2",
          5346 => x"39",
          5347 => x"51",
          5348 => x"d3",
          5349 => x"39",
          5350 => x"51",
          5351 => x"3f",
          5352 => x"04",
          5353 => x"77",
          5354 => x"74",
          5355 => x"8a",
          5356 => x"75",
          5357 => x"51",
          5358 => x"e8",
          5359 => x"fe",
          5360 => x"81",
          5361 => x"52",
          5362 => x"eb",
          5363 => x"de",
          5364 => x"79",
          5365 => x"81",
          5366 => x"ff",
          5367 => x"87",
          5368 => x"f5",
          5369 => x"7f",
          5370 => x"05",
          5371 => x"33",
          5372 => x"66",
          5373 => x"5a",
          5374 => x"78",
          5375 => x"dc",
          5376 => x"a0",
          5377 => x"e4",
          5378 => x"b4",
          5379 => x"74",
          5380 => x"fc",
          5381 => x"2e",
          5382 => x"a0",
          5383 => x"80",
          5384 => x"16",
          5385 => x"27",
          5386 => x"22",
          5387 => x"e8",
          5388 => x"f0",
          5389 => x"81",
          5390 => x"ff",
          5391 => x"82",
          5392 => x"c3",
          5393 => x"53",
          5394 => x"8e",
          5395 => x"52",
          5396 => x"51",
          5397 => x"3f",
          5398 => x"d3",
          5399 => x"85",
          5400 => x"15",
          5401 => x"74",
          5402 => x"78",
          5403 => x"72",
          5404 => x"d3",
          5405 => x"8b",
          5406 => x"39",
          5407 => x"51",
          5408 => x"3f",
          5409 => x"a0",
          5410 => x"af",
          5411 => x"39",
          5412 => x"51",
          5413 => x"3f",
          5414 => x"77",
          5415 => x"74",
          5416 => x"79",
          5417 => x"55",
          5418 => x"27",
          5419 => x"80",
          5420 => x"73",
          5421 => x"85",
          5422 => x"83",
          5423 => x"fe",
          5424 => x"81",
          5425 => x"39",
          5426 => x"51",
          5427 => x"3f",
          5428 => x"1a",
          5429 => x"f9",
          5430 => x"de",
          5431 => x"2b",
          5432 => x"51",
          5433 => x"2e",
          5434 => x"a5",
          5435 => x"9d",
          5436 => x"c0",
          5437 => x"70",
          5438 => x"a0",
          5439 => x"70",
          5440 => x"2a",
          5441 => x"51",
          5442 => x"2e",
          5443 => x"dd",
          5444 => x"2e",
          5445 => x"85",
          5446 => x"8c",
          5447 => x"53",
          5448 => x"fd",
          5449 => x"53",
          5450 => x"c0",
          5451 => x"0d",
          5452 => x"0d",
          5453 => x"05",
          5454 => x"33",
          5455 => x"70",
          5456 => x"25",
          5457 => x"74",
          5458 => x"51",
          5459 => x"56",
          5460 => x"80",
          5461 => x"53",
          5462 => x"3d",
          5463 => x"ff",
          5464 => x"81",
          5465 => x"56",
          5466 => x"08",
          5467 => x"de",
          5468 => x"c0",
          5469 => x"81",
          5470 => x"59",
          5471 => x"05",
          5472 => x"53",
          5473 => x"51",
          5474 => x"81",
          5475 => x"56",
          5476 => x"08",
          5477 => x"55",
          5478 => x"89",
          5479 => x"75",
          5480 => x"d8",
          5481 => x"d8",
          5482 => x"85",
          5483 => x"70",
          5484 => x"25",
          5485 => x"80",
          5486 => x"74",
          5487 => x"38",
          5488 => x"53",
          5489 => x"88",
          5490 => x"51",
          5491 => x"75",
          5492 => x"de",
          5493 => x"3d",
          5494 => x"3d",
          5495 => x"84",
          5496 => x"33",
          5497 => x"57",
          5498 => x"52",
          5499 => x"c1",
          5500 => x"c0",
          5501 => x"75",
          5502 => x"38",
          5503 => x"98",
          5504 => x"60",
          5505 => x"81",
          5506 => x"7e",
          5507 => x"77",
          5508 => x"c0",
          5509 => x"39",
          5510 => x"81",
          5511 => x"89",
          5512 => x"fc",
          5513 => x"9b",
          5514 => x"d4",
          5515 => x"d4",
          5516 => x"ff",
          5517 => x"81",
          5518 => x"51",
          5519 => x"3f",
          5520 => x"54",
          5521 => x"53",
          5522 => x"33",
          5523 => x"c0",
          5524 => x"d0",
          5525 => x"2e",
          5526 => x"fb",
          5527 => x"3d",
          5528 => x"3d",
          5529 => x"96",
          5530 => x"ff",
          5531 => x"81",
          5532 => x"ad",
          5533 => x"dc",
          5534 => x"a5",
          5535 => x"fe",
          5536 => x"72",
          5537 => x"81",
          5538 => x"71",
          5539 => x"38",
          5540 => x"f2",
          5541 => x"d4",
          5542 => x"f4",
          5543 => x"51",
          5544 => x"3f",
          5545 => x"70",
          5546 => x"52",
          5547 => x"95",
          5548 => x"fe",
          5549 => x"81",
          5550 => x"fe",
          5551 => x"80",
          5552 => x"dd",
          5553 => x"2a",
          5554 => x"51",
          5555 => x"2e",
          5556 => x"51",
          5557 => x"3f",
          5558 => x"51",
          5559 => x"3f",
          5560 => x"f1",
          5561 => x"84",
          5562 => x"06",
          5563 => x"80",
          5564 => x"81",
          5565 => x"a9",
          5566 => x"b0",
          5567 => x"a1",
          5568 => x"fe",
          5569 => x"72",
          5570 => x"81",
          5571 => x"71",
          5572 => x"38",
          5573 => x"f1",
          5574 => x"d5",
          5575 => x"f3",
          5576 => x"51",
          5577 => x"3f",
          5578 => x"70",
          5579 => x"52",
          5580 => x"95",
          5581 => x"fe",
          5582 => x"81",
          5583 => x"fe",
          5584 => x"80",
          5585 => x"d9",
          5586 => x"2a",
          5587 => x"51",
          5588 => x"2e",
          5589 => x"51",
          5590 => x"3f",
          5591 => x"51",
          5592 => x"3f",
          5593 => x"f0",
          5594 => x"88",
          5595 => x"06",
          5596 => x"80",
          5597 => x"81",
          5598 => x"a5",
          5599 => x"80",
          5600 => x"9d",
          5601 => x"fe",
          5602 => x"fe",
          5603 => x"84",
          5604 => x"fa",
          5605 => x"70",
          5606 => x"55",
          5607 => x"2e",
          5608 => x"8e",
          5609 => x"0c",
          5610 => x"53",
          5611 => x"81",
          5612 => x"74",
          5613 => x"ff",
          5614 => x"53",
          5615 => x"83",
          5616 => x"74",
          5617 => x"38",
          5618 => x"75",
          5619 => x"53",
          5620 => x"09",
          5621 => x"38",
          5622 => x"81",
          5623 => x"80",
          5624 => x"29",
          5625 => x"05",
          5626 => x"70",
          5627 => x"fe",
          5628 => x"81",
          5629 => x"8b",
          5630 => x"33",
          5631 => x"2e",
          5632 => x"81",
          5633 => x"ff",
          5634 => x"94",
          5635 => x"38",
          5636 => x"81",
          5637 => x"88",
          5638 => x"fb",
          5639 => x"79",
          5640 => x"56",
          5641 => x"51",
          5642 => x"3f",
          5643 => x"33",
          5644 => x"38",
          5645 => x"d6",
          5646 => x"f5",
          5647 => x"b9",
          5648 => x"de",
          5649 => x"70",
          5650 => x"08",
          5651 => x"82",
          5652 => x"51",
          5653 => x"db",
          5654 => x"db",
          5655 => x"73",
          5656 => x"81",
          5657 => x"81",
          5658 => x"74",
          5659 => x"f4",
          5660 => x"de",
          5661 => x"2e",
          5662 => x"de",
          5663 => x"fe",
          5664 => x"8e",
          5665 => x"c4",
          5666 => x"3f",
          5667 => x"db",
          5668 => x"db",
          5669 => x"73",
          5670 => x"81",
          5671 => x"74",
          5672 => x"ff",
          5673 => x"80",
          5674 => x"c0",
          5675 => x"0d",
          5676 => x"0d",
          5677 => x"81",
          5678 => x"40",
          5679 => x"7c",
          5680 => x"d7",
          5681 => x"c0",
          5682 => x"06",
          5683 => x"2e",
          5684 => x"a2",
          5685 => x"d0",
          5686 => x"70",
          5687 => x"82",
          5688 => x"53",
          5689 => x"df",
          5690 => x"b7",
          5691 => x"de",
          5692 => x"2e",
          5693 => x"d6",
          5694 => x"bc",
          5695 => x"40",
          5696 => x"8c",
          5697 => x"b8",
          5698 => x"70",
          5699 => x"f8",
          5700 => x"fe",
          5701 => x"3d",
          5702 => x"51",
          5703 => x"81",
          5704 => x"90",
          5705 => x"2c",
          5706 => x"80",
          5707 => x"ce",
          5708 => x"c3",
          5709 => x"38",
          5710 => x"83",
          5711 => x"ab",
          5712 => x"78",
          5713 => x"af",
          5714 => x"24",
          5715 => x"80",
          5716 => x"38",
          5717 => x"78",
          5718 => x"82",
          5719 => x"2e",
          5720 => x"8f",
          5721 => x"80",
          5722 => x"87",
          5723 => x"c0",
          5724 => x"78",
          5725 => x"a9",
          5726 => x"2e",
          5727 => x"8f",
          5728 => x"80",
          5729 => x"9e",
          5730 => x"c2",
          5731 => x"38",
          5732 => x"78",
          5733 => x"8d",
          5734 => x"80",
          5735 => x"38",
          5736 => x"2e",
          5737 => x"78",
          5738 => x"8b",
          5739 => x"c5",
          5740 => x"38",
          5741 => x"78",
          5742 => x"8d",
          5743 => x"80",
          5744 => x"ab",
          5745 => x"39",
          5746 => x"2e",
          5747 => x"78",
          5748 => x"92",
          5749 => x"f8",
          5750 => x"38",
          5751 => x"2e",
          5752 => x"8e",
          5753 => x"81",
          5754 => x"b4",
          5755 => x"85",
          5756 => x"38",
          5757 => x"b7",
          5758 => x"11",
          5759 => x"05",
          5760 => x"95",
          5761 => x"c0",
          5762 => x"81",
          5763 => x"90",
          5764 => x"3d",
          5765 => x"53",
          5766 => x"51",
          5767 => x"3f",
          5768 => x"08",
          5769 => x"38",
          5770 => x"83",
          5771 => x"02",
          5772 => x"33",
          5773 => x"cf",
          5774 => x"ff",
          5775 => x"81",
          5776 => x"81",
          5777 => x"78",
          5778 => x"d7",
          5779 => x"f9",
          5780 => x"5f",
          5781 => x"81",
          5782 => x"8c",
          5783 => x"3d",
          5784 => x"53",
          5785 => x"51",
          5786 => x"3f",
          5787 => x"08",
          5788 => x"8d",
          5789 => x"80",
          5790 => x"cf",
          5791 => x"ff",
          5792 => x"81",
          5793 => x"52",
          5794 => x"51",
          5795 => x"b7",
          5796 => x"11",
          5797 => x"05",
          5798 => x"fd",
          5799 => x"c0",
          5800 => x"87",
          5801 => x"26",
          5802 => x"b7",
          5803 => x"11",
          5804 => x"05",
          5805 => x"e1",
          5806 => x"c0",
          5807 => x"81",
          5808 => x"43",
          5809 => x"d7",
          5810 => x"51",
          5811 => x"3f",
          5812 => x"05",
          5813 => x"52",
          5814 => x"29",
          5815 => x"05",
          5816 => x"fb",
          5817 => x"c0",
          5818 => x"38",
          5819 => x"51",
          5820 => x"3f",
          5821 => x"89",
          5822 => x"fe",
          5823 => x"fe",
          5824 => x"81",
          5825 => x"b8",
          5826 => x"05",
          5827 => x"e6",
          5828 => x"53",
          5829 => x"08",
          5830 => x"f4",
          5831 => x"d5",
          5832 => x"fe",
          5833 => x"fe",
          5834 => x"81",
          5835 => x"b8",
          5836 => x"05",
          5837 => x"e5",
          5838 => x"de",
          5839 => x"3d",
          5840 => x"52",
          5841 => x"ec",
          5842 => x"c0",
          5843 => x"fe",
          5844 => x"59",
          5845 => x"3f",
          5846 => x"58",
          5847 => x"57",
          5848 => x"55",
          5849 => x"08",
          5850 => x"54",
          5851 => x"52",
          5852 => x"e6",
          5853 => x"c0",
          5854 => x"fb",
          5855 => x"de",
          5856 => x"ee",
          5857 => x"f9",
          5858 => x"fe",
          5859 => x"fe",
          5860 => x"fe",
          5861 => x"81",
          5862 => x"80",
          5863 => x"38",
          5864 => x"f0",
          5865 => x"f8",
          5866 => x"fe",
          5867 => x"de",
          5868 => x"2e",
          5869 => x"b7",
          5870 => x"11",
          5871 => x"05",
          5872 => x"d5",
          5873 => x"c0",
          5874 => x"81",
          5875 => x"42",
          5876 => x"51",
          5877 => x"3f",
          5878 => x"5a",
          5879 => x"88",
          5880 => x"59",
          5881 => x"84",
          5882 => x"7a",
          5883 => x"38",
          5884 => x"b7",
          5885 => x"11",
          5886 => x"05",
          5887 => x"99",
          5888 => x"c0",
          5889 => x"38",
          5890 => x"33",
          5891 => x"2e",
          5892 => x"db",
          5893 => x"80",
          5894 => x"db",
          5895 => x"78",
          5896 => x"38",
          5897 => x"08",
          5898 => x"81",
          5899 => x"59",
          5900 => x"88",
          5901 => x"9c",
          5902 => x"39",
          5903 => x"33",
          5904 => x"2e",
          5905 => x"db",
          5906 => x"9a",
          5907 => x"d2",
          5908 => x"80",
          5909 => x"81",
          5910 => x"44",
          5911 => x"db",
          5912 => x"80",
          5913 => x"3d",
          5914 => x"53",
          5915 => x"51",
          5916 => x"3f",
          5917 => x"08",
          5918 => x"81",
          5919 => x"59",
          5920 => x"89",
          5921 => x"90",
          5922 => x"cc",
          5923 => x"d5",
          5924 => x"80",
          5925 => x"81",
          5926 => x"43",
          5927 => x"db",
          5928 => x"78",
          5929 => x"38",
          5930 => x"08",
          5931 => x"81",
          5932 => x"59",
          5933 => x"88",
          5934 => x"a8",
          5935 => x"39",
          5936 => x"33",
          5937 => x"2e",
          5938 => x"db",
          5939 => x"88",
          5940 => x"bc",
          5941 => x"43",
          5942 => x"ec",
          5943 => x"f8",
          5944 => x"fc",
          5945 => x"de",
          5946 => x"2e",
          5947 => x"62",
          5948 => x"88",
          5949 => x"81",
          5950 => x"2e",
          5951 => x"80",
          5952 => x"79",
          5953 => x"38",
          5954 => x"d7",
          5955 => x"f4",
          5956 => x"55",
          5957 => x"53",
          5958 => x"51",
          5959 => x"81",
          5960 => x"86",
          5961 => x"3d",
          5962 => x"53",
          5963 => x"51",
          5964 => x"3f",
          5965 => x"08",
          5966 => x"c5",
          5967 => x"fe",
          5968 => x"fe",
          5969 => x"fe",
          5970 => x"81",
          5971 => x"80",
          5972 => x"63",
          5973 => x"cb",
          5974 => x"34",
          5975 => x"44",
          5976 => x"f0",
          5977 => x"f8",
          5978 => x"fb",
          5979 => x"de",
          5980 => x"38",
          5981 => x"63",
          5982 => x"52",
          5983 => x"51",
          5984 => x"3f",
          5985 => x"79",
          5986 => x"f2",
          5987 => x"79",
          5988 => x"ae",
          5989 => x"38",
          5990 => x"a0",
          5991 => x"fe",
          5992 => x"fe",
          5993 => x"fe",
          5994 => x"81",
          5995 => x"80",
          5996 => x"63",
          5997 => x"cb",
          5998 => x"34",
          5999 => x"44",
          6000 => x"81",
          6001 => x"fe",
          6002 => x"ff",
          6003 => x"3d",
          6004 => x"53",
          6005 => x"51",
          6006 => x"3f",
          6007 => x"08",
          6008 => x"9d",
          6009 => x"fe",
          6010 => x"fe",
          6011 => x"fe",
          6012 => x"81",
          6013 => x"80",
          6014 => x"60",
          6015 => x"05",
          6016 => x"82",
          6017 => x"78",
          6018 => x"fe",
          6019 => x"fe",
          6020 => x"fe",
          6021 => x"81",
          6022 => x"df",
          6023 => x"39",
          6024 => x"54",
          6025 => x"94",
          6026 => x"f8",
          6027 => x"52",
          6028 => x"f8",
          6029 => x"45",
          6030 => x"78",
          6031 => x"c1",
          6032 => x"26",
          6033 => x"82",
          6034 => x"39",
          6035 => x"e4",
          6036 => x"f8",
          6037 => x"fb",
          6038 => x"de",
          6039 => x"2e",
          6040 => x"59",
          6041 => x"22",
          6042 => x"05",
          6043 => x"41",
          6044 => x"81",
          6045 => x"fe",
          6046 => x"ff",
          6047 => x"3d",
          6048 => x"53",
          6049 => x"51",
          6050 => x"3f",
          6051 => x"08",
          6052 => x"ed",
          6053 => x"fe",
          6054 => x"fe",
          6055 => x"fe",
          6056 => x"81",
          6057 => x"80",
          6058 => x"60",
          6059 => x"59",
          6060 => x"41",
          6061 => x"e4",
          6062 => x"f8",
          6063 => x"fa",
          6064 => x"de",
          6065 => x"38",
          6066 => x"60",
          6067 => x"52",
          6068 => x"51",
          6069 => x"3f",
          6070 => x"79",
          6071 => x"9e",
          6072 => x"79",
          6073 => x"ae",
          6074 => x"38",
          6075 => x"9c",
          6076 => x"fe",
          6077 => x"fe",
          6078 => x"fe",
          6079 => x"81",
          6080 => x"80",
          6081 => x"60",
          6082 => x"59",
          6083 => x"41",
          6084 => x"81",
          6085 => x"fe",
          6086 => x"ff",
          6087 => x"3d",
          6088 => x"53",
          6089 => x"51",
          6090 => x"3f",
          6091 => x"08",
          6092 => x"81",
          6093 => x"59",
          6094 => x"89",
          6095 => x"8c",
          6096 => x"cd",
          6097 => x"d5",
          6098 => x"80",
          6099 => x"81",
          6100 => x"44",
          6101 => x"db",
          6102 => x"78",
          6103 => x"38",
          6104 => x"08",
          6105 => x"81",
          6106 => x"59",
          6107 => x"88",
          6108 => x"a4",
          6109 => x"39",
          6110 => x"33",
          6111 => x"2e",
          6112 => x"db",
          6113 => x"89",
          6114 => x"bc",
          6115 => x"05",
          6116 => x"fe",
          6117 => x"fe",
          6118 => x"fe",
          6119 => x"81",
          6120 => x"80",
          6121 => x"db",
          6122 => x"78",
          6123 => x"38",
          6124 => x"08",
          6125 => x"39",
          6126 => x"33",
          6127 => x"2e",
          6128 => x"db",
          6129 => x"bb",
          6130 => x"d6",
          6131 => x"80",
          6132 => x"81",
          6133 => x"43",
          6134 => x"db",
          6135 => x"78",
          6136 => x"38",
          6137 => x"08",
          6138 => x"81",
          6139 => x"59",
          6140 => x"88",
          6141 => x"b0",
          6142 => x"39",
          6143 => x"08",
          6144 => x"b7",
          6145 => x"11",
          6146 => x"05",
          6147 => x"89",
          6148 => x"c0",
          6149 => x"81",
          6150 => x"42",
          6151 => x"51",
          6152 => x"3f",
          6153 => x"63",
          6154 => x"79",
          6155 => x"62",
          6156 => x"06",
          6157 => x"53",
          6158 => x"d8",
          6159 => x"f3",
          6160 => x"1a",
          6161 => x"81",
          6162 => x"b9",
          6163 => x"cc",
          6164 => x"ec",
          6165 => x"fe",
          6166 => x"f1",
          6167 => x"d8",
          6168 => x"ed",
          6169 => x"51",
          6170 => x"3f",
          6171 => x"84",
          6172 => x"87",
          6173 => x"0c",
          6174 => x"0b",
          6175 => x"94",
          6176 => x"fc",
          6177 => x"b8",
          6178 => x"39",
          6179 => x"51",
          6180 => x"3f",
          6181 => x"0b",
          6182 => x"84",
          6183 => x"83",
          6184 => x"94",
          6185 => x"d9",
          6186 => x"fe",
          6187 => x"fe",
          6188 => x"fe",
          6189 => x"81",
          6190 => x"80",
          6191 => x"38",
          6192 => x"d9",
          6193 => x"f2",
          6194 => x"59",
          6195 => x"3d",
          6196 => x"53",
          6197 => x"51",
          6198 => x"3f",
          6199 => x"08",
          6200 => x"9d",
          6201 => x"81",
          6202 => x"fe",
          6203 => x"63",
          6204 => x"81",
          6205 => x"5e",
          6206 => x"08",
          6207 => x"81",
          6208 => x"c0",
          6209 => x"d9",
          6210 => x"f2",
          6211 => x"f1",
          6212 => x"f8",
          6213 => x"a8",
          6214 => x"e5",
          6215 => x"39",
          6216 => x"51",
          6217 => x"3f",
          6218 => x"a0",
          6219 => x"81",
          6220 => x"39",
          6221 => x"51",
          6222 => x"2e",
          6223 => x"7c",
          6224 => x"dc",
          6225 => x"60",
          6226 => x"78",
          6227 => x"d0",
          6228 => x"fe",
          6229 => x"fe",
          6230 => x"81",
          6231 => x"7a",
          6232 => x"82",
          6233 => x"7b",
          6234 => x"38",
          6235 => x"8c",
          6236 => x"39",
          6237 => x"b0",
          6238 => x"39",
          6239 => x"56",
          6240 => x"da",
          6241 => x"53",
          6242 => x"52",
          6243 => x"b0",
          6244 => x"f1",
          6245 => x"39",
          6246 => x"52",
          6247 => x"b0",
          6248 => x"f1",
          6249 => x"39",
          6250 => x"da",
          6251 => x"53",
          6252 => x"52",
          6253 => x"b0",
          6254 => x"f0",
          6255 => x"39",
          6256 => x"53",
          6257 => x"52",
          6258 => x"b0",
          6259 => x"f0",
          6260 => x"db",
          6261 => x"de",
          6262 => x"56",
          6263 => x"46",
          6264 => x"80",
          6265 => x"80",
          6266 => x"80",
          6267 => x"ff",
          6268 => x"e7",
          6269 => x"de",
          6270 => x"de",
          6271 => x"70",
          6272 => x"07",
          6273 => x"5b",
          6274 => x"83",
          6275 => x"78",
          6276 => x"38",
          6277 => x"81",
          6278 => x"59",
          6279 => x"38",
          6280 => x"7d",
          6281 => x"59",
          6282 => x"7d",
          6283 => x"81",
          6284 => x"38",
          6285 => x"51",
          6286 => x"3f",
          6287 => x"fc",
          6288 => x"0b",
          6289 => x"34",
          6290 => x"8c",
          6291 => x"55",
          6292 => x"52",
          6293 => x"ce",
          6294 => x"de",
          6295 => x"2b",
          6296 => x"53",
          6297 => x"52",
          6298 => x"ce",
          6299 => x"81",
          6300 => x"07",
          6301 => x"c0",
          6302 => x"08",
          6303 => x"84",
          6304 => x"51",
          6305 => x"3f",
          6306 => x"08",
          6307 => x"08",
          6308 => x"84",
          6309 => x"51",
          6310 => x"3f",
          6311 => x"c0",
          6312 => x"0c",
          6313 => x"0b",
          6314 => x"84",
          6315 => x"83",
          6316 => x"94",
          6317 => x"ba",
          6318 => x"d0",
          6319 => x"0b",
          6320 => x"0c",
          6321 => x"3f",
          6322 => x"3f",
          6323 => x"51",
          6324 => x"3f",
          6325 => x"51",
          6326 => x"3f",
          6327 => x"51",
          6328 => x"3f",
          6329 => x"bb",
          6330 => x"3f",
          6331 => x"00",
          6332 => x"ff",
          6333 => x"ff",
          6334 => x"00",
          6335 => x"ff",
          6336 => x"16",
          6337 => x"16",
          6338 => x"16",
          6339 => x"16",
          6340 => x"16",
          6341 => x"53",
          6342 => x"53",
          6343 => x"53",
          6344 => x"53",
          6345 => x"53",
          6346 => x"53",
          6347 => x"53",
          6348 => x"53",
          6349 => x"53",
          6350 => x"53",
          6351 => x"53",
          6352 => x"53",
          6353 => x"53",
          6354 => x"53",
          6355 => x"53",
          6356 => x"53",
          6357 => x"53",
          6358 => x"53",
          6359 => x"53",
          6360 => x"53",
          6361 => x"2f",
          6362 => x"25",
          6363 => x"64",
          6364 => x"3a",
          6365 => x"25",
          6366 => x"0a",
          6367 => x"43",
          6368 => x"6e",
          6369 => x"75",
          6370 => x"69",
          6371 => x"00",
          6372 => x"66",
          6373 => x"20",
          6374 => x"20",
          6375 => x"66",
          6376 => x"00",
          6377 => x"44",
          6378 => x"63",
          6379 => x"69",
          6380 => x"65",
          6381 => x"74",
          6382 => x"0a",
          6383 => x"20",
          6384 => x"20",
          6385 => x"41",
          6386 => x"28",
          6387 => x"58",
          6388 => x"38",
          6389 => x"0a",
          6390 => x"20",
          6391 => x"52",
          6392 => x"20",
          6393 => x"28",
          6394 => x"58",
          6395 => x"38",
          6396 => x"0a",
          6397 => x"20",
          6398 => x"53",
          6399 => x"52",
          6400 => x"28",
          6401 => x"58",
          6402 => x"38",
          6403 => x"0a",
          6404 => x"20",
          6405 => x"41",
          6406 => x"20",
          6407 => x"28",
          6408 => x"58",
          6409 => x"38",
          6410 => x"0a",
          6411 => x"20",
          6412 => x"4d",
          6413 => x"20",
          6414 => x"28",
          6415 => x"58",
          6416 => x"38",
          6417 => x"0a",
          6418 => x"20",
          6419 => x"20",
          6420 => x"44",
          6421 => x"28",
          6422 => x"69",
          6423 => x"20",
          6424 => x"32",
          6425 => x"0a",
          6426 => x"20",
          6427 => x"4d",
          6428 => x"20",
          6429 => x"28",
          6430 => x"65",
          6431 => x"20",
          6432 => x"32",
          6433 => x"0a",
          6434 => x"20",
          6435 => x"54",
          6436 => x"54",
          6437 => x"28",
          6438 => x"6e",
          6439 => x"73",
          6440 => x"32",
          6441 => x"0a",
          6442 => x"20",
          6443 => x"53",
          6444 => x"4e",
          6445 => x"55",
          6446 => x"00",
          6447 => x"20",
          6448 => x"20",
          6449 => x"0a",
          6450 => x"20",
          6451 => x"43",
          6452 => x"00",
          6453 => x"20",
          6454 => x"32",
          6455 => x"00",
          6456 => x"20",
          6457 => x"49",
          6458 => x"00",
          6459 => x"64",
          6460 => x"73",
          6461 => x"0a",
          6462 => x"20",
          6463 => x"55",
          6464 => x"73",
          6465 => x"56",
          6466 => x"6f",
          6467 => x"64",
          6468 => x"73",
          6469 => x"20",
          6470 => x"58",
          6471 => x"00",
          6472 => x"20",
          6473 => x"55",
          6474 => x"6d",
          6475 => x"20",
          6476 => x"72",
          6477 => x"64",
          6478 => x"73",
          6479 => x"20",
          6480 => x"58",
          6481 => x"00",
          6482 => x"20",
          6483 => x"61",
          6484 => x"53",
          6485 => x"74",
          6486 => x"64",
          6487 => x"73",
          6488 => x"20",
          6489 => x"20",
          6490 => x"58",
          6491 => x"00",
          6492 => x"73",
          6493 => x"00",
          6494 => x"20",
          6495 => x"55",
          6496 => x"20",
          6497 => x"20",
          6498 => x"20",
          6499 => x"20",
          6500 => x"20",
          6501 => x"20",
          6502 => x"58",
          6503 => x"00",
          6504 => x"20",
          6505 => x"73",
          6506 => x"20",
          6507 => x"63",
          6508 => x"72",
          6509 => x"20",
          6510 => x"20",
          6511 => x"20",
          6512 => x"25",
          6513 => x"4d",
          6514 => x"00",
          6515 => x"20",
          6516 => x"52",
          6517 => x"43",
          6518 => x"6b",
          6519 => x"65",
          6520 => x"20",
          6521 => x"20",
          6522 => x"20",
          6523 => x"25",
          6524 => x"4d",
          6525 => x"00",
          6526 => x"20",
          6527 => x"73",
          6528 => x"6e",
          6529 => x"44",
          6530 => x"20",
          6531 => x"63",
          6532 => x"72",
          6533 => x"20",
          6534 => x"25",
          6535 => x"4d",
          6536 => x"00",
          6537 => x"61",
          6538 => x"00",
          6539 => x"64",
          6540 => x"00",
          6541 => x"65",
          6542 => x"00",
          6543 => x"4f",
          6544 => x"4f",
          6545 => x"00",
          6546 => x"6b",
          6547 => x"6e",
          6548 => x"00",
          6549 => x"2b",
          6550 => x"3c",
          6551 => x"5b",
          6552 => x"00",
          6553 => x"54",
          6554 => x"54",
          6555 => x"00",
          6556 => x"90",
          6557 => x"4f",
          6558 => x"30",
          6559 => x"20",
          6560 => x"45",
          6561 => x"20",
          6562 => x"33",
          6563 => x"20",
          6564 => x"20",
          6565 => x"45",
          6566 => x"20",
          6567 => x"20",
          6568 => x"20",
          6569 => x"66",
          6570 => x"00",
          6571 => x"00",
          6572 => x"00",
          6573 => x"45",
          6574 => x"8f",
          6575 => x"45",
          6576 => x"8e",
          6577 => x"92",
          6578 => x"55",
          6579 => x"9a",
          6580 => x"9e",
          6581 => x"4f",
          6582 => x"a6",
          6583 => x"aa",
          6584 => x"ae",
          6585 => x"b2",
          6586 => x"b6",
          6587 => x"ba",
          6588 => x"be",
          6589 => x"c2",
          6590 => x"c6",
          6591 => x"ca",
          6592 => x"ce",
          6593 => x"d2",
          6594 => x"d6",
          6595 => x"da",
          6596 => x"de",
          6597 => x"e2",
          6598 => x"e6",
          6599 => x"ea",
          6600 => x"ee",
          6601 => x"f2",
          6602 => x"f6",
          6603 => x"fa",
          6604 => x"fe",
          6605 => x"2c",
          6606 => x"5d",
          6607 => x"2a",
          6608 => x"3f",
          6609 => x"00",
          6610 => x"00",
          6611 => x"00",
          6612 => x"02",
          6613 => x"00",
          6614 => x"00",
          6615 => x"00",
          6616 => x"00",
          6617 => x"00",
          6618 => x"6e",
          6619 => x"00",
          6620 => x"6f",
          6621 => x"00",
          6622 => x"6e",
          6623 => x"00",
          6624 => x"6f",
          6625 => x"00",
          6626 => x"78",
          6627 => x"00",
          6628 => x"6c",
          6629 => x"00",
          6630 => x"75",
          6631 => x"00",
          6632 => x"72",
          6633 => x"00",
          6634 => x"62",
          6635 => x"68",
          6636 => x"77",
          6637 => x"64",
          6638 => x"65",
          6639 => x"64",
          6640 => x"65",
          6641 => x"6c",
          6642 => x"00",
          6643 => x"70",
          6644 => x"73",
          6645 => x"74",
          6646 => x"73",
          6647 => x"00",
          6648 => x"66",
          6649 => x"00",
          6650 => x"73",
          6651 => x"00",
          6652 => x"73",
          6653 => x"72",
          6654 => x"0a",
          6655 => x"74",
          6656 => x"61",
          6657 => x"72",
          6658 => x"2e",
          6659 => x"00",
          6660 => x"73",
          6661 => x"6f",
          6662 => x"65",
          6663 => x"2e",
          6664 => x"00",
          6665 => x"20",
          6666 => x"65",
          6667 => x"75",
          6668 => x"0a",
          6669 => x"20",
          6670 => x"68",
          6671 => x"75",
          6672 => x"0a",
          6673 => x"76",
          6674 => x"64",
          6675 => x"6c",
          6676 => x"6d",
          6677 => x"00",
          6678 => x"63",
          6679 => x"20",
          6680 => x"69",
          6681 => x"0a",
          6682 => x"6c",
          6683 => x"6c",
          6684 => x"64",
          6685 => x"78",
          6686 => x"73",
          6687 => x"00",
          6688 => x"6c",
          6689 => x"61",
          6690 => x"65",
          6691 => x"76",
          6692 => x"64",
          6693 => x"00",
          6694 => x"20",
          6695 => x"77",
          6696 => x"65",
          6697 => x"6f",
          6698 => x"74",
          6699 => x"0a",
          6700 => x"69",
          6701 => x"6e",
          6702 => x"65",
          6703 => x"73",
          6704 => x"76",
          6705 => x"64",
          6706 => x"00",
          6707 => x"73",
          6708 => x"6f",
          6709 => x"6e",
          6710 => x"65",
          6711 => x"00",
          6712 => x"20",
          6713 => x"70",
          6714 => x"62",
          6715 => x"66",
          6716 => x"73",
          6717 => x"65",
          6718 => x"6f",
          6719 => x"20",
          6720 => x"64",
          6721 => x"2e",
          6722 => x"00",
          6723 => x"72",
          6724 => x"20",
          6725 => x"72",
          6726 => x"2e",
          6727 => x"00",
          6728 => x"6d",
          6729 => x"74",
          6730 => x"70",
          6731 => x"74",
          6732 => x"20",
          6733 => x"63",
          6734 => x"65",
          6735 => x"00",
          6736 => x"6c",
          6737 => x"73",
          6738 => x"63",
          6739 => x"2e",
          6740 => x"00",
          6741 => x"73",
          6742 => x"69",
          6743 => x"6e",
          6744 => x"65",
          6745 => x"79",
          6746 => x"00",
          6747 => x"6f",
          6748 => x"6e",
          6749 => x"70",
          6750 => x"66",
          6751 => x"73",
          6752 => x"00",
          6753 => x"72",
          6754 => x"74",
          6755 => x"20",
          6756 => x"6f",
          6757 => x"63",
          6758 => x"00",
          6759 => x"63",
          6760 => x"73",
          6761 => x"00",
          6762 => x"6b",
          6763 => x"6e",
          6764 => x"72",
          6765 => x"0a",
          6766 => x"6c",
          6767 => x"79",
          6768 => x"20",
          6769 => x"61",
          6770 => x"6c",
          6771 => x"79",
          6772 => x"2f",
          6773 => x"2e",
          6774 => x"00",
          6775 => x"38",
          6776 => x"00",
          6777 => x"20",
          6778 => x"34",
          6779 => x"00",
          6780 => x"20",
          6781 => x"20",
          6782 => x"00",
          6783 => x"32",
          6784 => x"00",
          6785 => x"00",
          6786 => x"00",
          6787 => x"0a",
          6788 => x"61",
          6789 => x"00",
          6790 => x"55",
          6791 => x"00",
          6792 => x"2a",
          6793 => x"20",
          6794 => x"00",
          6795 => x"2f",
          6796 => x"32",
          6797 => x"00",
          6798 => x"2e",
          6799 => x"00",
          6800 => x"50",
          6801 => x"72",
          6802 => x"25",
          6803 => x"29",
          6804 => x"20",
          6805 => x"2a",
          6806 => x"00",
          6807 => x"55",
          6808 => x"49",
          6809 => x"72",
          6810 => x"74",
          6811 => x"6e",
          6812 => x"72",
          6813 => x"00",
          6814 => x"6d",
          6815 => x"69",
          6816 => x"72",
          6817 => x"74",
          6818 => x"00",
          6819 => x"32",
          6820 => x"74",
          6821 => x"75",
          6822 => x"00",
          6823 => x"43",
          6824 => x"52",
          6825 => x"6e",
          6826 => x"72",
          6827 => x"0a",
          6828 => x"43",
          6829 => x"57",
          6830 => x"6e",
          6831 => x"72",
          6832 => x"0a",
          6833 => x"52",
          6834 => x"52",
          6835 => x"6e",
          6836 => x"72",
          6837 => x"0a",
          6838 => x"52",
          6839 => x"54",
          6840 => x"6e",
          6841 => x"72",
          6842 => x"0a",
          6843 => x"52",
          6844 => x"52",
          6845 => x"6e",
          6846 => x"72",
          6847 => x"0a",
          6848 => x"52",
          6849 => x"54",
          6850 => x"6e",
          6851 => x"72",
          6852 => x"0a",
          6853 => x"74",
          6854 => x"67",
          6855 => x"20",
          6856 => x"65",
          6857 => x"2e",
          6858 => x"00",
          6859 => x"61",
          6860 => x"6e",
          6861 => x"69",
          6862 => x"2e",
          6863 => x"00",
          6864 => x"74",
          6865 => x"65",
          6866 => x"61",
          6867 => x"00",
          6868 => x"00",
          6869 => x"69",
          6870 => x"20",
          6871 => x"69",
          6872 => x"69",
          6873 => x"73",
          6874 => x"64",
          6875 => x"72",
          6876 => x"2c",
          6877 => x"65",
          6878 => x"20",
          6879 => x"74",
          6880 => x"6e",
          6881 => x"6c",
          6882 => x"00",
          6883 => x"00",
          6884 => x"64",
          6885 => x"73",
          6886 => x"64",
          6887 => x"00",
          6888 => x"69",
          6889 => x"6c",
          6890 => x"64",
          6891 => x"00",
          6892 => x"69",
          6893 => x"20",
          6894 => x"69",
          6895 => x"69",
          6896 => x"73",
          6897 => x"00",
          6898 => x"3d",
          6899 => x"00",
          6900 => x"3a",
          6901 => x"65",
          6902 => x"6e",
          6903 => x"2e",
          6904 => x"00",
          6905 => x"6d",
          6906 => x"65",
          6907 => x"79",
          6908 => x"00",
          6909 => x"6f",
          6910 => x"65",
          6911 => x"0a",
          6912 => x"38",
          6913 => x"30",
          6914 => x"00",
          6915 => x"3f",
          6916 => x"00",
          6917 => x"38",
          6918 => x"30",
          6919 => x"00",
          6920 => x"38",
          6921 => x"30",
          6922 => x"00",
          6923 => x"61",
          6924 => x"69",
          6925 => x"2e",
          6926 => x"00",
          6927 => x"38",
          6928 => x"3e",
          6929 => x"6c",
          6930 => x"00",
          6931 => x"73",
          6932 => x"69",
          6933 => x"69",
          6934 => x"72",
          6935 => x"74",
          6936 => x"00",
          6937 => x"61",
          6938 => x"6e",
          6939 => x"6e",
          6940 => x"72",
          6941 => x"73",
          6942 => x"00",
          6943 => x"73",
          6944 => x"65",
          6945 => x"61",
          6946 => x"66",
          6947 => x"0a",
          6948 => x"61",
          6949 => x"6e",
          6950 => x"61",
          6951 => x"66",
          6952 => x"0a",
          6953 => x"65",
          6954 => x"69",
          6955 => x"63",
          6956 => x"20",
          6957 => x"30",
          6958 => x"2e",
          6959 => x"00",
          6960 => x"6c",
          6961 => x"67",
          6962 => x"64",
          6963 => x"20",
          6964 => x"78",
          6965 => x"2e",
          6966 => x"00",
          6967 => x"6c",
          6968 => x"65",
          6969 => x"6e",
          6970 => x"63",
          6971 => x"20",
          6972 => x"29",
          6973 => x"00",
          6974 => x"73",
          6975 => x"74",
          6976 => x"20",
          6977 => x"6c",
          6978 => x"74",
          6979 => x"2e",
          6980 => x"00",
          6981 => x"6c",
          6982 => x"65",
          6983 => x"74",
          6984 => x"2e",
          6985 => x"00",
          6986 => x"55",
          6987 => x"6e",
          6988 => x"3a",
          6989 => x"5c",
          6990 => x"25",
          6991 => x"00",
          6992 => x"3a",
          6993 => x"5c",
          6994 => x"00",
          6995 => x"3a",
          6996 => x"00",
          6997 => x"64",
          6998 => x"6d",
          6999 => x"64",
          7000 => x"00",
          7001 => x"6e",
          7002 => x"67",
          7003 => x"0a",
          7004 => x"61",
          7005 => x"6e",
          7006 => x"6e",
          7007 => x"72",
          7008 => x"73",
          7009 => x"0a",
          7010 => x"00",
          7011 => x"00",
          7012 => x"7f",
          7013 => x"00",
          7014 => x"7f",
          7015 => x"00",
          7016 => x"7f",
          7017 => x"00",
          7018 => x"00",
          7019 => x"00",
          7020 => x"ff",
          7021 => x"00",
          7022 => x"00",
          7023 => x"78",
          7024 => x"00",
          7025 => x"e1",
          7026 => x"e1",
          7027 => x"e1",
          7028 => x"00",
          7029 => x"01",
          7030 => x"01",
          7031 => x"10",
          7032 => x"00",
          7033 => x"00",
          7034 => x"00",
          7035 => x"00",
          7036 => x"67",
          7037 => x"01",
          7038 => x"00",
          7039 => x"00",
          7040 => x"67",
          7041 => x"01",
          7042 => x"00",
          7043 => x"00",
          7044 => x"67",
          7045 => x"03",
          7046 => x"00",
          7047 => x"00",
          7048 => x"67",
          7049 => x"03",
          7050 => x"00",
          7051 => x"00",
          7052 => x"67",
          7053 => x"03",
          7054 => x"00",
          7055 => x"00",
          7056 => x"67",
          7057 => x"04",
          7058 => x"00",
          7059 => x"00",
          7060 => x"67",
          7061 => x"04",
          7062 => x"00",
          7063 => x"00",
          7064 => x"67",
          7065 => x"04",
          7066 => x"00",
          7067 => x"00",
          7068 => x"67",
          7069 => x"04",
          7070 => x"00",
          7071 => x"00",
          7072 => x"67",
          7073 => x"04",
          7074 => x"00",
          7075 => x"00",
          7076 => x"67",
          7077 => x"04",
          7078 => x"00",
          7079 => x"00",
          7080 => x"67",
          7081 => x"05",
          7082 => x"00",
          7083 => x"00",
          7084 => x"67",
          7085 => x"05",
          7086 => x"00",
          7087 => x"00",
          7088 => x"67",
          7089 => x"05",
          7090 => x"00",
          7091 => x"00",
          7092 => x"67",
          7093 => x"05",
          7094 => x"00",
          7095 => x"00",
          7096 => x"67",
          7097 => x"07",
          7098 => x"00",
          7099 => x"00",
          7100 => x"67",
          7101 => x"07",
          7102 => x"00",
          7103 => x"00",
          7104 => x"67",
          7105 => x"08",
          7106 => x"00",
          7107 => x"00",
          7108 => x"67",
          7109 => x"08",
          7110 => x"00",
          7111 => x"00",
          7112 => x"67",
          7113 => x"08",
          7114 => x"00",
          7115 => x"00",
          7116 => x"67",
          7117 => x"08",
          7118 => x"00",
          7119 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"a4",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8c",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"81",
           386 => x"a0",
           387 => x"de",
           388 => x"80",
           389 => x"de",
           390 => x"e2",
           391 => x"cc",
           392 => x"90",
           393 => x"cc",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"81",
           399 => x"82",
           400 => x"81",
           401 => x"b4",
           402 => x"de",
           403 => x"80",
           404 => x"de",
           405 => x"fb",
           406 => x"cc",
           407 => x"90",
           408 => x"cc",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"81",
           414 => x"82",
           415 => x"81",
           416 => x"b8",
           417 => x"de",
           418 => x"80",
           419 => x"de",
           420 => x"a3",
           421 => x"cc",
           422 => x"90",
           423 => x"cc",
           424 => x"2d",
           425 => x"08",
           426 => x"04",
           427 => x"0c",
           428 => x"81",
           429 => x"82",
           430 => x"81",
           431 => x"a2",
           432 => x"de",
           433 => x"80",
           434 => x"de",
           435 => x"8c",
           436 => x"cc",
           437 => x"90",
           438 => x"cc",
           439 => x"2d",
           440 => x"08",
           441 => x"04",
           442 => x"0c",
           443 => x"81",
           444 => x"82",
           445 => x"81",
           446 => x"9e",
           447 => x"de",
           448 => x"80",
           449 => x"de",
           450 => x"ea",
           451 => x"de",
           452 => x"80",
           453 => x"de",
           454 => x"f7",
           455 => x"de",
           456 => x"80",
           457 => x"de",
           458 => x"ef",
           459 => x"de",
           460 => x"80",
           461 => x"de",
           462 => x"f2",
           463 => x"de",
           464 => x"80",
           465 => x"de",
           466 => x"fc",
           467 => x"de",
           468 => x"80",
           469 => x"de",
           470 => x"85",
           471 => x"de",
           472 => x"80",
           473 => x"de",
           474 => x"f6",
           475 => x"de",
           476 => x"80",
           477 => x"de",
           478 => x"ff",
           479 => x"de",
           480 => x"80",
           481 => x"de",
           482 => x"80",
           483 => x"de",
           484 => x"80",
           485 => x"de",
           486 => x"81",
           487 => x"de",
           488 => x"80",
           489 => x"de",
           490 => x"89",
           491 => x"de",
           492 => x"80",
           493 => x"de",
           494 => x"86",
           495 => x"de",
           496 => x"80",
           497 => x"de",
           498 => x"8b",
           499 => x"de",
           500 => x"80",
           501 => x"de",
           502 => x"82",
           503 => x"de",
           504 => x"80",
           505 => x"de",
           506 => x"8e",
           507 => x"de",
           508 => x"80",
           509 => x"de",
           510 => x"8f",
           511 => x"de",
           512 => x"80",
           513 => x"de",
           514 => x"f8",
           515 => x"de",
           516 => x"80",
           517 => x"de",
           518 => x"f7",
           519 => x"de",
           520 => x"80",
           521 => x"de",
           522 => x"f9",
           523 => x"de",
           524 => x"80",
           525 => x"de",
           526 => x"82",
           527 => x"de",
           528 => x"80",
           529 => x"de",
           530 => x"90",
           531 => x"de",
           532 => x"80",
           533 => x"de",
           534 => x"92",
           535 => x"de",
           536 => x"80",
           537 => x"de",
           538 => x"96",
           539 => x"de",
           540 => x"80",
           541 => x"de",
           542 => x"e9",
           543 => x"de",
           544 => x"80",
           545 => x"de",
           546 => x"99",
           547 => x"de",
           548 => x"80",
           549 => x"de",
           550 => x"99",
           551 => x"cc",
           552 => x"90",
           553 => x"cc",
           554 => x"2d",
           555 => x"08",
           556 => x"04",
           557 => x"0c",
           558 => x"81",
           559 => x"82",
           560 => x"81",
           561 => x"9b",
           562 => x"de",
           563 => x"80",
           564 => x"de",
           565 => x"b3",
           566 => x"cc",
           567 => x"90",
           568 => x"cc",
           569 => x"2d",
           570 => x"08",
           571 => x"04",
           572 => x"0c",
           573 => x"2d",
           574 => x"08",
           575 => x"04",
           576 => x"10",
           577 => x"10",
           578 => x"10",
           579 => x"10",
           580 => x"10",
           581 => x"10",
           582 => x"10",
           583 => x"10",
           584 => x"04",
           585 => x"81",
           586 => x"83",
           587 => x"05",
           588 => x"10",
           589 => x"72",
           590 => x"51",
           591 => x"72",
           592 => x"06",
           593 => x"72",
           594 => x"10",
           595 => x"10",
           596 => x"ed",
           597 => x"53",
           598 => x"de",
           599 => x"f5",
           600 => x"38",
           601 => x"84",
           602 => x"0b",
           603 => x"db",
           604 => x"51",
           605 => x"04",
           606 => x"cc",
           607 => x"de",
           608 => x"3d",
           609 => x"81",
           610 => x"8c",
           611 => x"81",
           612 => x"88",
           613 => x"83",
           614 => x"de",
           615 => x"81",
           616 => x"54",
           617 => x"81",
           618 => x"04",
           619 => x"08",
           620 => x"cc",
           621 => x"0d",
           622 => x"de",
           623 => x"05",
           624 => x"de",
           625 => x"05",
           626 => x"a1",
           627 => x"c0",
           628 => x"de",
           629 => x"85",
           630 => x"de",
           631 => x"81",
           632 => x"02",
           633 => x"0c",
           634 => x"80",
           635 => x"cc",
           636 => x"0c",
           637 => x"08",
           638 => x"80",
           639 => x"81",
           640 => x"88",
           641 => x"81",
           642 => x"88",
           643 => x"0b",
           644 => x"08",
           645 => x"81",
           646 => x"fc",
           647 => x"38",
           648 => x"de",
           649 => x"05",
           650 => x"cc",
           651 => x"08",
           652 => x"08",
           653 => x"81",
           654 => x"8c",
           655 => x"25",
           656 => x"de",
           657 => x"05",
           658 => x"de",
           659 => x"05",
           660 => x"81",
           661 => x"f0",
           662 => x"de",
           663 => x"05",
           664 => x"81",
           665 => x"cc",
           666 => x"0c",
           667 => x"08",
           668 => x"81",
           669 => x"fc",
           670 => x"53",
           671 => x"08",
           672 => x"52",
           673 => x"08",
           674 => x"51",
           675 => x"81",
           676 => x"70",
           677 => x"08",
           678 => x"54",
           679 => x"08",
           680 => x"80",
           681 => x"81",
           682 => x"f8",
           683 => x"81",
           684 => x"f8",
           685 => x"de",
           686 => x"05",
           687 => x"de",
           688 => x"89",
           689 => x"de",
           690 => x"81",
           691 => x"02",
           692 => x"0c",
           693 => x"80",
           694 => x"cc",
           695 => x"0c",
           696 => x"08",
           697 => x"80",
           698 => x"81",
           699 => x"88",
           700 => x"81",
           701 => x"88",
           702 => x"0b",
           703 => x"08",
           704 => x"81",
           705 => x"8c",
           706 => x"25",
           707 => x"de",
           708 => x"05",
           709 => x"de",
           710 => x"05",
           711 => x"81",
           712 => x"8c",
           713 => x"81",
           714 => x"88",
           715 => x"bd",
           716 => x"c0",
           717 => x"de",
           718 => x"05",
           719 => x"de",
           720 => x"05",
           721 => x"90",
           722 => x"cc",
           723 => x"08",
           724 => x"cc",
           725 => x"0c",
           726 => x"08",
           727 => x"70",
           728 => x"0c",
           729 => x"0d",
           730 => x"0c",
           731 => x"cc",
           732 => x"de",
           733 => x"3d",
           734 => x"81",
           735 => x"fc",
           736 => x"0b",
           737 => x"08",
           738 => x"81",
           739 => x"8c",
           740 => x"de",
           741 => x"05",
           742 => x"38",
           743 => x"08",
           744 => x"80",
           745 => x"80",
           746 => x"cc",
           747 => x"08",
           748 => x"81",
           749 => x"8c",
           750 => x"81",
           751 => x"8c",
           752 => x"de",
           753 => x"05",
           754 => x"de",
           755 => x"05",
           756 => x"39",
           757 => x"08",
           758 => x"80",
           759 => x"38",
           760 => x"08",
           761 => x"81",
           762 => x"88",
           763 => x"ad",
           764 => x"cc",
           765 => x"08",
           766 => x"08",
           767 => x"31",
           768 => x"08",
           769 => x"81",
           770 => x"f8",
           771 => x"de",
           772 => x"05",
           773 => x"de",
           774 => x"05",
           775 => x"cc",
           776 => x"08",
           777 => x"de",
           778 => x"05",
           779 => x"cc",
           780 => x"08",
           781 => x"de",
           782 => x"05",
           783 => x"39",
           784 => x"08",
           785 => x"80",
           786 => x"81",
           787 => x"88",
           788 => x"81",
           789 => x"f4",
           790 => x"91",
           791 => x"cc",
           792 => x"08",
           793 => x"cc",
           794 => x"0c",
           795 => x"cc",
           796 => x"08",
           797 => x"0c",
           798 => x"81",
           799 => x"04",
           800 => x"76",
           801 => x"8c",
           802 => x"33",
           803 => x"55",
           804 => x"8a",
           805 => x"06",
           806 => x"2e",
           807 => x"12",
           808 => x"2e",
           809 => x"73",
           810 => x"55",
           811 => x"52",
           812 => x"09",
           813 => x"38",
           814 => x"c0",
           815 => x"0d",
           816 => x"88",
           817 => x"70",
           818 => x"07",
           819 => x"8f",
           820 => x"38",
           821 => x"84",
           822 => x"72",
           823 => x"05",
           824 => x"71",
           825 => x"53",
           826 => x"70",
           827 => x"0c",
           828 => x"71",
           829 => x"38",
           830 => x"90",
           831 => x"70",
           832 => x"0c",
           833 => x"71",
           834 => x"38",
           835 => x"8e",
           836 => x"0d",
           837 => x"72",
           838 => x"53",
           839 => x"93",
           840 => x"73",
           841 => x"54",
           842 => x"2e",
           843 => x"73",
           844 => x"71",
           845 => x"ff",
           846 => x"70",
           847 => x"38",
           848 => x"70",
           849 => x"81",
           850 => x"81",
           851 => x"71",
           852 => x"ff",
           853 => x"54",
           854 => x"38",
           855 => x"73",
           856 => x"75",
           857 => x"71",
           858 => x"de",
           859 => x"52",
           860 => x"04",
           861 => x"f7",
           862 => x"14",
           863 => x"84",
           864 => x"06",
           865 => x"70",
           866 => x"14",
           867 => x"08",
           868 => x"71",
           869 => x"dc",
           870 => x"54",
           871 => x"39",
           872 => x"de",
           873 => x"3d",
           874 => x"3d",
           875 => x"83",
           876 => x"2b",
           877 => x"3f",
           878 => x"08",
           879 => x"72",
           880 => x"54",
           881 => x"25",
           882 => x"81",
           883 => x"84",
           884 => x"fb",
           885 => x"70",
           886 => x"53",
           887 => x"2e",
           888 => x"71",
           889 => x"a0",
           890 => x"06",
           891 => x"12",
           892 => x"71",
           893 => x"81",
           894 => x"73",
           895 => x"ff",
           896 => x"55",
           897 => x"83",
           898 => x"70",
           899 => x"38",
           900 => x"73",
           901 => x"51",
           902 => x"09",
           903 => x"38",
           904 => x"81",
           905 => x"72",
           906 => x"51",
           907 => x"c0",
           908 => x"0d",
           909 => x"0d",
           910 => x"08",
           911 => x"38",
           912 => x"05",
           913 => x"9b",
           914 => x"de",
           915 => x"38",
           916 => x"39",
           917 => x"81",
           918 => x"86",
           919 => x"fc",
           920 => x"82",
           921 => x"05",
           922 => x"52",
           923 => x"81",
           924 => x"13",
           925 => x"51",
           926 => x"9e",
           927 => x"38",
           928 => x"51",
           929 => x"97",
           930 => x"38",
           931 => x"51",
           932 => x"bb",
           933 => x"38",
           934 => x"51",
           935 => x"bb",
           936 => x"38",
           937 => x"55",
           938 => x"87",
           939 => x"d9",
           940 => x"22",
           941 => x"73",
           942 => x"80",
           943 => x"0b",
           944 => x"9c",
           945 => x"87",
           946 => x"0c",
           947 => x"87",
           948 => x"0c",
           949 => x"87",
           950 => x"0c",
           951 => x"87",
           952 => x"0c",
           953 => x"87",
           954 => x"0c",
           955 => x"87",
           956 => x"0c",
           957 => x"98",
           958 => x"87",
           959 => x"0c",
           960 => x"c0",
           961 => x"80",
           962 => x"de",
           963 => x"3d",
           964 => x"3d",
           965 => x"87",
           966 => x"5d",
           967 => x"87",
           968 => x"08",
           969 => x"23",
           970 => x"b8",
           971 => x"82",
           972 => x"c0",
           973 => x"5a",
           974 => x"34",
           975 => x"b0",
           976 => x"84",
           977 => x"c0",
           978 => x"5a",
           979 => x"34",
           980 => x"a8",
           981 => x"86",
           982 => x"c0",
           983 => x"5c",
           984 => x"23",
           985 => x"a0",
           986 => x"8a",
           987 => x"7d",
           988 => x"ff",
           989 => x"7b",
           990 => x"06",
           991 => x"33",
           992 => x"33",
           993 => x"33",
           994 => x"33",
           995 => x"33",
           996 => x"ff",
           997 => x"81",
           998 => x"95",
           999 => x"3d",
          1000 => x"3d",
          1001 => x"05",
          1002 => x"70",
          1003 => x"52",
          1004 => x"0b",
          1005 => x"34",
          1006 => x"04",
          1007 => x"77",
          1008 => x"db",
          1009 => x"81",
          1010 => x"55",
          1011 => x"94",
          1012 => x"80",
          1013 => x"87",
          1014 => x"51",
          1015 => x"96",
          1016 => x"06",
          1017 => x"70",
          1018 => x"38",
          1019 => x"70",
          1020 => x"51",
          1021 => x"72",
          1022 => x"81",
          1023 => x"70",
          1024 => x"38",
          1025 => x"70",
          1026 => x"51",
          1027 => x"38",
          1028 => x"06",
          1029 => x"94",
          1030 => x"80",
          1031 => x"87",
          1032 => x"52",
          1033 => x"75",
          1034 => x"0c",
          1035 => x"04",
          1036 => x"02",
          1037 => x"0b",
          1038 => x"88",
          1039 => x"ff",
          1040 => x"56",
          1041 => x"84",
          1042 => x"2e",
          1043 => x"c0",
          1044 => x"70",
          1045 => x"2a",
          1046 => x"53",
          1047 => x"80",
          1048 => x"71",
          1049 => x"81",
          1050 => x"70",
          1051 => x"81",
          1052 => x"06",
          1053 => x"80",
          1054 => x"71",
          1055 => x"81",
          1056 => x"70",
          1057 => x"73",
          1058 => x"51",
          1059 => x"80",
          1060 => x"2e",
          1061 => x"c0",
          1062 => x"75",
          1063 => x"3d",
          1064 => x"3d",
          1065 => x"80",
          1066 => x"81",
          1067 => x"53",
          1068 => x"2e",
          1069 => x"71",
          1070 => x"81",
          1071 => x"81",
          1072 => x"70",
          1073 => x"59",
          1074 => x"87",
          1075 => x"51",
          1076 => x"86",
          1077 => x"94",
          1078 => x"08",
          1079 => x"70",
          1080 => x"54",
          1081 => x"2e",
          1082 => x"91",
          1083 => x"06",
          1084 => x"d7",
          1085 => x"32",
          1086 => x"51",
          1087 => x"2e",
          1088 => x"93",
          1089 => x"06",
          1090 => x"ff",
          1091 => x"81",
          1092 => x"87",
          1093 => x"52",
          1094 => x"86",
          1095 => x"94",
          1096 => x"72",
          1097 => x"74",
          1098 => x"ff",
          1099 => x"57",
          1100 => x"38",
          1101 => x"c0",
          1102 => x"0d",
          1103 => x"0d",
          1104 => x"db",
          1105 => x"81",
          1106 => x"52",
          1107 => x"84",
          1108 => x"2e",
          1109 => x"c0",
          1110 => x"70",
          1111 => x"2a",
          1112 => x"51",
          1113 => x"80",
          1114 => x"71",
          1115 => x"51",
          1116 => x"80",
          1117 => x"2e",
          1118 => x"c0",
          1119 => x"71",
          1120 => x"ff",
          1121 => x"c0",
          1122 => x"3d",
          1123 => x"3d",
          1124 => x"81",
          1125 => x"70",
          1126 => x"52",
          1127 => x"94",
          1128 => x"80",
          1129 => x"87",
          1130 => x"52",
          1131 => x"82",
          1132 => x"06",
          1133 => x"ff",
          1134 => x"2e",
          1135 => x"81",
          1136 => x"87",
          1137 => x"52",
          1138 => x"86",
          1139 => x"94",
          1140 => x"08",
          1141 => x"70",
          1142 => x"53",
          1143 => x"de",
          1144 => x"3d",
          1145 => x"3d",
          1146 => x"9e",
          1147 => x"9c",
          1148 => x"51",
          1149 => x"2e",
          1150 => x"87",
          1151 => x"08",
          1152 => x"0c",
          1153 => x"a8",
          1154 => x"90",
          1155 => x"9e",
          1156 => x"db",
          1157 => x"c0",
          1158 => x"81",
          1159 => x"87",
          1160 => x"08",
          1161 => x"0c",
          1162 => x"a0",
          1163 => x"a0",
          1164 => x"9e",
          1165 => x"db",
          1166 => x"c0",
          1167 => x"81",
          1168 => x"87",
          1169 => x"08",
          1170 => x"0c",
          1171 => x"b8",
          1172 => x"b0",
          1173 => x"9e",
          1174 => x"db",
          1175 => x"c0",
          1176 => x"81",
          1177 => x"87",
          1178 => x"08",
          1179 => x"0c",
          1180 => x"80",
          1181 => x"81",
          1182 => x"87",
          1183 => x"08",
          1184 => x"0c",
          1185 => x"88",
          1186 => x"c8",
          1187 => x"9e",
          1188 => x"db",
          1189 => x"0b",
          1190 => x"34",
          1191 => x"c0",
          1192 => x"70",
          1193 => x"06",
          1194 => x"70",
          1195 => x"38",
          1196 => x"81",
          1197 => x"80",
          1198 => x"9e",
          1199 => x"88",
          1200 => x"51",
          1201 => x"80",
          1202 => x"81",
          1203 => x"db",
          1204 => x"0b",
          1205 => x"90",
          1206 => x"80",
          1207 => x"52",
          1208 => x"2e",
          1209 => x"52",
          1210 => x"d3",
          1211 => x"87",
          1212 => x"08",
          1213 => x"80",
          1214 => x"52",
          1215 => x"83",
          1216 => x"71",
          1217 => x"34",
          1218 => x"c0",
          1219 => x"70",
          1220 => x"06",
          1221 => x"70",
          1222 => x"38",
          1223 => x"81",
          1224 => x"80",
          1225 => x"9e",
          1226 => x"90",
          1227 => x"51",
          1228 => x"80",
          1229 => x"81",
          1230 => x"db",
          1231 => x"0b",
          1232 => x"90",
          1233 => x"80",
          1234 => x"52",
          1235 => x"2e",
          1236 => x"52",
          1237 => x"d7",
          1238 => x"87",
          1239 => x"08",
          1240 => x"80",
          1241 => x"52",
          1242 => x"83",
          1243 => x"71",
          1244 => x"34",
          1245 => x"c0",
          1246 => x"70",
          1247 => x"06",
          1248 => x"70",
          1249 => x"38",
          1250 => x"81",
          1251 => x"80",
          1252 => x"9e",
          1253 => x"80",
          1254 => x"51",
          1255 => x"80",
          1256 => x"81",
          1257 => x"db",
          1258 => x"0b",
          1259 => x"90",
          1260 => x"80",
          1261 => x"52",
          1262 => x"83",
          1263 => x"71",
          1264 => x"34",
          1265 => x"90",
          1266 => x"80",
          1267 => x"2a",
          1268 => x"70",
          1269 => x"34",
          1270 => x"c0",
          1271 => x"70",
          1272 => x"51",
          1273 => x"80",
          1274 => x"81",
          1275 => x"db",
          1276 => x"c0",
          1277 => x"70",
          1278 => x"70",
          1279 => x"51",
          1280 => x"db",
          1281 => x"0b",
          1282 => x"90",
          1283 => x"06",
          1284 => x"70",
          1285 => x"38",
          1286 => x"81",
          1287 => x"87",
          1288 => x"08",
          1289 => x"51",
          1290 => x"db",
          1291 => x"3d",
          1292 => x"3d",
          1293 => x"fc",
          1294 => x"3f",
          1295 => x"33",
          1296 => x"2e",
          1297 => x"c7",
          1298 => x"f5",
          1299 => x"a4",
          1300 => x"3f",
          1301 => x"33",
          1302 => x"2e",
          1303 => x"db",
          1304 => x"db",
          1305 => x"54",
          1306 => x"bc",
          1307 => x"3f",
          1308 => x"33",
          1309 => x"2e",
          1310 => x"db",
          1311 => x"db",
          1312 => x"54",
          1313 => x"d8",
          1314 => x"3f",
          1315 => x"33",
          1316 => x"2e",
          1317 => x"db",
          1318 => x"db",
          1319 => x"54",
          1320 => x"f4",
          1321 => x"3f",
          1322 => x"33",
          1323 => x"2e",
          1324 => x"db",
          1325 => x"db",
          1326 => x"54",
          1327 => x"90",
          1328 => x"3f",
          1329 => x"33",
          1330 => x"2e",
          1331 => x"db",
          1332 => x"db",
          1333 => x"54",
          1334 => x"ac",
          1335 => x"3f",
          1336 => x"33",
          1337 => x"2e",
          1338 => x"db",
          1339 => x"81",
          1340 => x"8a",
          1341 => x"db",
          1342 => x"73",
          1343 => x"38",
          1344 => x"33",
          1345 => x"e8",
          1346 => x"3f",
          1347 => x"33",
          1348 => x"2e",
          1349 => x"db",
          1350 => x"81",
          1351 => x"8a",
          1352 => x"db",
          1353 => x"73",
          1354 => x"38",
          1355 => x"51",
          1356 => x"81",
          1357 => x"54",
          1358 => x"88",
          1359 => x"bc",
          1360 => x"3f",
          1361 => x"33",
          1362 => x"2e",
          1363 => x"c9",
          1364 => x"ed",
          1365 => x"d9",
          1366 => x"80",
          1367 => x"81",
          1368 => x"83",
          1369 => x"db",
          1370 => x"73",
          1371 => x"38",
          1372 => x"51",
          1373 => x"81",
          1374 => x"83",
          1375 => x"db",
          1376 => x"81",
          1377 => x"89",
          1378 => x"db",
          1379 => x"81",
          1380 => x"89",
          1381 => x"db",
          1382 => x"81",
          1383 => x"89",
          1384 => x"ca",
          1385 => x"fa",
          1386 => x"c0",
          1387 => x"ca",
          1388 => x"f1",
          1389 => x"c4",
          1390 => x"84",
          1391 => x"51",
          1392 => x"81",
          1393 => x"bd",
          1394 => x"76",
          1395 => x"54",
          1396 => x"08",
          1397 => x"a0",
          1398 => x"3f",
          1399 => x"33",
          1400 => x"2e",
          1401 => x"db",
          1402 => x"bd",
          1403 => x"75",
          1404 => x"3f",
          1405 => x"08",
          1406 => x"29",
          1407 => x"54",
          1408 => x"c0",
          1409 => x"cb",
          1410 => x"99",
          1411 => x"d2",
          1412 => x"80",
          1413 => x"81",
          1414 => x"56",
          1415 => x"52",
          1416 => x"d5",
          1417 => x"c0",
          1418 => x"c0",
          1419 => x"31",
          1420 => x"de",
          1421 => x"81",
          1422 => x"87",
          1423 => x"d7",
          1424 => x"fd",
          1425 => x"0d",
          1426 => x"0d",
          1427 => x"33",
          1428 => x"71",
          1429 => x"38",
          1430 => x"81",
          1431 => x"52",
          1432 => x"81",
          1433 => x"9d",
          1434 => x"ac",
          1435 => x"81",
          1436 => x"91",
          1437 => x"bc",
          1438 => x"81",
          1439 => x"85",
          1440 => x"c8",
          1441 => x"3f",
          1442 => x"04",
          1443 => x"0c",
          1444 => x"87",
          1445 => x"0c",
          1446 => x"0d",
          1447 => x"84",
          1448 => x"52",
          1449 => x"70",
          1450 => x"81",
          1451 => x"72",
          1452 => x"0d",
          1453 => x"0d",
          1454 => x"84",
          1455 => x"db",
          1456 => x"80",
          1457 => x"09",
          1458 => x"e4",
          1459 => x"81",
          1460 => x"73",
          1461 => x"3d",
          1462 => x"db",
          1463 => x"c0",
          1464 => x"04",
          1465 => x"02",
          1466 => x"53",
          1467 => x"09",
          1468 => x"38",
          1469 => x"3f",
          1470 => x"08",
          1471 => x"2e",
          1472 => x"72",
          1473 => x"d8",
          1474 => x"81",
          1475 => x"8f",
          1476 => x"d0",
          1477 => x"80",
          1478 => x"72",
          1479 => x"84",
          1480 => x"fe",
          1481 => x"97",
          1482 => x"de",
          1483 => x"81",
          1484 => x"54",
          1485 => x"3f",
          1486 => x"d0",
          1487 => x"0d",
          1488 => x"0d",
          1489 => x"33",
          1490 => x"06",
          1491 => x"80",
          1492 => x"72",
          1493 => x"51",
          1494 => x"ff",
          1495 => x"39",
          1496 => x"04",
          1497 => x"77",
          1498 => x"08",
          1499 => x"d0",
          1500 => x"73",
          1501 => x"ff",
          1502 => x"71",
          1503 => x"38",
          1504 => x"06",
          1505 => x"54",
          1506 => x"e7",
          1507 => x"de",
          1508 => x"3d",
          1509 => x"3d",
          1510 => x"59",
          1511 => x"81",
          1512 => x"56",
          1513 => x"84",
          1514 => x"a5",
          1515 => x"06",
          1516 => x"80",
          1517 => x"81",
          1518 => x"58",
          1519 => x"b0",
          1520 => x"06",
          1521 => x"5a",
          1522 => x"ad",
          1523 => x"06",
          1524 => x"5a",
          1525 => x"05",
          1526 => x"75",
          1527 => x"81",
          1528 => x"77",
          1529 => x"08",
          1530 => x"05",
          1531 => x"5d",
          1532 => x"39",
          1533 => x"72",
          1534 => x"38",
          1535 => x"7b",
          1536 => x"05",
          1537 => x"70",
          1538 => x"33",
          1539 => x"39",
          1540 => x"32",
          1541 => x"72",
          1542 => x"78",
          1543 => x"70",
          1544 => x"07",
          1545 => x"07",
          1546 => x"51",
          1547 => x"80",
          1548 => x"79",
          1549 => x"70",
          1550 => x"33",
          1551 => x"80",
          1552 => x"38",
          1553 => x"e0",
          1554 => x"38",
          1555 => x"81",
          1556 => x"53",
          1557 => x"2e",
          1558 => x"73",
          1559 => x"a2",
          1560 => x"c3",
          1561 => x"38",
          1562 => x"24",
          1563 => x"80",
          1564 => x"8c",
          1565 => x"39",
          1566 => x"2e",
          1567 => x"81",
          1568 => x"80",
          1569 => x"80",
          1570 => x"d5",
          1571 => x"73",
          1572 => x"8e",
          1573 => x"39",
          1574 => x"2e",
          1575 => x"80",
          1576 => x"84",
          1577 => x"56",
          1578 => x"74",
          1579 => x"72",
          1580 => x"38",
          1581 => x"15",
          1582 => x"54",
          1583 => x"38",
          1584 => x"56",
          1585 => x"81",
          1586 => x"72",
          1587 => x"38",
          1588 => x"90",
          1589 => x"06",
          1590 => x"2e",
          1591 => x"51",
          1592 => x"74",
          1593 => x"53",
          1594 => x"fd",
          1595 => x"51",
          1596 => x"ef",
          1597 => x"19",
          1598 => x"53",
          1599 => x"39",
          1600 => x"39",
          1601 => x"39",
          1602 => x"39",
          1603 => x"39",
          1604 => x"d0",
          1605 => x"39",
          1606 => x"70",
          1607 => x"53",
          1608 => x"88",
          1609 => x"19",
          1610 => x"39",
          1611 => x"54",
          1612 => x"74",
          1613 => x"70",
          1614 => x"07",
          1615 => x"55",
          1616 => x"80",
          1617 => x"72",
          1618 => x"38",
          1619 => x"90",
          1620 => x"80",
          1621 => x"5e",
          1622 => x"74",
          1623 => x"3f",
          1624 => x"08",
          1625 => x"7c",
          1626 => x"54",
          1627 => x"81",
          1628 => x"55",
          1629 => x"92",
          1630 => x"53",
          1631 => x"2e",
          1632 => x"14",
          1633 => x"ff",
          1634 => x"14",
          1635 => x"70",
          1636 => x"34",
          1637 => x"30",
          1638 => x"9f",
          1639 => x"57",
          1640 => x"85",
          1641 => x"b1",
          1642 => x"2a",
          1643 => x"51",
          1644 => x"2e",
          1645 => x"3d",
          1646 => x"05",
          1647 => x"34",
          1648 => x"76",
          1649 => x"54",
          1650 => x"72",
          1651 => x"54",
          1652 => x"70",
          1653 => x"56",
          1654 => x"81",
          1655 => x"7b",
          1656 => x"73",
          1657 => x"3f",
          1658 => x"53",
          1659 => x"74",
          1660 => x"53",
          1661 => x"eb",
          1662 => x"77",
          1663 => x"53",
          1664 => x"14",
          1665 => x"54",
          1666 => x"3f",
          1667 => x"74",
          1668 => x"53",
          1669 => x"fb",
          1670 => x"51",
          1671 => x"ef",
          1672 => x"0d",
          1673 => x"0d",
          1674 => x"70",
          1675 => x"08",
          1676 => x"51",
          1677 => x"85",
          1678 => x"fe",
          1679 => x"81",
          1680 => x"85",
          1681 => x"52",
          1682 => x"ca",
          1683 => x"d8",
          1684 => x"73",
          1685 => x"81",
          1686 => x"84",
          1687 => x"fd",
          1688 => x"de",
          1689 => x"81",
          1690 => x"87",
          1691 => x"53",
          1692 => x"fa",
          1693 => x"81",
          1694 => x"85",
          1695 => x"fb",
          1696 => x"79",
          1697 => x"08",
          1698 => x"57",
          1699 => x"71",
          1700 => x"e0",
          1701 => x"d4",
          1702 => x"2d",
          1703 => x"08",
          1704 => x"53",
          1705 => x"80",
          1706 => x"8d",
          1707 => x"72",
          1708 => x"30",
          1709 => x"51",
          1710 => x"80",
          1711 => x"71",
          1712 => x"38",
          1713 => x"97",
          1714 => x"25",
          1715 => x"16",
          1716 => x"25",
          1717 => x"14",
          1718 => x"34",
          1719 => x"72",
          1720 => x"3f",
          1721 => x"73",
          1722 => x"72",
          1723 => x"f7",
          1724 => x"53",
          1725 => x"c0",
          1726 => x"0d",
          1727 => x"0d",
          1728 => x"08",
          1729 => x"d4",
          1730 => x"76",
          1731 => x"ef",
          1732 => x"de",
          1733 => x"3d",
          1734 => x"3d",
          1735 => x"5a",
          1736 => x"7a",
          1737 => x"08",
          1738 => x"53",
          1739 => x"09",
          1740 => x"38",
          1741 => x"0c",
          1742 => x"ad",
          1743 => x"06",
          1744 => x"76",
          1745 => x"0c",
          1746 => x"33",
          1747 => x"73",
          1748 => x"81",
          1749 => x"38",
          1750 => x"05",
          1751 => x"08",
          1752 => x"53",
          1753 => x"2e",
          1754 => x"57",
          1755 => x"2e",
          1756 => x"39",
          1757 => x"13",
          1758 => x"08",
          1759 => x"53",
          1760 => x"55",
          1761 => x"80",
          1762 => x"14",
          1763 => x"88",
          1764 => x"27",
          1765 => x"eb",
          1766 => x"53",
          1767 => x"89",
          1768 => x"38",
          1769 => x"55",
          1770 => x"8a",
          1771 => x"a0",
          1772 => x"c2",
          1773 => x"74",
          1774 => x"e0",
          1775 => x"ff",
          1776 => x"d0",
          1777 => x"ff",
          1778 => x"90",
          1779 => x"38",
          1780 => x"81",
          1781 => x"53",
          1782 => x"ca",
          1783 => x"27",
          1784 => x"77",
          1785 => x"08",
          1786 => x"0c",
          1787 => x"33",
          1788 => x"ff",
          1789 => x"80",
          1790 => x"74",
          1791 => x"79",
          1792 => x"74",
          1793 => x"0c",
          1794 => x"04",
          1795 => x"7a",
          1796 => x"80",
          1797 => x"58",
          1798 => x"33",
          1799 => x"a0",
          1800 => x"06",
          1801 => x"13",
          1802 => x"39",
          1803 => x"09",
          1804 => x"38",
          1805 => x"11",
          1806 => x"08",
          1807 => x"54",
          1808 => x"2e",
          1809 => x"80",
          1810 => x"08",
          1811 => x"0c",
          1812 => x"33",
          1813 => x"80",
          1814 => x"38",
          1815 => x"80",
          1816 => x"38",
          1817 => x"57",
          1818 => x"0c",
          1819 => x"33",
          1820 => x"39",
          1821 => x"74",
          1822 => x"38",
          1823 => x"80",
          1824 => x"89",
          1825 => x"38",
          1826 => x"d0",
          1827 => x"55",
          1828 => x"80",
          1829 => x"39",
          1830 => x"d9",
          1831 => x"80",
          1832 => x"27",
          1833 => x"80",
          1834 => x"89",
          1835 => x"70",
          1836 => x"55",
          1837 => x"70",
          1838 => x"55",
          1839 => x"27",
          1840 => x"14",
          1841 => x"06",
          1842 => x"74",
          1843 => x"73",
          1844 => x"38",
          1845 => x"14",
          1846 => x"05",
          1847 => x"08",
          1848 => x"54",
          1849 => x"39",
          1850 => x"84",
          1851 => x"55",
          1852 => x"81",
          1853 => x"de",
          1854 => x"3d",
          1855 => x"3d",
          1856 => x"05",
          1857 => x"52",
          1858 => x"87",
          1859 => x"e8",
          1860 => x"71",
          1861 => x"0c",
          1862 => x"04",
          1863 => x"02",
          1864 => x"02",
          1865 => x"05",
          1866 => x"83",
          1867 => x"26",
          1868 => x"72",
          1869 => x"c0",
          1870 => x"53",
          1871 => x"74",
          1872 => x"38",
          1873 => x"73",
          1874 => x"c0",
          1875 => x"51",
          1876 => x"85",
          1877 => x"98",
          1878 => x"52",
          1879 => x"82",
          1880 => x"70",
          1881 => x"38",
          1882 => x"8c",
          1883 => x"ec",
          1884 => x"fc",
          1885 => x"52",
          1886 => x"87",
          1887 => x"08",
          1888 => x"2e",
          1889 => x"81",
          1890 => x"34",
          1891 => x"13",
          1892 => x"81",
          1893 => x"86",
          1894 => x"f3",
          1895 => x"62",
          1896 => x"05",
          1897 => x"57",
          1898 => x"83",
          1899 => x"fe",
          1900 => x"de",
          1901 => x"06",
          1902 => x"71",
          1903 => x"71",
          1904 => x"2b",
          1905 => x"80",
          1906 => x"92",
          1907 => x"c0",
          1908 => x"41",
          1909 => x"5a",
          1910 => x"87",
          1911 => x"0c",
          1912 => x"84",
          1913 => x"08",
          1914 => x"70",
          1915 => x"53",
          1916 => x"2e",
          1917 => x"08",
          1918 => x"70",
          1919 => x"34",
          1920 => x"80",
          1921 => x"53",
          1922 => x"2e",
          1923 => x"53",
          1924 => x"26",
          1925 => x"80",
          1926 => x"87",
          1927 => x"08",
          1928 => x"38",
          1929 => x"8c",
          1930 => x"80",
          1931 => x"78",
          1932 => x"99",
          1933 => x"0c",
          1934 => x"8c",
          1935 => x"08",
          1936 => x"51",
          1937 => x"38",
          1938 => x"8d",
          1939 => x"17",
          1940 => x"81",
          1941 => x"53",
          1942 => x"2e",
          1943 => x"fc",
          1944 => x"52",
          1945 => x"7d",
          1946 => x"ed",
          1947 => x"80",
          1948 => x"71",
          1949 => x"38",
          1950 => x"53",
          1951 => x"c0",
          1952 => x"0d",
          1953 => x"0d",
          1954 => x"02",
          1955 => x"05",
          1956 => x"58",
          1957 => x"80",
          1958 => x"fc",
          1959 => x"de",
          1960 => x"06",
          1961 => x"71",
          1962 => x"81",
          1963 => x"38",
          1964 => x"2b",
          1965 => x"80",
          1966 => x"92",
          1967 => x"c0",
          1968 => x"40",
          1969 => x"5a",
          1970 => x"c0",
          1971 => x"76",
          1972 => x"76",
          1973 => x"75",
          1974 => x"2a",
          1975 => x"51",
          1976 => x"80",
          1977 => x"7a",
          1978 => x"5c",
          1979 => x"81",
          1980 => x"81",
          1981 => x"06",
          1982 => x"80",
          1983 => x"87",
          1984 => x"08",
          1985 => x"38",
          1986 => x"8c",
          1987 => x"80",
          1988 => x"77",
          1989 => x"99",
          1990 => x"0c",
          1991 => x"8c",
          1992 => x"08",
          1993 => x"51",
          1994 => x"38",
          1995 => x"8d",
          1996 => x"70",
          1997 => x"84",
          1998 => x"5b",
          1999 => x"2e",
          2000 => x"fc",
          2001 => x"52",
          2002 => x"7d",
          2003 => x"f8",
          2004 => x"80",
          2005 => x"71",
          2006 => x"38",
          2007 => x"53",
          2008 => x"c0",
          2009 => x"0d",
          2010 => x"0d",
          2011 => x"05",
          2012 => x"02",
          2013 => x"05",
          2014 => x"54",
          2015 => x"fe",
          2016 => x"c0",
          2017 => x"53",
          2018 => x"80",
          2019 => x"0b",
          2020 => x"8c",
          2021 => x"71",
          2022 => x"dc",
          2023 => x"24",
          2024 => x"84",
          2025 => x"92",
          2026 => x"54",
          2027 => x"8d",
          2028 => x"39",
          2029 => x"80",
          2030 => x"cb",
          2031 => x"70",
          2032 => x"81",
          2033 => x"52",
          2034 => x"8a",
          2035 => x"98",
          2036 => x"71",
          2037 => x"c0",
          2038 => x"52",
          2039 => x"81",
          2040 => x"c0",
          2041 => x"53",
          2042 => x"82",
          2043 => x"71",
          2044 => x"39",
          2045 => x"39",
          2046 => x"77",
          2047 => x"81",
          2048 => x"72",
          2049 => x"84",
          2050 => x"73",
          2051 => x"0c",
          2052 => x"04",
          2053 => x"74",
          2054 => x"71",
          2055 => x"2b",
          2056 => x"c0",
          2057 => x"84",
          2058 => x"fd",
          2059 => x"83",
          2060 => x"12",
          2061 => x"2b",
          2062 => x"07",
          2063 => x"70",
          2064 => x"2b",
          2065 => x"07",
          2066 => x"0c",
          2067 => x"56",
          2068 => x"3d",
          2069 => x"3d",
          2070 => x"84",
          2071 => x"22",
          2072 => x"72",
          2073 => x"54",
          2074 => x"2a",
          2075 => x"34",
          2076 => x"04",
          2077 => x"73",
          2078 => x"70",
          2079 => x"05",
          2080 => x"88",
          2081 => x"72",
          2082 => x"54",
          2083 => x"2a",
          2084 => x"70",
          2085 => x"34",
          2086 => x"51",
          2087 => x"83",
          2088 => x"fe",
          2089 => x"75",
          2090 => x"51",
          2091 => x"92",
          2092 => x"81",
          2093 => x"73",
          2094 => x"55",
          2095 => x"51",
          2096 => x"3d",
          2097 => x"3d",
          2098 => x"76",
          2099 => x"72",
          2100 => x"05",
          2101 => x"11",
          2102 => x"38",
          2103 => x"04",
          2104 => x"78",
          2105 => x"56",
          2106 => x"81",
          2107 => x"74",
          2108 => x"56",
          2109 => x"31",
          2110 => x"52",
          2111 => x"80",
          2112 => x"71",
          2113 => x"38",
          2114 => x"c0",
          2115 => x"0d",
          2116 => x"0d",
          2117 => x"51",
          2118 => x"73",
          2119 => x"81",
          2120 => x"33",
          2121 => x"38",
          2122 => x"de",
          2123 => x"3d",
          2124 => x"0b",
          2125 => x"0c",
          2126 => x"81",
          2127 => x"04",
          2128 => x"7b",
          2129 => x"83",
          2130 => x"5a",
          2131 => x"80",
          2132 => x"54",
          2133 => x"53",
          2134 => x"53",
          2135 => x"52",
          2136 => x"3f",
          2137 => x"08",
          2138 => x"81",
          2139 => x"81",
          2140 => x"83",
          2141 => x"16",
          2142 => x"18",
          2143 => x"18",
          2144 => x"58",
          2145 => x"9f",
          2146 => x"33",
          2147 => x"2e",
          2148 => x"93",
          2149 => x"76",
          2150 => x"52",
          2151 => x"51",
          2152 => x"83",
          2153 => x"79",
          2154 => x"0c",
          2155 => x"04",
          2156 => x"78",
          2157 => x"80",
          2158 => x"17",
          2159 => x"38",
          2160 => x"fc",
          2161 => x"c0",
          2162 => x"de",
          2163 => x"38",
          2164 => x"53",
          2165 => x"81",
          2166 => x"f7",
          2167 => x"de",
          2168 => x"2e",
          2169 => x"55",
          2170 => x"b0",
          2171 => x"81",
          2172 => x"88",
          2173 => x"f8",
          2174 => x"70",
          2175 => x"c0",
          2176 => x"c0",
          2177 => x"de",
          2178 => x"91",
          2179 => x"55",
          2180 => x"09",
          2181 => x"f0",
          2182 => x"33",
          2183 => x"2e",
          2184 => x"80",
          2185 => x"80",
          2186 => x"c0",
          2187 => x"17",
          2188 => x"fd",
          2189 => x"d4",
          2190 => x"b2",
          2191 => x"96",
          2192 => x"85",
          2193 => x"75",
          2194 => x"3f",
          2195 => x"e4",
          2196 => x"98",
          2197 => x"9c",
          2198 => x"08",
          2199 => x"17",
          2200 => x"3f",
          2201 => x"52",
          2202 => x"51",
          2203 => x"a0",
          2204 => x"05",
          2205 => x"0c",
          2206 => x"75",
          2207 => x"33",
          2208 => x"3f",
          2209 => x"34",
          2210 => x"52",
          2211 => x"51",
          2212 => x"81",
          2213 => x"80",
          2214 => x"81",
          2215 => x"de",
          2216 => x"3d",
          2217 => x"3d",
          2218 => x"1a",
          2219 => x"fe",
          2220 => x"54",
          2221 => x"73",
          2222 => x"8a",
          2223 => x"71",
          2224 => x"08",
          2225 => x"75",
          2226 => x"0c",
          2227 => x"04",
          2228 => x"7a",
          2229 => x"56",
          2230 => x"77",
          2231 => x"38",
          2232 => x"08",
          2233 => x"38",
          2234 => x"54",
          2235 => x"2e",
          2236 => x"72",
          2237 => x"38",
          2238 => x"8d",
          2239 => x"39",
          2240 => x"81",
          2241 => x"b6",
          2242 => x"2a",
          2243 => x"2a",
          2244 => x"05",
          2245 => x"55",
          2246 => x"81",
          2247 => x"81",
          2248 => x"83",
          2249 => x"b4",
          2250 => x"17",
          2251 => x"a4",
          2252 => x"55",
          2253 => x"57",
          2254 => x"3f",
          2255 => x"08",
          2256 => x"74",
          2257 => x"14",
          2258 => x"70",
          2259 => x"07",
          2260 => x"71",
          2261 => x"52",
          2262 => x"72",
          2263 => x"75",
          2264 => x"58",
          2265 => x"76",
          2266 => x"15",
          2267 => x"73",
          2268 => x"3f",
          2269 => x"08",
          2270 => x"76",
          2271 => x"06",
          2272 => x"05",
          2273 => x"3f",
          2274 => x"08",
          2275 => x"06",
          2276 => x"76",
          2277 => x"15",
          2278 => x"73",
          2279 => x"3f",
          2280 => x"08",
          2281 => x"82",
          2282 => x"06",
          2283 => x"05",
          2284 => x"3f",
          2285 => x"08",
          2286 => x"58",
          2287 => x"58",
          2288 => x"c0",
          2289 => x"0d",
          2290 => x"0d",
          2291 => x"5a",
          2292 => x"59",
          2293 => x"82",
          2294 => x"98",
          2295 => x"82",
          2296 => x"33",
          2297 => x"2e",
          2298 => x"72",
          2299 => x"38",
          2300 => x"8d",
          2301 => x"39",
          2302 => x"81",
          2303 => x"f7",
          2304 => x"2a",
          2305 => x"2a",
          2306 => x"05",
          2307 => x"55",
          2308 => x"81",
          2309 => x"59",
          2310 => x"08",
          2311 => x"74",
          2312 => x"16",
          2313 => x"16",
          2314 => x"59",
          2315 => x"53",
          2316 => x"8f",
          2317 => x"2b",
          2318 => x"74",
          2319 => x"71",
          2320 => x"72",
          2321 => x"0b",
          2322 => x"74",
          2323 => x"17",
          2324 => x"75",
          2325 => x"3f",
          2326 => x"08",
          2327 => x"c0",
          2328 => x"38",
          2329 => x"06",
          2330 => x"78",
          2331 => x"54",
          2332 => x"77",
          2333 => x"33",
          2334 => x"71",
          2335 => x"51",
          2336 => x"34",
          2337 => x"76",
          2338 => x"17",
          2339 => x"75",
          2340 => x"3f",
          2341 => x"08",
          2342 => x"c0",
          2343 => x"38",
          2344 => x"ff",
          2345 => x"10",
          2346 => x"76",
          2347 => x"51",
          2348 => x"be",
          2349 => x"2a",
          2350 => x"05",
          2351 => x"f9",
          2352 => x"de",
          2353 => x"81",
          2354 => x"ab",
          2355 => x"0a",
          2356 => x"2b",
          2357 => x"70",
          2358 => x"70",
          2359 => x"54",
          2360 => x"81",
          2361 => x"8f",
          2362 => x"07",
          2363 => x"f7",
          2364 => x"0b",
          2365 => x"78",
          2366 => x"0c",
          2367 => x"04",
          2368 => x"7a",
          2369 => x"08",
          2370 => x"59",
          2371 => x"a4",
          2372 => x"17",
          2373 => x"38",
          2374 => x"aa",
          2375 => x"73",
          2376 => x"fd",
          2377 => x"de",
          2378 => x"81",
          2379 => x"80",
          2380 => x"39",
          2381 => x"eb",
          2382 => x"80",
          2383 => x"de",
          2384 => x"80",
          2385 => x"52",
          2386 => x"84",
          2387 => x"c0",
          2388 => x"de",
          2389 => x"2e",
          2390 => x"81",
          2391 => x"81",
          2392 => x"81",
          2393 => x"ff",
          2394 => x"80",
          2395 => x"75",
          2396 => x"3f",
          2397 => x"08",
          2398 => x"16",
          2399 => x"90",
          2400 => x"55",
          2401 => x"27",
          2402 => x"15",
          2403 => x"84",
          2404 => x"07",
          2405 => x"17",
          2406 => x"76",
          2407 => x"a6",
          2408 => x"73",
          2409 => x"0c",
          2410 => x"04",
          2411 => x"7c",
          2412 => x"59",
          2413 => x"95",
          2414 => x"08",
          2415 => x"2e",
          2416 => x"17",
          2417 => x"b2",
          2418 => x"ae",
          2419 => x"7a",
          2420 => x"3f",
          2421 => x"81",
          2422 => x"27",
          2423 => x"81",
          2424 => x"55",
          2425 => x"08",
          2426 => x"d2",
          2427 => x"08",
          2428 => x"08",
          2429 => x"38",
          2430 => x"17",
          2431 => x"54",
          2432 => x"82",
          2433 => x"7a",
          2434 => x"06",
          2435 => x"81",
          2436 => x"17",
          2437 => x"83",
          2438 => x"75",
          2439 => x"f9",
          2440 => x"59",
          2441 => x"08",
          2442 => x"81",
          2443 => x"81",
          2444 => x"59",
          2445 => x"08",
          2446 => x"70",
          2447 => x"25",
          2448 => x"81",
          2449 => x"54",
          2450 => x"55",
          2451 => x"38",
          2452 => x"08",
          2453 => x"38",
          2454 => x"54",
          2455 => x"90",
          2456 => x"18",
          2457 => x"38",
          2458 => x"39",
          2459 => x"38",
          2460 => x"16",
          2461 => x"08",
          2462 => x"38",
          2463 => x"78",
          2464 => x"38",
          2465 => x"51",
          2466 => x"81",
          2467 => x"80",
          2468 => x"80",
          2469 => x"c0",
          2470 => x"09",
          2471 => x"38",
          2472 => x"08",
          2473 => x"c0",
          2474 => x"30",
          2475 => x"80",
          2476 => x"07",
          2477 => x"55",
          2478 => x"38",
          2479 => x"09",
          2480 => x"ae",
          2481 => x"80",
          2482 => x"53",
          2483 => x"51",
          2484 => x"81",
          2485 => x"81",
          2486 => x"30",
          2487 => x"c0",
          2488 => x"25",
          2489 => x"79",
          2490 => x"38",
          2491 => x"8f",
          2492 => x"79",
          2493 => x"f9",
          2494 => x"de",
          2495 => x"74",
          2496 => x"8c",
          2497 => x"17",
          2498 => x"90",
          2499 => x"54",
          2500 => x"86",
          2501 => x"90",
          2502 => x"17",
          2503 => x"54",
          2504 => x"34",
          2505 => x"56",
          2506 => x"90",
          2507 => x"80",
          2508 => x"81",
          2509 => x"55",
          2510 => x"56",
          2511 => x"81",
          2512 => x"8c",
          2513 => x"f8",
          2514 => x"70",
          2515 => x"f0",
          2516 => x"c0",
          2517 => x"56",
          2518 => x"08",
          2519 => x"7b",
          2520 => x"f6",
          2521 => x"de",
          2522 => x"de",
          2523 => x"17",
          2524 => x"80",
          2525 => x"b4",
          2526 => x"57",
          2527 => x"77",
          2528 => x"81",
          2529 => x"15",
          2530 => x"78",
          2531 => x"81",
          2532 => x"53",
          2533 => x"15",
          2534 => x"e9",
          2535 => x"c0",
          2536 => x"df",
          2537 => x"22",
          2538 => x"30",
          2539 => x"70",
          2540 => x"51",
          2541 => x"81",
          2542 => x"8a",
          2543 => x"f8",
          2544 => x"7c",
          2545 => x"56",
          2546 => x"80",
          2547 => x"f1",
          2548 => x"06",
          2549 => x"e9",
          2550 => x"18",
          2551 => x"08",
          2552 => x"38",
          2553 => x"82",
          2554 => x"38",
          2555 => x"54",
          2556 => x"74",
          2557 => x"82",
          2558 => x"22",
          2559 => x"79",
          2560 => x"38",
          2561 => x"98",
          2562 => x"cd",
          2563 => x"22",
          2564 => x"54",
          2565 => x"26",
          2566 => x"52",
          2567 => x"b0",
          2568 => x"c0",
          2569 => x"de",
          2570 => x"2e",
          2571 => x"0b",
          2572 => x"08",
          2573 => x"98",
          2574 => x"de",
          2575 => x"85",
          2576 => x"bd",
          2577 => x"31",
          2578 => x"73",
          2579 => x"f4",
          2580 => x"de",
          2581 => x"18",
          2582 => x"18",
          2583 => x"08",
          2584 => x"72",
          2585 => x"38",
          2586 => x"58",
          2587 => x"89",
          2588 => x"18",
          2589 => x"ff",
          2590 => x"05",
          2591 => x"80",
          2592 => x"de",
          2593 => x"3d",
          2594 => x"3d",
          2595 => x"08",
          2596 => x"a0",
          2597 => x"54",
          2598 => x"77",
          2599 => x"80",
          2600 => x"0c",
          2601 => x"53",
          2602 => x"80",
          2603 => x"38",
          2604 => x"06",
          2605 => x"b5",
          2606 => x"98",
          2607 => x"14",
          2608 => x"92",
          2609 => x"2a",
          2610 => x"56",
          2611 => x"26",
          2612 => x"80",
          2613 => x"16",
          2614 => x"77",
          2615 => x"53",
          2616 => x"38",
          2617 => x"51",
          2618 => x"81",
          2619 => x"53",
          2620 => x"0b",
          2621 => x"08",
          2622 => x"38",
          2623 => x"de",
          2624 => x"2e",
          2625 => x"98",
          2626 => x"de",
          2627 => x"80",
          2628 => x"8a",
          2629 => x"15",
          2630 => x"80",
          2631 => x"14",
          2632 => x"51",
          2633 => x"81",
          2634 => x"53",
          2635 => x"de",
          2636 => x"2e",
          2637 => x"82",
          2638 => x"c0",
          2639 => x"ba",
          2640 => x"81",
          2641 => x"ff",
          2642 => x"81",
          2643 => x"52",
          2644 => x"f3",
          2645 => x"c0",
          2646 => x"72",
          2647 => x"72",
          2648 => x"f2",
          2649 => x"de",
          2650 => x"15",
          2651 => x"15",
          2652 => x"b4",
          2653 => x"0c",
          2654 => x"81",
          2655 => x"8a",
          2656 => x"f7",
          2657 => x"7d",
          2658 => x"5b",
          2659 => x"76",
          2660 => x"3f",
          2661 => x"08",
          2662 => x"c0",
          2663 => x"38",
          2664 => x"08",
          2665 => x"08",
          2666 => x"f0",
          2667 => x"de",
          2668 => x"81",
          2669 => x"80",
          2670 => x"de",
          2671 => x"18",
          2672 => x"51",
          2673 => x"81",
          2674 => x"81",
          2675 => x"81",
          2676 => x"c0",
          2677 => x"83",
          2678 => x"77",
          2679 => x"72",
          2680 => x"38",
          2681 => x"75",
          2682 => x"81",
          2683 => x"a5",
          2684 => x"c0",
          2685 => x"52",
          2686 => x"8e",
          2687 => x"c0",
          2688 => x"de",
          2689 => x"2e",
          2690 => x"73",
          2691 => x"81",
          2692 => x"87",
          2693 => x"de",
          2694 => x"3d",
          2695 => x"3d",
          2696 => x"11",
          2697 => x"ec",
          2698 => x"c0",
          2699 => x"ff",
          2700 => x"33",
          2701 => x"71",
          2702 => x"81",
          2703 => x"94",
          2704 => x"d0",
          2705 => x"c0",
          2706 => x"73",
          2707 => x"81",
          2708 => x"85",
          2709 => x"fc",
          2710 => x"79",
          2711 => x"ff",
          2712 => x"12",
          2713 => x"eb",
          2714 => x"70",
          2715 => x"72",
          2716 => x"81",
          2717 => x"73",
          2718 => x"94",
          2719 => x"d6",
          2720 => x"0d",
          2721 => x"0d",
          2722 => x"55",
          2723 => x"5a",
          2724 => x"08",
          2725 => x"8a",
          2726 => x"08",
          2727 => x"ee",
          2728 => x"de",
          2729 => x"81",
          2730 => x"80",
          2731 => x"15",
          2732 => x"55",
          2733 => x"38",
          2734 => x"e6",
          2735 => x"33",
          2736 => x"70",
          2737 => x"58",
          2738 => x"86",
          2739 => x"de",
          2740 => x"73",
          2741 => x"83",
          2742 => x"73",
          2743 => x"38",
          2744 => x"06",
          2745 => x"80",
          2746 => x"75",
          2747 => x"38",
          2748 => x"08",
          2749 => x"54",
          2750 => x"2e",
          2751 => x"83",
          2752 => x"73",
          2753 => x"38",
          2754 => x"51",
          2755 => x"81",
          2756 => x"58",
          2757 => x"08",
          2758 => x"15",
          2759 => x"38",
          2760 => x"0b",
          2761 => x"77",
          2762 => x"0c",
          2763 => x"04",
          2764 => x"77",
          2765 => x"54",
          2766 => x"51",
          2767 => x"81",
          2768 => x"55",
          2769 => x"08",
          2770 => x"14",
          2771 => x"51",
          2772 => x"81",
          2773 => x"55",
          2774 => x"08",
          2775 => x"53",
          2776 => x"08",
          2777 => x"08",
          2778 => x"3f",
          2779 => x"14",
          2780 => x"08",
          2781 => x"3f",
          2782 => x"17",
          2783 => x"de",
          2784 => x"3d",
          2785 => x"3d",
          2786 => x"08",
          2787 => x"54",
          2788 => x"53",
          2789 => x"81",
          2790 => x"8d",
          2791 => x"08",
          2792 => x"34",
          2793 => x"15",
          2794 => x"0d",
          2795 => x"0d",
          2796 => x"57",
          2797 => x"17",
          2798 => x"08",
          2799 => x"82",
          2800 => x"89",
          2801 => x"55",
          2802 => x"14",
          2803 => x"16",
          2804 => x"71",
          2805 => x"38",
          2806 => x"09",
          2807 => x"38",
          2808 => x"73",
          2809 => x"81",
          2810 => x"ae",
          2811 => x"05",
          2812 => x"15",
          2813 => x"70",
          2814 => x"34",
          2815 => x"8a",
          2816 => x"38",
          2817 => x"05",
          2818 => x"81",
          2819 => x"17",
          2820 => x"12",
          2821 => x"34",
          2822 => x"9c",
          2823 => x"e8",
          2824 => x"de",
          2825 => x"0c",
          2826 => x"e7",
          2827 => x"de",
          2828 => x"17",
          2829 => x"51",
          2830 => x"81",
          2831 => x"84",
          2832 => x"3d",
          2833 => x"3d",
          2834 => x"08",
          2835 => x"61",
          2836 => x"55",
          2837 => x"2e",
          2838 => x"55",
          2839 => x"2e",
          2840 => x"80",
          2841 => x"94",
          2842 => x"1c",
          2843 => x"81",
          2844 => x"61",
          2845 => x"56",
          2846 => x"2e",
          2847 => x"83",
          2848 => x"73",
          2849 => x"70",
          2850 => x"25",
          2851 => x"51",
          2852 => x"38",
          2853 => x"0c",
          2854 => x"51",
          2855 => x"26",
          2856 => x"80",
          2857 => x"34",
          2858 => x"51",
          2859 => x"81",
          2860 => x"55",
          2861 => x"91",
          2862 => x"1d",
          2863 => x"8b",
          2864 => x"79",
          2865 => x"3f",
          2866 => x"57",
          2867 => x"55",
          2868 => x"2e",
          2869 => x"80",
          2870 => x"18",
          2871 => x"1a",
          2872 => x"70",
          2873 => x"2a",
          2874 => x"07",
          2875 => x"5a",
          2876 => x"8c",
          2877 => x"54",
          2878 => x"81",
          2879 => x"39",
          2880 => x"70",
          2881 => x"2a",
          2882 => x"75",
          2883 => x"8c",
          2884 => x"2e",
          2885 => x"a0",
          2886 => x"38",
          2887 => x"0c",
          2888 => x"76",
          2889 => x"38",
          2890 => x"b8",
          2891 => x"70",
          2892 => x"5a",
          2893 => x"76",
          2894 => x"38",
          2895 => x"70",
          2896 => x"dc",
          2897 => x"72",
          2898 => x"80",
          2899 => x"51",
          2900 => x"73",
          2901 => x"38",
          2902 => x"18",
          2903 => x"1a",
          2904 => x"55",
          2905 => x"2e",
          2906 => x"83",
          2907 => x"73",
          2908 => x"70",
          2909 => x"25",
          2910 => x"51",
          2911 => x"38",
          2912 => x"75",
          2913 => x"81",
          2914 => x"81",
          2915 => x"27",
          2916 => x"73",
          2917 => x"38",
          2918 => x"70",
          2919 => x"32",
          2920 => x"80",
          2921 => x"2a",
          2922 => x"56",
          2923 => x"81",
          2924 => x"57",
          2925 => x"f5",
          2926 => x"2b",
          2927 => x"25",
          2928 => x"80",
          2929 => x"cd",
          2930 => x"57",
          2931 => x"e6",
          2932 => x"de",
          2933 => x"2e",
          2934 => x"18",
          2935 => x"1a",
          2936 => x"56",
          2937 => x"3f",
          2938 => x"08",
          2939 => x"e8",
          2940 => x"54",
          2941 => x"80",
          2942 => x"17",
          2943 => x"34",
          2944 => x"11",
          2945 => x"74",
          2946 => x"75",
          2947 => x"d4",
          2948 => x"3f",
          2949 => x"08",
          2950 => x"9f",
          2951 => x"99",
          2952 => x"e0",
          2953 => x"ff",
          2954 => x"79",
          2955 => x"74",
          2956 => x"57",
          2957 => x"77",
          2958 => x"76",
          2959 => x"38",
          2960 => x"73",
          2961 => x"09",
          2962 => x"38",
          2963 => x"84",
          2964 => x"27",
          2965 => x"39",
          2966 => x"f2",
          2967 => x"80",
          2968 => x"54",
          2969 => x"34",
          2970 => x"58",
          2971 => x"f2",
          2972 => x"de",
          2973 => x"81",
          2974 => x"80",
          2975 => x"1b",
          2976 => x"51",
          2977 => x"81",
          2978 => x"56",
          2979 => x"08",
          2980 => x"9c",
          2981 => x"33",
          2982 => x"80",
          2983 => x"38",
          2984 => x"bf",
          2985 => x"86",
          2986 => x"15",
          2987 => x"2a",
          2988 => x"51",
          2989 => x"92",
          2990 => x"79",
          2991 => x"e4",
          2992 => x"de",
          2993 => x"2e",
          2994 => x"52",
          2995 => x"ba",
          2996 => x"39",
          2997 => x"33",
          2998 => x"80",
          2999 => x"74",
          3000 => x"81",
          3001 => x"38",
          3002 => x"70",
          3003 => x"82",
          3004 => x"54",
          3005 => x"96",
          3006 => x"06",
          3007 => x"2e",
          3008 => x"ff",
          3009 => x"1c",
          3010 => x"80",
          3011 => x"81",
          3012 => x"ba",
          3013 => x"b6",
          3014 => x"2a",
          3015 => x"51",
          3016 => x"38",
          3017 => x"70",
          3018 => x"81",
          3019 => x"55",
          3020 => x"e1",
          3021 => x"08",
          3022 => x"1d",
          3023 => x"7c",
          3024 => x"3f",
          3025 => x"08",
          3026 => x"fa",
          3027 => x"81",
          3028 => x"8f",
          3029 => x"f6",
          3030 => x"5b",
          3031 => x"70",
          3032 => x"59",
          3033 => x"73",
          3034 => x"c6",
          3035 => x"81",
          3036 => x"70",
          3037 => x"52",
          3038 => x"8d",
          3039 => x"38",
          3040 => x"09",
          3041 => x"a5",
          3042 => x"d0",
          3043 => x"ff",
          3044 => x"53",
          3045 => x"91",
          3046 => x"73",
          3047 => x"d0",
          3048 => x"71",
          3049 => x"f7",
          3050 => x"81",
          3051 => x"55",
          3052 => x"55",
          3053 => x"81",
          3054 => x"74",
          3055 => x"56",
          3056 => x"12",
          3057 => x"70",
          3058 => x"38",
          3059 => x"81",
          3060 => x"51",
          3061 => x"51",
          3062 => x"89",
          3063 => x"70",
          3064 => x"53",
          3065 => x"70",
          3066 => x"51",
          3067 => x"09",
          3068 => x"38",
          3069 => x"38",
          3070 => x"77",
          3071 => x"70",
          3072 => x"2a",
          3073 => x"07",
          3074 => x"51",
          3075 => x"8f",
          3076 => x"84",
          3077 => x"83",
          3078 => x"94",
          3079 => x"74",
          3080 => x"38",
          3081 => x"0c",
          3082 => x"86",
          3083 => x"f0",
          3084 => x"81",
          3085 => x"8c",
          3086 => x"fa",
          3087 => x"56",
          3088 => x"17",
          3089 => x"b0",
          3090 => x"52",
          3091 => x"e0",
          3092 => x"81",
          3093 => x"81",
          3094 => x"b2",
          3095 => x"b4",
          3096 => x"c0",
          3097 => x"ff",
          3098 => x"55",
          3099 => x"d5",
          3100 => x"06",
          3101 => x"80",
          3102 => x"33",
          3103 => x"81",
          3104 => x"81",
          3105 => x"81",
          3106 => x"eb",
          3107 => x"70",
          3108 => x"07",
          3109 => x"73",
          3110 => x"81",
          3111 => x"81",
          3112 => x"83",
          3113 => x"e4",
          3114 => x"16",
          3115 => x"3f",
          3116 => x"08",
          3117 => x"c0",
          3118 => x"9d",
          3119 => x"81",
          3120 => x"81",
          3121 => x"e0",
          3122 => x"de",
          3123 => x"81",
          3124 => x"80",
          3125 => x"82",
          3126 => x"de",
          3127 => x"3d",
          3128 => x"3d",
          3129 => x"84",
          3130 => x"05",
          3131 => x"80",
          3132 => x"51",
          3133 => x"81",
          3134 => x"58",
          3135 => x"0b",
          3136 => x"08",
          3137 => x"38",
          3138 => x"08",
          3139 => x"de",
          3140 => x"08",
          3141 => x"56",
          3142 => x"86",
          3143 => x"75",
          3144 => x"fe",
          3145 => x"54",
          3146 => x"2e",
          3147 => x"14",
          3148 => x"ca",
          3149 => x"c0",
          3150 => x"06",
          3151 => x"54",
          3152 => x"38",
          3153 => x"86",
          3154 => x"82",
          3155 => x"06",
          3156 => x"56",
          3157 => x"38",
          3158 => x"80",
          3159 => x"81",
          3160 => x"52",
          3161 => x"51",
          3162 => x"81",
          3163 => x"81",
          3164 => x"81",
          3165 => x"83",
          3166 => x"87",
          3167 => x"2e",
          3168 => x"82",
          3169 => x"06",
          3170 => x"56",
          3171 => x"38",
          3172 => x"74",
          3173 => x"a3",
          3174 => x"c0",
          3175 => x"06",
          3176 => x"2e",
          3177 => x"80",
          3178 => x"3d",
          3179 => x"83",
          3180 => x"15",
          3181 => x"53",
          3182 => x"8d",
          3183 => x"15",
          3184 => x"3f",
          3185 => x"08",
          3186 => x"70",
          3187 => x"0c",
          3188 => x"16",
          3189 => x"80",
          3190 => x"80",
          3191 => x"54",
          3192 => x"84",
          3193 => x"5b",
          3194 => x"80",
          3195 => x"7a",
          3196 => x"fc",
          3197 => x"de",
          3198 => x"ff",
          3199 => x"77",
          3200 => x"81",
          3201 => x"76",
          3202 => x"81",
          3203 => x"2e",
          3204 => x"8d",
          3205 => x"26",
          3206 => x"bf",
          3207 => x"f4",
          3208 => x"c0",
          3209 => x"ff",
          3210 => x"84",
          3211 => x"81",
          3212 => x"38",
          3213 => x"51",
          3214 => x"81",
          3215 => x"83",
          3216 => x"58",
          3217 => x"80",
          3218 => x"db",
          3219 => x"de",
          3220 => x"77",
          3221 => x"80",
          3222 => x"82",
          3223 => x"c4",
          3224 => x"11",
          3225 => x"06",
          3226 => x"8d",
          3227 => x"26",
          3228 => x"74",
          3229 => x"78",
          3230 => x"c1",
          3231 => x"59",
          3232 => x"15",
          3233 => x"2e",
          3234 => x"13",
          3235 => x"72",
          3236 => x"38",
          3237 => x"eb",
          3238 => x"14",
          3239 => x"3f",
          3240 => x"08",
          3241 => x"c0",
          3242 => x"23",
          3243 => x"57",
          3244 => x"83",
          3245 => x"c7",
          3246 => x"d8",
          3247 => x"c0",
          3248 => x"ff",
          3249 => x"8d",
          3250 => x"14",
          3251 => x"3f",
          3252 => x"08",
          3253 => x"14",
          3254 => x"3f",
          3255 => x"08",
          3256 => x"06",
          3257 => x"72",
          3258 => x"97",
          3259 => x"22",
          3260 => x"84",
          3261 => x"5a",
          3262 => x"83",
          3263 => x"14",
          3264 => x"79",
          3265 => x"ac",
          3266 => x"de",
          3267 => x"81",
          3268 => x"80",
          3269 => x"38",
          3270 => x"08",
          3271 => x"ff",
          3272 => x"38",
          3273 => x"83",
          3274 => x"83",
          3275 => x"74",
          3276 => x"85",
          3277 => x"89",
          3278 => x"76",
          3279 => x"c3",
          3280 => x"70",
          3281 => x"7b",
          3282 => x"73",
          3283 => x"17",
          3284 => x"ac",
          3285 => x"55",
          3286 => x"09",
          3287 => x"38",
          3288 => x"51",
          3289 => x"81",
          3290 => x"83",
          3291 => x"53",
          3292 => x"82",
          3293 => x"82",
          3294 => x"e0",
          3295 => x"ab",
          3296 => x"c0",
          3297 => x"0c",
          3298 => x"53",
          3299 => x"56",
          3300 => x"81",
          3301 => x"13",
          3302 => x"74",
          3303 => x"82",
          3304 => x"74",
          3305 => x"81",
          3306 => x"06",
          3307 => x"83",
          3308 => x"2a",
          3309 => x"72",
          3310 => x"26",
          3311 => x"ff",
          3312 => x"0c",
          3313 => x"15",
          3314 => x"0b",
          3315 => x"76",
          3316 => x"81",
          3317 => x"38",
          3318 => x"51",
          3319 => x"81",
          3320 => x"83",
          3321 => x"53",
          3322 => x"09",
          3323 => x"f9",
          3324 => x"52",
          3325 => x"b8",
          3326 => x"c0",
          3327 => x"38",
          3328 => x"08",
          3329 => x"84",
          3330 => x"d8",
          3331 => x"de",
          3332 => x"ff",
          3333 => x"72",
          3334 => x"2e",
          3335 => x"80",
          3336 => x"14",
          3337 => x"3f",
          3338 => x"08",
          3339 => x"a4",
          3340 => x"81",
          3341 => x"84",
          3342 => x"d7",
          3343 => x"de",
          3344 => x"8a",
          3345 => x"2e",
          3346 => x"9d",
          3347 => x"14",
          3348 => x"3f",
          3349 => x"08",
          3350 => x"84",
          3351 => x"d7",
          3352 => x"de",
          3353 => x"15",
          3354 => x"34",
          3355 => x"22",
          3356 => x"72",
          3357 => x"23",
          3358 => x"23",
          3359 => x"15",
          3360 => x"75",
          3361 => x"0c",
          3362 => x"04",
          3363 => x"77",
          3364 => x"73",
          3365 => x"38",
          3366 => x"72",
          3367 => x"38",
          3368 => x"71",
          3369 => x"38",
          3370 => x"84",
          3371 => x"52",
          3372 => x"09",
          3373 => x"38",
          3374 => x"51",
          3375 => x"81",
          3376 => x"81",
          3377 => x"88",
          3378 => x"08",
          3379 => x"39",
          3380 => x"73",
          3381 => x"74",
          3382 => x"0c",
          3383 => x"04",
          3384 => x"02",
          3385 => x"7a",
          3386 => x"fc",
          3387 => x"f4",
          3388 => x"54",
          3389 => x"de",
          3390 => x"bc",
          3391 => x"c0",
          3392 => x"81",
          3393 => x"70",
          3394 => x"73",
          3395 => x"38",
          3396 => x"78",
          3397 => x"2e",
          3398 => x"74",
          3399 => x"0c",
          3400 => x"80",
          3401 => x"80",
          3402 => x"70",
          3403 => x"51",
          3404 => x"81",
          3405 => x"54",
          3406 => x"c0",
          3407 => x"0d",
          3408 => x"0d",
          3409 => x"05",
          3410 => x"33",
          3411 => x"54",
          3412 => x"84",
          3413 => x"bf",
          3414 => x"98",
          3415 => x"53",
          3416 => x"05",
          3417 => x"fa",
          3418 => x"c0",
          3419 => x"de",
          3420 => x"a4",
          3421 => x"68",
          3422 => x"70",
          3423 => x"c6",
          3424 => x"c0",
          3425 => x"de",
          3426 => x"38",
          3427 => x"05",
          3428 => x"2b",
          3429 => x"80",
          3430 => x"86",
          3431 => x"06",
          3432 => x"2e",
          3433 => x"74",
          3434 => x"38",
          3435 => x"09",
          3436 => x"38",
          3437 => x"f8",
          3438 => x"c0",
          3439 => x"39",
          3440 => x"33",
          3441 => x"73",
          3442 => x"77",
          3443 => x"81",
          3444 => x"73",
          3445 => x"38",
          3446 => x"bc",
          3447 => x"07",
          3448 => x"b4",
          3449 => x"2a",
          3450 => x"51",
          3451 => x"2e",
          3452 => x"62",
          3453 => x"e8",
          3454 => x"de",
          3455 => x"82",
          3456 => x"52",
          3457 => x"51",
          3458 => x"62",
          3459 => x"8b",
          3460 => x"53",
          3461 => x"51",
          3462 => x"80",
          3463 => x"05",
          3464 => x"3f",
          3465 => x"0b",
          3466 => x"75",
          3467 => x"f1",
          3468 => x"11",
          3469 => x"80",
          3470 => x"97",
          3471 => x"51",
          3472 => x"81",
          3473 => x"55",
          3474 => x"08",
          3475 => x"b7",
          3476 => x"c4",
          3477 => x"05",
          3478 => x"2a",
          3479 => x"51",
          3480 => x"80",
          3481 => x"84",
          3482 => x"39",
          3483 => x"70",
          3484 => x"54",
          3485 => x"a9",
          3486 => x"06",
          3487 => x"2e",
          3488 => x"55",
          3489 => x"73",
          3490 => x"d6",
          3491 => x"de",
          3492 => x"ff",
          3493 => x"0c",
          3494 => x"de",
          3495 => x"f8",
          3496 => x"2a",
          3497 => x"51",
          3498 => x"2e",
          3499 => x"80",
          3500 => x"7a",
          3501 => x"a0",
          3502 => x"a4",
          3503 => x"53",
          3504 => x"e6",
          3505 => x"de",
          3506 => x"de",
          3507 => x"1b",
          3508 => x"05",
          3509 => x"d3",
          3510 => x"c0",
          3511 => x"c0",
          3512 => x"0c",
          3513 => x"56",
          3514 => x"84",
          3515 => x"90",
          3516 => x"0b",
          3517 => x"80",
          3518 => x"0c",
          3519 => x"1a",
          3520 => x"2a",
          3521 => x"51",
          3522 => x"2e",
          3523 => x"81",
          3524 => x"80",
          3525 => x"38",
          3526 => x"08",
          3527 => x"8a",
          3528 => x"89",
          3529 => x"59",
          3530 => x"76",
          3531 => x"d7",
          3532 => x"de",
          3533 => x"81",
          3534 => x"81",
          3535 => x"82",
          3536 => x"c0",
          3537 => x"09",
          3538 => x"38",
          3539 => x"78",
          3540 => x"30",
          3541 => x"80",
          3542 => x"77",
          3543 => x"38",
          3544 => x"06",
          3545 => x"c3",
          3546 => x"1a",
          3547 => x"38",
          3548 => x"06",
          3549 => x"2e",
          3550 => x"52",
          3551 => x"a6",
          3552 => x"c0",
          3553 => x"82",
          3554 => x"75",
          3555 => x"de",
          3556 => x"9c",
          3557 => x"39",
          3558 => x"74",
          3559 => x"de",
          3560 => x"3d",
          3561 => x"3d",
          3562 => x"65",
          3563 => x"5d",
          3564 => x"0c",
          3565 => x"05",
          3566 => x"f9",
          3567 => x"de",
          3568 => x"81",
          3569 => x"8a",
          3570 => x"33",
          3571 => x"2e",
          3572 => x"56",
          3573 => x"90",
          3574 => x"06",
          3575 => x"74",
          3576 => x"b6",
          3577 => x"82",
          3578 => x"34",
          3579 => x"aa",
          3580 => x"91",
          3581 => x"56",
          3582 => x"8c",
          3583 => x"1a",
          3584 => x"74",
          3585 => x"38",
          3586 => x"80",
          3587 => x"38",
          3588 => x"70",
          3589 => x"56",
          3590 => x"b2",
          3591 => x"11",
          3592 => x"77",
          3593 => x"5b",
          3594 => x"38",
          3595 => x"88",
          3596 => x"8f",
          3597 => x"08",
          3598 => x"d5",
          3599 => x"de",
          3600 => x"81",
          3601 => x"9f",
          3602 => x"2e",
          3603 => x"74",
          3604 => x"98",
          3605 => x"7e",
          3606 => x"3f",
          3607 => x"08",
          3608 => x"83",
          3609 => x"c0",
          3610 => x"89",
          3611 => x"77",
          3612 => x"d6",
          3613 => x"7f",
          3614 => x"58",
          3615 => x"75",
          3616 => x"75",
          3617 => x"77",
          3618 => x"7c",
          3619 => x"33",
          3620 => x"3f",
          3621 => x"08",
          3622 => x"7e",
          3623 => x"56",
          3624 => x"2e",
          3625 => x"16",
          3626 => x"55",
          3627 => x"94",
          3628 => x"53",
          3629 => x"b0",
          3630 => x"31",
          3631 => x"05",
          3632 => x"3f",
          3633 => x"56",
          3634 => x"9c",
          3635 => x"19",
          3636 => x"06",
          3637 => x"31",
          3638 => x"76",
          3639 => x"7b",
          3640 => x"08",
          3641 => x"d1",
          3642 => x"de",
          3643 => x"81",
          3644 => x"94",
          3645 => x"ff",
          3646 => x"05",
          3647 => x"cf",
          3648 => x"76",
          3649 => x"17",
          3650 => x"1e",
          3651 => x"18",
          3652 => x"5e",
          3653 => x"39",
          3654 => x"81",
          3655 => x"90",
          3656 => x"f2",
          3657 => x"63",
          3658 => x"40",
          3659 => x"7e",
          3660 => x"fc",
          3661 => x"51",
          3662 => x"81",
          3663 => x"55",
          3664 => x"08",
          3665 => x"18",
          3666 => x"80",
          3667 => x"74",
          3668 => x"39",
          3669 => x"70",
          3670 => x"81",
          3671 => x"56",
          3672 => x"80",
          3673 => x"38",
          3674 => x"0b",
          3675 => x"82",
          3676 => x"39",
          3677 => x"19",
          3678 => x"83",
          3679 => x"18",
          3680 => x"56",
          3681 => x"27",
          3682 => x"09",
          3683 => x"2e",
          3684 => x"94",
          3685 => x"83",
          3686 => x"56",
          3687 => x"38",
          3688 => x"22",
          3689 => x"89",
          3690 => x"55",
          3691 => x"75",
          3692 => x"18",
          3693 => x"9c",
          3694 => x"85",
          3695 => x"08",
          3696 => x"d7",
          3697 => x"de",
          3698 => x"81",
          3699 => x"80",
          3700 => x"38",
          3701 => x"ff",
          3702 => x"ff",
          3703 => x"38",
          3704 => x"0c",
          3705 => x"85",
          3706 => x"19",
          3707 => x"b0",
          3708 => x"19",
          3709 => x"81",
          3710 => x"74",
          3711 => x"3f",
          3712 => x"08",
          3713 => x"98",
          3714 => x"7e",
          3715 => x"3f",
          3716 => x"08",
          3717 => x"d2",
          3718 => x"c0",
          3719 => x"89",
          3720 => x"78",
          3721 => x"d5",
          3722 => x"7f",
          3723 => x"58",
          3724 => x"75",
          3725 => x"75",
          3726 => x"78",
          3727 => x"7c",
          3728 => x"33",
          3729 => x"3f",
          3730 => x"08",
          3731 => x"7e",
          3732 => x"78",
          3733 => x"74",
          3734 => x"38",
          3735 => x"b0",
          3736 => x"31",
          3737 => x"05",
          3738 => x"51",
          3739 => x"7e",
          3740 => x"83",
          3741 => x"89",
          3742 => x"db",
          3743 => x"08",
          3744 => x"26",
          3745 => x"51",
          3746 => x"81",
          3747 => x"fd",
          3748 => x"77",
          3749 => x"55",
          3750 => x"0c",
          3751 => x"83",
          3752 => x"80",
          3753 => x"55",
          3754 => x"83",
          3755 => x"9c",
          3756 => x"7e",
          3757 => x"3f",
          3758 => x"08",
          3759 => x"75",
          3760 => x"94",
          3761 => x"ff",
          3762 => x"05",
          3763 => x"3f",
          3764 => x"0b",
          3765 => x"7b",
          3766 => x"08",
          3767 => x"76",
          3768 => x"08",
          3769 => x"1c",
          3770 => x"08",
          3771 => x"5c",
          3772 => x"83",
          3773 => x"74",
          3774 => x"fd",
          3775 => x"18",
          3776 => x"07",
          3777 => x"19",
          3778 => x"75",
          3779 => x"0c",
          3780 => x"04",
          3781 => x"7a",
          3782 => x"05",
          3783 => x"56",
          3784 => x"81",
          3785 => x"57",
          3786 => x"08",
          3787 => x"90",
          3788 => x"86",
          3789 => x"06",
          3790 => x"73",
          3791 => x"e9",
          3792 => x"08",
          3793 => x"cc",
          3794 => x"de",
          3795 => x"81",
          3796 => x"80",
          3797 => x"16",
          3798 => x"33",
          3799 => x"55",
          3800 => x"34",
          3801 => x"53",
          3802 => x"08",
          3803 => x"3f",
          3804 => x"52",
          3805 => x"c9",
          3806 => x"88",
          3807 => x"96",
          3808 => x"f0",
          3809 => x"92",
          3810 => x"ca",
          3811 => x"81",
          3812 => x"34",
          3813 => x"df",
          3814 => x"c0",
          3815 => x"33",
          3816 => x"55",
          3817 => x"17",
          3818 => x"de",
          3819 => x"3d",
          3820 => x"3d",
          3821 => x"52",
          3822 => x"3f",
          3823 => x"08",
          3824 => x"c0",
          3825 => x"86",
          3826 => x"52",
          3827 => x"bc",
          3828 => x"c0",
          3829 => x"de",
          3830 => x"38",
          3831 => x"08",
          3832 => x"81",
          3833 => x"86",
          3834 => x"ff",
          3835 => x"3d",
          3836 => x"3f",
          3837 => x"0b",
          3838 => x"08",
          3839 => x"81",
          3840 => x"81",
          3841 => x"80",
          3842 => x"de",
          3843 => x"3d",
          3844 => x"3d",
          3845 => x"93",
          3846 => x"52",
          3847 => x"e9",
          3848 => x"de",
          3849 => x"81",
          3850 => x"80",
          3851 => x"58",
          3852 => x"3d",
          3853 => x"e0",
          3854 => x"de",
          3855 => x"81",
          3856 => x"bc",
          3857 => x"c7",
          3858 => x"98",
          3859 => x"73",
          3860 => x"38",
          3861 => x"12",
          3862 => x"39",
          3863 => x"33",
          3864 => x"70",
          3865 => x"55",
          3866 => x"2e",
          3867 => x"7f",
          3868 => x"54",
          3869 => x"81",
          3870 => x"94",
          3871 => x"39",
          3872 => x"08",
          3873 => x"81",
          3874 => x"85",
          3875 => x"de",
          3876 => x"3d",
          3877 => x"3d",
          3878 => x"5b",
          3879 => x"34",
          3880 => x"3d",
          3881 => x"52",
          3882 => x"e8",
          3883 => x"de",
          3884 => x"81",
          3885 => x"82",
          3886 => x"43",
          3887 => x"11",
          3888 => x"58",
          3889 => x"80",
          3890 => x"38",
          3891 => x"3d",
          3892 => x"d5",
          3893 => x"de",
          3894 => x"81",
          3895 => x"82",
          3896 => x"52",
          3897 => x"c8",
          3898 => x"c0",
          3899 => x"de",
          3900 => x"c1",
          3901 => x"7b",
          3902 => x"3f",
          3903 => x"08",
          3904 => x"74",
          3905 => x"3f",
          3906 => x"08",
          3907 => x"c0",
          3908 => x"38",
          3909 => x"51",
          3910 => x"81",
          3911 => x"57",
          3912 => x"08",
          3913 => x"52",
          3914 => x"f2",
          3915 => x"de",
          3916 => x"a6",
          3917 => x"74",
          3918 => x"3f",
          3919 => x"08",
          3920 => x"c0",
          3921 => x"cc",
          3922 => x"2e",
          3923 => x"86",
          3924 => x"81",
          3925 => x"81",
          3926 => x"3d",
          3927 => x"52",
          3928 => x"c9",
          3929 => x"3d",
          3930 => x"11",
          3931 => x"5a",
          3932 => x"2e",
          3933 => x"b9",
          3934 => x"16",
          3935 => x"33",
          3936 => x"73",
          3937 => x"16",
          3938 => x"26",
          3939 => x"75",
          3940 => x"38",
          3941 => x"05",
          3942 => x"6f",
          3943 => x"ff",
          3944 => x"55",
          3945 => x"74",
          3946 => x"38",
          3947 => x"11",
          3948 => x"74",
          3949 => x"39",
          3950 => x"09",
          3951 => x"38",
          3952 => x"11",
          3953 => x"74",
          3954 => x"81",
          3955 => x"70",
          3956 => x"cd",
          3957 => x"08",
          3958 => x"5c",
          3959 => x"73",
          3960 => x"38",
          3961 => x"1a",
          3962 => x"55",
          3963 => x"38",
          3964 => x"73",
          3965 => x"38",
          3966 => x"76",
          3967 => x"74",
          3968 => x"33",
          3969 => x"05",
          3970 => x"15",
          3971 => x"ba",
          3972 => x"05",
          3973 => x"ff",
          3974 => x"06",
          3975 => x"57",
          3976 => x"18",
          3977 => x"54",
          3978 => x"70",
          3979 => x"34",
          3980 => x"ee",
          3981 => x"34",
          3982 => x"c0",
          3983 => x"0d",
          3984 => x"0d",
          3985 => x"3d",
          3986 => x"71",
          3987 => x"ec",
          3988 => x"de",
          3989 => x"81",
          3990 => x"82",
          3991 => x"15",
          3992 => x"82",
          3993 => x"15",
          3994 => x"76",
          3995 => x"90",
          3996 => x"81",
          3997 => x"06",
          3998 => x"72",
          3999 => x"56",
          4000 => x"54",
          4001 => x"17",
          4002 => x"78",
          4003 => x"38",
          4004 => x"22",
          4005 => x"59",
          4006 => x"78",
          4007 => x"76",
          4008 => x"51",
          4009 => x"3f",
          4010 => x"08",
          4011 => x"54",
          4012 => x"53",
          4013 => x"3f",
          4014 => x"08",
          4015 => x"38",
          4016 => x"75",
          4017 => x"18",
          4018 => x"31",
          4019 => x"57",
          4020 => x"b1",
          4021 => x"08",
          4022 => x"38",
          4023 => x"51",
          4024 => x"81",
          4025 => x"54",
          4026 => x"08",
          4027 => x"9a",
          4028 => x"c0",
          4029 => x"81",
          4030 => x"de",
          4031 => x"16",
          4032 => x"16",
          4033 => x"2e",
          4034 => x"76",
          4035 => x"dc",
          4036 => x"31",
          4037 => x"18",
          4038 => x"90",
          4039 => x"81",
          4040 => x"06",
          4041 => x"56",
          4042 => x"9a",
          4043 => x"74",
          4044 => x"3f",
          4045 => x"08",
          4046 => x"c0",
          4047 => x"81",
          4048 => x"56",
          4049 => x"52",
          4050 => x"84",
          4051 => x"c0",
          4052 => x"ff",
          4053 => x"81",
          4054 => x"38",
          4055 => x"98",
          4056 => x"a6",
          4057 => x"16",
          4058 => x"39",
          4059 => x"16",
          4060 => x"75",
          4061 => x"53",
          4062 => x"aa",
          4063 => x"79",
          4064 => x"3f",
          4065 => x"08",
          4066 => x"0b",
          4067 => x"82",
          4068 => x"39",
          4069 => x"16",
          4070 => x"bb",
          4071 => x"2a",
          4072 => x"08",
          4073 => x"15",
          4074 => x"15",
          4075 => x"90",
          4076 => x"16",
          4077 => x"33",
          4078 => x"53",
          4079 => x"34",
          4080 => x"06",
          4081 => x"2e",
          4082 => x"9c",
          4083 => x"85",
          4084 => x"16",
          4085 => x"72",
          4086 => x"0c",
          4087 => x"04",
          4088 => x"79",
          4089 => x"75",
          4090 => x"8a",
          4091 => x"89",
          4092 => x"52",
          4093 => x"05",
          4094 => x"3f",
          4095 => x"08",
          4096 => x"c0",
          4097 => x"38",
          4098 => x"7a",
          4099 => x"d8",
          4100 => x"de",
          4101 => x"81",
          4102 => x"80",
          4103 => x"16",
          4104 => x"2b",
          4105 => x"74",
          4106 => x"86",
          4107 => x"84",
          4108 => x"06",
          4109 => x"73",
          4110 => x"38",
          4111 => x"52",
          4112 => x"da",
          4113 => x"c0",
          4114 => x"0c",
          4115 => x"14",
          4116 => x"23",
          4117 => x"51",
          4118 => x"81",
          4119 => x"55",
          4120 => x"09",
          4121 => x"38",
          4122 => x"39",
          4123 => x"84",
          4124 => x"0c",
          4125 => x"81",
          4126 => x"89",
          4127 => x"fc",
          4128 => x"87",
          4129 => x"53",
          4130 => x"e7",
          4131 => x"de",
          4132 => x"38",
          4133 => x"08",
          4134 => x"3d",
          4135 => x"3d",
          4136 => x"89",
          4137 => x"54",
          4138 => x"54",
          4139 => x"81",
          4140 => x"53",
          4141 => x"08",
          4142 => x"74",
          4143 => x"de",
          4144 => x"73",
          4145 => x"3f",
          4146 => x"08",
          4147 => x"39",
          4148 => x"08",
          4149 => x"d3",
          4150 => x"de",
          4151 => x"81",
          4152 => x"84",
          4153 => x"06",
          4154 => x"53",
          4155 => x"de",
          4156 => x"38",
          4157 => x"51",
          4158 => x"72",
          4159 => x"cf",
          4160 => x"de",
          4161 => x"32",
          4162 => x"72",
          4163 => x"70",
          4164 => x"08",
          4165 => x"54",
          4166 => x"de",
          4167 => x"3d",
          4168 => x"3d",
          4169 => x"80",
          4170 => x"70",
          4171 => x"52",
          4172 => x"3f",
          4173 => x"08",
          4174 => x"c0",
          4175 => x"64",
          4176 => x"d6",
          4177 => x"de",
          4178 => x"81",
          4179 => x"a0",
          4180 => x"cb",
          4181 => x"98",
          4182 => x"73",
          4183 => x"38",
          4184 => x"39",
          4185 => x"88",
          4186 => x"75",
          4187 => x"3f",
          4188 => x"c0",
          4189 => x"0d",
          4190 => x"0d",
          4191 => x"5c",
          4192 => x"3d",
          4193 => x"93",
          4194 => x"d6",
          4195 => x"c0",
          4196 => x"de",
          4197 => x"80",
          4198 => x"0c",
          4199 => x"11",
          4200 => x"90",
          4201 => x"56",
          4202 => x"74",
          4203 => x"75",
          4204 => x"e4",
          4205 => x"81",
          4206 => x"5b",
          4207 => x"81",
          4208 => x"75",
          4209 => x"73",
          4210 => x"81",
          4211 => x"82",
          4212 => x"76",
          4213 => x"f0",
          4214 => x"f4",
          4215 => x"c0",
          4216 => x"d1",
          4217 => x"c0",
          4218 => x"ce",
          4219 => x"c0",
          4220 => x"81",
          4221 => x"07",
          4222 => x"05",
          4223 => x"53",
          4224 => x"98",
          4225 => x"26",
          4226 => x"f9",
          4227 => x"08",
          4228 => x"08",
          4229 => x"98",
          4230 => x"81",
          4231 => x"58",
          4232 => x"3f",
          4233 => x"08",
          4234 => x"c0",
          4235 => x"38",
          4236 => x"77",
          4237 => x"5d",
          4238 => x"74",
          4239 => x"81",
          4240 => x"b4",
          4241 => x"bb",
          4242 => x"de",
          4243 => x"ff",
          4244 => x"30",
          4245 => x"1b",
          4246 => x"5b",
          4247 => x"39",
          4248 => x"ff",
          4249 => x"81",
          4250 => x"f0",
          4251 => x"30",
          4252 => x"1b",
          4253 => x"5b",
          4254 => x"83",
          4255 => x"58",
          4256 => x"92",
          4257 => x"0c",
          4258 => x"12",
          4259 => x"33",
          4260 => x"54",
          4261 => x"34",
          4262 => x"c0",
          4263 => x"0d",
          4264 => x"0d",
          4265 => x"fc",
          4266 => x"52",
          4267 => x"3f",
          4268 => x"08",
          4269 => x"c0",
          4270 => x"38",
          4271 => x"56",
          4272 => x"38",
          4273 => x"70",
          4274 => x"81",
          4275 => x"55",
          4276 => x"80",
          4277 => x"38",
          4278 => x"54",
          4279 => x"08",
          4280 => x"38",
          4281 => x"81",
          4282 => x"53",
          4283 => x"52",
          4284 => x"8c",
          4285 => x"c0",
          4286 => x"19",
          4287 => x"c9",
          4288 => x"08",
          4289 => x"ff",
          4290 => x"81",
          4291 => x"ff",
          4292 => x"06",
          4293 => x"56",
          4294 => x"08",
          4295 => x"81",
          4296 => x"82",
          4297 => x"75",
          4298 => x"54",
          4299 => x"08",
          4300 => x"27",
          4301 => x"17",
          4302 => x"de",
          4303 => x"76",
          4304 => x"3f",
          4305 => x"08",
          4306 => x"08",
          4307 => x"90",
          4308 => x"c0",
          4309 => x"90",
          4310 => x"80",
          4311 => x"75",
          4312 => x"75",
          4313 => x"de",
          4314 => x"3d",
          4315 => x"3d",
          4316 => x"a0",
          4317 => x"05",
          4318 => x"51",
          4319 => x"81",
          4320 => x"55",
          4321 => x"08",
          4322 => x"78",
          4323 => x"08",
          4324 => x"70",
          4325 => x"ae",
          4326 => x"c0",
          4327 => x"de",
          4328 => x"db",
          4329 => x"fb",
          4330 => x"85",
          4331 => x"06",
          4332 => x"86",
          4333 => x"c7",
          4334 => x"2b",
          4335 => x"24",
          4336 => x"02",
          4337 => x"33",
          4338 => x"58",
          4339 => x"76",
          4340 => x"6b",
          4341 => x"cc",
          4342 => x"de",
          4343 => x"84",
          4344 => x"06",
          4345 => x"73",
          4346 => x"d4",
          4347 => x"81",
          4348 => x"94",
          4349 => x"81",
          4350 => x"5a",
          4351 => x"08",
          4352 => x"8a",
          4353 => x"54",
          4354 => x"81",
          4355 => x"55",
          4356 => x"08",
          4357 => x"81",
          4358 => x"52",
          4359 => x"e5",
          4360 => x"c0",
          4361 => x"de",
          4362 => x"38",
          4363 => x"cf",
          4364 => x"c0",
          4365 => x"88",
          4366 => x"c0",
          4367 => x"38",
          4368 => x"c2",
          4369 => x"c0",
          4370 => x"c0",
          4371 => x"81",
          4372 => x"07",
          4373 => x"55",
          4374 => x"2e",
          4375 => x"80",
          4376 => x"80",
          4377 => x"77",
          4378 => x"3f",
          4379 => x"08",
          4380 => x"38",
          4381 => x"ba",
          4382 => x"de",
          4383 => x"74",
          4384 => x"0c",
          4385 => x"04",
          4386 => x"82",
          4387 => x"c0",
          4388 => x"3d",
          4389 => x"3f",
          4390 => x"08",
          4391 => x"c0",
          4392 => x"38",
          4393 => x"52",
          4394 => x"52",
          4395 => x"3f",
          4396 => x"08",
          4397 => x"c0",
          4398 => x"88",
          4399 => x"39",
          4400 => x"08",
          4401 => x"81",
          4402 => x"38",
          4403 => x"05",
          4404 => x"2a",
          4405 => x"55",
          4406 => x"81",
          4407 => x"5a",
          4408 => x"3d",
          4409 => x"c1",
          4410 => x"de",
          4411 => x"55",
          4412 => x"c0",
          4413 => x"87",
          4414 => x"c0",
          4415 => x"09",
          4416 => x"38",
          4417 => x"de",
          4418 => x"2e",
          4419 => x"86",
          4420 => x"81",
          4421 => x"81",
          4422 => x"de",
          4423 => x"78",
          4424 => x"3f",
          4425 => x"08",
          4426 => x"c0",
          4427 => x"38",
          4428 => x"52",
          4429 => x"ff",
          4430 => x"78",
          4431 => x"b4",
          4432 => x"54",
          4433 => x"15",
          4434 => x"b2",
          4435 => x"ca",
          4436 => x"b6",
          4437 => x"53",
          4438 => x"53",
          4439 => x"3f",
          4440 => x"b4",
          4441 => x"d4",
          4442 => x"b6",
          4443 => x"54",
          4444 => x"d5",
          4445 => x"53",
          4446 => x"11",
          4447 => x"d7",
          4448 => x"81",
          4449 => x"34",
          4450 => x"a4",
          4451 => x"c0",
          4452 => x"de",
          4453 => x"38",
          4454 => x"0a",
          4455 => x"05",
          4456 => x"d0",
          4457 => x"64",
          4458 => x"c9",
          4459 => x"54",
          4460 => x"15",
          4461 => x"81",
          4462 => x"34",
          4463 => x"b8",
          4464 => x"de",
          4465 => x"8b",
          4466 => x"75",
          4467 => x"ff",
          4468 => x"73",
          4469 => x"0c",
          4470 => x"04",
          4471 => x"a9",
          4472 => x"51",
          4473 => x"82",
          4474 => x"ff",
          4475 => x"a9",
          4476 => x"ee",
          4477 => x"c0",
          4478 => x"de",
          4479 => x"d3",
          4480 => x"a9",
          4481 => x"9d",
          4482 => x"58",
          4483 => x"81",
          4484 => x"55",
          4485 => x"08",
          4486 => x"02",
          4487 => x"33",
          4488 => x"54",
          4489 => x"82",
          4490 => x"53",
          4491 => x"52",
          4492 => x"88",
          4493 => x"b4",
          4494 => x"53",
          4495 => x"3d",
          4496 => x"ff",
          4497 => x"aa",
          4498 => x"73",
          4499 => x"3f",
          4500 => x"08",
          4501 => x"c0",
          4502 => x"63",
          4503 => x"81",
          4504 => x"65",
          4505 => x"2e",
          4506 => x"55",
          4507 => x"81",
          4508 => x"84",
          4509 => x"06",
          4510 => x"73",
          4511 => x"3f",
          4512 => x"08",
          4513 => x"c0",
          4514 => x"38",
          4515 => x"53",
          4516 => x"95",
          4517 => x"16",
          4518 => x"87",
          4519 => x"05",
          4520 => x"34",
          4521 => x"70",
          4522 => x"81",
          4523 => x"55",
          4524 => x"74",
          4525 => x"73",
          4526 => x"78",
          4527 => x"83",
          4528 => x"16",
          4529 => x"2a",
          4530 => x"51",
          4531 => x"80",
          4532 => x"38",
          4533 => x"80",
          4534 => x"52",
          4535 => x"be",
          4536 => x"c0",
          4537 => x"51",
          4538 => x"3f",
          4539 => x"de",
          4540 => x"2e",
          4541 => x"81",
          4542 => x"52",
          4543 => x"b5",
          4544 => x"de",
          4545 => x"80",
          4546 => x"58",
          4547 => x"c0",
          4548 => x"38",
          4549 => x"54",
          4550 => x"09",
          4551 => x"38",
          4552 => x"52",
          4553 => x"af",
          4554 => x"81",
          4555 => x"34",
          4556 => x"de",
          4557 => x"38",
          4558 => x"ca",
          4559 => x"c0",
          4560 => x"de",
          4561 => x"38",
          4562 => x"b5",
          4563 => x"de",
          4564 => x"74",
          4565 => x"0c",
          4566 => x"04",
          4567 => x"02",
          4568 => x"33",
          4569 => x"80",
          4570 => x"57",
          4571 => x"95",
          4572 => x"52",
          4573 => x"d2",
          4574 => x"de",
          4575 => x"81",
          4576 => x"80",
          4577 => x"5a",
          4578 => x"3d",
          4579 => x"c9",
          4580 => x"de",
          4581 => x"81",
          4582 => x"b8",
          4583 => x"cf",
          4584 => x"a0",
          4585 => x"55",
          4586 => x"75",
          4587 => x"71",
          4588 => x"33",
          4589 => x"74",
          4590 => x"57",
          4591 => x"8b",
          4592 => x"54",
          4593 => x"15",
          4594 => x"ff",
          4595 => x"81",
          4596 => x"55",
          4597 => x"c0",
          4598 => x"0d",
          4599 => x"0d",
          4600 => x"53",
          4601 => x"05",
          4602 => x"51",
          4603 => x"81",
          4604 => x"55",
          4605 => x"08",
          4606 => x"76",
          4607 => x"93",
          4608 => x"51",
          4609 => x"81",
          4610 => x"55",
          4611 => x"08",
          4612 => x"80",
          4613 => x"81",
          4614 => x"86",
          4615 => x"38",
          4616 => x"86",
          4617 => x"90",
          4618 => x"54",
          4619 => x"ff",
          4620 => x"76",
          4621 => x"83",
          4622 => x"51",
          4623 => x"3f",
          4624 => x"08",
          4625 => x"de",
          4626 => x"3d",
          4627 => x"3d",
          4628 => x"5c",
          4629 => x"98",
          4630 => x"52",
          4631 => x"d1",
          4632 => x"de",
          4633 => x"de",
          4634 => x"70",
          4635 => x"08",
          4636 => x"51",
          4637 => x"80",
          4638 => x"38",
          4639 => x"06",
          4640 => x"80",
          4641 => x"38",
          4642 => x"5f",
          4643 => x"3d",
          4644 => x"ff",
          4645 => x"81",
          4646 => x"57",
          4647 => x"08",
          4648 => x"74",
          4649 => x"c3",
          4650 => x"de",
          4651 => x"81",
          4652 => x"bf",
          4653 => x"c0",
          4654 => x"c0",
          4655 => x"59",
          4656 => x"81",
          4657 => x"56",
          4658 => x"33",
          4659 => x"16",
          4660 => x"27",
          4661 => x"56",
          4662 => x"80",
          4663 => x"80",
          4664 => x"ff",
          4665 => x"70",
          4666 => x"56",
          4667 => x"e8",
          4668 => x"76",
          4669 => x"81",
          4670 => x"80",
          4671 => x"57",
          4672 => x"78",
          4673 => x"51",
          4674 => x"2e",
          4675 => x"73",
          4676 => x"38",
          4677 => x"08",
          4678 => x"b1",
          4679 => x"de",
          4680 => x"81",
          4681 => x"a7",
          4682 => x"33",
          4683 => x"c3",
          4684 => x"2e",
          4685 => x"e4",
          4686 => x"2e",
          4687 => x"56",
          4688 => x"05",
          4689 => x"e3",
          4690 => x"c0",
          4691 => x"76",
          4692 => x"0c",
          4693 => x"04",
          4694 => x"82",
          4695 => x"ff",
          4696 => x"9d",
          4697 => x"fa",
          4698 => x"c0",
          4699 => x"c0",
          4700 => x"81",
          4701 => x"83",
          4702 => x"53",
          4703 => x"3d",
          4704 => x"ff",
          4705 => x"73",
          4706 => x"70",
          4707 => x"52",
          4708 => x"9f",
          4709 => x"bc",
          4710 => x"74",
          4711 => x"6d",
          4712 => x"70",
          4713 => x"af",
          4714 => x"de",
          4715 => x"2e",
          4716 => x"70",
          4717 => x"57",
          4718 => x"fd",
          4719 => x"c0",
          4720 => x"8d",
          4721 => x"2b",
          4722 => x"81",
          4723 => x"86",
          4724 => x"c0",
          4725 => x"9f",
          4726 => x"ff",
          4727 => x"54",
          4728 => x"8a",
          4729 => x"70",
          4730 => x"06",
          4731 => x"ff",
          4732 => x"38",
          4733 => x"15",
          4734 => x"80",
          4735 => x"74",
          4736 => x"b4",
          4737 => x"89",
          4738 => x"c0",
          4739 => x"81",
          4740 => x"88",
          4741 => x"26",
          4742 => x"39",
          4743 => x"86",
          4744 => x"81",
          4745 => x"ff",
          4746 => x"38",
          4747 => x"54",
          4748 => x"81",
          4749 => x"81",
          4750 => x"78",
          4751 => x"5a",
          4752 => x"6d",
          4753 => x"81",
          4754 => x"57",
          4755 => x"9f",
          4756 => x"38",
          4757 => x"54",
          4758 => x"81",
          4759 => x"b1",
          4760 => x"2e",
          4761 => x"a7",
          4762 => x"15",
          4763 => x"54",
          4764 => x"09",
          4765 => x"38",
          4766 => x"76",
          4767 => x"41",
          4768 => x"52",
          4769 => x"52",
          4770 => x"b3",
          4771 => x"c0",
          4772 => x"de",
          4773 => x"f7",
          4774 => x"74",
          4775 => x"e5",
          4776 => x"c0",
          4777 => x"de",
          4778 => x"38",
          4779 => x"38",
          4780 => x"74",
          4781 => x"39",
          4782 => x"08",
          4783 => x"81",
          4784 => x"38",
          4785 => x"74",
          4786 => x"38",
          4787 => x"51",
          4788 => x"3f",
          4789 => x"08",
          4790 => x"c0",
          4791 => x"a0",
          4792 => x"c0",
          4793 => x"51",
          4794 => x"3f",
          4795 => x"0b",
          4796 => x"8b",
          4797 => x"67",
          4798 => x"a7",
          4799 => x"81",
          4800 => x"34",
          4801 => x"ad",
          4802 => x"de",
          4803 => x"73",
          4804 => x"de",
          4805 => x"3d",
          4806 => x"3d",
          4807 => x"02",
          4808 => x"cb",
          4809 => x"3d",
          4810 => x"72",
          4811 => x"5a",
          4812 => x"81",
          4813 => x"58",
          4814 => x"08",
          4815 => x"91",
          4816 => x"77",
          4817 => x"7c",
          4818 => x"38",
          4819 => x"59",
          4820 => x"90",
          4821 => x"81",
          4822 => x"06",
          4823 => x"73",
          4824 => x"54",
          4825 => x"82",
          4826 => x"39",
          4827 => x"8b",
          4828 => x"11",
          4829 => x"2b",
          4830 => x"54",
          4831 => x"fe",
          4832 => x"ff",
          4833 => x"70",
          4834 => x"07",
          4835 => x"de",
          4836 => x"8c",
          4837 => x"40",
          4838 => x"55",
          4839 => x"88",
          4840 => x"08",
          4841 => x"38",
          4842 => x"77",
          4843 => x"56",
          4844 => x"51",
          4845 => x"3f",
          4846 => x"55",
          4847 => x"08",
          4848 => x"38",
          4849 => x"de",
          4850 => x"2e",
          4851 => x"81",
          4852 => x"ff",
          4853 => x"38",
          4854 => x"08",
          4855 => x"16",
          4856 => x"2e",
          4857 => x"87",
          4858 => x"74",
          4859 => x"74",
          4860 => x"81",
          4861 => x"38",
          4862 => x"ff",
          4863 => x"2e",
          4864 => x"7b",
          4865 => x"80",
          4866 => x"81",
          4867 => x"81",
          4868 => x"06",
          4869 => x"56",
          4870 => x"52",
          4871 => x"af",
          4872 => x"de",
          4873 => x"81",
          4874 => x"80",
          4875 => x"81",
          4876 => x"56",
          4877 => x"d3",
          4878 => x"ff",
          4879 => x"7c",
          4880 => x"55",
          4881 => x"b3",
          4882 => x"1b",
          4883 => x"1b",
          4884 => x"33",
          4885 => x"54",
          4886 => x"34",
          4887 => x"fe",
          4888 => x"08",
          4889 => x"74",
          4890 => x"75",
          4891 => x"16",
          4892 => x"33",
          4893 => x"73",
          4894 => x"77",
          4895 => x"de",
          4896 => x"3d",
          4897 => x"3d",
          4898 => x"02",
          4899 => x"eb",
          4900 => x"3d",
          4901 => x"59",
          4902 => x"8b",
          4903 => x"81",
          4904 => x"24",
          4905 => x"81",
          4906 => x"84",
          4907 => x"dc",
          4908 => x"51",
          4909 => x"2e",
          4910 => x"75",
          4911 => x"c0",
          4912 => x"06",
          4913 => x"7e",
          4914 => x"d0",
          4915 => x"c0",
          4916 => x"06",
          4917 => x"56",
          4918 => x"74",
          4919 => x"76",
          4920 => x"81",
          4921 => x"8a",
          4922 => x"b2",
          4923 => x"fc",
          4924 => x"52",
          4925 => x"a4",
          4926 => x"de",
          4927 => x"38",
          4928 => x"80",
          4929 => x"74",
          4930 => x"26",
          4931 => x"15",
          4932 => x"74",
          4933 => x"38",
          4934 => x"80",
          4935 => x"84",
          4936 => x"92",
          4937 => x"80",
          4938 => x"38",
          4939 => x"06",
          4940 => x"2e",
          4941 => x"56",
          4942 => x"78",
          4943 => x"89",
          4944 => x"2b",
          4945 => x"43",
          4946 => x"38",
          4947 => x"30",
          4948 => x"77",
          4949 => x"91",
          4950 => x"c2",
          4951 => x"f8",
          4952 => x"52",
          4953 => x"a4",
          4954 => x"56",
          4955 => x"08",
          4956 => x"77",
          4957 => x"77",
          4958 => x"c0",
          4959 => x"45",
          4960 => x"bf",
          4961 => x"8e",
          4962 => x"26",
          4963 => x"74",
          4964 => x"48",
          4965 => x"75",
          4966 => x"38",
          4967 => x"81",
          4968 => x"fa",
          4969 => x"2a",
          4970 => x"56",
          4971 => x"2e",
          4972 => x"87",
          4973 => x"82",
          4974 => x"38",
          4975 => x"55",
          4976 => x"83",
          4977 => x"81",
          4978 => x"56",
          4979 => x"80",
          4980 => x"38",
          4981 => x"83",
          4982 => x"06",
          4983 => x"78",
          4984 => x"91",
          4985 => x"0b",
          4986 => x"22",
          4987 => x"80",
          4988 => x"74",
          4989 => x"38",
          4990 => x"56",
          4991 => x"17",
          4992 => x"57",
          4993 => x"2e",
          4994 => x"75",
          4995 => x"79",
          4996 => x"fe",
          4997 => x"81",
          4998 => x"84",
          4999 => x"05",
          5000 => x"5e",
          5001 => x"80",
          5002 => x"c0",
          5003 => x"8a",
          5004 => x"fd",
          5005 => x"75",
          5006 => x"38",
          5007 => x"78",
          5008 => x"8c",
          5009 => x"0b",
          5010 => x"22",
          5011 => x"80",
          5012 => x"74",
          5013 => x"38",
          5014 => x"56",
          5015 => x"17",
          5016 => x"57",
          5017 => x"2e",
          5018 => x"75",
          5019 => x"79",
          5020 => x"fe",
          5021 => x"81",
          5022 => x"10",
          5023 => x"81",
          5024 => x"9f",
          5025 => x"38",
          5026 => x"de",
          5027 => x"81",
          5028 => x"05",
          5029 => x"2a",
          5030 => x"56",
          5031 => x"17",
          5032 => x"81",
          5033 => x"60",
          5034 => x"65",
          5035 => x"12",
          5036 => x"30",
          5037 => x"74",
          5038 => x"59",
          5039 => x"7d",
          5040 => x"81",
          5041 => x"76",
          5042 => x"41",
          5043 => x"76",
          5044 => x"90",
          5045 => x"62",
          5046 => x"51",
          5047 => x"26",
          5048 => x"75",
          5049 => x"31",
          5050 => x"65",
          5051 => x"fe",
          5052 => x"81",
          5053 => x"58",
          5054 => x"09",
          5055 => x"38",
          5056 => x"08",
          5057 => x"26",
          5058 => x"78",
          5059 => x"79",
          5060 => x"78",
          5061 => x"86",
          5062 => x"82",
          5063 => x"06",
          5064 => x"83",
          5065 => x"81",
          5066 => x"27",
          5067 => x"8f",
          5068 => x"55",
          5069 => x"26",
          5070 => x"59",
          5071 => x"62",
          5072 => x"74",
          5073 => x"38",
          5074 => x"88",
          5075 => x"c0",
          5076 => x"26",
          5077 => x"86",
          5078 => x"1a",
          5079 => x"79",
          5080 => x"38",
          5081 => x"80",
          5082 => x"2e",
          5083 => x"83",
          5084 => x"9f",
          5085 => x"8b",
          5086 => x"06",
          5087 => x"74",
          5088 => x"84",
          5089 => x"52",
          5090 => x"a2",
          5091 => x"53",
          5092 => x"52",
          5093 => x"a2",
          5094 => x"80",
          5095 => x"51",
          5096 => x"3f",
          5097 => x"34",
          5098 => x"ff",
          5099 => x"1b",
          5100 => x"a2",
          5101 => x"90",
          5102 => x"83",
          5103 => x"70",
          5104 => x"80",
          5105 => x"55",
          5106 => x"ff",
          5107 => x"66",
          5108 => x"ff",
          5109 => x"38",
          5110 => x"ff",
          5111 => x"1b",
          5112 => x"f2",
          5113 => x"74",
          5114 => x"51",
          5115 => x"3f",
          5116 => x"1c",
          5117 => x"98",
          5118 => x"a0",
          5119 => x"ff",
          5120 => x"51",
          5121 => x"3f",
          5122 => x"1b",
          5123 => x"e4",
          5124 => x"2e",
          5125 => x"80",
          5126 => x"88",
          5127 => x"80",
          5128 => x"ff",
          5129 => x"7c",
          5130 => x"51",
          5131 => x"3f",
          5132 => x"1b",
          5133 => x"bc",
          5134 => x"b0",
          5135 => x"a0",
          5136 => x"52",
          5137 => x"ff",
          5138 => x"ff",
          5139 => x"c0",
          5140 => x"0b",
          5141 => x"34",
          5142 => x"cc",
          5143 => x"c7",
          5144 => x"39",
          5145 => x"0a",
          5146 => x"51",
          5147 => x"3f",
          5148 => x"ff",
          5149 => x"1b",
          5150 => x"da",
          5151 => x"0b",
          5152 => x"a9",
          5153 => x"34",
          5154 => x"cd",
          5155 => x"1b",
          5156 => x"8f",
          5157 => x"d5",
          5158 => x"1b",
          5159 => x"ff",
          5160 => x"81",
          5161 => x"7a",
          5162 => x"ff",
          5163 => x"81",
          5164 => x"c0",
          5165 => x"38",
          5166 => x"09",
          5167 => x"ee",
          5168 => x"60",
          5169 => x"7a",
          5170 => x"ff",
          5171 => x"84",
          5172 => x"52",
          5173 => x"9f",
          5174 => x"8b",
          5175 => x"52",
          5176 => x"9f",
          5177 => x"8a",
          5178 => x"52",
          5179 => x"51",
          5180 => x"3f",
          5181 => x"83",
          5182 => x"ff",
          5183 => x"82",
          5184 => x"1b",
          5185 => x"ec",
          5186 => x"d5",
          5187 => x"ff",
          5188 => x"75",
          5189 => x"05",
          5190 => x"7e",
          5191 => x"e5",
          5192 => x"60",
          5193 => x"52",
          5194 => x"9a",
          5195 => x"53",
          5196 => x"51",
          5197 => x"3f",
          5198 => x"58",
          5199 => x"09",
          5200 => x"38",
          5201 => x"51",
          5202 => x"3f",
          5203 => x"1b",
          5204 => x"a0",
          5205 => x"52",
          5206 => x"91",
          5207 => x"ff",
          5208 => x"81",
          5209 => x"f8",
          5210 => x"7a",
          5211 => x"84",
          5212 => x"61",
          5213 => x"26",
          5214 => x"57",
          5215 => x"53",
          5216 => x"51",
          5217 => x"3f",
          5218 => x"08",
          5219 => x"84",
          5220 => x"de",
          5221 => x"7a",
          5222 => x"aa",
          5223 => x"75",
          5224 => x"56",
          5225 => x"81",
          5226 => x"80",
          5227 => x"38",
          5228 => x"83",
          5229 => x"63",
          5230 => x"74",
          5231 => x"38",
          5232 => x"54",
          5233 => x"52",
          5234 => x"99",
          5235 => x"de",
          5236 => x"c1",
          5237 => x"75",
          5238 => x"56",
          5239 => x"8c",
          5240 => x"2e",
          5241 => x"56",
          5242 => x"ff",
          5243 => x"84",
          5244 => x"2e",
          5245 => x"56",
          5246 => x"58",
          5247 => x"38",
          5248 => x"77",
          5249 => x"ff",
          5250 => x"82",
          5251 => x"78",
          5252 => x"c2",
          5253 => x"1b",
          5254 => x"34",
          5255 => x"16",
          5256 => x"82",
          5257 => x"83",
          5258 => x"84",
          5259 => x"67",
          5260 => x"fd",
          5261 => x"51",
          5262 => x"3f",
          5263 => x"16",
          5264 => x"c0",
          5265 => x"bf",
          5266 => x"86",
          5267 => x"de",
          5268 => x"16",
          5269 => x"83",
          5270 => x"ff",
          5271 => x"66",
          5272 => x"1b",
          5273 => x"8c",
          5274 => x"77",
          5275 => x"7e",
          5276 => x"91",
          5277 => x"81",
          5278 => x"a2",
          5279 => x"80",
          5280 => x"ff",
          5281 => x"81",
          5282 => x"c0",
          5283 => x"89",
          5284 => x"8a",
          5285 => x"86",
          5286 => x"c0",
          5287 => x"81",
          5288 => x"99",
          5289 => x"f5",
          5290 => x"60",
          5291 => x"79",
          5292 => x"5a",
          5293 => x"78",
          5294 => x"8d",
          5295 => x"55",
          5296 => x"fc",
          5297 => x"51",
          5298 => x"7a",
          5299 => x"81",
          5300 => x"8c",
          5301 => x"74",
          5302 => x"38",
          5303 => x"81",
          5304 => x"81",
          5305 => x"8a",
          5306 => x"06",
          5307 => x"76",
          5308 => x"76",
          5309 => x"55",
          5310 => x"c0",
          5311 => x"0d",
          5312 => x"0d",
          5313 => x"93",
          5314 => x"38",
          5315 => x"81",
          5316 => x"52",
          5317 => x"81",
          5318 => x"81",
          5319 => x"cf",
          5320 => x"f9",
          5321 => x"90",
          5322 => x"39",
          5323 => x"51",
          5324 => x"81",
          5325 => x"80",
          5326 => x"d0",
          5327 => x"dd",
          5328 => x"d8",
          5329 => x"39",
          5330 => x"51",
          5331 => x"81",
          5332 => x"80",
          5333 => x"d1",
          5334 => x"c1",
          5335 => x"b0",
          5336 => x"81",
          5337 => x"b5",
          5338 => x"e0",
          5339 => x"81",
          5340 => x"a9",
          5341 => x"a0",
          5342 => x"81",
          5343 => x"9d",
          5344 => x"d4",
          5345 => x"81",
          5346 => x"91",
          5347 => x"84",
          5348 => x"81",
          5349 => x"85",
          5350 => x"a8",
          5351 => x"a1",
          5352 => x"0d",
          5353 => x"0d",
          5354 => x"56",
          5355 => x"26",
          5356 => x"52",
          5357 => x"29",
          5358 => x"87",
          5359 => x"51",
          5360 => x"3f",
          5361 => x"08",
          5362 => x"fe",
          5363 => x"81",
          5364 => x"54",
          5365 => x"52",
          5366 => x"51",
          5367 => x"3f",
          5368 => x"04",
          5369 => x"7d",
          5370 => x"8c",
          5371 => x"05",
          5372 => x"15",
          5373 => x"5a",
          5374 => x"5c",
          5375 => x"d3",
          5376 => x"8c",
          5377 => x"d3",
          5378 => x"86",
          5379 => x"55",
          5380 => x"80",
          5381 => x"90",
          5382 => x"79",
          5383 => x"38",
          5384 => x"74",
          5385 => x"78",
          5386 => x"72",
          5387 => x"d3",
          5388 => x"8b",
          5389 => x"39",
          5390 => x"51",
          5391 => x"3f",
          5392 => x"80",
          5393 => x"16",
          5394 => x"27",
          5395 => x"08",
          5396 => x"dc",
          5397 => x"cd",
          5398 => x"81",
          5399 => x"ff",
          5400 => x"84",
          5401 => x"39",
          5402 => x"72",
          5403 => x"38",
          5404 => x"81",
          5405 => x"ff",
          5406 => x"89",
          5407 => x"84",
          5408 => x"bd",
          5409 => x"55",
          5410 => x"f6",
          5411 => x"80",
          5412 => x"88",
          5413 => x"a9",
          5414 => x"74",
          5415 => x"38",
          5416 => x"33",
          5417 => x"52",
          5418 => x"74",
          5419 => x"72",
          5420 => x"38",
          5421 => x"26",
          5422 => x"51",
          5423 => x"51",
          5424 => x"3f",
          5425 => x"d3",
          5426 => x"8c",
          5427 => x"f1",
          5428 => x"77",
          5429 => x"fe",
          5430 => x"81",
          5431 => x"98",
          5432 => x"2c",
          5433 => x"a0",
          5434 => x"06",
          5435 => x"f9",
          5436 => x"de",
          5437 => x"2b",
          5438 => x"70",
          5439 => x"30",
          5440 => x"9f",
          5441 => x"56",
          5442 => x"9b",
          5443 => x"72",
          5444 => x"9b",
          5445 => x"06",
          5446 => x"53",
          5447 => x"1c",
          5448 => x"26",
          5449 => x"ff",
          5450 => x"de",
          5451 => x"3d",
          5452 => x"3d",
          5453 => x"84",
          5454 => x"05",
          5455 => x"30",
          5456 => x"80",
          5457 => x"ff",
          5458 => x"51",
          5459 => x"5b",
          5460 => x"74",
          5461 => x"81",
          5462 => x"8c",
          5463 => x"57",
          5464 => x"3f",
          5465 => x"08",
          5466 => x"c0",
          5467 => x"81",
          5468 => x"87",
          5469 => x"0c",
          5470 => x"08",
          5471 => x"d4",
          5472 => x"80",
          5473 => x"76",
          5474 => x"3f",
          5475 => x"08",
          5476 => x"c0",
          5477 => x"7a",
          5478 => x"2e",
          5479 => x"19",
          5480 => x"59",
          5481 => x"3d",
          5482 => x"cc",
          5483 => x"30",
          5484 => x"80",
          5485 => x"79",
          5486 => x"38",
          5487 => x"90",
          5488 => x"90",
          5489 => x"98",
          5490 => x"78",
          5491 => x"3f",
          5492 => x"81",
          5493 => x"96",
          5494 => x"f9",
          5495 => x"02",
          5496 => x"05",
          5497 => x"ff",
          5498 => x"7a",
          5499 => x"fe",
          5500 => x"de",
          5501 => x"38",
          5502 => x"88",
          5503 => x"2e",
          5504 => x"39",
          5505 => x"54",
          5506 => x"53",
          5507 => x"51",
          5508 => x"de",
          5509 => x"83",
          5510 => x"76",
          5511 => x"0c",
          5512 => x"04",
          5513 => x"02",
          5514 => x"81",
          5515 => x"81",
          5516 => x"55",
          5517 => x"3f",
          5518 => x"22",
          5519 => x"89",
          5520 => x"ac",
          5521 => x"b8",
          5522 => x"c1",
          5523 => x"d4",
          5524 => x"87",
          5525 => x"80",
          5526 => x"fe",
          5527 => x"86",
          5528 => x"fe",
          5529 => x"c0",
          5530 => x"53",
          5531 => x"3f",
          5532 => x"f2",
          5533 => x"d4",
          5534 => x"f4",
          5535 => x"51",
          5536 => x"3f",
          5537 => x"70",
          5538 => x"52",
          5539 => x"95",
          5540 => x"fe",
          5541 => x"81",
          5542 => x"fe",
          5543 => x"80",
          5544 => x"fe",
          5545 => x"2a",
          5546 => x"51",
          5547 => x"2e",
          5548 => x"51",
          5549 => x"3f",
          5550 => x"51",
          5551 => x"3f",
          5552 => x"f1",
          5553 => x"83",
          5554 => x"06",
          5555 => x"80",
          5556 => x"81",
          5557 => x"ca",
          5558 => x"9c",
          5559 => x"c2",
          5560 => x"fe",
          5561 => x"72",
          5562 => x"81",
          5563 => x"71",
          5564 => x"38",
          5565 => x"f1",
          5566 => x"d5",
          5567 => x"f3",
          5568 => x"51",
          5569 => x"3f",
          5570 => x"70",
          5571 => x"52",
          5572 => x"95",
          5573 => x"fe",
          5574 => x"81",
          5575 => x"fe",
          5576 => x"80",
          5577 => x"fa",
          5578 => x"2a",
          5579 => x"51",
          5580 => x"2e",
          5581 => x"51",
          5582 => x"3f",
          5583 => x"51",
          5584 => x"3f",
          5585 => x"f0",
          5586 => x"87",
          5587 => x"06",
          5588 => x"80",
          5589 => x"81",
          5590 => x"c6",
          5591 => x"ec",
          5592 => x"be",
          5593 => x"fe",
          5594 => x"72",
          5595 => x"81",
          5596 => x"71",
          5597 => x"38",
          5598 => x"f0",
          5599 => x"d6",
          5600 => x"f2",
          5601 => x"51",
          5602 => x"3f",
          5603 => x"3f",
          5604 => x"04",
          5605 => x"78",
          5606 => x"55",
          5607 => x"80",
          5608 => x"38",
          5609 => x"77",
          5610 => x"33",
          5611 => x"39",
          5612 => x"80",
          5613 => x"81",
          5614 => x"57",
          5615 => x"2e",
          5616 => x"53",
          5617 => x"84",
          5618 => x"38",
          5619 => x"06",
          5620 => x"2e",
          5621 => x"88",
          5622 => x"70",
          5623 => x"34",
          5624 => x"90",
          5625 => x"f0",
          5626 => x"53",
          5627 => x"55",
          5628 => x"3f",
          5629 => x"08",
          5630 => x"15",
          5631 => x"81",
          5632 => x"38",
          5633 => x"81",
          5634 => x"53",
          5635 => x"d2",
          5636 => x"72",
          5637 => x"0c",
          5638 => x"04",
          5639 => x"77",
          5640 => x"56",
          5641 => x"75",
          5642 => x"d4",
          5643 => x"ec",
          5644 => x"a7",
          5645 => x"81",
          5646 => x"81",
          5647 => x"ff",
          5648 => x"81",
          5649 => x"30",
          5650 => x"c0",
          5651 => x"25",
          5652 => x"51",
          5653 => x"81",
          5654 => x"81",
          5655 => x"54",
          5656 => x"09",
          5657 => x"38",
          5658 => x"53",
          5659 => x"51",
          5660 => x"81",
          5661 => x"80",
          5662 => x"81",
          5663 => x"51",
          5664 => x"3f",
          5665 => x"f5",
          5666 => x"a6",
          5667 => x"81",
          5668 => x"81",
          5669 => x"54",
          5670 => x"09",
          5671 => x"38",
          5672 => x"51",
          5673 => x"3f",
          5674 => x"de",
          5675 => x"3d",
          5676 => x"3d",
          5677 => x"71",
          5678 => x"0c",
          5679 => x"52",
          5680 => x"88",
          5681 => x"de",
          5682 => x"ff",
          5683 => x"7d",
          5684 => x"06",
          5685 => x"d6",
          5686 => x"3d",
          5687 => x"ff",
          5688 => x"7c",
          5689 => x"81",
          5690 => x"ff",
          5691 => x"81",
          5692 => x"7d",
          5693 => x"81",
          5694 => x"92",
          5695 => x"70",
          5696 => x"d7",
          5697 => x"fc",
          5698 => x"3d",
          5699 => x"80",
          5700 => x"51",
          5701 => x"b7",
          5702 => x"05",
          5703 => x"3f",
          5704 => x"08",
          5705 => x"90",
          5706 => x"78",
          5707 => x"8a",
          5708 => x"80",
          5709 => x"dc",
          5710 => x"2e",
          5711 => x"78",
          5712 => x"38",
          5713 => x"81",
          5714 => x"82",
          5715 => x"78",
          5716 => x"ae",
          5717 => x"39",
          5718 => x"82",
          5719 => x"94",
          5720 => x"38",
          5721 => x"78",
          5722 => x"85",
          5723 => x"80",
          5724 => x"38",
          5725 => x"83",
          5726 => x"bc",
          5727 => x"38",
          5728 => x"78",
          5729 => x"87",
          5730 => x"80",
          5731 => x"bf",
          5732 => x"39",
          5733 => x"2e",
          5734 => x"78",
          5735 => x"a9",
          5736 => x"d0",
          5737 => x"38",
          5738 => x"24",
          5739 => x"80",
          5740 => x"eb",
          5741 => x"39",
          5742 => x"2e",
          5743 => x"78",
          5744 => x"8d",
          5745 => x"ed",
          5746 => x"82",
          5747 => x"38",
          5748 => x"24",
          5749 => x"80",
          5750 => x"ce",
          5751 => x"f9",
          5752 => x"38",
          5753 => x"78",
          5754 => x"8e",
          5755 => x"81",
          5756 => x"ba",
          5757 => x"39",
          5758 => x"f4",
          5759 => x"f8",
          5760 => x"82",
          5761 => x"de",
          5762 => x"38",
          5763 => x"51",
          5764 => x"b7",
          5765 => x"11",
          5766 => x"05",
          5767 => x"fa",
          5768 => x"c0",
          5769 => x"88",
          5770 => x"25",
          5771 => x"43",
          5772 => x"05",
          5773 => x"80",
          5774 => x"51",
          5775 => x"3f",
          5776 => x"08",
          5777 => x"59",
          5778 => x"81",
          5779 => x"fe",
          5780 => x"81",
          5781 => x"39",
          5782 => x"51",
          5783 => x"b7",
          5784 => x"11",
          5785 => x"05",
          5786 => x"ae",
          5787 => x"c0",
          5788 => x"fd",
          5789 => x"53",
          5790 => x"80",
          5791 => x"51",
          5792 => x"3f",
          5793 => x"08",
          5794 => x"c8",
          5795 => x"39",
          5796 => x"f4",
          5797 => x"f8",
          5798 => x"80",
          5799 => x"de",
          5800 => x"2e",
          5801 => x"89",
          5802 => x"38",
          5803 => x"f0",
          5804 => x"f8",
          5805 => x"80",
          5806 => x"de",
          5807 => x"38",
          5808 => x"08",
          5809 => x"81",
          5810 => x"79",
          5811 => x"eb",
          5812 => x"cb",
          5813 => x"79",
          5814 => x"b4",
          5815 => x"f0",
          5816 => x"b3",
          5817 => x"de",
          5818 => x"93",
          5819 => x"a0",
          5820 => x"cd",
          5821 => x"fc",
          5822 => x"3d",
          5823 => x"51",
          5824 => x"3f",
          5825 => x"08",
          5826 => x"f8",
          5827 => x"fe",
          5828 => x"81",
          5829 => x"c0",
          5830 => x"51",
          5831 => x"80",
          5832 => x"3d",
          5833 => x"51",
          5834 => x"3f",
          5835 => x"08",
          5836 => x"f8",
          5837 => x"fe",
          5838 => x"81",
          5839 => x"b8",
          5840 => x"05",
          5841 => x"e5",
          5842 => x"de",
          5843 => x"3d",
          5844 => x"52",
          5845 => x"dd",
          5846 => x"8c",
          5847 => x"f4",
          5848 => x"80",
          5849 => x"c0",
          5850 => x"06",
          5851 => x"79",
          5852 => x"f4",
          5853 => x"de",
          5854 => x"2e",
          5855 => x"81",
          5856 => x"51",
          5857 => x"fa",
          5858 => x"3d",
          5859 => x"53",
          5860 => x"51",
          5861 => x"3f",
          5862 => x"08",
          5863 => x"e2",
          5864 => x"fe",
          5865 => x"fe",
          5866 => x"fe",
          5867 => x"81",
          5868 => x"80",
          5869 => x"38",
          5870 => x"ec",
          5871 => x"f8",
          5872 => x"fe",
          5873 => x"de",
          5874 => x"38",
          5875 => x"08",
          5876 => x"d4",
          5877 => x"e9",
          5878 => x"5c",
          5879 => x"27",
          5880 => x"61",
          5881 => x"70",
          5882 => x"0c",
          5883 => x"f5",
          5884 => x"39",
          5885 => x"f4",
          5886 => x"f8",
          5887 => x"fe",
          5888 => x"de",
          5889 => x"df",
          5890 => x"d4",
          5891 => x"80",
          5892 => x"81",
          5893 => x"44",
          5894 => x"81",
          5895 => x"59",
          5896 => x"88",
          5897 => x"94",
          5898 => x"39",
          5899 => x"33",
          5900 => x"2e",
          5901 => x"db",
          5902 => x"ab",
          5903 => x"d7",
          5904 => x"80",
          5905 => x"81",
          5906 => x"44",
          5907 => x"db",
          5908 => x"78",
          5909 => x"38",
          5910 => x"08",
          5911 => x"81",
          5912 => x"fc",
          5913 => x"b7",
          5914 => x"11",
          5915 => x"05",
          5916 => x"a6",
          5917 => x"c0",
          5918 => x"38",
          5919 => x"33",
          5920 => x"2e",
          5921 => x"db",
          5922 => x"80",
          5923 => x"db",
          5924 => x"78",
          5925 => x"38",
          5926 => x"08",
          5927 => x"81",
          5928 => x"59",
          5929 => x"88",
          5930 => x"a0",
          5931 => x"39",
          5932 => x"33",
          5933 => x"2e",
          5934 => x"db",
          5935 => x"99",
          5936 => x"d2",
          5937 => x"80",
          5938 => x"81",
          5939 => x"43",
          5940 => x"db",
          5941 => x"05",
          5942 => x"fe",
          5943 => x"fe",
          5944 => x"fe",
          5945 => x"81",
          5946 => x"80",
          5947 => x"80",
          5948 => x"79",
          5949 => x"38",
          5950 => x"90",
          5951 => x"78",
          5952 => x"38",
          5953 => x"83",
          5954 => x"81",
          5955 => x"fe",
          5956 => x"a0",
          5957 => x"61",
          5958 => x"63",
          5959 => x"3f",
          5960 => x"51",
          5961 => x"b7",
          5962 => x"11",
          5963 => x"05",
          5964 => x"e6",
          5965 => x"c0",
          5966 => x"f7",
          5967 => x"3d",
          5968 => x"53",
          5969 => x"51",
          5970 => x"3f",
          5971 => x"08",
          5972 => x"38",
          5973 => x"80",
          5974 => x"79",
          5975 => x"05",
          5976 => x"fe",
          5977 => x"fe",
          5978 => x"fe",
          5979 => x"81",
          5980 => x"e0",
          5981 => x"39",
          5982 => x"54",
          5983 => x"80",
          5984 => x"a1",
          5985 => x"52",
          5986 => x"f9",
          5987 => x"45",
          5988 => x"78",
          5989 => x"ea",
          5990 => x"27",
          5991 => x"3d",
          5992 => x"53",
          5993 => x"51",
          5994 => x"3f",
          5995 => x"08",
          5996 => x"38",
          5997 => x"80",
          5998 => x"79",
          5999 => x"05",
          6000 => x"39",
          6001 => x"51",
          6002 => x"3f",
          6003 => x"b7",
          6004 => x"11",
          6005 => x"05",
          6006 => x"b0",
          6007 => x"c0",
          6008 => x"f6",
          6009 => x"3d",
          6010 => x"53",
          6011 => x"51",
          6012 => x"3f",
          6013 => x"08",
          6014 => x"38",
          6015 => x"be",
          6016 => x"70",
          6017 => x"23",
          6018 => x"3d",
          6019 => x"53",
          6020 => x"51",
          6021 => x"3f",
          6022 => x"08",
          6023 => x"e2",
          6024 => x"22",
          6025 => x"d8",
          6026 => x"f7",
          6027 => x"f8",
          6028 => x"fe",
          6029 => x"79",
          6030 => x"59",
          6031 => x"f5",
          6032 => x"9f",
          6033 => x"60",
          6034 => x"d5",
          6035 => x"fe",
          6036 => x"fe",
          6037 => x"fe",
          6038 => x"81",
          6039 => x"80",
          6040 => x"60",
          6041 => x"05",
          6042 => x"82",
          6043 => x"78",
          6044 => x"39",
          6045 => x"51",
          6046 => x"3f",
          6047 => x"b7",
          6048 => x"11",
          6049 => x"05",
          6050 => x"80",
          6051 => x"c0",
          6052 => x"f4",
          6053 => x"3d",
          6054 => x"53",
          6055 => x"51",
          6056 => x"3f",
          6057 => x"08",
          6058 => x"38",
          6059 => x"0c",
          6060 => x"05",
          6061 => x"fe",
          6062 => x"fe",
          6063 => x"fe",
          6064 => x"81",
          6065 => x"e4",
          6066 => x"39",
          6067 => x"54",
          6068 => x"a0",
          6069 => x"cd",
          6070 => x"52",
          6071 => x"f7",
          6072 => x"45",
          6073 => x"78",
          6074 => x"96",
          6075 => x"27",
          6076 => x"3d",
          6077 => x"53",
          6078 => x"51",
          6079 => x"3f",
          6080 => x"08",
          6081 => x"38",
          6082 => x"0c",
          6083 => x"05",
          6084 => x"39",
          6085 => x"51",
          6086 => x"3f",
          6087 => x"b7",
          6088 => x"11",
          6089 => x"05",
          6090 => x"ee",
          6091 => x"c0",
          6092 => x"38",
          6093 => x"33",
          6094 => x"2e",
          6095 => x"db",
          6096 => x"80",
          6097 => x"db",
          6098 => x"78",
          6099 => x"38",
          6100 => x"08",
          6101 => x"81",
          6102 => x"59",
          6103 => x"88",
          6104 => x"9c",
          6105 => x"39",
          6106 => x"33",
          6107 => x"2e",
          6108 => x"db",
          6109 => x"9a",
          6110 => x"d2",
          6111 => x"80",
          6112 => x"81",
          6113 => x"44",
          6114 => x"db",
          6115 => x"80",
          6116 => x"3d",
          6117 => x"53",
          6118 => x"51",
          6119 => x"3f",
          6120 => x"08",
          6121 => x"81",
          6122 => x"59",
          6123 => x"89",
          6124 => x"90",
          6125 => x"cc",
          6126 => x"d5",
          6127 => x"80",
          6128 => x"81",
          6129 => x"43",
          6130 => x"db",
          6131 => x"78",
          6132 => x"38",
          6133 => x"08",
          6134 => x"81",
          6135 => x"59",
          6136 => x"88",
          6137 => x"a8",
          6138 => x"39",
          6139 => x"33",
          6140 => x"2e",
          6141 => x"db",
          6142 => x"88",
          6143 => x"bc",
          6144 => x"43",
          6145 => x"ec",
          6146 => x"f8",
          6147 => x"f6",
          6148 => x"de",
          6149 => x"38",
          6150 => x"08",
          6151 => x"ac",
          6152 => x"9d",
          6153 => x"79",
          6154 => x"38",
          6155 => x"78",
          6156 => x"81",
          6157 => x"78",
          6158 => x"81",
          6159 => x"fe",
          6160 => x"84",
          6161 => x"39",
          6162 => x"51",
          6163 => x"d8",
          6164 => x"ed",
          6165 => x"51",
          6166 => x"3f",
          6167 => x"81",
          6168 => x"fe",
          6169 => x"a2",
          6170 => x"ad",
          6171 => x"39",
          6172 => x"0b",
          6173 => x"84",
          6174 => x"81",
          6175 => x"94",
          6176 => x"d8",
          6177 => x"ed",
          6178 => x"f6",
          6179 => x"90",
          6180 => x"ad",
          6181 => x"83",
          6182 => x"94",
          6183 => x"80",
          6184 => x"c0",
          6185 => x"f0",
          6186 => x"3d",
          6187 => x"53",
          6188 => x"51",
          6189 => x"3f",
          6190 => x"08",
          6191 => x"c2",
          6192 => x"81",
          6193 => x"fe",
          6194 => x"63",
          6195 => x"b7",
          6196 => x"11",
          6197 => x"05",
          6198 => x"be",
          6199 => x"c0",
          6200 => x"f0",
          6201 => x"52",
          6202 => x"51",
          6203 => x"3f",
          6204 => x"2d",
          6205 => x"08",
          6206 => x"c0",
          6207 => x"f0",
          6208 => x"de",
          6209 => x"81",
          6210 => x"fe",
          6211 => x"ef",
          6212 => x"d9",
          6213 => x"ec",
          6214 => x"bd",
          6215 => x"e2",
          6216 => x"94",
          6217 => x"99",
          6218 => x"ff",
          6219 => x"e6",
          6220 => x"ce",
          6221 => x"33",
          6222 => x"80",
          6223 => x"38",
          6224 => x"81",
          6225 => x"70",
          6226 => x"5a",
          6227 => x"81",
          6228 => x"3d",
          6229 => x"51",
          6230 => x"3f",
          6231 => x"08",
          6232 => x"7b",
          6233 => x"38",
          6234 => x"89",
          6235 => x"2e",
          6236 => x"cd",
          6237 => x"2e",
          6238 => x"c5",
          6239 => x"a8",
          6240 => x"81",
          6241 => x"80",
          6242 => x"b0",
          6243 => x"ff",
          6244 => x"fe",
          6245 => x"bb",
          6246 => x"d0",
          6247 => x"ff",
          6248 => x"fe",
          6249 => x"ab",
          6250 => x"81",
          6251 => x"80",
          6252 => x"c0",
          6253 => x"ff",
          6254 => x"fe",
          6255 => x"93",
          6256 => x"80",
          6257 => x"cc",
          6258 => x"ff",
          6259 => x"fe",
          6260 => x"81",
          6261 => x"81",
          6262 => x"80",
          6263 => x"11",
          6264 => x"55",
          6265 => x"80",
          6266 => x"80",
          6267 => x"3d",
          6268 => x"51",
          6269 => x"81",
          6270 => x"81",
          6271 => x"09",
          6272 => x"72",
          6273 => x"51",
          6274 => x"7b",
          6275 => x"38",
          6276 => x"8d",
          6277 => x"70",
          6278 => x"5d",
          6279 => x"c3",
          6280 => x"32",
          6281 => x"07",
          6282 => x"38",
          6283 => x"09",
          6284 => x"ce",
          6285 => x"d4",
          6286 => x"e9",
          6287 => x"39",
          6288 => x"80",
          6289 => x"f4",
          6290 => x"94",
          6291 => x"54",
          6292 => x"80",
          6293 => x"fe",
          6294 => x"81",
          6295 => x"90",
          6296 => x"55",
          6297 => x"80",
          6298 => x"fe",
          6299 => x"72",
          6300 => x"08",
          6301 => x"87",
          6302 => x"70",
          6303 => x"87",
          6304 => x"72",
          6305 => x"f1",
          6306 => x"c0",
          6307 => x"75",
          6308 => x"87",
          6309 => x"73",
          6310 => x"dd",
          6311 => x"de",
          6312 => x"75",
          6313 => x"83",
          6314 => x"94",
          6315 => x"80",
          6316 => x"c0",
          6317 => x"9f",
          6318 => x"de",
          6319 => x"bb",
          6320 => x"d4",
          6321 => x"9e",
          6322 => x"c5",
          6323 => x"e4",
          6324 => x"ce",
          6325 => x"f0",
          6326 => x"e5",
          6327 => x"e1",
          6328 => x"a8",
          6329 => x"e6",
          6330 => x"c6",
          6331 => x"00",
          6332 => x"ff",
          6333 => x"00",
          6334 => x"ff",
          6335 => x"ff",
          6336 => x"00",
          6337 => x"00",
          6338 => x"00",
          6339 => x"00",
          6340 => x"00",
          6341 => x"00",
          6342 => x"00",
          6343 => x"00",
          6344 => x"00",
          6345 => x"00",
          6346 => x"00",
          6347 => x"00",
          6348 => x"00",
          6349 => x"00",
          6350 => x"00",
          6351 => x"00",
          6352 => x"00",
          6353 => x"00",
          6354 => x"00",
          6355 => x"00",
          6356 => x"00",
          6357 => x"00",
          6358 => x"00",
          6359 => x"00",
          6360 => x"00",
          6361 => x"64",
          6362 => x"2f",
          6363 => x"25",
          6364 => x"64",
          6365 => x"2e",
          6366 => x"64",
          6367 => x"6f",
          6368 => x"6f",
          6369 => x"67",
          6370 => x"74",
          6371 => x"00",
          6372 => x"28",
          6373 => x"6d",
          6374 => x"43",
          6375 => x"6e",
          6376 => x"29",
          6377 => x"0a",
          6378 => x"69",
          6379 => x"20",
          6380 => x"6c",
          6381 => x"6e",
          6382 => x"3a",
          6383 => x"20",
          6384 => x"42",
          6385 => x"52",
          6386 => x"20",
          6387 => x"38",
          6388 => x"30",
          6389 => x"2e",
          6390 => x"20",
          6391 => x"44",
          6392 => x"20",
          6393 => x"20",
          6394 => x"38",
          6395 => x"30",
          6396 => x"2e",
          6397 => x"20",
          6398 => x"4e",
          6399 => x"42",
          6400 => x"20",
          6401 => x"38",
          6402 => x"30",
          6403 => x"2e",
          6404 => x"20",
          6405 => x"52",
          6406 => x"20",
          6407 => x"20",
          6408 => x"38",
          6409 => x"30",
          6410 => x"2e",
          6411 => x"20",
          6412 => x"41",
          6413 => x"20",
          6414 => x"20",
          6415 => x"38",
          6416 => x"30",
          6417 => x"2e",
          6418 => x"20",
          6419 => x"44",
          6420 => x"52",
          6421 => x"20",
          6422 => x"76",
          6423 => x"73",
          6424 => x"30",
          6425 => x"2e",
          6426 => x"20",
          6427 => x"49",
          6428 => x"31",
          6429 => x"20",
          6430 => x"6d",
          6431 => x"20",
          6432 => x"30",
          6433 => x"2e",
          6434 => x"20",
          6435 => x"4e",
          6436 => x"43",
          6437 => x"20",
          6438 => x"61",
          6439 => x"6c",
          6440 => x"30",
          6441 => x"2e",
          6442 => x"20",
          6443 => x"49",
          6444 => x"4f",
          6445 => x"42",
          6446 => x"00",
          6447 => x"20",
          6448 => x"42",
          6449 => x"43",
          6450 => x"20",
          6451 => x"4f",
          6452 => x"0a",
          6453 => x"20",
          6454 => x"53",
          6455 => x"00",
          6456 => x"20",
          6457 => x"50",
          6458 => x"00",
          6459 => x"64",
          6460 => x"73",
          6461 => x"3a",
          6462 => x"20",
          6463 => x"50",
          6464 => x"65",
          6465 => x"20",
          6466 => x"74",
          6467 => x"41",
          6468 => x"65",
          6469 => x"3d",
          6470 => x"38",
          6471 => x"00",
          6472 => x"20",
          6473 => x"50",
          6474 => x"65",
          6475 => x"79",
          6476 => x"61",
          6477 => x"41",
          6478 => x"65",
          6479 => x"3d",
          6480 => x"38",
          6481 => x"00",
          6482 => x"20",
          6483 => x"74",
          6484 => x"20",
          6485 => x"72",
          6486 => x"64",
          6487 => x"73",
          6488 => x"20",
          6489 => x"3d",
          6490 => x"38",
          6491 => x"00",
          6492 => x"69",
          6493 => x"0a",
          6494 => x"20",
          6495 => x"50",
          6496 => x"64",
          6497 => x"20",
          6498 => x"20",
          6499 => x"20",
          6500 => x"20",
          6501 => x"3d",
          6502 => x"34",
          6503 => x"00",
          6504 => x"20",
          6505 => x"79",
          6506 => x"6d",
          6507 => x"6f",
          6508 => x"46",
          6509 => x"20",
          6510 => x"20",
          6511 => x"3d",
          6512 => x"2e",
          6513 => x"64",
          6514 => x"0a",
          6515 => x"20",
          6516 => x"44",
          6517 => x"20",
          6518 => x"63",
          6519 => x"72",
          6520 => x"20",
          6521 => x"20",
          6522 => x"3d",
          6523 => x"2e",
          6524 => x"64",
          6525 => x"0a",
          6526 => x"20",
          6527 => x"69",
          6528 => x"6f",
          6529 => x"53",
          6530 => x"4d",
          6531 => x"6f",
          6532 => x"46",
          6533 => x"3d",
          6534 => x"2e",
          6535 => x"64",
          6536 => x"0a",
          6537 => x"6d",
          6538 => x"00",
          6539 => x"65",
          6540 => x"6d",
          6541 => x"6c",
          6542 => x"00",
          6543 => x"56",
          6544 => x"56",
          6545 => x"6e",
          6546 => x"6e",
          6547 => x"77",
          6548 => x"44",
          6549 => x"2a",
          6550 => x"3b",
          6551 => x"3f",
          6552 => x"7f",
          6553 => x"41",
          6554 => x"41",
          6555 => x"00",
          6556 => x"fe",
          6557 => x"44",
          6558 => x"2e",
          6559 => x"4f",
          6560 => x"4d",
          6561 => x"20",
          6562 => x"54",
          6563 => x"20",
          6564 => x"4f",
          6565 => x"4d",
          6566 => x"20",
          6567 => x"54",
          6568 => x"20",
          6569 => x"00",
          6570 => x"00",
          6571 => x"00",
          6572 => x"00",
          6573 => x"9a",
          6574 => x"41",
          6575 => x"45",
          6576 => x"49",
          6577 => x"92",
          6578 => x"4f",
          6579 => x"99",
          6580 => x"9d",
          6581 => x"49",
          6582 => x"a5",
          6583 => x"a9",
          6584 => x"ad",
          6585 => x"b1",
          6586 => x"b5",
          6587 => x"b9",
          6588 => x"bd",
          6589 => x"c1",
          6590 => x"c5",
          6591 => x"c9",
          6592 => x"cd",
          6593 => x"d1",
          6594 => x"d5",
          6595 => x"d9",
          6596 => x"dd",
          6597 => x"e1",
          6598 => x"e5",
          6599 => x"e9",
          6600 => x"ed",
          6601 => x"f1",
          6602 => x"f5",
          6603 => x"f9",
          6604 => x"fd",
          6605 => x"2e",
          6606 => x"5b",
          6607 => x"22",
          6608 => x"3e",
          6609 => x"00",
          6610 => x"01",
          6611 => x"10",
          6612 => x"00",
          6613 => x"00",
          6614 => x"01",
          6615 => x"04",
          6616 => x"10",
          6617 => x"00",
          6618 => x"69",
          6619 => x"00",
          6620 => x"69",
          6621 => x"6c",
          6622 => x"69",
          6623 => x"00",
          6624 => x"6c",
          6625 => x"00",
          6626 => x"65",
          6627 => x"00",
          6628 => x"63",
          6629 => x"72",
          6630 => x"64",
          6631 => x"00",
          6632 => x"73",
          6633 => x"00",
          6634 => x"65",
          6635 => x"65",
          6636 => x"65",
          6637 => x"69",
          6638 => x"69",
          6639 => x"66",
          6640 => x"66",
          6641 => x"61",
          6642 => x"00",
          6643 => x"6d",
          6644 => x"65",
          6645 => x"72",
          6646 => x"65",
          6647 => x"00",
          6648 => x"6e",
          6649 => x"00",
          6650 => x"65",
          6651 => x"00",
          6652 => x"69",
          6653 => x"45",
          6654 => x"72",
          6655 => x"6e",
          6656 => x"6e",
          6657 => x"65",
          6658 => x"72",
          6659 => x"00",
          6660 => x"69",
          6661 => x"6e",
          6662 => x"72",
          6663 => x"79",
          6664 => x"00",
          6665 => x"6f",
          6666 => x"6c",
          6667 => x"6f",
          6668 => x"2e",
          6669 => x"6f",
          6670 => x"74",
          6671 => x"6f",
          6672 => x"2e",
          6673 => x"6e",
          6674 => x"69",
          6675 => x"69",
          6676 => x"61",
          6677 => x"0a",
          6678 => x"63",
          6679 => x"73",
          6680 => x"6e",
          6681 => x"2e",
          6682 => x"69",
          6683 => x"61",
          6684 => x"61",
          6685 => x"65",
          6686 => x"74",
          6687 => x"00",
          6688 => x"69",
          6689 => x"68",
          6690 => x"6c",
          6691 => x"6e",
          6692 => x"69",
          6693 => x"00",
          6694 => x"44",
          6695 => x"20",
          6696 => x"74",
          6697 => x"72",
          6698 => x"63",
          6699 => x"2e",
          6700 => x"72",
          6701 => x"20",
          6702 => x"62",
          6703 => x"69",
          6704 => x"6e",
          6705 => x"69",
          6706 => x"00",
          6707 => x"69",
          6708 => x"6e",
          6709 => x"65",
          6710 => x"6c",
          6711 => x"0a",
          6712 => x"6f",
          6713 => x"6d",
          6714 => x"69",
          6715 => x"20",
          6716 => x"65",
          6717 => x"74",
          6718 => x"66",
          6719 => x"64",
          6720 => x"20",
          6721 => x"6b",
          6722 => x"00",
          6723 => x"6f",
          6724 => x"74",
          6725 => x"6f",
          6726 => x"64",
          6727 => x"00",
          6728 => x"69",
          6729 => x"75",
          6730 => x"6f",
          6731 => x"61",
          6732 => x"6e",
          6733 => x"6e",
          6734 => x"6c",
          6735 => x"0a",
          6736 => x"69",
          6737 => x"69",
          6738 => x"6f",
          6739 => x"64",
          6740 => x"00",
          6741 => x"6e",
          6742 => x"66",
          6743 => x"65",
          6744 => x"6d",
          6745 => x"72",
          6746 => x"00",
          6747 => x"6f",
          6748 => x"61",
          6749 => x"6f",
          6750 => x"20",
          6751 => x"65",
          6752 => x"00",
          6753 => x"61",
          6754 => x"65",
          6755 => x"73",
          6756 => x"63",
          6757 => x"65",
          6758 => x"0a",
          6759 => x"75",
          6760 => x"73",
          6761 => x"00",
          6762 => x"6e",
          6763 => x"77",
          6764 => x"72",
          6765 => x"2e",
          6766 => x"25",
          6767 => x"62",
          6768 => x"73",
          6769 => x"20",
          6770 => x"25",
          6771 => x"62",
          6772 => x"73",
          6773 => x"63",
          6774 => x"00",
          6775 => x"30",
          6776 => x"00",
          6777 => x"20",
          6778 => x"30",
          6779 => x"00",
          6780 => x"20",
          6781 => x"20",
          6782 => x"00",
          6783 => x"30",
          6784 => x"00",
          6785 => x"20",
          6786 => x"7c",
          6787 => x"0d",
          6788 => x"65",
          6789 => x"00",
          6790 => x"50",
          6791 => x"00",
          6792 => x"2a",
          6793 => x"73",
          6794 => x"00",
          6795 => x"39",
          6796 => x"2f",
          6797 => x"39",
          6798 => x"31",
          6799 => x"00",
          6800 => x"5a",
          6801 => x"20",
          6802 => x"20",
          6803 => x"78",
          6804 => x"73",
          6805 => x"20",
          6806 => x"0a",
          6807 => x"50",
          6808 => x"20",
          6809 => x"65",
          6810 => x"70",
          6811 => x"61",
          6812 => x"65",
          6813 => x"00",
          6814 => x"69",
          6815 => x"20",
          6816 => x"65",
          6817 => x"70",
          6818 => x"00",
          6819 => x"53",
          6820 => x"6e",
          6821 => x"72",
          6822 => x"0a",
          6823 => x"4f",
          6824 => x"20",
          6825 => x"69",
          6826 => x"72",
          6827 => x"74",
          6828 => x"4f",
          6829 => x"20",
          6830 => x"69",
          6831 => x"72",
          6832 => x"74",
          6833 => x"41",
          6834 => x"20",
          6835 => x"69",
          6836 => x"72",
          6837 => x"74",
          6838 => x"41",
          6839 => x"20",
          6840 => x"69",
          6841 => x"72",
          6842 => x"74",
          6843 => x"41",
          6844 => x"20",
          6845 => x"69",
          6846 => x"72",
          6847 => x"74",
          6848 => x"41",
          6849 => x"20",
          6850 => x"69",
          6851 => x"72",
          6852 => x"74",
          6853 => x"65",
          6854 => x"6e",
          6855 => x"70",
          6856 => x"6d",
          6857 => x"2e",
          6858 => x"00",
          6859 => x"6e",
          6860 => x"69",
          6861 => x"74",
          6862 => x"72",
          6863 => x"0a",
          6864 => x"75",
          6865 => x"78",
          6866 => x"62",
          6867 => x"00",
          6868 => x"3a",
          6869 => x"61",
          6870 => x"64",
          6871 => x"20",
          6872 => x"74",
          6873 => x"69",
          6874 => x"73",
          6875 => x"61",
          6876 => x"30",
          6877 => x"6c",
          6878 => x"65",
          6879 => x"69",
          6880 => x"61",
          6881 => x"6c",
          6882 => x"0a",
          6883 => x"20",
          6884 => x"61",
          6885 => x"69",
          6886 => x"69",
          6887 => x"00",
          6888 => x"6e",
          6889 => x"61",
          6890 => x"65",
          6891 => x"00",
          6892 => x"61",
          6893 => x"64",
          6894 => x"20",
          6895 => x"74",
          6896 => x"69",
          6897 => x"0a",
          6898 => x"63",
          6899 => x"0a",
          6900 => x"75",
          6901 => x"6c",
          6902 => x"69",
          6903 => x"2e",
          6904 => x"00",
          6905 => x"75",
          6906 => x"4d",
          6907 => x"72",
          6908 => x"00",
          6909 => x"43",
          6910 => x"6c",
          6911 => x"2e",
          6912 => x"30",
          6913 => x"25",
          6914 => x"2d",
          6915 => x"3f",
          6916 => x"00",
          6917 => x"30",
          6918 => x"25",
          6919 => x"2d",
          6920 => x"30",
          6921 => x"25",
          6922 => x"2d",
          6923 => x"65",
          6924 => x"68",
          6925 => x"2e",
          6926 => x"00",
          6927 => x"30",
          6928 => x"2d",
          6929 => x"38",
          6930 => x"00",
          6931 => x"69",
          6932 => x"6c",
          6933 => x"20",
          6934 => x"65",
          6935 => x"70",
          6936 => x"00",
          6937 => x"6e",
          6938 => x"69",
          6939 => x"69",
          6940 => x"72",
          6941 => x"74",
          6942 => x"00",
          6943 => x"69",
          6944 => x"6c",
          6945 => x"75",
          6946 => x"20",
          6947 => x"6f",
          6948 => x"6e",
          6949 => x"69",
          6950 => x"75",
          6951 => x"20",
          6952 => x"6f",
          6953 => x"78",
          6954 => x"74",
          6955 => x"20",
          6956 => x"65",
          6957 => x"25",
          6958 => x"20",
          6959 => x"0a",
          6960 => x"61",
          6961 => x"6e",
          6962 => x"6f",
          6963 => x"40",
          6964 => x"38",
          6965 => x"2e",
          6966 => x"00",
          6967 => x"61",
          6968 => x"72",
          6969 => x"72",
          6970 => x"20",
          6971 => x"65",
          6972 => x"64",
          6973 => x"00",
          6974 => x"65",
          6975 => x"72",
          6976 => x"67",
          6977 => x"70",
          6978 => x"61",
          6979 => x"6e",
          6980 => x"0a",
          6981 => x"6f",
          6982 => x"72",
          6983 => x"6f",
          6984 => x"67",
          6985 => x"0a",
          6986 => x"50",
          6987 => x"69",
          6988 => x"64",
          6989 => x"73",
          6990 => x"2e",
          6991 => x"00",
          6992 => x"64",
          6993 => x"73",
          6994 => x"00",
          6995 => x"64",
          6996 => x"73",
          6997 => x"61",
          6998 => x"6f",
          6999 => x"6e",
          7000 => x"00",
          7001 => x"75",
          7002 => x"6e",
          7003 => x"2e",
          7004 => x"6e",
          7005 => x"69",
          7006 => x"69",
          7007 => x"72",
          7008 => x"74",
          7009 => x"2e",
          7010 => x"00",
          7011 => x"00",
          7012 => x"00",
          7013 => x"00",
          7014 => x"00",
          7015 => x"01",
          7016 => x"00",
          7017 => x"01",
          7018 => x"81",
          7019 => x"00",
          7020 => x"7f",
          7021 => x"00",
          7022 => x"00",
          7023 => x"00",
          7024 => x"00",
          7025 => x"f5",
          7026 => x"f5",
          7027 => x"f5",
          7028 => x"00",
          7029 => x"01",
          7030 => x"01",
          7031 => x"01",
          7032 => x"00",
          7033 => x"00",
          7034 => x"00",
          7035 => x"00",
          7036 => x"00",
          7037 => x"02",
          7038 => x"00",
          7039 => x"00",
          7040 => x"00",
          7041 => x"04",
          7042 => x"00",
          7043 => x"00",
          7044 => x"00",
          7045 => x"14",
          7046 => x"00",
          7047 => x"00",
          7048 => x"00",
          7049 => x"2b",
          7050 => x"00",
          7051 => x"00",
          7052 => x"00",
          7053 => x"30",
          7054 => x"00",
          7055 => x"00",
          7056 => x"00",
          7057 => x"3c",
          7058 => x"00",
          7059 => x"00",
          7060 => x"00",
          7061 => x"40",
          7062 => x"00",
          7063 => x"00",
          7064 => x"00",
          7065 => x"45",
          7066 => x"00",
          7067 => x"00",
          7068 => x"00",
          7069 => x"41",
          7070 => x"00",
          7071 => x"00",
          7072 => x"00",
          7073 => x"42",
          7074 => x"00",
          7075 => x"00",
          7076 => x"00",
          7077 => x"43",
          7078 => x"00",
          7079 => x"00",
          7080 => x"00",
          7081 => x"50",
          7082 => x"00",
          7083 => x"00",
          7084 => x"00",
          7085 => x"51",
          7086 => x"00",
          7087 => x"00",
          7088 => x"00",
          7089 => x"54",
          7090 => x"00",
          7091 => x"00",
          7092 => x"00",
          7093 => x"55",
          7094 => x"00",
          7095 => x"00",
          7096 => x"00",
          7097 => x"79",
          7098 => x"00",
          7099 => x"00",
          7100 => x"00",
          7101 => x"78",
          7102 => x"00",
          7103 => x"00",
          7104 => x"00",
          7105 => x"82",
          7106 => x"00",
          7107 => x"00",
          7108 => x"00",
          7109 => x"83",
          7110 => x"00",
          7111 => x"00",
          7112 => x"00",
          7113 => x"85",
          7114 => x"00",
          7115 => x"00",
          7116 => x"00",
          7117 => x"87",
          7118 => x"00",
          7119 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"d8",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"bc",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"f0",
           163 => x"10",
           164 => x"06",
           165 => x"92",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"dd",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"c9",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"94",
           269 => x"0b",
           270 => x"0b",
           271 => x"b2",
           272 => x"0b",
           273 => x"0b",
           274 => x"d0",
           275 => x"0b",
           276 => x"0b",
           277 => x"ee",
           278 => x"0b",
           279 => x"0b",
           280 => x"8c",
           281 => x"0b",
           282 => x"0b",
           283 => x"aa",
           284 => x"0b",
           285 => x"0b",
           286 => x"c8",
           287 => x"0b",
           288 => x"0b",
           289 => x"e6",
           290 => x"0b",
           291 => x"0b",
           292 => x"84",
           293 => x"0b",
           294 => x"0b",
           295 => x"a4",
           296 => x"0b",
           297 => x"0b",
           298 => x"c4",
           299 => x"0b",
           300 => x"0b",
           301 => x"e4",
           302 => x"0b",
           303 => x"0b",
           304 => x"84",
           305 => x"0b",
           306 => x"0b",
           307 => x"a4",
           308 => x"0b",
           309 => x"0b",
           310 => x"c4",
           311 => x"0b",
           312 => x"0b",
           313 => x"e4",
           314 => x"0b",
           315 => x"0b",
           316 => x"84",
           317 => x"0b",
           318 => x"0b",
           319 => x"a4",
           320 => x"0b",
           321 => x"0b",
           322 => x"c4",
           323 => x"0b",
           324 => x"0b",
           325 => x"e4",
           326 => x"0b",
           327 => x"0b",
           328 => x"84",
           329 => x"0b",
           330 => x"0b",
           331 => x"a3",
           332 => x"0b",
           333 => x"0b",
           334 => x"c1",
           335 => x"0b",
           336 => x"0b",
           337 => x"df",
           338 => x"0b",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"81",
           388 => x"82",
           389 => x"81",
           390 => x"ad",
           391 => x"de",
           392 => x"80",
           393 => x"de",
           394 => x"a1",
           395 => x"cc",
           396 => x"90",
           397 => x"cc",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"81",
           403 => x"82",
           404 => x"81",
           405 => x"b5",
           406 => x"de",
           407 => x"80",
           408 => x"de",
           409 => x"e2",
           410 => x"cc",
           411 => x"90",
           412 => x"cc",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"81",
           418 => x"82",
           419 => x"81",
           420 => x"b4",
           421 => x"de",
           422 => x"80",
           423 => x"de",
           424 => x"b9",
           425 => x"cc",
           426 => x"90",
           427 => x"cc",
           428 => x"2d",
           429 => x"08",
           430 => x"04",
           431 => x"0c",
           432 => x"81",
           433 => x"82",
           434 => x"81",
           435 => x"a3",
           436 => x"de",
           437 => x"80",
           438 => x"de",
           439 => x"a8",
           440 => x"cc",
           441 => x"90",
           442 => x"cc",
           443 => x"2d",
           444 => x"08",
           445 => x"04",
           446 => x"0c",
           447 => x"81",
           448 => x"82",
           449 => x"81",
           450 => x"80",
           451 => x"81",
           452 => x"82",
           453 => x"81",
           454 => x"80",
           455 => x"81",
           456 => x"82",
           457 => x"81",
           458 => x"80",
           459 => x"81",
           460 => x"82",
           461 => x"81",
           462 => x"80",
           463 => x"81",
           464 => x"82",
           465 => x"81",
           466 => x"80",
           467 => x"81",
           468 => x"82",
           469 => x"81",
           470 => x"81",
           471 => x"81",
           472 => x"82",
           473 => x"81",
           474 => x"80",
           475 => x"81",
           476 => x"82",
           477 => x"81",
           478 => x"80",
           479 => x"81",
           480 => x"82",
           481 => x"81",
           482 => x"81",
           483 => x"81",
           484 => x"82",
           485 => x"81",
           486 => x"81",
           487 => x"81",
           488 => x"82",
           489 => x"81",
           490 => x"81",
           491 => x"81",
           492 => x"82",
           493 => x"81",
           494 => x"81",
           495 => x"81",
           496 => x"82",
           497 => x"81",
           498 => x"81",
           499 => x"81",
           500 => x"82",
           501 => x"81",
           502 => x"81",
           503 => x"81",
           504 => x"82",
           505 => x"81",
           506 => x"81",
           507 => x"81",
           508 => x"82",
           509 => x"81",
           510 => x"81",
           511 => x"81",
           512 => x"82",
           513 => x"81",
           514 => x"80",
           515 => x"81",
           516 => x"82",
           517 => x"81",
           518 => x"80",
           519 => x"81",
           520 => x"82",
           521 => x"81",
           522 => x"80",
           523 => x"81",
           524 => x"82",
           525 => x"81",
           526 => x"81",
           527 => x"81",
           528 => x"82",
           529 => x"81",
           530 => x"81",
           531 => x"81",
           532 => x"82",
           533 => x"81",
           534 => x"81",
           535 => x"81",
           536 => x"82",
           537 => x"81",
           538 => x"81",
           539 => x"81",
           540 => x"82",
           541 => x"81",
           542 => x"80",
           543 => x"81",
           544 => x"82",
           545 => x"81",
           546 => x"81",
           547 => x"81",
           548 => x"82",
           549 => x"81",
           550 => x"bb",
           551 => x"de",
           552 => x"80",
           553 => x"de",
           554 => x"83",
           555 => x"cc",
           556 => x"90",
           557 => x"cc",
           558 => x"2d",
           559 => x"08",
           560 => x"04",
           561 => x"0c",
           562 => x"81",
           563 => x"82",
           564 => x"81",
           565 => x"9c",
           566 => x"de",
           567 => x"80",
           568 => x"de",
           569 => x"a0",
           570 => x"cc",
           571 => x"90",
           572 => x"cc",
           573 => x"ff",
           574 => x"cc",
           575 => x"90",
           576 => x"10",
           577 => x"10",
           578 => x"10",
           579 => x"10",
           580 => x"10",
           581 => x"10",
           582 => x"10",
           583 => x"10",
           584 => x"51",
           585 => x"73",
           586 => x"73",
           587 => x"81",
           588 => x"10",
           589 => x"07",
           590 => x"0c",
           591 => x"72",
           592 => x"81",
           593 => x"09",
           594 => x"71",
           595 => x"0a",
           596 => x"72",
           597 => x"51",
           598 => x"81",
           599 => x"81",
           600 => x"8e",
           601 => x"70",
           602 => x"0c",
           603 => x"92",
           604 => x"81",
           605 => x"be",
           606 => x"de",
           607 => x"81",
           608 => x"fd",
           609 => x"53",
           610 => x"08",
           611 => x"52",
           612 => x"08",
           613 => x"51",
           614 => x"81",
           615 => x"70",
           616 => x"0c",
           617 => x"0d",
           618 => x"0c",
           619 => x"cc",
           620 => x"de",
           621 => x"3d",
           622 => x"81",
           623 => x"8c",
           624 => x"81",
           625 => x"88",
           626 => x"83",
           627 => x"de",
           628 => x"81",
           629 => x"54",
           630 => x"81",
           631 => x"04",
           632 => x"08",
           633 => x"cc",
           634 => x"0d",
           635 => x"de",
           636 => x"05",
           637 => x"cc",
           638 => x"08",
           639 => x"38",
           640 => x"08",
           641 => x"30",
           642 => x"08",
           643 => x"80",
           644 => x"cc",
           645 => x"0c",
           646 => x"08",
           647 => x"8a",
           648 => x"81",
           649 => x"f4",
           650 => x"de",
           651 => x"05",
           652 => x"cc",
           653 => x"0c",
           654 => x"08",
           655 => x"80",
           656 => x"81",
           657 => x"8c",
           658 => x"81",
           659 => x"8c",
           660 => x"0b",
           661 => x"08",
           662 => x"81",
           663 => x"fc",
           664 => x"38",
           665 => x"de",
           666 => x"05",
           667 => x"cc",
           668 => x"08",
           669 => x"08",
           670 => x"80",
           671 => x"cc",
           672 => x"08",
           673 => x"cc",
           674 => x"08",
           675 => x"3f",
           676 => x"08",
           677 => x"cc",
           678 => x"0c",
           679 => x"cc",
           680 => x"08",
           681 => x"38",
           682 => x"08",
           683 => x"30",
           684 => x"08",
           685 => x"81",
           686 => x"f8",
           687 => x"81",
           688 => x"54",
           689 => x"81",
           690 => x"04",
           691 => x"08",
           692 => x"cc",
           693 => x"0d",
           694 => x"de",
           695 => x"05",
           696 => x"cc",
           697 => x"08",
           698 => x"38",
           699 => x"08",
           700 => x"30",
           701 => x"08",
           702 => x"81",
           703 => x"cc",
           704 => x"0c",
           705 => x"08",
           706 => x"80",
           707 => x"81",
           708 => x"8c",
           709 => x"81",
           710 => x"8c",
           711 => x"53",
           712 => x"08",
           713 => x"52",
           714 => x"08",
           715 => x"51",
           716 => x"de",
           717 => x"81",
           718 => x"f8",
           719 => x"81",
           720 => x"fc",
           721 => x"2e",
           722 => x"de",
           723 => x"05",
           724 => x"de",
           725 => x"05",
           726 => x"cc",
           727 => x"08",
           728 => x"c0",
           729 => x"3d",
           730 => x"cc",
           731 => x"de",
           732 => x"81",
           733 => x"fd",
           734 => x"0b",
           735 => x"08",
           736 => x"80",
           737 => x"cc",
           738 => x"0c",
           739 => x"08",
           740 => x"81",
           741 => x"88",
           742 => x"b9",
           743 => x"cc",
           744 => x"08",
           745 => x"38",
           746 => x"de",
           747 => x"05",
           748 => x"38",
           749 => x"08",
           750 => x"10",
           751 => x"08",
           752 => x"81",
           753 => x"fc",
           754 => x"81",
           755 => x"fc",
           756 => x"b8",
           757 => x"cc",
           758 => x"08",
           759 => x"e1",
           760 => x"cc",
           761 => x"08",
           762 => x"08",
           763 => x"26",
           764 => x"de",
           765 => x"05",
           766 => x"cc",
           767 => x"08",
           768 => x"cc",
           769 => x"0c",
           770 => x"08",
           771 => x"81",
           772 => x"fc",
           773 => x"81",
           774 => x"f8",
           775 => x"de",
           776 => x"05",
           777 => x"81",
           778 => x"fc",
           779 => x"de",
           780 => x"05",
           781 => x"81",
           782 => x"8c",
           783 => x"95",
           784 => x"cc",
           785 => x"08",
           786 => x"38",
           787 => x"08",
           788 => x"70",
           789 => x"08",
           790 => x"51",
           791 => x"de",
           792 => x"05",
           793 => x"de",
           794 => x"05",
           795 => x"de",
           796 => x"05",
           797 => x"c0",
           798 => x"0d",
           799 => x"0c",
           800 => x"0d",
           801 => x"02",
           802 => x"05",
           803 => x"53",
           804 => x"27",
           805 => x"83",
           806 => x"80",
           807 => x"ff",
           808 => x"ff",
           809 => x"73",
           810 => x"05",
           811 => x"12",
           812 => x"2e",
           813 => x"ef",
           814 => x"de",
           815 => x"3d",
           816 => x"74",
           817 => x"07",
           818 => x"2b",
           819 => x"51",
           820 => x"a5",
           821 => x"70",
           822 => x"0c",
           823 => x"84",
           824 => x"72",
           825 => x"05",
           826 => x"71",
           827 => x"53",
           828 => x"52",
           829 => x"dd",
           830 => x"27",
           831 => x"71",
           832 => x"53",
           833 => x"52",
           834 => x"f2",
           835 => x"ff",
           836 => x"3d",
           837 => x"70",
           838 => x"06",
           839 => x"70",
           840 => x"73",
           841 => x"56",
           842 => x"08",
           843 => x"38",
           844 => x"52",
           845 => x"81",
           846 => x"54",
           847 => x"9d",
           848 => x"55",
           849 => x"09",
           850 => x"38",
           851 => x"14",
           852 => x"81",
           853 => x"56",
           854 => x"e5",
           855 => x"55",
           856 => x"06",
           857 => x"06",
           858 => x"81",
           859 => x"52",
           860 => x"0d",
           861 => x"70",
           862 => x"ff",
           863 => x"f8",
           864 => x"80",
           865 => x"51",
           866 => x"84",
           867 => x"71",
           868 => x"54",
           869 => x"2e",
           870 => x"75",
           871 => x"94",
           872 => x"81",
           873 => x"87",
           874 => x"fe",
           875 => x"52",
           876 => x"88",
           877 => x"86",
           878 => x"c0",
           879 => x"06",
           880 => x"14",
           881 => x"80",
           882 => x"71",
           883 => x"0c",
           884 => x"04",
           885 => x"77",
           886 => x"53",
           887 => x"80",
           888 => x"38",
           889 => x"70",
           890 => x"81",
           891 => x"81",
           892 => x"39",
           893 => x"39",
           894 => x"80",
           895 => x"81",
           896 => x"55",
           897 => x"2e",
           898 => x"55",
           899 => x"84",
           900 => x"38",
           901 => x"06",
           902 => x"2e",
           903 => x"88",
           904 => x"70",
           905 => x"34",
           906 => x"71",
           907 => x"de",
           908 => x"3d",
           909 => x"3d",
           910 => x"72",
           911 => x"91",
           912 => x"fc",
           913 => x"51",
           914 => x"81",
           915 => x"85",
           916 => x"83",
           917 => x"72",
           918 => x"0c",
           919 => x"04",
           920 => x"76",
           921 => x"ff",
           922 => x"81",
           923 => x"26",
           924 => x"83",
           925 => x"05",
           926 => x"70",
           927 => x"8a",
           928 => x"33",
           929 => x"70",
           930 => x"fe",
           931 => x"33",
           932 => x"70",
           933 => x"f2",
           934 => x"33",
           935 => x"70",
           936 => x"e6",
           937 => x"22",
           938 => x"74",
           939 => x"80",
           940 => x"13",
           941 => x"52",
           942 => x"26",
           943 => x"81",
           944 => x"98",
           945 => x"22",
           946 => x"bc",
           947 => x"33",
           948 => x"b8",
           949 => x"33",
           950 => x"b4",
           951 => x"33",
           952 => x"b0",
           953 => x"33",
           954 => x"ac",
           955 => x"33",
           956 => x"a8",
           957 => x"c0",
           958 => x"73",
           959 => x"a0",
           960 => x"87",
           961 => x"0c",
           962 => x"81",
           963 => x"86",
           964 => x"f3",
           965 => x"5b",
           966 => x"9c",
           967 => x"0c",
           968 => x"bc",
           969 => x"7b",
           970 => x"98",
           971 => x"79",
           972 => x"87",
           973 => x"08",
           974 => x"1c",
           975 => x"98",
           976 => x"79",
           977 => x"87",
           978 => x"08",
           979 => x"1c",
           980 => x"98",
           981 => x"79",
           982 => x"87",
           983 => x"08",
           984 => x"1c",
           985 => x"98",
           986 => x"79",
           987 => x"80",
           988 => x"83",
           989 => x"59",
           990 => x"ff",
           991 => x"1b",
           992 => x"1b",
           993 => x"1b",
           994 => x"1b",
           995 => x"1b",
           996 => x"83",
           997 => x"52",
           998 => x"51",
           999 => x"8f",
          1000 => x"ff",
          1001 => x"8f",
          1002 => x"30",
          1003 => x"51",
          1004 => x"0b",
          1005 => x"88",
          1006 => x"0d",
          1007 => x"0d",
          1008 => x"81",
          1009 => x"70",
          1010 => x"57",
          1011 => x"c0",
          1012 => x"74",
          1013 => x"38",
          1014 => x"94",
          1015 => x"70",
          1016 => x"81",
          1017 => x"52",
          1018 => x"8c",
          1019 => x"2a",
          1020 => x"51",
          1021 => x"38",
          1022 => x"70",
          1023 => x"51",
          1024 => x"8d",
          1025 => x"2a",
          1026 => x"51",
          1027 => x"be",
          1028 => x"ff",
          1029 => x"c0",
          1030 => x"70",
          1031 => x"38",
          1032 => x"90",
          1033 => x"0c",
          1034 => x"c0",
          1035 => x"0d",
          1036 => x"0d",
          1037 => x"33",
          1038 => x"db",
          1039 => x"81",
          1040 => x"55",
          1041 => x"94",
          1042 => x"80",
          1043 => x"87",
          1044 => x"51",
          1045 => x"96",
          1046 => x"06",
          1047 => x"70",
          1048 => x"38",
          1049 => x"70",
          1050 => x"51",
          1051 => x"72",
          1052 => x"81",
          1053 => x"70",
          1054 => x"38",
          1055 => x"70",
          1056 => x"51",
          1057 => x"38",
          1058 => x"06",
          1059 => x"94",
          1060 => x"80",
          1061 => x"87",
          1062 => x"52",
          1063 => x"87",
          1064 => x"f9",
          1065 => x"54",
          1066 => x"70",
          1067 => x"53",
          1068 => x"77",
          1069 => x"38",
          1070 => x"06",
          1071 => x"0b",
          1072 => x"33",
          1073 => x"06",
          1074 => x"58",
          1075 => x"84",
          1076 => x"2e",
          1077 => x"c0",
          1078 => x"70",
          1079 => x"2a",
          1080 => x"53",
          1081 => x"80",
          1082 => x"71",
          1083 => x"81",
          1084 => x"70",
          1085 => x"81",
          1086 => x"06",
          1087 => x"80",
          1088 => x"71",
          1089 => x"81",
          1090 => x"70",
          1091 => x"74",
          1092 => x"51",
          1093 => x"80",
          1094 => x"2e",
          1095 => x"c0",
          1096 => x"77",
          1097 => x"17",
          1098 => x"81",
          1099 => x"53",
          1100 => x"84",
          1101 => x"de",
          1102 => x"3d",
          1103 => x"3d",
          1104 => x"81",
          1105 => x"70",
          1106 => x"54",
          1107 => x"94",
          1108 => x"80",
          1109 => x"87",
          1110 => x"51",
          1111 => x"82",
          1112 => x"06",
          1113 => x"70",
          1114 => x"38",
          1115 => x"06",
          1116 => x"94",
          1117 => x"80",
          1118 => x"87",
          1119 => x"52",
          1120 => x"81",
          1121 => x"de",
          1122 => x"84",
          1123 => x"fe",
          1124 => x"0b",
          1125 => x"33",
          1126 => x"06",
          1127 => x"c0",
          1128 => x"70",
          1129 => x"38",
          1130 => x"94",
          1131 => x"70",
          1132 => x"81",
          1133 => x"51",
          1134 => x"80",
          1135 => x"72",
          1136 => x"51",
          1137 => x"80",
          1138 => x"2e",
          1139 => x"c0",
          1140 => x"71",
          1141 => x"2b",
          1142 => x"51",
          1143 => x"81",
          1144 => x"84",
          1145 => x"ff",
          1146 => x"c0",
          1147 => x"70",
          1148 => x"06",
          1149 => x"80",
          1150 => x"38",
          1151 => x"a4",
          1152 => x"8c",
          1153 => x"9e",
          1154 => x"db",
          1155 => x"c0",
          1156 => x"81",
          1157 => x"87",
          1158 => x"08",
          1159 => x"0c",
          1160 => x"9c",
          1161 => x"9c",
          1162 => x"9e",
          1163 => x"db",
          1164 => x"c0",
          1165 => x"81",
          1166 => x"87",
          1167 => x"08",
          1168 => x"0c",
          1169 => x"b4",
          1170 => x"ac",
          1171 => x"9e",
          1172 => x"db",
          1173 => x"c0",
          1174 => x"81",
          1175 => x"87",
          1176 => x"08",
          1177 => x"0c",
          1178 => x"c4",
          1179 => x"bc",
          1180 => x"9e",
          1181 => x"70",
          1182 => x"23",
          1183 => x"84",
          1184 => x"c4",
          1185 => x"9e",
          1186 => x"db",
          1187 => x"c0",
          1188 => x"81",
          1189 => x"81",
          1190 => x"d0",
          1191 => x"87",
          1192 => x"08",
          1193 => x"0a",
          1194 => x"52",
          1195 => x"83",
          1196 => x"71",
          1197 => x"34",
          1198 => x"c0",
          1199 => x"70",
          1200 => x"06",
          1201 => x"70",
          1202 => x"38",
          1203 => x"81",
          1204 => x"80",
          1205 => x"9e",
          1206 => x"90",
          1207 => x"51",
          1208 => x"80",
          1209 => x"81",
          1210 => x"db",
          1211 => x"0b",
          1212 => x"90",
          1213 => x"80",
          1214 => x"52",
          1215 => x"2e",
          1216 => x"52",
          1217 => x"d4",
          1218 => x"87",
          1219 => x"08",
          1220 => x"80",
          1221 => x"52",
          1222 => x"83",
          1223 => x"71",
          1224 => x"34",
          1225 => x"c0",
          1226 => x"70",
          1227 => x"06",
          1228 => x"70",
          1229 => x"38",
          1230 => x"81",
          1231 => x"80",
          1232 => x"9e",
          1233 => x"84",
          1234 => x"51",
          1235 => x"80",
          1236 => x"81",
          1237 => x"db",
          1238 => x"0b",
          1239 => x"90",
          1240 => x"80",
          1241 => x"52",
          1242 => x"2e",
          1243 => x"52",
          1244 => x"d8",
          1245 => x"87",
          1246 => x"08",
          1247 => x"80",
          1248 => x"52",
          1249 => x"83",
          1250 => x"71",
          1251 => x"34",
          1252 => x"c0",
          1253 => x"70",
          1254 => x"06",
          1255 => x"70",
          1256 => x"38",
          1257 => x"81",
          1258 => x"80",
          1259 => x"9e",
          1260 => x"a0",
          1261 => x"52",
          1262 => x"2e",
          1263 => x"52",
          1264 => x"db",
          1265 => x"9e",
          1266 => x"98",
          1267 => x"8a",
          1268 => x"51",
          1269 => x"dc",
          1270 => x"87",
          1271 => x"08",
          1272 => x"06",
          1273 => x"70",
          1274 => x"38",
          1275 => x"81",
          1276 => x"87",
          1277 => x"08",
          1278 => x"06",
          1279 => x"51",
          1280 => x"81",
          1281 => x"80",
          1282 => x"9e",
          1283 => x"88",
          1284 => x"52",
          1285 => x"83",
          1286 => x"71",
          1287 => x"34",
          1288 => x"90",
          1289 => x"06",
          1290 => x"81",
          1291 => x"83",
          1292 => x"fb",
          1293 => x"c6",
          1294 => x"86",
          1295 => x"d0",
          1296 => x"80",
          1297 => x"81",
          1298 => x"85",
          1299 => x"c7",
          1300 => x"ee",
          1301 => x"d2",
          1302 => x"80",
          1303 => x"81",
          1304 => x"81",
          1305 => x"11",
          1306 => x"c7",
          1307 => x"b6",
          1308 => x"d7",
          1309 => x"80",
          1310 => x"81",
          1311 => x"81",
          1312 => x"11",
          1313 => x"c7",
          1314 => x"9a",
          1315 => x"d4",
          1316 => x"80",
          1317 => x"81",
          1318 => x"81",
          1319 => x"11",
          1320 => x"c7",
          1321 => x"fe",
          1322 => x"d5",
          1323 => x"80",
          1324 => x"81",
          1325 => x"81",
          1326 => x"11",
          1327 => x"c8",
          1328 => x"e2",
          1329 => x"d6",
          1330 => x"80",
          1331 => x"81",
          1332 => x"81",
          1333 => x"11",
          1334 => x"c8",
          1335 => x"c6",
          1336 => x"db",
          1337 => x"80",
          1338 => x"81",
          1339 => x"52",
          1340 => x"51",
          1341 => x"81",
          1342 => x"54",
          1343 => x"8d",
          1344 => x"e0",
          1345 => x"c8",
          1346 => x"9a",
          1347 => x"dd",
          1348 => x"80",
          1349 => x"81",
          1350 => x"52",
          1351 => x"51",
          1352 => x"81",
          1353 => x"54",
          1354 => x"88",
          1355 => x"a8",
          1356 => x"3f",
          1357 => x"33",
          1358 => x"2e",
          1359 => x"c9",
          1360 => x"fe",
          1361 => x"d8",
          1362 => x"80",
          1363 => x"81",
          1364 => x"83",
          1365 => x"db",
          1366 => x"73",
          1367 => x"38",
          1368 => x"51",
          1369 => x"81",
          1370 => x"54",
          1371 => x"88",
          1372 => x"e0",
          1373 => x"3f",
          1374 => x"51",
          1375 => x"81",
          1376 => x"52",
          1377 => x"51",
          1378 => x"81",
          1379 => x"52",
          1380 => x"51",
          1381 => x"81",
          1382 => x"52",
          1383 => x"51",
          1384 => x"81",
          1385 => x"f5",
          1386 => x"db",
          1387 => x"81",
          1388 => x"88",
          1389 => x"db",
          1390 => x"bd",
          1391 => x"75",
          1392 => x"3f",
          1393 => x"08",
          1394 => x"29",
          1395 => x"54",
          1396 => x"c0",
          1397 => x"cb",
          1398 => x"ca",
          1399 => x"d7",
          1400 => x"80",
          1401 => x"81",
          1402 => x"56",
          1403 => x"52",
          1404 => x"86",
          1405 => x"c0",
          1406 => x"c0",
          1407 => x"31",
          1408 => x"de",
          1409 => x"81",
          1410 => x"88",
          1411 => x"db",
          1412 => x"73",
          1413 => x"38",
          1414 => x"08",
          1415 => x"c0",
          1416 => x"e6",
          1417 => x"de",
          1418 => x"84",
          1419 => x"71",
          1420 => x"81",
          1421 => x"52",
          1422 => x"51",
          1423 => x"81",
          1424 => x"81",
          1425 => x"3d",
          1426 => x"3d",
          1427 => x"05",
          1428 => x"52",
          1429 => x"aa",
          1430 => x"29",
          1431 => x"05",
          1432 => x"04",
          1433 => x"51",
          1434 => x"cc",
          1435 => x"39",
          1436 => x"51",
          1437 => x"cc",
          1438 => x"39",
          1439 => x"51",
          1440 => x"cc",
          1441 => x"9b",
          1442 => x"0d",
          1443 => x"80",
          1444 => x"0b",
          1445 => x"84",
          1446 => x"3d",
          1447 => x"96",
          1448 => x"52",
          1449 => x"0c",
          1450 => x"70",
          1451 => x"0c",
          1452 => x"3d",
          1453 => x"3d",
          1454 => x"96",
          1455 => x"81",
          1456 => x"52",
          1457 => x"73",
          1458 => x"db",
          1459 => x"70",
          1460 => x"0c",
          1461 => x"83",
          1462 => x"81",
          1463 => x"87",
          1464 => x"0c",
          1465 => x"0d",
          1466 => x"33",
          1467 => x"2e",
          1468 => x"85",
          1469 => x"ed",
          1470 => x"d8",
          1471 => x"80",
          1472 => x"72",
          1473 => x"de",
          1474 => x"05",
          1475 => x"0c",
          1476 => x"de",
          1477 => x"71",
          1478 => x"38",
          1479 => x"2d",
          1480 => x"04",
          1481 => x"02",
          1482 => x"81",
          1483 => x"76",
          1484 => x"0c",
          1485 => x"ad",
          1486 => x"de",
          1487 => x"3d",
          1488 => x"3d",
          1489 => x"73",
          1490 => x"ff",
          1491 => x"71",
          1492 => x"38",
          1493 => x"06",
          1494 => x"54",
          1495 => x"e7",
          1496 => x"0d",
          1497 => x"0d",
          1498 => x"d0",
          1499 => x"de",
          1500 => x"54",
          1501 => x"81",
          1502 => x"53",
          1503 => x"8e",
          1504 => x"ff",
          1505 => x"14",
          1506 => x"3f",
          1507 => x"81",
          1508 => x"86",
          1509 => x"ec",
          1510 => x"68",
          1511 => x"70",
          1512 => x"33",
          1513 => x"2e",
          1514 => x"75",
          1515 => x"81",
          1516 => x"38",
          1517 => x"70",
          1518 => x"33",
          1519 => x"75",
          1520 => x"81",
          1521 => x"81",
          1522 => x"75",
          1523 => x"81",
          1524 => x"82",
          1525 => x"81",
          1526 => x"56",
          1527 => x"09",
          1528 => x"38",
          1529 => x"71",
          1530 => x"81",
          1531 => x"59",
          1532 => x"9d",
          1533 => x"53",
          1534 => x"95",
          1535 => x"29",
          1536 => x"76",
          1537 => x"79",
          1538 => x"5b",
          1539 => x"e5",
          1540 => x"ec",
          1541 => x"70",
          1542 => x"25",
          1543 => x"32",
          1544 => x"72",
          1545 => x"73",
          1546 => x"58",
          1547 => x"73",
          1548 => x"38",
          1549 => x"79",
          1550 => x"5b",
          1551 => x"75",
          1552 => x"de",
          1553 => x"80",
          1554 => x"89",
          1555 => x"70",
          1556 => x"55",
          1557 => x"cf",
          1558 => x"38",
          1559 => x"24",
          1560 => x"80",
          1561 => x"8e",
          1562 => x"c3",
          1563 => x"73",
          1564 => x"81",
          1565 => x"99",
          1566 => x"c4",
          1567 => x"38",
          1568 => x"73",
          1569 => x"81",
          1570 => x"80",
          1571 => x"38",
          1572 => x"2e",
          1573 => x"f9",
          1574 => x"d8",
          1575 => x"38",
          1576 => x"77",
          1577 => x"08",
          1578 => x"80",
          1579 => x"55",
          1580 => x"8d",
          1581 => x"70",
          1582 => x"51",
          1583 => x"f5",
          1584 => x"2a",
          1585 => x"74",
          1586 => x"53",
          1587 => x"8f",
          1588 => x"fc",
          1589 => x"81",
          1590 => x"80",
          1591 => x"73",
          1592 => x"3f",
          1593 => x"56",
          1594 => x"27",
          1595 => x"a0",
          1596 => x"3f",
          1597 => x"84",
          1598 => x"33",
          1599 => x"93",
          1600 => x"95",
          1601 => x"91",
          1602 => x"8d",
          1603 => x"89",
          1604 => x"fb",
          1605 => x"86",
          1606 => x"2a",
          1607 => x"51",
          1608 => x"2e",
          1609 => x"84",
          1610 => x"86",
          1611 => x"78",
          1612 => x"08",
          1613 => x"32",
          1614 => x"72",
          1615 => x"51",
          1616 => x"74",
          1617 => x"38",
          1618 => x"88",
          1619 => x"7a",
          1620 => x"55",
          1621 => x"3d",
          1622 => x"52",
          1623 => x"cd",
          1624 => x"c0",
          1625 => x"06",
          1626 => x"52",
          1627 => x"3f",
          1628 => x"08",
          1629 => x"27",
          1630 => x"14",
          1631 => x"f8",
          1632 => x"87",
          1633 => x"81",
          1634 => x"b0",
          1635 => x"7d",
          1636 => x"5f",
          1637 => x"75",
          1638 => x"07",
          1639 => x"54",
          1640 => x"26",
          1641 => x"ff",
          1642 => x"84",
          1643 => x"06",
          1644 => x"80",
          1645 => x"96",
          1646 => x"e0",
          1647 => x"73",
          1648 => x"57",
          1649 => x"06",
          1650 => x"54",
          1651 => x"a0",
          1652 => x"2a",
          1653 => x"54",
          1654 => x"38",
          1655 => x"76",
          1656 => x"38",
          1657 => x"fd",
          1658 => x"06",
          1659 => x"38",
          1660 => x"56",
          1661 => x"26",
          1662 => x"3d",
          1663 => x"05",
          1664 => x"ff",
          1665 => x"53",
          1666 => x"d9",
          1667 => x"38",
          1668 => x"56",
          1669 => x"27",
          1670 => x"a0",
          1671 => x"3f",
          1672 => x"3d",
          1673 => x"3d",
          1674 => x"70",
          1675 => x"52",
          1676 => x"73",
          1677 => x"3f",
          1678 => x"04",
          1679 => x"74",
          1680 => x"0c",
          1681 => x"05",
          1682 => x"fa",
          1683 => x"de",
          1684 => x"80",
          1685 => x"0b",
          1686 => x"0c",
          1687 => x"04",
          1688 => x"81",
          1689 => x"76",
          1690 => x"0c",
          1691 => x"05",
          1692 => x"53",
          1693 => x"72",
          1694 => x"0c",
          1695 => x"04",
          1696 => x"77",
          1697 => x"d4",
          1698 => x"54",
          1699 => x"54",
          1700 => x"80",
          1701 => x"de",
          1702 => x"71",
          1703 => x"c0",
          1704 => x"06",
          1705 => x"2e",
          1706 => x"72",
          1707 => x"38",
          1708 => x"70",
          1709 => x"25",
          1710 => x"73",
          1711 => x"38",
          1712 => x"86",
          1713 => x"54",
          1714 => x"73",
          1715 => x"ff",
          1716 => x"72",
          1717 => x"74",
          1718 => x"72",
          1719 => x"54",
          1720 => x"81",
          1721 => x"39",
          1722 => x"80",
          1723 => x"51",
          1724 => x"81",
          1725 => x"de",
          1726 => x"3d",
          1727 => x"3d",
          1728 => x"d4",
          1729 => x"de",
          1730 => x"53",
          1731 => x"fe",
          1732 => x"81",
          1733 => x"84",
          1734 => x"f8",
          1735 => x"7c",
          1736 => x"70",
          1737 => x"75",
          1738 => x"55",
          1739 => x"2e",
          1740 => x"87",
          1741 => x"76",
          1742 => x"73",
          1743 => x"81",
          1744 => x"81",
          1745 => x"77",
          1746 => x"70",
          1747 => x"58",
          1748 => x"09",
          1749 => x"c2",
          1750 => x"81",
          1751 => x"75",
          1752 => x"55",
          1753 => x"e2",
          1754 => x"90",
          1755 => x"f8",
          1756 => x"8f",
          1757 => x"81",
          1758 => x"75",
          1759 => x"55",
          1760 => x"81",
          1761 => x"27",
          1762 => x"d0",
          1763 => x"55",
          1764 => x"73",
          1765 => x"80",
          1766 => x"14",
          1767 => x"72",
          1768 => x"e0",
          1769 => x"80",
          1770 => x"39",
          1771 => x"55",
          1772 => x"80",
          1773 => x"e0",
          1774 => x"38",
          1775 => x"81",
          1776 => x"53",
          1777 => x"81",
          1778 => x"53",
          1779 => x"8e",
          1780 => x"70",
          1781 => x"55",
          1782 => x"27",
          1783 => x"77",
          1784 => x"74",
          1785 => x"76",
          1786 => x"77",
          1787 => x"70",
          1788 => x"55",
          1789 => x"77",
          1790 => x"38",
          1791 => x"74",
          1792 => x"55",
          1793 => x"c0",
          1794 => x"0d",
          1795 => x"0d",
          1796 => x"56",
          1797 => x"0c",
          1798 => x"70",
          1799 => x"73",
          1800 => x"81",
          1801 => x"81",
          1802 => x"ed",
          1803 => x"2e",
          1804 => x"8e",
          1805 => x"08",
          1806 => x"76",
          1807 => x"56",
          1808 => x"b0",
          1809 => x"06",
          1810 => x"75",
          1811 => x"76",
          1812 => x"70",
          1813 => x"73",
          1814 => x"8b",
          1815 => x"73",
          1816 => x"85",
          1817 => x"82",
          1818 => x"76",
          1819 => x"70",
          1820 => x"ac",
          1821 => x"a0",
          1822 => x"fa",
          1823 => x"53",
          1824 => x"57",
          1825 => x"98",
          1826 => x"39",
          1827 => x"80",
          1828 => x"26",
          1829 => x"86",
          1830 => x"80",
          1831 => x"57",
          1832 => x"74",
          1833 => x"38",
          1834 => x"27",
          1835 => x"14",
          1836 => x"06",
          1837 => x"14",
          1838 => x"06",
          1839 => x"74",
          1840 => x"f9",
          1841 => x"ff",
          1842 => x"89",
          1843 => x"38",
          1844 => x"c5",
          1845 => x"29",
          1846 => x"81",
          1847 => x"76",
          1848 => x"56",
          1849 => x"ba",
          1850 => x"2e",
          1851 => x"30",
          1852 => x"0c",
          1853 => x"81",
          1854 => x"8a",
          1855 => x"ff",
          1856 => x"8f",
          1857 => x"81",
          1858 => x"26",
          1859 => x"db",
          1860 => x"52",
          1861 => x"c0",
          1862 => x"0d",
          1863 => x"0d",
          1864 => x"33",
          1865 => x"9f",
          1866 => x"53",
          1867 => x"81",
          1868 => x"38",
          1869 => x"87",
          1870 => x"11",
          1871 => x"54",
          1872 => x"84",
          1873 => x"54",
          1874 => x"87",
          1875 => x"11",
          1876 => x"0c",
          1877 => x"c0",
          1878 => x"70",
          1879 => x"70",
          1880 => x"51",
          1881 => x"8a",
          1882 => x"98",
          1883 => x"70",
          1884 => x"08",
          1885 => x"06",
          1886 => x"38",
          1887 => x"8c",
          1888 => x"80",
          1889 => x"71",
          1890 => x"14",
          1891 => x"e8",
          1892 => x"70",
          1893 => x"0c",
          1894 => x"04",
          1895 => x"60",
          1896 => x"8c",
          1897 => x"33",
          1898 => x"5b",
          1899 => x"5a",
          1900 => x"81",
          1901 => x"81",
          1902 => x"52",
          1903 => x"38",
          1904 => x"84",
          1905 => x"92",
          1906 => x"c0",
          1907 => x"87",
          1908 => x"13",
          1909 => x"57",
          1910 => x"0b",
          1911 => x"8c",
          1912 => x"0c",
          1913 => x"75",
          1914 => x"2a",
          1915 => x"51",
          1916 => x"80",
          1917 => x"7b",
          1918 => x"7b",
          1919 => x"5d",
          1920 => x"59",
          1921 => x"06",
          1922 => x"73",
          1923 => x"81",
          1924 => x"ff",
          1925 => x"72",
          1926 => x"38",
          1927 => x"8c",
          1928 => x"c3",
          1929 => x"98",
          1930 => x"71",
          1931 => x"38",
          1932 => x"2e",
          1933 => x"76",
          1934 => x"92",
          1935 => x"72",
          1936 => x"06",
          1937 => x"f7",
          1938 => x"5a",
          1939 => x"80",
          1940 => x"70",
          1941 => x"5a",
          1942 => x"80",
          1943 => x"73",
          1944 => x"06",
          1945 => x"38",
          1946 => x"fe",
          1947 => x"fc",
          1948 => x"52",
          1949 => x"83",
          1950 => x"71",
          1951 => x"de",
          1952 => x"3d",
          1953 => x"3d",
          1954 => x"64",
          1955 => x"bf",
          1956 => x"40",
          1957 => x"59",
          1958 => x"58",
          1959 => x"81",
          1960 => x"81",
          1961 => x"52",
          1962 => x"09",
          1963 => x"b1",
          1964 => x"84",
          1965 => x"92",
          1966 => x"c0",
          1967 => x"87",
          1968 => x"13",
          1969 => x"56",
          1970 => x"87",
          1971 => x"0c",
          1972 => x"82",
          1973 => x"58",
          1974 => x"84",
          1975 => x"06",
          1976 => x"71",
          1977 => x"38",
          1978 => x"05",
          1979 => x"0c",
          1980 => x"73",
          1981 => x"81",
          1982 => x"71",
          1983 => x"38",
          1984 => x"8c",
          1985 => x"d0",
          1986 => x"98",
          1987 => x"71",
          1988 => x"38",
          1989 => x"2e",
          1990 => x"76",
          1991 => x"92",
          1992 => x"72",
          1993 => x"06",
          1994 => x"f7",
          1995 => x"59",
          1996 => x"1a",
          1997 => x"06",
          1998 => x"59",
          1999 => x"80",
          2000 => x"73",
          2001 => x"06",
          2002 => x"38",
          2003 => x"fe",
          2004 => x"fc",
          2005 => x"52",
          2006 => x"83",
          2007 => x"71",
          2008 => x"de",
          2009 => x"3d",
          2010 => x"3d",
          2011 => x"84",
          2012 => x"33",
          2013 => x"b7",
          2014 => x"54",
          2015 => x"fa",
          2016 => x"de",
          2017 => x"06",
          2018 => x"72",
          2019 => x"85",
          2020 => x"98",
          2021 => x"56",
          2022 => x"80",
          2023 => x"76",
          2024 => x"74",
          2025 => x"c0",
          2026 => x"54",
          2027 => x"2e",
          2028 => x"d4",
          2029 => x"2e",
          2030 => x"80",
          2031 => x"08",
          2032 => x"70",
          2033 => x"51",
          2034 => x"2e",
          2035 => x"c0",
          2036 => x"52",
          2037 => x"87",
          2038 => x"08",
          2039 => x"38",
          2040 => x"87",
          2041 => x"14",
          2042 => x"70",
          2043 => x"52",
          2044 => x"96",
          2045 => x"92",
          2046 => x"0a",
          2047 => x"39",
          2048 => x"0c",
          2049 => x"39",
          2050 => x"54",
          2051 => x"c0",
          2052 => x"0d",
          2053 => x"0d",
          2054 => x"33",
          2055 => x"88",
          2056 => x"de",
          2057 => x"51",
          2058 => x"04",
          2059 => x"75",
          2060 => x"82",
          2061 => x"90",
          2062 => x"2b",
          2063 => x"33",
          2064 => x"88",
          2065 => x"71",
          2066 => x"c0",
          2067 => x"54",
          2068 => x"85",
          2069 => x"ff",
          2070 => x"02",
          2071 => x"05",
          2072 => x"70",
          2073 => x"05",
          2074 => x"88",
          2075 => x"72",
          2076 => x"0d",
          2077 => x"0d",
          2078 => x"52",
          2079 => x"81",
          2080 => x"70",
          2081 => x"70",
          2082 => x"05",
          2083 => x"88",
          2084 => x"72",
          2085 => x"54",
          2086 => x"2a",
          2087 => x"34",
          2088 => x"04",
          2089 => x"76",
          2090 => x"54",
          2091 => x"2e",
          2092 => x"70",
          2093 => x"33",
          2094 => x"05",
          2095 => x"11",
          2096 => x"84",
          2097 => x"fe",
          2098 => x"77",
          2099 => x"53",
          2100 => x"81",
          2101 => x"ff",
          2102 => x"f4",
          2103 => x"0d",
          2104 => x"0d",
          2105 => x"56",
          2106 => x"70",
          2107 => x"33",
          2108 => x"05",
          2109 => x"71",
          2110 => x"56",
          2111 => x"72",
          2112 => x"38",
          2113 => x"e2",
          2114 => x"de",
          2115 => x"3d",
          2116 => x"3d",
          2117 => x"54",
          2118 => x"71",
          2119 => x"38",
          2120 => x"70",
          2121 => x"f3",
          2122 => x"81",
          2123 => x"84",
          2124 => x"80",
          2125 => x"c0",
          2126 => x"0b",
          2127 => x"0c",
          2128 => x"0d",
          2129 => x"0b",
          2130 => x"56",
          2131 => x"2e",
          2132 => x"81",
          2133 => x"08",
          2134 => x"70",
          2135 => x"33",
          2136 => x"a2",
          2137 => x"c0",
          2138 => x"09",
          2139 => x"38",
          2140 => x"08",
          2141 => x"b0",
          2142 => x"a4",
          2143 => x"9c",
          2144 => x"56",
          2145 => x"27",
          2146 => x"16",
          2147 => x"82",
          2148 => x"06",
          2149 => x"54",
          2150 => x"78",
          2151 => x"33",
          2152 => x"3f",
          2153 => x"5a",
          2154 => x"c0",
          2155 => x"0d",
          2156 => x"0d",
          2157 => x"56",
          2158 => x"b0",
          2159 => x"af",
          2160 => x"fe",
          2161 => x"de",
          2162 => x"81",
          2163 => x"9f",
          2164 => x"74",
          2165 => x"52",
          2166 => x"51",
          2167 => x"81",
          2168 => x"80",
          2169 => x"ff",
          2170 => x"74",
          2171 => x"76",
          2172 => x"0c",
          2173 => x"04",
          2174 => x"7a",
          2175 => x"fe",
          2176 => x"de",
          2177 => x"81",
          2178 => x"81",
          2179 => x"33",
          2180 => x"2e",
          2181 => x"80",
          2182 => x"17",
          2183 => x"81",
          2184 => x"06",
          2185 => x"84",
          2186 => x"de",
          2187 => x"b4",
          2188 => x"56",
          2189 => x"82",
          2190 => x"84",
          2191 => x"fc",
          2192 => x"8b",
          2193 => x"52",
          2194 => x"a9",
          2195 => x"85",
          2196 => x"84",
          2197 => x"fc",
          2198 => x"17",
          2199 => x"9c",
          2200 => x"91",
          2201 => x"08",
          2202 => x"17",
          2203 => x"3f",
          2204 => x"81",
          2205 => x"19",
          2206 => x"53",
          2207 => x"17",
          2208 => x"82",
          2209 => x"18",
          2210 => x"80",
          2211 => x"33",
          2212 => x"3f",
          2213 => x"08",
          2214 => x"38",
          2215 => x"81",
          2216 => x"8a",
          2217 => x"fb",
          2218 => x"fe",
          2219 => x"08",
          2220 => x"56",
          2221 => x"74",
          2222 => x"38",
          2223 => x"75",
          2224 => x"16",
          2225 => x"53",
          2226 => x"c0",
          2227 => x"0d",
          2228 => x"0d",
          2229 => x"08",
          2230 => x"81",
          2231 => x"df",
          2232 => x"15",
          2233 => x"d7",
          2234 => x"33",
          2235 => x"82",
          2236 => x"38",
          2237 => x"89",
          2238 => x"2e",
          2239 => x"bf",
          2240 => x"2e",
          2241 => x"81",
          2242 => x"81",
          2243 => x"89",
          2244 => x"08",
          2245 => x"52",
          2246 => x"3f",
          2247 => x"08",
          2248 => x"74",
          2249 => x"14",
          2250 => x"81",
          2251 => x"2a",
          2252 => x"05",
          2253 => x"57",
          2254 => x"f5",
          2255 => x"c0",
          2256 => x"38",
          2257 => x"06",
          2258 => x"33",
          2259 => x"78",
          2260 => x"06",
          2261 => x"5c",
          2262 => x"53",
          2263 => x"38",
          2264 => x"06",
          2265 => x"39",
          2266 => x"a4",
          2267 => x"52",
          2268 => x"bd",
          2269 => x"c0",
          2270 => x"38",
          2271 => x"fe",
          2272 => x"b4",
          2273 => x"8d",
          2274 => x"c0",
          2275 => x"ff",
          2276 => x"39",
          2277 => x"a4",
          2278 => x"52",
          2279 => x"91",
          2280 => x"c0",
          2281 => x"76",
          2282 => x"fc",
          2283 => x"b4",
          2284 => x"f8",
          2285 => x"c0",
          2286 => x"06",
          2287 => x"81",
          2288 => x"de",
          2289 => x"3d",
          2290 => x"3d",
          2291 => x"7e",
          2292 => x"82",
          2293 => x"27",
          2294 => x"76",
          2295 => x"27",
          2296 => x"75",
          2297 => x"79",
          2298 => x"38",
          2299 => x"89",
          2300 => x"2e",
          2301 => x"80",
          2302 => x"2e",
          2303 => x"81",
          2304 => x"81",
          2305 => x"89",
          2306 => x"08",
          2307 => x"52",
          2308 => x"3f",
          2309 => x"08",
          2310 => x"c0",
          2311 => x"38",
          2312 => x"06",
          2313 => x"81",
          2314 => x"06",
          2315 => x"77",
          2316 => x"2e",
          2317 => x"84",
          2318 => x"06",
          2319 => x"06",
          2320 => x"53",
          2321 => x"81",
          2322 => x"34",
          2323 => x"a4",
          2324 => x"52",
          2325 => x"d9",
          2326 => x"c0",
          2327 => x"de",
          2328 => x"94",
          2329 => x"ff",
          2330 => x"05",
          2331 => x"54",
          2332 => x"38",
          2333 => x"74",
          2334 => x"06",
          2335 => x"07",
          2336 => x"74",
          2337 => x"39",
          2338 => x"a4",
          2339 => x"52",
          2340 => x"9d",
          2341 => x"c0",
          2342 => x"de",
          2343 => x"d8",
          2344 => x"ff",
          2345 => x"76",
          2346 => x"06",
          2347 => x"05",
          2348 => x"3f",
          2349 => x"87",
          2350 => x"08",
          2351 => x"51",
          2352 => x"81",
          2353 => x"59",
          2354 => x"08",
          2355 => x"f0",
          2356 => x"82",
          2357 => x"06",
          2358 => x"05",
          2359 => x"54",
          2360 => x"3f",
          2361 => x"08",
          2362 => x"74",
          2363 => x"51",
          2364 => x"81",
          2365 => x"34",
          2366 => x"c0",
          2367 => x"0d",
          2368 => x"0d",
          2369 => x"72",
          2370 => x"56",
          2371 => x"27",
          2372 => x"98",
          2373 => x"9d",
          2374 => x"2e",
          2375 => x"53",
          2376 => x"51",
          2377 => x"81",
          2378 => x"54",
          2379 => x"08",
          2380 => x"93",
          2381 => x"80",
          2382 => x"54",
          2383 => x"81",
          2384 => x"54",
          2385 => x"74",
          2386 => x"fb",
          2387 => x"de",
          2388 => x"81",
          2389 => x"80",
          2390 => x"38",
          2391 => x"08",
          2392 => x"38",
          2393 => x"08",
          2394 => x"38",
          2395 => x"52",
          2396 => x"d6",
          2397 => x"c0",
          2398 => x"98",
          2399 => x"11",
          2400 => x"57",
          2401 => x"74",
          2402 => x"81",
          2403 => x"0c",
          2404 => x"81",
          2405 => x"84",
          2406 => x"55",
          2407 => x"ff",
          2408 => x"54",
          2409 => x"c0",
          2410 => x"0d",
          2411 => x"0d",
          2412 => x"08",
          2413 => x"79",
          2414 => x"17",
          2415 => x"80",
          2416 => x"98",
          2417 => x"26",
          2418 => x"58",
          2419 => x"52",
          2420 => x"fd",
          2421 => x"74",
          2422 => x"08",
          2423 => x"38",
          2424 => x"08",
          2425 => x"c0",
          2426 => x"82",
          2427 => x"17",
          2428 => x"c0",
          2429 => x"c7",
          2430 => x"90",
          2431 => x"56",
          2432 => x"2e",
          2433 => x"77",
          2434 => x"81",
          2435 => x"38",
          2436 => x"98",
          2437 => x"26",
          2438 => x"56",
          2439 => x"51",
          2440 => x"80",
          2441 => x"c0",
          2442 => x"09",
          2443 => x"38",
          2444 => x"08",
          2445 => x"c0",
          2446 => x"30",
          2447 => x"80",
          2448 => x"07",
          2449 => x"08",
          2450 => x"55",
          2451 => x"ef",
          2452 => x"c0",
          2453 => x"95",
          2454 => x"08",
          2455 => x"27",
          2456 => x"98",
          2457 => x"89",
          2458 => x"85",
          2459 => x"db",
          2460 => x"81",
          2461 => x"17",
          2462 => x"89",
          2463 => x"75",
          2464 => x"ac",
          2465 => x"7a",
          2466 => x"3f",
          2467 => x"08",
          2468 => x"38",
          2469 => x"de",
          2470 => x"2e",
          2471 => x"86",
          2472 => x"c0",
          2473 => x"de",
          2474 => x"70",
          2475 => x"07",
          2476 => x"7c",
          2477 => x"55",
          2478 => x"f8",
          2479 => x"2e",
          2480 => x"ff",
          2481 => x"55",
          2482 => x"ff",
          2483 => x"76",
          2484 => x"3f",
          2485 => x"08",
          2486 => x"08",
          2487 => x"de",
          2488 => x"80",
          2489 => x"55",
          2490 => x"94",
          2491 => x"2e",
          2492 => x"53",
          2493 => x"51",
          2494 => x"81",
          2495 => x"55",
          2496 => x"75",
          2497 => x"98",
          2498 => x"05",
          2499 => x"56",
          2500 => x"26",
          2501 => x"15",
          2502 => x"84",
          2503 => x"07",
          2504 => x"18",
          2505 => x"ff",
          2506 => x"2e",
          2507 => x"39",
          2508 => x"39",
          2509 => x"08",
          2510 => x"81",
          2511 => x"74",
          2512 => x"0c",
          2513 => x"04",
          2514 => x"7a",
          2515 => x"f3",
          2516 => x"de",
          2517 => x"81",
          2518 => x"c0",
          2519 => x"38",
          2520 => x"51",
          2521 => x"81",
          2522 => x"81",
          2523 => x"b0",
          2524 => x"84",
          2525 => x"52",
          2526 => x"52",
          2527 => x"3f",
          2528 => x"39",
          2529 => x"8a",
          2530 => x"75",
          2531 => x"38",
          2532 => x"19",
          2533 => x"81",
          2534 => x"ed",
          2535 => x"de",
          2536 => x"2e",
          2537 => x"15",
          2538 => x"70",
          2539 => x"07",
          2540 => x"53",
          2541 => x"75",
          2542 => x"0c",
          2543 => x"04",
          2544 => x"7a",
          2545 => x"58",
          2546 => x"f0",
          2547 => x"80",
          2548 => x"9f",
          2549 => x"80",
          2550 => x"90",
          2551 => x"17",
          2552 => x"aa",
          2553 => x"53",
          2554 => x"88",
          2555 => x"08",
          2556 => x"38",
          2557 => x"53",
          2558 => x"17",
          2559 => x"72",
          2560 => x"fe",
          2561 => x"08",
          2562 => x"80",
          2563 => x"16",
          2564 => x"2b",
          2565 => x"75",
          2566 => x"73",
          2567 => x"f5",
          2568 => x"de",
          2569 => x"81",
          2570 => x"ff",
          2571 => x"81",
          2572 => x"c0",
          2573 => x"38",
          2574 => x"81",
          2575 => x"26",
          2576 => x"58",
          2577 => x"73",
          2578 => x"39",
          2579 => x"51",
          2580 => x"81",
          2581 => x"98",
          2582 => x"94",
          2583 => x"17",
          2584 => x"58",
          2585 => x"9a",
          2586 => x"81",
          2587 => x"74",
          2588 => x"98",
          2589 => x"83",
          2590 => x"b4",
          2591 => x"0c",
          2592 => x"81",
          2593 => x"8a",
          2594 => x"f8",
          2595 => x"70",
          2596 => x"08",
          2597 => x"57",
          2598 => x"0a",
          2599 => x"38",
          2600 => x"15",
          2601 => x"08",
          2602 => x"72",
          2603 => x"cb",
          2604 => x"ff",
          2605 => x"81",
          2606 => x"13",
          2607 => x"94",
          2608 => x"74",
          2609 => x"85",
          2610 => x"22",
          2611 => x"73",
          2612 => x"38",
          2613 => x"8a",
          2614 => x"05",
          2615 => x"06",
          2616 => x"8a",
          2617 => x"73",
          2618 => x"3f",
          2619 => x"08",
          2620 => x"81",
          2621 => x"c0",
          2622 => x"ff",
          2623 => x"81",
          2624 => x"ff",
          2625 => x"38",
          2626 => x"81",
          2627 => x"26",
          2628 => x"7b",
          2629 => x"98",
          2630 => x"55",
          2631 => x"94",
          2632 => x"73",
          2633 => x"3f",
          2634 => x"08",
          2635 => x"81",
          2636 => x"80",
          2637 => x"38",
          2638 => x"de",
          2639 => x"2e",
          2640 => x"55",
          2641 => x"08",
          2642 => x"38",
          2643 => x"08",
          2644 => x"fb",
          2645 => x"de",
          2646 => x"38",
          2647 => x"0c",
          2648 => x"51",
          2649 => x"81",
          2650 => x"98",
          2651 => x"90",
          2652 => x"16",
          2653 => x"15",
          2654 => x"74",
          2655 => x"0c",
          2656 => x"04",
          2657 => x"7b",
          2658 => x"5b",
          2659 => x"52",
          2660 => x"ac",
          2661 => x"c0",
          2662 => x"de",
          2663 => x"ec",
          2664 => x"c0",
          2665 => x"17",
          2666 => x"51",
          2667 => x"81",
          2668 => x"54",
          2669 => x"08",
          2670 => x"81",
          2671 => x"9c",
          2672 => x"33",
          2673 => x"72",
          2674 => x"09",
          2675 => x"38",
          2676 => x"de",
          2677 => x"72",
          2678 => x"55",
          2679 => x"53",
          2680 => x"8e",
          2681 => x"56",
          2682 => x"09",
          2683 => x"38",
          2684 => x"de",
          2685 => x"81",
          2686 => x"fd",
          2687 => x"de",
          2688 => x"81",
          2689 => x"80",
          2690 => x"38",
          2691 => x"09",
          2692 => x"38",
          2693 => x"81",
          2694 => x"8b",
          2695 => x"fd",
          2696 => x"9a",
          2697 => x"eb",
          2698 => x"de",
          2699 => x"ff",
          2700 => x"70",
          2701 => x"53",
          2702 => x"09",
          2703 => x"38",
          2704 => x"eb",
          2705 => x"de",
          2706 => x"2b",
          2707 => x"72",
          2708 => x"0c",
          2709 => x"04",
          2710 => x"77",
          2711 => x"ff",
          2712 => x"9a",
          2713 => x"55",
          2714 => x"76",
          2715 => x"53",
          2716 => x"09",
          2717 => x"38",
          2718 => x"52",
          2719 => x"eb",
          2720 => x"3d",
          2721 => x"3d",
          2722 => x"5b",
          2723 => x"08",
          2724 => x"15",
          2725 => x"81",
          2726 => x"15",
          2727 => x"51",
          2728 => x"81",
          2729 => x"58",
          2730 => x"08",
          2731 => x"9c",
          2732 => x"33",
          2733 => x"86",
          2734 => x"80",
          2735 => x"13",
          2736 => x"06",
          2737 => x"06",
          2738 => x"72",
          2739 => x"81",
          2740 => x"53",
          2741 => x"2e",
          2742 => x"53",
          2743 => x"a9",
          2744 => x"74",
          2745 => x"72",
          2746 => x"38",
          2747 => x"99",
          2748 => x"c0",
          2749 => x"06",
          2750 => x"88",
          2751 => x"06",
          2752 => x"54",
          2753 => x"a0",
          2754 => x"74",
          2755 => x"3f",
          2756 => x"08",
          2757 => x"c0",
          2758 => x"98",
          2759 => x"fa",
          2760 => x"80",
          2761 => x"0c",
          2762 => x"c0",
          2763 => x"0d",
          2764 => x"0d",
          2765 => x"57",
          2766 => x"73",
          2767 => x"3f",
          2768 => x"08",
          2769 => x"c0",
          2770 => x"98",
          2771 => x"75",
          2772 => x"3f",
          2773 => x"08",
          2774 => x"c0",
          2775 => x"a0",
          2776 => x"c0",
          2777 => x"14",
          2778 => x"db",
          2779 => x"a0",
          2780 => x"14",
          2781 => x"ac",
          2782 => x"83",
          2783 => x"81",
          2784 => x"87",
          2785 => x"fd",
          2786 => x"70",
          2787 => x"08",
          2788 => x"55",
          2789 => x"3f",
          2790 => x"08",
          2791 => x"13",
          2792 => x"73",
          2793 => x"83",
          2794 => x"3d",
          2795 => x"3d",
          2796 => x"57",
          2797 => x"89",
          2798 => x"17",
          2799 => x"81",
          2800 => x"70",
          2801 => x"55",
          2802 => x"08",
          2803 => x"81",
          2804 => x"52",
          2805 => x"a8",
          2806 => x"2e",
          2807 => x"84",
          2808 => x"52",
          2809 => x"09",
          2810 => x"38",
          2811 => x"81",
          2812 => x"81",
          2813 => x"73",
          2814 => x"55",
          2815 => x"55",
          2816 => x"c5",
          2817 => x"88",
          2818 => x"0b",
          2819 => x"9c",
          2820 => x"8b",
          2821 => x"17",
          2822 => x"08",
          2823 => x"52",
          2824 => x"81",
          2825 => x"76",
          2826 => x"51",
          2827 => x"81",
          2828 => x"86",
          2829 => x"12",
          2830 => x"3f",
          2831 => x"08",
          2832 => x"88",
          2833 => x"f3",
          2834 => x"70",
          2835 => x"80",
          2836 => x"51",
          2837 => x"af",
          2838 => x"81",
          2839 => x"dc",
          2840 => x"74",
          2841 => x"38",
          2842 => x"88",
          2843 => x"39",
          2844 => x"80",
          2845 => x"56",
          2846 => x"af",
          2847 => x"06",
          2848 => x"56",
          2849 => x"32",
          2850 => x"80",
          2851 => x"51",
          2852 => x"dc",
          2853 => x"1c",
          2854 => x"33",
          2855 => x"9f",
          2856 => x"ff",
          2857 => x"1c",
          2858 => x"7a",
          2859 => x"3f",
          2860 => x"08",
          2861 => x"39",
          2862 => x"a0",
          2863 => x"5e",
          2864 => x"52",
          2865 => x"ff",
          2866 => x"59",
          2867 => x"33",
          2868 => x"ae",
          2869 => x"06",
          2870 => x"78",
          2871 => x"81",
          2872 => x"32",
          2873 => x"9f",
          2874 => x"26",
          2875 => x"53",
          2876 => x"73",
          2877 => x"17",
          2878 => x"34",
          2879 => x"db",
          2880 => x"32",
          2881 => x"9f",
          2882 => x"54",
          2883 => x"2e",
          2884 => x"80",
          2885 => x"75",
          2886 => x"bd",
          2887 => x"7e",
          2888 => x"a0",
          2889 => x"bd",
          2890 => x"82",
          2891 => x"18",
          2892 => x"1a",
          2893 => x"a0",
          2894 => x"fc",
          2895 => x"32",
          2896 => x"80",
          2897 => x"30",
          2898 => x"71",
          2899 => x"51",
          2900 => x"55",
          2901 => x"ac",
          2902 => x"81",
          2903 => x"78",
          2904 => x"51",
          2905 => x"af",
          2906 => x"06",
          2907 => x"55",
          2908 => x"32",
          2909 => x"80",
          2910 => x"51",
          2911 => x"db",
          2912 => x"39",
          2913 => x"09",
          2914 => x"38",
          2915 => x"7c",
          2916 => x"54",
          2917 => x"a2",
          2918 => x"32",
          2919 => x"ae",
          2920 => x"72",
          2921 => x"9f",
          2922 => x"51",
          2923 => x"74",
          2924 => x"88",
          2925 => x"fe",
          2926 => x"98",
          2927 => x"80",
          2928 => x"75",
          2929 => x"81",
          2930 => x"33",
          2931 => x"51",
          2932 => x"81",
          2933 => x"80",
          2934 => x"78",
          2935 => x"81",
          2936 => x"5a",
          2937 => x"d2",
          2938 => x"c0",
          2939 => x"80",
          2940 => x"1c",
          2941 => x"27",
          2942 => x"79",
          2943 => x"74",
          2944 => x"7a",
          2945 => x"74",
          2946 => x"39",
          2947 => x"cc",
          2948 => x"fe",
          2949 => x"c0",
          2950 => x"ff",
          2951 => x"73",
          2952 => x"38",
          2953 => x"81",
          2954 => x"54",
          2955 => x"75",
          2956 => x"17",
          2957 => x"39",
          2958 => x"0c",
          2959 => x"99",
          2960 => x"54",
          2961 => x"2e",
          2962 => x"84",
          2963 => x"34",
          2964 => x"76",
          2965 => x"8b",
          2966 => x"81",
          2967 => x"56",
          2968 => x"80",
          2969 => x"1b",
          2970 => x"08",
          2971 => x"51",
          2972 => x"81",
          2973 => x"56",
          2974 => x"08",
          2975 => x"98",
          2976 => x"76",
          2977 => x"3f",
          2978 => x"08",
          2979 => x"c0",
          2980 => x"38",
          2981 => x"70",
          2982 => x"73",
          2983 => x"be",
          2984 => x"33",
          2985 => x"73",
          2986 => x"8b",
          2987 => x"83",
          2988 => x"06",
          2989 => x"73",
          2990 => x"53",
          2991 => x"51",
          2992 => x"81",
          2993 => x"80",
          2994 => x"75",
          2995 => x"f3",
          2996 => x"9f",
          2997 => x"1c",
          2998 => x"74",
          2999 => x"38",
          3000 => x"09",
          3001 => x"e7",
          3002 => x"2a",
          3003 => x"77",
          3004 => x"51",
          3005 => x"2e",
          3006 => x"81",
          3007 => x"80",
          3008 => x"38",
          3009 => x"ab",
          3010 => x"55",
          3011 => x"75",
          3012 => x"73",
          3013 => x"55",
          3014 => x"82",
          3015 => x"06",
          3016 => x"ab",
          3017 => x"33",
          3018 => x"70",
          3019 => x"55",
          3020 => x"2e",
          3021 => x"1b",
          3022 => x"06",
          3023 => x"52",
          3024 => x"db",
          3025 => x"c0",
          3026 => x"0c",
          3027 => x"74",
          3028 => x"0c",
          3029 => x"04",
          3030 => x"7c",
          3031 => x"08",
          3032 => x"55",
          3033 => x"59",
          3034 => x"81",
          3035 => x"70",
          3036 => x"33",
          3037 => x"52",
          3038 => x"2e",
          3039 => x"ee",
          3040 => x"2e",
          3041 => x"81",
          3042 => x"33",
          3043 => x"81",
          3044 => x"52",
          3045 => x"26",
          3046 => x"14",
          3047 => x"06",
          3048 => x"52",
          3049 => x"80",
          3050 => x"0b",
          3051 => x"59",
          3052 => x"7a",
          3053 => x"70",
          3054 => x"33",
          3055 => x"05",
          3056 => x"9f",
          3057 => x"53",
          3058 => x"89",
          3059 => x"70",
          3060 => x"54",
          3061 => x"12",
          3062 => x"26",
          3063 => x"12",
          3064 => x"06",
          3065 => x"30",
          3066 => x"51",
          3067 => x"2e",
          3068 => x"85",
          3069 => x"be",
          3070 => x"74",
          3071 => x"30",
          3072 => x"9f",
          3073 => x"2a",
          3074 => x"54",
          3075 => x"2e",
          3076 => x"15",
          3077 => x"55",
          3078 => x"ff",
          3079 => x"39",
          3080 => x"86",
          3081 => x"7c",
          3082 => x"51",
          3083 => x"de",
          3084 => x"70",
          3085 => x"0c",
          3086 => x"04",
          3087 => x"78",
          3088 => x"83",
          3089 => x"0b",
          3090 => x"79",
          3091 => x"e2",
          3092 => x"55",
          3093 => x"08",
          3094 => x"84",
          3095 => x"df",
          3096 => x"de",
          3097 => x"ff",
          3098 => x"83",
          3099 => x"d4",
          3100 => x"81",
          3101 => x"38",
          3102 => x"17",
          3103 => x"74",
          3104 => x"09",
          3105 => x"38",
          3106 => x"81",
          3107 => x"30",
          3108 => x"79",
          3109 => x"54",
          3110 => x"74",
          3111 => x"09",
          3112 => x"38",
          3113 => x"cc",
          3114 => x"ea",
          3115 => x"b1",
          3116 => x"c0",
          3117 => x"de",
          3118 => x"2e",
          3119 => x"53",
          3120 => x"52",
          3121 => x"51",
          3122 => x"81",
          3123 => x"55",
          3124 => x"08",
          3125 => x"38",
          3126 => x"81",
          3127 => x"88",
          3128 => x"f2",
          3129 => x"02",
          3130 => x"cb",
          3131 => x"55",
          3132 => x"60",
          3133 => x"3f",
          3134 => x"08",
          3135 => x"80",
          3136 => x"c0",
          3137 => x"fc",
          3138 => x"c0",
          3139 => x"81",
          3140 => x"70",
          3141 => x"8c",
          3142 => x"2e",
          3143 => x"73",
          3144 => x"81",
          3145 => x"33",
          3146 => x"80",
          3147 => x"81",
          3148 => x"d7",
          3149 => x"de",
          3150 => x"ff",
          3151 => x"06",
          3152 => x"98",
          3153 => x"2e",
          3154 => x"74",
          3155 => x"81",
          3156 => x"8a",
          3157 => x"ac",
          3158 => x"39",
          3159 => x"77",
          3160 => x"81",
          3161 => x"33",
          3162 => x"3f",
          3163 => x"08",
          3164 => x"70",
          3165 => x"55",
          3166 => x"86",
          3167 => x"80",
          3168 => x"74",
          3169 => x"81",
          3170 => x"8a",
          3171 => x"f4",
          3172 => x"53",
          3173 => x"fd",
          3174 => x"de",
          3175 => x"ff",
          3176 => x"82",
          3177 => x"06",
          3178 => x"8c",
          3179 => x"58",
          3180 => x"f6",
          3181 => x"58",
          3182 => x"2e",
          3183 => x"fa",
          3184 => x"e8",
          3185 => x"c0",
          3186 => x"78",
          3187 => x"5a",
          3188 => x"90",
          3189 => x"75",
          3190 => x"38",
          3191 => x"3d",
          3192 => x"70",
          3193 => x"08",
          3194 => x"7a",
          3195 => x"38",
          3196 => x"51",
          3197 => x"81",
          3198 => x"81",
          3199 => x"81",
          3200 => x"38",
          3201 => x"83",
          3202 => x"38",
          3203 => x"84",
          3204 => x"38",
          3205 => x"81",
          3206 => x"38",
          3207 => x"db",
          3208 => x"de",
          3209 => x"ff",
          3210 => x"72",
          3211 => x"09",
          3212 => x"d0",
          3213 => x"14",
          3214 => x"3f",
          3215 => x"08",
          3216 => x"06",
          3217 => x"38",
          3218 => x"51",
          3219 => x"81",
          3220 => x"58",
          3221 => x"0c",
          3222 => x"33",
          3223 => x"80",
          3224 => x"ff",
          3225 => x"ff",
          3226 => x"55",
          3227 => x"81",
          3228 => x"38",
          3229 => x"06",
          3230 => x"80",
          3231 => x"52",
          3232 => x"8a",
          3233 => x"80",
          3234 => x"ff",
          3235 => x"53",
          3236 => x"86",
          3237 => x"83",
          3238 => x"c5",
          3239 => x"f5",
          3240 => x"c0",
          3241 => x"de",
          3242 => x"15",
          3243 => x"06",
          3244 => x"76",
          3245 => x"80",
          3246 => x"da",
          3247 => x"de",
          3248 => x"ff",
          3249 => x"74",
          3250 => x"d4",
          3251 => x"dc",
          3252 => x"c0",
          3253 => x"c2",
          3254 => x"b9",
          3255 => x"c0",
          3256 => x"ff",
          3257 => x"56",
          3258 => x"83",
          3259 => x"14",
          3260 => x"71",
          3261 => x"5a",
          3262 => x"26",
          3263 => x"8a",
          3264 => x"74",
          3265 => x"ff",
          3266 => x"81",
          3267 => x"55",
          3268 => x"08",
          3269 => x"ec",
          3270 => x"c0",
          3271 => x"ff",
          3272 => x"83",
          3273 => x"74",
          3274 => x"26",
          3275 => x"57",
          3276 => x"26",
          3277 => x"57",
          3278 => x"56",
          3279 => x"82",
          3280 => x"15",
          3281 => x"0c",
          3282 => x"0c",
          3283 => x"a4",
          3284 => x"1d",
          3285 => x"54",
          3286 => x"2e",
          3287 => x"af",
          3288 => x"14",
          3289 => x"3f",
          3290 => x"08",
          3291 => x"06",
          3292 => x"72",
          3293 => x"79",
          3294 => x"80",
          3295 => x"d9",
          3296 => x"de",
          3297 => x"15",
          3298 => x"2b",
          3299 => x"8d",
          3300 => x"2e",
          3301 => x"77",
          3302 => x"0c",
          3303 => x"76",
          3304 => x"38",
          3305 => x"70",
          3306 => x"81",
          3307 => x"53",
          3308 => x"89",
          3309 => x"56",
          3310 => x"08",
          3311 => x"38",
          3312 => x"15",
          3313 => x"8c",
          3314 => x"80",
          3315 => x"34",
          3316 => x"09",
          3317 => x"92",
          3318 => x"14",
          3319 => x"3f",
          3320 => x"08",
          3321 => x"06",
          3322 => x"2e",
          3323 => x"80",
          3324 => x"1b",
          3325 => x"db",
          3326 => x"de",
          3327 => x"ea",
          3328 => x"c0",
          3329 => x"34",
          3330 => x"51",
          3331 => x"81",
          3332 => x"83",
          3333 => x"53",
          3334 => x"d5",
          3335 => x"06",
          3336 => x"b4",
          3337 => x"84",
          3338 => x"c0",
          3339 => x"85",
          3340 => x"09",
          3341 => x"38",
          3342 => x"51",
          3343 => x"81",
          3344 => x"86",
          3345 => x"f2",
          3346 => x"06",
          3347 => x"9c",
          3348 => x"d8",
          3349 => x"c0",
          3350 => x"0c",
          3351 => x"51",
          3352 => x"81",
          3353 => x"8c",
          3354 => x"74",
          3355 => x"ec",
          3356 => x"53",
          3357 => x"ec",
          3358 => x"15",
          3359 => x"94",
          3360 => x"56",
          3361 => x"c0",
          3362 => x"0d",
          3363 => x"0d",
          3364 => x"55",
          3365 => x"b9",
          3366 => x"53",
          3367 => x"b1",
          3368 => x"52",
          3369 => x"a9",
          3370 => x"22",
          3371 => x"57",
          3372 => x"2e",
          3373 => x"99",
          3374 => x"33",
          3375 => x"3f",
          3376 => x"08",
          3377 => x"71",
          3378 => x"74",
          3379 => x"83",
          3380 => x"78",
          3381 => x"52",
          3382 => x"c0",
          3383 => x"0d",
          3384 => x"0d",
          3385 => x"33",
          3386 => x"3d",
          3387 => x"56",
          3388 => x"8b",
          3389 => x"81",
          3390 => x"24",
          3391 => x"de",
          3392 => x"29",
          3393 => x"05",
          3394 => x"55",
          3395 => x"84",
          3396 => x"34",
          3397 => x"80",
          3398 => x"80",
          3399 => x"75",
          3400 => x"75",
          3401 => x"38",
          3402 => x"3d",
          3403 => x"05",
          3404 => x"3f",
          3405 => x"08",
          3406 => x"de",
          3407 => x"3d",
          3408 => x"3d",
          3409 => x"84",
          3410 => x"05",
          3411 => x"89",
          3412 => x"2e",
          3413 => x"77",
          3414 => x"54",
          3415 => x"05",
          3416 => x"84",
          3417 => x"f6",
          3418 => x"de",
          3419 => x"81",
          3420 => x"84",
          3421 => x"5c",
          3422 => x"3d",
          3423 => x"ed",
          3424 => x"de",
          3425 => x"81",
          3426 => x"92",
          3427 => x"d7",
          3428 => x"98",
          3429 => x"73",
          3430 => x"38",
          3431 => x"9c",
          3432 => x"80",
          3433 => x"38",
          3434 => x"95",
          3435 => x"2e",
          3436 => x"aa",
          3437 => x"ea",
          3438 => x"de",
          3439 => x"9e",
          3440 => x"05",
          3441 => x"54",
          3442 => x"38",
          3443 => x"70",
          3444 => x"54",
          3445 => x"8e",
          3446 => x"83",
          3447 => x"88",
          3448 => x"83",
          3449 => x"83",
          3450 => x"06",
          3451 => x"80",
          3452 => x"38",
          3453 => x"51",
          3454 => x"81",
          3455 => x"56",
          3456 => x"0a",
          3457 => x"05",
          3458 => x"3f",
          3459 => x"0b",
          3460 => x"80",
          3461 => x"7a",
          3462 => x"3f",
          3463 => x"9c",
          3464 => x"d1",
          3465 => x"81",
          3466 => x"34",
          3467 => x"80",
          3468 => x"b0",
          3469 => x"54",
          3470 => x"52",
          3471 => x"05",
          3472 => x"3f",
          3473 => x"08",
          3474 => x"c0",
          3475 => x"38",
          3476 => x"82",
          3477 => x"b2",
          3478 => x"84",
          3479 => x"06",
          3480 => x"73",
          3481 => x"38",
          3482 => x"ad",
          3483 => x"2a",
          3484 => x"51",
          3485 => x"2e",
          3486 => x"81",
          3487 => x"80",
          3488 => x"87",
          3489 => x"39",
          3490 => x"51",
          3491 => x"81",
          3492 => x"7b",
          3493 => x"12",
          3494 => x"81",
          3495 => x"81",
          3496 => x"83",
          3497 => x"06",
          3498 => x"80",
          3499 => x"77",
          3500 => x"58",
          3501 => x"08",
          3502 => x"63",
          3503 => x"63",
          3504 => x"57",
          3505 => x"81",
          3506 => x"81",
          3507 => x"88",
          3508 => x"9c",
          3509 => x"d2",
          3510 => x"de",
          3511 => x"de",
          3512 => x"1b",
          3513 => x"0c",
          3514 => x"22",
          3515 => x"77",
          3516 => x"80",
          3517 => x"34",
          3518 => x"1a",
          3519 => x"94",
          3520 => x"85",
          3521 => x"06",
          3522 => x"80",
          3523 => x"38",
          3524 => x"08",
          3525 => x"84",
          3526 => x"c0",
          3527 => x"0c",
          3528 => x"70",
          3529 => x"52",
          3530 => x"39",
          3531 => x"51",
          3532 => x"81",
          3533 => x"57",
          3534 => x"08",
          3535 => x"38",
          3536 => x"de",
          3537 => x"2e",
          3538 => x"83",
          3539 => x"75",
          3540 => x"74",
          3541 => x"07",
          3542 => x"54",
          3543 => x"8a",
          3544 => x"75",
          3545 => x"73",
          3546 => x"98",
          3547 => x"a9",
          3548 => x"ff",
          3549 => x"80",
          3550 => x"76",
          3551 => x"d6",
          3552 => x"de",
          3553 => x"38",
          3554 => x"39",
          3555 => x"81",
          3556 => x"05",
          3557 => x"84",
          3558 => x"0c",
          3559 => x"81",
          3560 => x"97",
          3561 => x"f2",
          3562 => x"63",
          3563 => x"40",
          3564 => x"7e",
          3565 => x"fc",
          3566 => x"51",
          3567 => x"81",
          3568 => x"55",
          3569 => x"08",
          3570 => x"19",
          3571 => x"80",
          3572 => x"74",
          3573 => x"39",
          3574 => x"81",
          3575 => x"56",
          3576 => x"82",
          3577 => x"39",
          3578 => x"1a",
          3579 => x"82",
          3580 => x"0b",
          3581 => x"81",
          3582 => x"39",
          3583 => x"94",
          3584 => x"55",
          3585 => x"83",
          3586 => x"7b",
          3587 => x"89",
          3588 => x"08",
          3589 => x"06",
          3590 => x"81",
          3591 => x"8a",
          3592 => x"05",
          3593 => x"06",
          3594 => x"a8",
          3595 => x"38",
          3596 => x"55",
          3597 => x"19",
          3598 => x"51",
          3599 => x"81",
          3600 => x"55",
          3601 => x"ff",
          3602 => x"ff",
          3603 => x"38",
          3604 => x"0c",
          3605 => x"52",
          3606 => x"cb",
          3607 => x"c0",
          3608 => x"ff",
          3609 => x"de",
          3610 => x"7c",
          3611 => x"57",
          3612 => x"80",
          3613 => x"1a",
          3614 => x"22",
          3615 => x"75",
          3616 => x"38",
          3617 => x"58",
          3618 => x"53",
          3619 => x"1b",
          3620 => x"88",
          3621 => x"c0",
          3622 => x"38",
          3623 => x"33",
          3624 => x"80",
          3625 => x"b0",
          3626 => x"31",
          3627 => x"27",
          3628 => x"80",
          3629 => x"52",
          3630 => x"77",
          3631 => x"7d",
          3632 => x"e0",
          3633 => x"2b",
          3634 => x"76",
          3635 => x"94",
          3636 => x"ff",
          3637 => x"71",
          3638 => x"7b",
          3639 => x"38",
          3640 => x"19",
          3641 => x"51",
          3642 => x"81",
          3643 => x"fe",
          3644 => x"53",
          3645 => x"83",
          3646 => x"b4",
          3647 => x"51",
          3648 => x"7b",
          3649 => x"08",
          3650 => x"76",
          3651 => x"08",
          3652 => x"0c",
          3653 => x"f3",
          3654 => x"75",
          3655 => x"0c",
          3656 => x"04",
          3657 => x"60",
          3658 => x"40",
          3659 => x"80",
          3660 => x"3d",
          3661 => x"77",
          3662 => x"3f",
          3663 => x"08",
          3664 => x"c0",
          3665 => x"91",
          3666 => x"74",
          3667 => x"38",
          3668 => x"b8",
          3669 => x"33",
          3670 => x"70",
          3671 => x"56",
          3672 => x"74",
          3673 => x"a4",
          3674 => x"82",
          3675 => x"34",
          3676 => x"98",
          3677 => x"91",
          3678 => x"56",
          3679 => x"94",
          3680 => x"11",
          3681 => x"76",
          3682 => x"75",
          3683 => x"80",
          3684 => x"38",
          3685 => x"70",
          3686 => x"56",
          3687 => x"fd",
          3688 => x"11",
          3689 => x"77",
          3690 => x"5c",
          3691 => x"38",
          3692 => x"88",
          3693 => x"74",
          3694 => x"52",
          3695 => x"18",
          3696 => x"51",
          3697 => x"81",
          3698 => x"55",
          3699 => x"08",
          3700 => x"ab",
          3701 => x"2e",
          3702 => x"74",
          3703 => x"95",
          3704 => x"19",
          3705 => x"08",
          3706 => x"88",
          3707 => x"55",
          3708 => x"9c",
          3709 => x"09",
          3710 => x"38",
          3711 => x"c1",
          3712 => x"c0",
          3713 => x"38",
          3714 => x"52",
          3715 => x"97",
          3716 => x"c0",
          3717 => x"fe",
          3718 => x"de",
          3719 => x"7c",
          3720 => x"57",
          3721 => x"80",
          3722 => x"1b",
          3723 => x"22",
          3724 => x"75",
          3725 => x"38",
          3726 => x"59",
          3727 => x"53",
          3728 => x"1a",
          3729 => x"be",
          3730 => x"c0",
          3731 => x"38",
          3732 => x"08",
          3733 => x"56",
          3734 => x"9b",
          3735 => x"53",
          3736 => x"77",
          3737 => x"7d",
          3738 => x"16",
          3739 => x"3f",
          3740 => x"0b",
          3741 => x"78",
          3742 => x"80",
          3743 => x"18",
          3744 => x"08",
          3745 => x"7e",
          3746 => x"3f",
          3747 => x"08",
          3748 => x"7e",
          3749 => x"0c",
          3750 => x"19",
          3751 => x"08",
          3752 => x"84",
          3753 => x"57",
          3754 => x"27",
          3755 => x"56",
          3756 => x"52",
          3757 => x"f9",
          3758 => x"c0",
          3759 => x"38",
          3760 => x"52",
          3761 => x"83",
          3762 => x"b4",
          3763 => x"d4",
          3764 => x"81",
          3765 => x"34",
          3766 => x"7e",
          3767 => x"0c",
          3768 => x"1a",
          3769 => x"94",
          3770 => x"1b",
          3771 => x"5e",
          3772 => x"27",
          3773 => x"55",
          3774 => x"0c",
          3775 => x"90",
          3776 => x"c0",
          3777 => x"90",
          3778 => x"56",
          3779 => x"c0",
          3780 => x"0d",
          3781 => x"0d",
          3782 => x"fc",
          3783 => x"52",
          3784 => x"3f",
          3785 => x"08",
          3786 => x"c0",
          3787 => x"38",
          3788 => x"70",
          3789 => x"81",
          3790 => x"55",
          3791 => x"80",
          3792 => x"16",
          3793 => x"51",
          3794 => x"81",
          3795 => x"57",
          3796 => x"08",
          3797 => x"a4",
          3798 => x"11",
          3799 => x"55",
          3800 => x"16",
          3801 => x"08",
          3802 => x"75",
          3803 => x"e8",
          3804 => x"08",
          3805 => x"51",
          3806 => x"82",
          3807 => x"52",
          3808 => x"c9",
          3809 => x"52",
          3810 => x"c9",
          3811 => x"54",
          3812 => x"15",
          3813 => x"cc",
          3814 => x"de",
          3815 => x"17",
          3816 => x"06",
          3817 => x"90",
          3818 => x"81",
          3819 => x"8a",
          3820 => x"fc",
          3821 => x"70",
          3822 => x"d9",
          3823 => x"c0",
          3824 => x"de",
          3825 => x"38",
          3826 => x"05",
          3827 => x"f1",
          3828 => x"de",
          3829 => x"81",
          3830 => x"87",
          3831 => x"c0",
          3832 => x"72",
          3833 => x"0c",
          3834 => x"04",
          3835 => x"84",
          3836 => x"e4",
          3837 => x"80",
          3838 => x"c0",
          3839 => x"38",
          3840 => x"08",
          3841 => x"34",
          3842 => x"81",
          3843 => x"83",
          3844 => x"ef",
          3845 => x"53",
          3846 => x"05",
          3847 => x"51",
          3848 => x"81",
          3849 => x"55",
          3850 => x"08",
          3851 => x"76",
          3852 => x"93",
          3853 => x"51",
          3854 => x"81",
          3855 => x"55",
          3856 => x"08",
          3857 => x"80",
          3858 => x"70",
          3859 => x"56",
          3860 => x"89",
          3861 => x"94",
          3862 => x"b2",
          3863 => x"05",
          3864 => x"2a",
          3865 => x"51",
          3866 => x"80",
          3867 => x"76",
          3868 => x"52",
          3869 => x"3f",
          3870 => x"08",
          3871 => x"8e",
          3872 => x"c0",
          3873 => x"09",
          3874 => x"38",
          3875 => x"81",
          3876 => x"93",
          3877 => x"e4",
          3878 => x"6f",
          3879 => x"7a",
          3880 => x"9e",
          3881 => x"05",
          3882 => x"51",
          3883 => x"81",
          3884 => x"57",
          3885 => x"08",
          3886 => x"7b",
          3887 => x"94",
          3888 => x"55",
          3889 => x"73",
          3890 => x"ed",
          3891 => x"93",
          3892 => x"55",
          3893 => x"81",
          3894 => x"57",
          3895 => x"08",
          3896 => x"68",
          3897 => x"c9",
          3898 => x"de",
          3899 => x"81",
          3900 => x"82",
          3901 => x"52",
          3902 => x"a3",
          3903 => x"c0",
          3904 => x"52",
          3905 => x"b8",
          3906 => x"c0",
          3907 => x"de",
          3908 => x"a2",
          3909 => x"74",
          3910 => x"3f",
          3911 => x"08",
          3912 => x"c0",
          3913 => x"69",
          3914 => x"d9",
          3915 => x"81",
          3916 => x"2e",
          3917 => x"52",
          3918 => x"cf",
          3919 => x"c0",
          3920 => x"de",
          3921 => x"2e",
          3922 => x"84",
          3923 => x"06",
          3924 => x"57",
          3925 => x"76",
          3926 => x"9e",
          3927 => x"05",
          3928 => x"dc",
          3929 => x"90",
          3930 => x"81",
          3931 => x"56",
          3932 => x"80",
          3933 => x"02",
          3934 => x"81",
          3935 => x"70",
          3936 => x"56",
          3937 => x"81",
          3938 => x"78",
          3939 => x"38",
          3940 => x"99",
          3941 => x"81",
          3942 => x"18",
          3943 => x"18",
          3944 => x"58",
          3945 => x"33",
          3946 => x"ee",
          3947 => x"6f",
          3948 => x"af",
          3949 => x"8d",
          3950 => x"2e",
          3951 => x"8a",
          3952 => x"6f",
          3953 => x"af",
          3954 => x"0b",
          3955 => x"33",
          3956 => x"81",
          3957 => x"70",
          3958 => x"52",
          3959 => x"56",
          3960 => x"8d",
          3961 => x"70",
          3962 => x"51",
          3963 => x"f5",
          3964 => x"54",
          3965 => x"a7",
          3966 => x"74",
          3967 => x"38",
          3968 => x"73",
          3969 => x"81",
          3970 => x"81",
          3971 => x"39",
          3972 => x"81",
          3973 => x"74",
          3974 => x"81",
          3975 => x"91",
          3976 => x"6e",
          3977 => x"59",
          3978 => x"7a",
          3979 => x"5c",
          3980 => x"26",
          3981 => x"7a",
          3982 => x"de",
          3983 => x"3d",
          3984 => x"3d",
          3985 => x"8d",
          3986 => x"54",
          3987 => x"55",
          3988 => x"81",
          3989 => x"53",
          3990 => x"08",
          3991 => x"91",
          3992 => x"72",
          3993 => x"8c",
          3994 => x"73",
          3995 => x"38",
          3996 => x"70",
          3997 => x"81",
          3998 => x"57",
          3999 => x"73",
          4000 => x"08",
          4001 => x"94",
          4002 => x"75",
          4003 => x"97",
          4004 => x"11",
          4005 => x"2b",
          4006 => x"73",
          4007 => x"38",
          4008 => x"16",
          4009 => x"d2",
          4010 => x"c0",
          4011 => x"78",
          4012 => x"55",
          4013 => x"c2",
          4014 => x"c0",
          4015 => x"96",
          4016 => x"70",
          4017 => x"94",
          4018 => x"71",
          4019 => x"08",
          4020 => x"53",
          4021 => x"15",
          4022 => x"a6",
          4023 => x"74",
          4024 => x"3f",
          4025 => x"08",
          4026 => x"c0",
          4027 => x"81",
          4028 => x"de",
          4029 => x"2e",
          4030 => x"81",
          4031 => x"88",
          4032 => x"98",
          4033 => x"80",
          4034 => x"38",
          4035 => x"80",
          4036 => x"77",
          4037 => x"08",
          4038 => x"0c",
          4039 => x"70",
          4040 => x"81",
          4041 => x"5a",
          4042 => x"2e",
          4043 => x"52",
          4044 => x"f9",
          4045 => x"c0",
          4046 => x"de",
          4047 => x"38",
          4048 => x"08",
          4049 => x"73",
          4050 => x"c7",
          4051 => x"de",
          4052 => x"73",
          4053 => x"38",
          4054 => x"af",
          4055 => x"73",
          4056 => x"27",
          4057 => x"98",
          4058 => x"a0",
          4059 => x"08",
          4060 => x"0c",
          4061 => x"06",
          4062 => x"2e",
          4063 => x"52",
          4064 => x"a3",
          4065 => x"c0",
          4066 => x"82",
          4067 => x"34",
          4068 => x"c4",
          4069 => x"91",
          4070 => x"53",
          4071 => x"89",
          4072 => x"c0",
          4073 => x"94",
          4074 => x"8c",
          4075 => x"27",
          4076 => x"8c",
          4077 => x"15",
          4078 => x"07",
          4079 => x"16",
          4080 => x"ff",
          4081 => x"80",
          4082 => x"77",
          4083 => x"2e",
          4084 => x"9c",
          4085 => x"53",
          4086 => x"c0",
          4087 => x"0d",
          4088 => x"0d",
          4089 => x"54",
          4090 => x"81",
          4091 => x"53",
          4092 => x"05",
          4093 => x"84",
          4094 => x"e7",
          4095 => x"c0",
          4096 => x"de",
          4097 => x"ea",
          4098 => x"0c",
          4099 => x"51",
          4100 => x"81",
          4101 => x"55",
          4102 => x"08",
          4103 => x"ab",
          4104 => x"98",
          4105 => x"80",
          4106 => x"38",
          4107 => x"70",
          4108 => x"81",
          4109 => x"57",
          4110 => x"ad",
          4111 => x"08",
          4112 => x"d3",
          4113 => x"de",
          4114 => x"17",
          4115 => x"86",
          4116 => x"17",
          4117 => x"75",
          4118 => x"3f",
          4119 => x"08",
          4120 => x"2e",
          4121 => x"85",
          4122 => x"86",
          4123 => x"2e",
          4124 => x"76",
          4125 => x"73",
          4126 => x"0c",
          4127 => x"04",
          4128 => x"76",
          4129 => x"05",
          4130 => x"53",
          4131 => x"81",
          4132 => x"87",
          4133 => x"c0",
          4134 => x"86",
          4135 => x"fb",
          4136 => x"79",
          4137 => x"05",
          4138 => x"56",
          4139 => x"3f",
          4140 => x"08",
          4141 => x"c0",
          4142 => x"38",
          4143 => x"81",
          4144 => x"52",
          4145 => x"f8",
          4146 => x"c0",
          4147 => x"ca",
          4148 => x"c0",
          4149 => x"51",
          4150 => x"81",
          4151 => x"53",
          4152 => x"08",
          4153 => x"81",
          4154 => x"80",
          4155 => x"81",
          4156 => x"a6",
          4157 => x"73",
          4158 => x"3f",
          4159 => x"51",
          4160 => x"81",
          4161 => x"84",
          4162 => x"70",
          4163 => x"2c",
          4164 => x"c0",
          4165 => x"51",
          4166 => x"81",
          4167 => x"87",
          4168 => x"ee",
          4169 => x"57",
          4170 => x"3d",
          4171 => x"3d",
          4172 => x"af",
          4173 => x"c0",
          4174 => x"de",
          4175 => x"38",
          4176 => x"51",
          4177 => x"81",
          4178 => x"55",
          4179 => x"08",
          4180 => x"80",
          4181 => x"70",
          4182 => x"58",
          4183 => x"85",
          4184 => x"8d",
          4185 => x"2e",
          4186 => x"52",
          4187 => x"be",
          4188 => x"de",
          4189 => x"3d",
          4190 => x"3d",
          4191 => x"55",
          4192 => x"92",
          4193 => x"52",
          4194 => x"de",
          4195 => x"de",
          4196 => x"81",
          4197 => x"82",
          4198 => x"74",
          4199 => x"98",
          4200 => x"11",
          4201 => x"59",
          4202 => x"75",
          4203 => x"38",
          4204 => x"81",
          4205 => x"5b",
          4206 => x"82",
          4207 => x"39",
          4208 => x"08",
          4209 => x"59",
          4210 => x"09",
          4211 => x"38",
          4212 => x"57",
          4213 => x"3d",
          4214 => x"c1",
          4215 => x"de",
          4216 => x"2e",
          4217 => x"de",
          4218 => x"2e",
          4219 => x"de",
          4220 => x"70",
          4221 => x"08",
          4222 => x"7a",
          4223 => x"7f",
          4224 => x"54",
          4225 => x"77",
          4226 => x"80",
          4227 => x"15",
          4228 => x"c0",
          4229 => x"75",
          4230 => x"52",
          4231 => x"52",
          4232 => x"8d",
          4233 => x"c0",
          4234 => x"de",
          4235 => x"d6",
          4236 => x"33",
          4237 => x"1a",
          4238 => x"54",
          4239 => x"09",
          4240 => x"38",
          4241 => x"ff",
          4242 => x"81",
          4243 => x"83",
          4244 => x"70",
          4245 => x"25",
          4246 => x"59",
          4247 => x"9b",
          4248 => x"51",
          4249 => x"3f",
          4250 => x"08",
          4251 => x"70",
          4252 => x"25",
          4253 => x"59",
          4254 => x"75",
          4255 => x"7a",
          4256 => x"ff",
          4257 => x"7c",
          4258 => x"90",
          4259 => x"11",
          4260 => x"56",
          4261 => x"15",
          4262 => x"de",
          4263 => x"3d",
          4264 => x"3d",
          4265 => x"3d",
          4266 => x"70",
          4267 => x"dd",
          4268 => x"c0",
          4269 => x"de",
          4270 => x"a8",
          4271 => x"33",
          4272 => x"a0",
          4273 => x"33",
          4274 => x"70",
          4275 => x"55",
          4276 => x"73",
          4277 => x"8e",
          4278 => x"08",
          4279 => x"18",
          4280 => x"80",
          4281 => x"38",
          4282 => x"08",
          4283 => x"08",
          4284 => x"c4",
          4285 => x"de",
          4286 => x"88",
          4287 => x"80",
          4288 => x"17",
          4289 => x"51",
          4290 => x"3f",
          4291 => x"08",
          4292 => x"81",
          4293 => x"81",
          4294 => x"c0",
          4295 => x"09",
          4296 => x"38",
          4297 => x"39",
          4298 => x"77",
          4299 => x"c0",
          4300 => x"08",
          4301 => x"98",
          4302 => x"81",
          4303 => x"52",
          4304 => x"bd",
          4305 => x"c0",
          4306 => x"17",
          4307 => x"0c",
          4308 => x"80",
          4309 => x"73",
          4310 => x"75",
          4311 => x"38",
          4312 => x"34",
          4313 => x"81",
          4314 => x"89",
          4315 => x"e2",
          4316 => x"53",
          4317 => x"a4",
          4318 => x"3d",
          4319 => x"3f",
          4320 => x"08",
          4321 => x"c0",
          4322 => x"38",
          4323 => x"3d",
          4324 => x"3d",
          4325 => x"d1",
          4326 => x"de",
          4327 => x"81",
          4328 => x"81",
          4329 => x"80",
          4330 => x"70",
          4331 => x"81",
          4332 => x"56",
          4333 => x"81",
          4334 => x"98",
          4335 => x"74",
          4336 => x"38",
          4337 => x"05",
          4338 => x"06",
          4339 => x"55",
          4340 => x"38",
          4341 => x"51",
          4342 => x"81",
          4343 => x"74",
          4344 => x"81",
          4345 => x"56",
          4346 => x"80",
          4347 => x"54",
          4348 => x"08",
          4349 => x"2e",
          4350 => x"73",
          4351 => x"c0",
          4352 => x"52",
          4353 => x"52",
          4354 => x"3f",
          4355 => x"08",
          4356 => x"c0",
          4357 => x"38",
          4358 => x"08",
          4359 => x"cc",
          4360 => x"de",
          4361 => x"81",
          4362 => x"86",
          4363 => x"80",
          4364 => x"de",
          4365 => x"2e",
          4366 => x"de",
          4367 => x"c0",
          4368 => x"ce",
          4369 => x"de",
          4370 => x"de",
          4371 => x"70",
          4372 => x"08",
          4373 => x"51",
          4374 => x"80",
          4375 => x"73",
          4376 => x"38",
          4377 => x"52",
          4378 => x"95",
          4379 => x"c0",
          4380 => x"8c",
          4381 => x"ff",
          4382 => x"81",
          4383 => x"55",
          4384 => x"c0",
          4385 => x"0d",
          4386 => x"0d",
          4387 => x"3d",
          4388 => x"9a",
          4389 => x"cb",
          4390 => x"c0",
          4391 => x"de",
          4392 => x"b0",
          4393 => x"69",
          4394 => x"70",
          4395 => x"97",
          4396 => x"c0",
          4397 => x"de",
          4398 => x"38",
          4399 => x"94",
          4400 => x"c0",
          4401 => x"09",
          4402 => x"88",
          4403 => x"df",
          4404 => x"85",
          4405 => x"51",
          4406 => x"74",
          4407 => x"78",
          4408 => x"8a",
          4409 => x"57",
          4410 => x"81",
          4411 => x"75",
          4412 => x"de",
          4413 => x"38",
          4414 => x"de",
          4415 => x"2e",
          4416 => x"83",
          4417 => x"81",
          4418 => x"ff",
          4419 => x"06",
          4420 => x"54",
          4421 => x"73",
          4422 => x"81",
          4423 => x"52",
          4424 => x"a4",
          4425 => x"c0",
          4426 => x"de",
          4427 => x"9a",
          4428 => x"a0",
          4429 => x"51",
          4430 => x"3f",
          4431 => x"0b",
          4432 => x"78",
          4433 => x"bf",
          4434 => x"88",
          4435 => x"80",
          4436 => x"ff",
          4437 => x"75",
          4438 => x"11",
          4439 => x"f8",
          4440 => x"78",
          4441 => x"80",
          4442 => x"ff",
          4443 => x"78",
          4444 => x"80",
          4445 => x"7f",
          4446 => x"d4",
          4447 => x"c9",
          4448 => x"54",
          4449 => x"15",
          4450 => x"cb",
          4451 => x"de",
          4452 => x"81",
          4453 => x"b2",
          4454 => x"b2",
          4455 => x"96",
          4456 => x"b5",
          4457 => x"53",
          4458 => x"51",
          4459 => x"64",
          4460 => x"8b",
          4461 => x"54",
          4462 => x"15",
          4463 => x"ff",
          4464 => x"81",
          4465 => x"54",
          4466 => x"53",
          4467 => x"51",
          4468 => x"3f",
          4469 => x"c0",
          4470 => x"0d",
          4471 => x"0d",
          4472 => x"05",
          4473 => x"3f",
          4474 => x"3d",
          4475 => x"52",
          4476 => x"d5",
          4477 => x"de",
          4478 => x"81",
          4479 => x"82",
          4480 => x"4d",
          4481 => x"52",
          4482 => x"52",
          4483 => x"3f",
          4484 => x"08",
          4485 => x"c0",
          4486 => x"38",
          4487 => x"05",
          4488 => x"06",
          4489 => x"73",
          4490 => x"a0",
          4491 => x"08",
          4492 => x"ff",
          4493 => x"ff",
          4494 => x"ac",
          4495 => x"92",
          4496 => x"54",
          4497 => x"3f",
          4498 => x"52",
          4499 => x"f7",
          4500 => x"c0",
          4501 => x"de",
          4502 => x"38",
          4503 => x"09",
          4504 => x"38",
          4505 => x"08",
          4506 => x"88",
          4507 => x"39",
          4508 => x"08",
          4509 => x"81",
          4510 => x"38",
          4511 => x"b1",
          4512 => x"c0",
          4513 => x"de",
          4514 => x"c8",
          4515 => x"93",
          4516 => x"ff",
          4517 => x"8d",
          4518 => x"b4",
          4519 => x"af",
          4520 => x"17",
          4521 => x"33",
          4522 => x"70",
          4523 => x"55",
          4524 => x"38",
          4525 => x"54",
          4526 => x"34",
          4527 => x"0b",
          4528 => x"8b",
          4529 => x"84",
          4530 => x"06",
          4531 => x"73",
          4532 => x"e5",
          4533 => x"2e",
          4534 => x"75",
          4535 => x"c6",
          4536 => x"de",
          4537 => x"78",
          4538 => x"bb",
          4539 => x"81",
          4540 => x"80",
          4541 => x"38",
          4542 => x"08",
          4543 => x"ff",
          4544 => x"81",
          4545 => x"79",
          4546 => x"58",
          4547 => x"de",
          4548 => x"c0",
          4549 => x"33",
          4550 => x"2e",
          4551 => x"99",
          4552 => x"75",
          4553 => x"c6",
          4554 => x"54",
          4555 => x"15",
          4556 => x"81",
          4557 => x"9c",
          4558 => x"c8",
          4559 => x"de",
          4560 => x"81",
          4561 => x"8c",
          4562 => x"ff",
          4563 => x"81",
          4564 => x"55",
          4565 => x"c0",
          4566 => x"0d",
          4567 => x"0d",
          4568 => x"05",
          4569 => x"05",
          4570 => x"33",
          4571 => x"53",
          4572 => x"05",
          4573 => x"51",
          4574 => x"81",
          4575 => x"55",
          4576 => x"08",
          4577 => x"78",
          4578 => x"95",
          4579 => x"51",
          4580 => x"81",
          4581 => x"55",
          4582 => x"08",
          4583 => x"80",
          4584 => x"81",
          4585 => x"86",
          4586 => x"38",
          4587 => x"61",
          4588 => x"12",
          4589 => x"7a",
          4590 => x"51",
          4591 => x"74",
          4592 => x"78",
          4593 => x"83",
          4594 => x"51",
          4595 => x"3f",
          4596 => x"08",
          4597 => x"de",
          4598 => x"3d",
          4599 => x"3d",
          4600 => x"82",
          4601 => x"d0",
          4602 => x"3d",
          4603 => x"3f",
          4604 => x"08",
          4605 => x"c0",
          4606 => x"38",
          4607 => x"52",
          4608 => x"05",
          4609 => x"3f",
          4610 => x"08",
          4611 => x"c0",
          4612 => x"02",
          4613 => x"33",
          4614 => x"54",
          4615 => x"a6",
          4616 => x"22",
          4617 => x"71",
          4618 => x"53",
          4619 => x"51",
          4620 => x"3f",
          4621 => x"0b",
          4622 => x"76",
          4623 => x"b8",
          4624 => x"c0",
          4625 => x"81",
          4626 => x"93",
          4627 => x"ea",
          4628 => x"6b",
          4629 => x"53",
          4630 => x"05",
          4631 => x"51",
          4632 => x"81",
          4633 => x"81",
          4634 => x"30",
          4635 => x"c0",
          4636 => x"25",
          4637 => x"79",
          4638 => x"85",
          4639 => x"75",
          4640 => x"73",
          4641 => x"f9",
          4642 => x"80",
          4643 => x"8d",
          4644 => x"54",
          4645 => x"3f",
          4646 => x"08",
          4647 => x"c0",
          4648 => x"38",
          4649 => x"51",
          4650 => x"81",
          4651 => x"57",
          4652 => x"08",
          4653 => x"de",
          4654 => x"de",
          4655 => x"5b",
          4656 => x"18",
          4657 => x"18",
          4658 => x"74",
          4659 => x"81",
          4660 => x"78",
          4661 => x"8b",
          4662 => x"54",
          4663 => x"75",
          4664 => x"38",
          4665 => x"1b",
          4666 => x"55",
          4667 => x"2e",
          4668 => x"39",
          4669 => x"09",
          4670 => x"38",
          4671 => x"80",
          4672 => x"70",
          4673 => x"25",
          4674 => x"80",
          4675 => x"38",
          4676 => x"bc",
          4677 => x"11",
          4678 => x"ff",
          4679 => x"81",
          4680 => x"57",
          4681 => x"08",
          4682 => x"70",
          4683 => x"80",
          4684 => x"83",
          4685 => x"80",
          4686 => x"84",
          4687 => x"a7",
          4688 => x"b4",
          4689 => x"ad",
          4690 => x"de",
          4691 => x"0c",
          4692 => x"c0",
          4693 => x"0d",
          4694 => x"0d",
          4695 => x"3d",
          4696 => x"52",
          4697 => x"ce",
          4698 => x"de",
          4699 => x"de",
          4700 => x"54",
          4701 => x"08",
          4702 => x"8b",
          4703 => x"8b",
          4704 => x"59",
          4705 => x"3f",
          4706 => x"33",
          4707 => x"06",
          4708 => x"57",
          4709 => x"81",
          4710 => x"58",
          4711 => x"06",
          4712 => x"4e",
          4713 => x"ff",
          4714 => x"81",
          4715 => x"80",
          4716 => x"6c",
          4717 => x"53",
          4718 => x"ae",
          4719 => x"de",
          4720 => x"2e",
          4721 => x"88",
          4722 => x"6d",
          4723 => x"55",
          4724 => x"de",
          4725 => x"ff",
          4726 => x"83",
          4727 => x"51",
          4728 => x"26",
          4729 => x"15",
          4730 => x"ff",
          4731 => x"80",
          4732 => x"87",
          4733 => x"b4",
          4734 => x"74",
          4735 => x"38",
          4736 => x"ce",
          4737 => x"ae",
          4738 => x"de",
          4739 => x"38",
          4740 => x"27",
          4741 => x"89",
          4742 => x"8b",
          4743 => x"27",
          4744 => x"55",
          4745 => x"81",
          4746 => x"8f",
          4747 => x"2a",
          4748 => x"70",
          4749 => x"34",
          4750 => x"74",
          4751 => x"05",
          4752 => x"17",
          4753 => x"70",
          4754 => x"52",
          4755 => x"73",
          4756 => x"c8",
          4757 => x"33",
          4758 => x"73",
          4759 => x"81",
          4760 => x"80",
          4761 => x"02",
          4762 => x"76",
          4763 => x"51",
          4764 => x"2e",
          4765 => x"87",
          4766 => x"57",
          4767 => x"79",
          4768 => x"80",
          4769 => x"70",
          4770 => x"ba",
          4771 => x"de",
          4772 => x"81",
          4773 => x"80",
          4774 => x"52",
          4775 => x"bf",
          4776 => x"de",
          4777 => x"81",
          4778 => x"8d",
          4779 => x"c4",
          4780 => x"e5",
          4781 => x"c6",
          4782 => x"c0",
          4783 => x"09",
          4784 => x"cc",
          4785 => x"76",
          4786 => x"c4",
          4787 => x"74",
          4788 => x"b0",
          4789 => x"c0",
          4790 => x"de",
          4791 => x"38",
          4792 => x"de",
          4793 => x"67",
          4794 => x"db",
          4795 => x"88",
          4796 => x"34",
          4797 => x"52",
          4798 => x"ab",
          4799 => x"54",
          4800 => x"15",
          4801 => x"ff",
          4802 => x"81",
          4803 => x"54",
          4804 => x"81",
          4805 => x"9c",
          4806 => x"f2",
          4807 => x"62",
          4808 => x"80",
          4809 => x"93",
          4810 => x"55",
          4811 => x"5e",
          4812 => x"3f",
          4813 => x"08",
          4814 => x"c0",
          4815 => x"38",
          4816 => x"58",
          4817 => x"38",
          4818 => x"97",
          4819 => x"08",
          4820 => x"38",
          4821 => x"70",
          4822 => x"81",
          4823 => x"55",
          4824 => x"87",
          4825 => x"39",
          4826 => x"90",
          4827 => x"82",
          4828 => x"8a",
          4829 => x"89",
          4830 => x"7f",
          4831 => x"56",
          4832 => x"3f",
          4833 => x"06",
          4834 => x"72",
          4835 => x"81",
          4836 => x"05",
          4837 => x"7c",
          4838 => x"55",
          4839 => x"27",
          4840 => x"16",
          4841 => x"83",
          4842 => x"76",
          4843 => x"80",
          4844 => x"79",
          4845 => x"99",
          4846 => x"7f",
          4847 => x"14",
          4848 => x"83",
          4849 => x"81",
          4850 => x"81",
          4851 => x"38",
          4852 => x"08",
          4853 => x"95",
          4854 => x"c0",
          4855 => x"81",
          4856 => x"7b",
          4857 => x"06",
          4858 => x"39",
          4859 => x"56",
          4860 => x"09",
          4861 => x"b9",
          4862 => x"80",
          4863 => x"80",
          4864 => x"78",
          4865 => x"7a",
          4866 => x"38",
          4867 => x"73",
          4868 => x"81",
          4869 => x"ff",
          4870 => x"74",
          4871 => x"ff",
          4872 => x"81",
          4873 => x"58",
          4874 => x"08",
          4875 => x"74",
          4876 => x"16",
          4877 => x"73",
          4878 => x"39",
          4879 => x"7e",
          4880 => x"0c",
          4881 => x"2e",
          4882 => x"88",
          4883 => x"8c",
          4884 => x"1a",
          4885 => x"07",
          4886 => x"1b",
          4887 => x"08",
          4888 => x"16",
          4889 => x"75",
          4890 => x"38",
          4891 => x"90",
          4892 => x"15",
          4893 => x"54",
          4894 => x"34",
          4895 => x"81",
          4896 => x"90",
          4897 => x"e9",
          4898 => x"6d",
          4899 => x"80",
          4900 => x"9d",
          4901 => x"5c",
          4902 => x"3f",
          4903 => x"0b",
          4904 => x"08",
          4905 => x"38",
          4906 => x"08",
          4907 => x"de",
          4908 => x"08",
          4909 => x"80",
          4910 => x"80",
          4911 => x"de",
          4912 => x"ff",
          4913 => x"52",
          4914 => x"a0",
          4915 => x"de",
          4916 => x"ff",
          4917 => x"06",
          4918 => x"56",
          4919 => x"38",
          4920 => x"70",
          4921 => x"55",
          4922 => x"8b",
          4923 => x"3d",
          4924 => x"83",
          4925 => x"ff",
          4926 => x"81",
          4927 => x"99",
          4928 => x"74",
          4929 => x"38",
          4930 => x"80",
          4931 => x"ff",
          4932 => x"55",
          4933 => x"83",
          4934 => x"78",
          4935 => x"38",
          4936 => x"26",
          4937 => x"81",
          4938 => x"8b",
          4939 => x"79",
          4940 => x"80",
          4941 => x"93",
          4942 => x"39",
          4943 => x"6e",
          4944 => x"89",
          4945 => x"48",
          4946 => x"83",
          4947 => x"61",
          4948 => x"25",
          4949 => x"55",
          4950 => x"8a",
          4951 => x"3d",
          4952 => x"81",
          4953 => x"ff",
          4954 => x"81",
          4955 => x"c0",
          4956 => x"38",
          4957 => x"70",
          4958 => x"de",
          4959 => x"56",
          4960 => x"38",
          4961 => x"55",
          4962 => x"75",
          4963 => x"38",
          4964 => x"70",
          4965 => x"ff",
          4966 => x"83",
          4967 => x"78",
          4968 => x"89",
          4969 => x"81",
          4970 => x"06",
          4971 => x"80",
          4972 => x"77",
          4973 => x"74",
          4974 => x"8d",
          4975 => x"06",
          4976 => x"2e",
          4977 => x"77",
          4978 => x"93",
          4979 => x"74",
          4980 => x"cb",
          4981 => x"7d",
          4982 => x"81",
          4983 => x"38",
          4984 => x"66",
          4985 => x"81",
          4986 => x"d8",
          4987 => x"74",
          4988 => x"38",
          4989 => x"98",
          4990 => x"d8",
          4991 => x"82",
          4992 => x"57",
          4993 => x"80",
          4994 => x"76",
          4995 => x"38",
          4996 => x"51",
          4997 => x"3f",
          4998 => x"08",
          4999 => x"87",
          5000 => x"2a",
          5001 => x"5c",
          5002 => x"de",
          5003 => x"80",
          5004 => x"44",
          5005 => x"0a",
          5006 => x"ec",
          5007 => x"39",
          5008 => x"66",
          5009 => x"81",
          5010 => x"c8",
          5011 => x"74",
          5012 => x"38",
          5013 => x"98",
          5014 => x"c8",
          5015 => x"82",
          5016 => x"57",
          5017 => x"80",
          5018 => x"76",
          5019 => x"38",
          5020 => x"51",
          5021 => x"3f",
          5022 => x"08",
          5023 => x"57",
          5024 => x"08",
          5025 => x"96",
          5026 => x"81",
          5027 => x"10",
          5028 => x"08",
          5029 => x"72",
          5030 => x"59",
          5031 => x"ff",
          5032 => x"5d",
          5033 => x"44",
          5034 => x"11",
          5035 => x"70",
          5036 => x"71",
          5037 => x"06",
          5038 => x"52",
          5039 => x"40",
          5040 => x"09",
          5041 => x"38",
          5042 => x"18",
          5043 => x"39",
          5044 => x"79",
          5045 => x"70",
          5046 => x"58",
          5047 => x"76",
          5048 => x"38",
          5049 => x"7d",
          5050 => x"70",
          5051 => x"55",
          5052 => x"3f",
          5053 => x"08",
          5054 => x"2e",
          5055 => x"9b",
          5056 => x"c0",
          5057 => x"f5",
          5058 => x"38",
          5059 => x"38",
          5060 => x"59",
          5061 => x"38",
          5062 => x"7d",
          5063 => x"81",
          5064 => x"38",
          5065 => x"0b",
          5066 => x"08",
          5067 => x"78",
          5068 => x"1a",
          5069 => x"c0",
          5070 => x"74",
          5071 => x"39",
          5072 => x"55",
          5073 => x"8f",
          5074 => x"fd",
          5075 => x"de",
          5076 => x"f5",
          5077 => x"78",
          5078 => x"79",
          5079 => x"80",
          5080 => x"f1",
          5081 => x"39",
          5082 => x"81",
          5083 => x"06",
          5084 => x"55",
          5085 => x"27",
          5086 => x"81",
          5087 => x"56",
          5088 => x"38",
          5089 => x"80",
          5090 => x"ff",
          5091 => x"8b",
          5092 => x"f0",
          5093 => x"ff",
          5094 => x"84",
          5095 => x"1b",
          5096 => x"b3",
          5097 => x"1c",
          5098 => x"ff",
          5099 => x"8e",
          5100 => x"a1",
          5101 => x"0b",
          5102 => x"7d",
          5103 => x"30",
          5104 => x"84",
          5105 => x"51",
          5106 => x"51",
          5107 => x"3f",
          5108 => x"83",
          5109 => x"90",
          5110 => x"ff",
          5111 => x"93",
          5112 => x"a0",
          5113 => x"39",
          5114 => x"1b",
          5115 => x"85",
          5116 => x"95",
          5117 => x"52",
          5118 => x"ff",
          5119 => x"81",
          5120 => x"1b",
          5121 => x"cf",
          5122 => x"9c",
          5123 => x"a0",
          5124 => x"83",
          5125 => x"06",
          5126 => x"82",
          5127 => x"52",
          5128 => x"51",
          5129 => x"3f",
          5130 => x"1b",
          5131 => x"c5",
          5132 => x"ac",
          5133 => x"a0",
          5134 => x"52",
          5135 => x"ff",
          5136 => x"86",
          5137 => x"51",
          5138 => x"3f",
          5139 => x"80",
          5140 => x"a9",
          5141 => x"1c",
          5142 => x"81",
          5143 => x"80",
          5144 => x"ae",
          5145 => x"b2",
          5146 => x"1b",
          5147 => x"85",
          5148 => x"ff",
          5149 => x"96",
          5150 => x"9f",
          5151 => x"80",
          5152 => x"34",
          5153 => x"1c",
          5154 => x"81",
          5155 => x"ab",
          5156 => x"a0",
          5157 => x"d4",
          5158 => x"fe",
          5159 => x"59",
          5160 => x"3f",
          5161 => x"53",
          5162 => x"51",
          5163 => x"3f",
          5164 => x"de",
          5165 => x"e7",
          5166 => x"2e",
          5167 => x"80",
          5168 => x"54",
          5169 => x"53",
          5170 => x"51",
          5171 => x"3f",
          5172 => x"80",
          5173 => x"ff",
          5174 => x"84",
          5175 => x"d2",
          5176 => x"ff",
          5177 => x"86",
          5178 => x"f2",
          5179 => x"1b",
          5180 => x"81",
          5181 => x"52",
          5182 => x"51",
          5183 => x"3f",
          5184 => x"ec",
          5185 => x"9e",
          5186 => x"d4",
          5187 => x"51",
          5188 => x"3f",
          5189 => x"87",
          5190 => x"52",
          5191 => x"9a",
          5192 => x"54",
          5193 => x"7a",
          5194 => x"ff",
          5195 => x"65",
          5196 => x"7a",
          5197 => x"8f",
          5198 => x"80",
          5199 => x"2e",
          5200 => x"9a",
          5201 => x"7a",
          5202 => x"a9",
          5203 => x"84",
          5204 => x"9e",
          5205 => x"0a",
          5206 => x"51",
          5207 => x"ff",
          5208 => x"7d",
          5209 => x"38",
          5210 => x"52",
          5211 => x"9e",
          5212 => x"55",
          5213 => x"62",
          5214 => x"74",
          5215 => x"75",
          5216 => x"7e",
          5217 => x"fe",
          5218 => x"c0",
          5219 => x"38",
          5220 => x"81",
          5221 => x"52",
          5222 => x"9e",
          5223 => x"16",
          5224 => x"56",
          5225 => x"38",
          5226 => x"77",
          5227 => x"8d",
          5228 => x"7d",
          5229 => x"38",
          5230 => x"57",
          5231 => x"83",
          5232 => x"76",
          5233 => x"7a",
          5234 => x"ff",
          5235 => x"81",
          5236 => x"81",
          5237 => x"16",
          5238 => x"56",
          5239 => x"38",
          5240 => x"83",
          5241 => x"86",
          5242 => x"ff",
          5243 => x"38",
          5244 => x"82",
          5245 => x"81",
          5246 => x"06",
          5247 => x"fe",
          5248 => x"53",
          5249 => x"51",
          5250 => x"3f",
          5251 => x"52",
          5252 => x"9c",
          5253 => x"be",
          5254 => x"75",
          5255 => x"81",
          5256 => x"0b",
          5257 => x"77",
          5258 => x"75",
          5259 => x"60",
          5260 => x"80",
          5261 => x"75",
          5262 => x"be",
          5263 => x"85",
          5264 => x"de",
          5265 => x"2a",
          5266 => x"75",
          5267 => x"81",
          5268 => x"87",
          5269 => x"52",
          5270 => x"51",
          5271 => x"3f",
          5272 => x"ca",
          5273 => x"9c",
          5274 => x"54",
          5275 => x"52",
          5276 => x"98",
          5277 => x"56",
          5278 => x"08",
          5279 => x"53",
          5280 => x"51",
          5281 => x"3f",
          5282 => x"de",
          5283 => x"38",
          5284 => x"56",
          5285 => x"56",
          5286 => x"de",
          5287 => x"75",
          5288 => x"0c",
          5289 => x"04",
          5290 => x"7d",
          5291 => x"80",
          5292 => x"05",
          5293 => x"76",
          5294 => x"38",
          5295 => x"11",
          5296 => x"53",
          5297 => x"79",
          5298 => x"3f",
          5299 => x"09",
          5300 => x"38",
          5301 => x"55",
          5302 => x"db",
          5303 => x"70",
          5304 => x"34",
          5305 => x"74",
          5306 => x"81",
          5307 => x"80",
          5308 => x"55",
          5309 => x"76",
          5310 => x"de",
          5311 => x"3d",
          5312 => x"3d",
          5313 => x"71",
          5314 => x"8e",
          5315 => x"29",
          5316 => x"05",
          5317 => x"04",
          5318 => x"51",
          5319 => x"81",
          5320 => x"80",
          5321 => x"d0",
          5322 => x"f2",
          5323 => x"a4",
          5324 => x"39",
          5325 => x"51",
          5326 => x"81",
          5327 => x"80",
          5328 => x"d0",
          5329 => x"d6",
          5330 => x"e8",
          5331 => x"39",
          5332 => x"51",
          5333 => x"81",
          5334 => x"80",
          5335 => x"d1",
          5336 => x"39",
          5337 => x"51",
          5338 => x"d1",
          5339 => x"39",
          5340 => x"51",
          5341 => x"d2",
          5342 => x"39",
          5343 => x"51",
          5344 => x"d2",
          5345 => x"39",
          5346 => x"51",
          5347 => x"d3",
          5348 => x"39",
          5349 => x"51",
          5350 => x"d3",
          5351 => x"87",
          5352 => x"3d",
          5353 => x"3d",
          5354 => x"56",
          5355 => x"e7",
          5356 => x"74",
          5357 => x"e8",
          5358 => x"39",
          5359 => x"74",
          5360 => x"b6",
          5361 => x"c0",
          5362 => x"51",
          5363 => x"3f",
          5364 => x"08",
          5365 => x"75",
          5366 => x"b8",
          5367 => x"c6",
          5368 => x"0d",
          5369 => x"0d",
          5370 => x"02",
          5371 => x"c7",
          5372 => x"73",
          5373 => x"5d",
          5374 => x"5c",
          5375 => x"81",
          5376 => x"ff",
          5377 => x"81",
          5378 => x"ff",
          5379 => x"80",
          5380 => x"27",
          5381 => x"79",
          5382 => x"38",
          5383 => x"a7",
          5384 => x"39",
          5385 => x"72",
          5386 => x"38",
          5387 => x"81",
          5388 => x"ff",
          5389 => x"89",
          5390 => x"f4",
          5391 => x"82",
          5392 => x"55",
          5393 => x"74",
          5394 => x"78",
          5395 => x"72",
          5396 => x"d3",
          5397 => x"8b",
          5398 => x"39",
          5399 => x"51",
          5400 => x"3f",
          5401 => x"a1",
          5402 => x"53",
          5403 => x"8e",
          5404 => x"52",
          5405 => x"51",
          5406 => x"3f",
          5407 => x"d4",
          5408 => x"85",
          5409 => x"15",
          5410 => x"fe",
          5411 => x"ff",
          5412 => x"d4",
          5413 => x"85",
          5414 => x"55",
          5415 => x"aa",
          5416 => x"70",
          5417 => x"26",
          5418 => x"9f",
          5419 => x"38",
          5420 => x"8b",
          5421 => x"fe",
          5422 => x"73",
          5423 => x"a0",
          5424 => x"f9",
          5425 => x"55",
          5426 => x"d4",
          5427 => x"84",
          5428 => x"16",
          5429 => x"56",
          5430 => x"3f",
          5431 => x"08",
          5432 => x"98",
          5433 => x"74",
          5434 => x"81",
          5435 => x"fe",
          5436 => x"81",
          5437 => x"98",
          5438 => x"2c",
          5439 => x"70",
          5440 => x"07",
          5441 => x"56",
          5442 => x"74",
          5443 => x"38",
          5444 => x"74",
          5445 => x"81",
          5446 => x"80",
          5447 => x"7a",
          5448 => x"76",
          5449 => x"38",
          5450 => x"81",
          5451 => x"8d",
          5452 => x"ec",
          5453 => x"02",
          5454 => x"e3",
          5455 => x"72",
          5456 => x"07",
          5457 => x"87",
          5458 => x"07",
          5459 => x"5a",
          5460 => x"57",
          5461 => x"38",
          5462 => x"52",
          5463 => x"52",
          5464 => x"de",
          5465 => x"c0",
          5466 => x"de",
          5467 => x"38",
          5468 => x"08",
          5469 => x"88",
          5470 => x"c0",
          5471 => x"3d",
          5472 => x"84",
          5473 => x"52",
          5474 => x"9b",
          5475 => x"c0",
          5476 => x"de",
          5477 => x"38",
          5478 => x"80",
          5479 => x"74",
          5480 => x"59",
          5481 => x"96",
          5482 => x"51",
          5483 => x"75",
          5484 => x"07",
          5485 => x"55",
          5486 => x"95",
          5487 => x"2e",
          5488 => x"d4",
          5489 => x"c0",
          5490 => x"52",
          5491 => x"d6",
          5492 => x"76",
          5493 => x"0c",
          5494 => x"04",
          5495 => x"7b",
          5496 => x"b3",
          5497 => x"58",
          5498 => x"53",
          5499 => x"51",
          5500 => x"81",
          5501 => x"a4",
          5502 => x"2e",
          5503 => x"81",
          5504 => x"98",
          5505 => x"7f",
          5506 => x"c0",
          5507 => x"7d",
          5508 => x"81",
          5509 => x"57",
          5510 => x"04",
          5511 => x"c0",
          5512 => x"0d",
          5513 => x"0d",
          5514 => x"33",
          5515 => x"53",
          5516 => x"52",
          5517 => x"ee",
          5518 => x"c0",
          5519 => x"80",
          5520 => x"d4",
          5521 => x"d4",
          5522 => x"db",
          5523 => x"81",
          5524 => x"ff",
          5525 => x"74",
          5526 => x"38",
          5527 => x"3f",
          5528 => x"04",
          5529 => x"87",
          5530 => x"08",
          5531 => x"a2",
          5532 => x"fe",
          5533 => x"81",
          5534 => x"fe",
          5535 => x"80",
          5536 => x"9f",
          5537 => x"2a",
          5538 => x"51",
          5539 => x"2e",
          5540 => x"51",
          5541 => x"3f",
          5542 => x"51",
          5543 => x"3f",
          5544 => x"f1",
          5545 => x"82",
          5546 => x"06",
          5547 => x"80",
          5548 => x"81",
          5549 => x"eb",
          5550 => x"8c",
          5551 => x"e3",
          5552 => x"fe",
          5553 => x"72",
          5554 => x"81",
          5555 => x"71",
          5556 => x"38",
          5557 => x"f1",
          5558 => x"d5",
          5559 => x"f3",
          5560 => x"51",
          5561 => x"3f",
          5562 => x"70",
          5563 => x"52",
          5564 => x"95",
          5565 => x"fe",
          5566 => x"81",
          5567 => x"fe",
          5568 => x"80",
          5569 => x"9b",
          5570 => x"2a",
          5571 => x"51",
          5572 => x"2e",
          5573 => x"51",
          5574 => x"3f",
          5575 => x"51",
          5576 => x"3f",
          5577 => x"f0",
          5578 => x"86",
          5579 => x"06",
          5580 => x"80",
          5581 => x"81",
          5582 => x"e7",
          5583 => x"d8",
          5584 => x"df",
          5585 => x"fe",
          5586 => x"72",
          5587 => x"81",
          5588 => x"71",
          5589 => x"38",
          5590 => x"f0",
          5591 => x"d5",
          5592 => x"f2",
          5593 => x"51",
          5594 => x"3f",
          5595 => x"70",
          5596 => x"52",
          5597 => x"95",
          5598 => x"fe",
          5599 => x"81",
          5600 => x"fe",
          5601 => x"80",
          5602 => x"97",
          5603 => x"cb",
          5604 => x"0d",
          5605 => x"0d",
          5606 => x"70",
          5607 => x"73",
          5608 => x"f0",
          5609 => x"73",
          5610 => x"15",
          5611 => x"e4",
          5612 => x"54",
          5613 => x"70",
          5614 => x"57",
          5615 => x"a0",
          5616 => x"81",
          5617 => x"2e",
          5618 => x"e5",
          5619 => x"ff",
          5620 => x"a0",
          5621 => x"06",
          5622 => x"74",
          5623 => x"56",
          5624 => x"75",
          5625 => x"db",
          5626 => x"08",
          5627 => x"52",
          5628 => x"9e",
          5629 => x"c0",
          5630 => x"84",
          5631 => x"72",
          5632 => x"a3",
          5633 => x"70",
          5634 => x"57",
          5635 => x"27",
          5636 => x"53",
          5637 => x"c0",
          5638 => x"0d",
          5639 => x"0d",
          5640 => x"55",
          5641 => x"52",
          5642 => x"e8",
          5643 => x"db",
          5644 => x"73",
          5645 => x"53",
          5646 => x"52",
          5647 => x"51",
          5648 => x"3f",
          5649 => x"08",
          5650 => x"de",
          5651 => x"80",
          5652 => x"31",
          5653 => x"73",
          5654 => x"34",
          5655 => x"33",
          5656 => x"2e",
          5657 => x"ac",
          5658 => x"c4",
          5659 => x"75",
          5660 => x"3f",
          5661 => x"08",
          5662 => x"38",
          5663 => x"08",
          5664 => x"be",
          5665 => x"81",
          5666 => x"c6",
          5667 => x"0b",
          5668 => x"34",
          5669 => x"33",
          5670 => x"2e",
          5671 => x"89",
          5672 => x"75",
          5673 => x"d8",
          5674 => x"81",
          5675 => x"87",
          5676 => x"cb",
          5677 => x"70",
          5678 => x"c0",
          5679 => x"81",
          5680 => x"ff",
          5681 => x"81",
          5682 => x"81",
          5683 => x"78",
          5684 => x"81",
          5685 => x"81",
          5686 => x"99",
          5687 => x"59",
          5688 => x"3f",
          5689 => x"52",
          5690 => x"51",
          5691 => x"3f",
          5692 => x"08",
          5693 => x"38",
          5694 => x"51",
          5695 => x"81",
          5696 => x"81",
          5697 => x"fe",
          5698 => x"99",
          5699 => x"5a",
          5700 => x"79",
          5701 => x"3f",
          5702 => x"f8",
          5703 => x"f5",
          5704 => x"c0",
          5705 => x"70",
          5706 => x"59",
          5707 => x"2e",
          5708 => x"78",
          5709 => x"80",
          5710 => x"ab",
          5711 => x"38",
          5712 => x"a4",
          5713 => x"2e",
          5714 => x"78",
          5715 => x"38",
          5716 => x"ff",
          5717 => x"de",
          5718 => x"2e",
          5719 => x"78",
          5720 => x"ad",
          5721 => x"39",
          5722 => x"2e",
          5723 => x"78",
          5724 => x"90",
          5725 => x"2e",
          5726 => x"78",
          5727 => x"8b",
          5728 => x"39",
          5729 => x"2e",
          5730 => x"78",
          5731 => x"88",
          5732 => x"a2",
          5733 => x"d5",
          5734 => x"38",
          5735 => x"24",
          5736 => x"80",
          5737 => x"a7",
          5738 => x"d0",
          5739 => x"78",
          5740 => x"8a",
          5741 => x"fe",
          5742 => x"d1",
          5743 => x"38",
          5744 => x"2e",
          5745 => x"8e",
          5746 => x"81",
          5747 => x"c3",
          5748 => x"82",
          5749 => x"78",
          5750 => x"8d",
          5751 => x"80",
          5752 => x"ec",
          5753 => x"39",
          5754 => x"2e",
          5755 => x"78",
          5756 => x"8e",
          5757 => x"be",
          5758 => x"fe",
          5759 => x"fe",
          5760 => x"ff",
          5761 => x"81",
          5762 => x"88",
          5763 => x"90",
          5764 => x"39",
          5765 => x"f0",
          5766 => x"f8",
          5767 => x"81",
          5768 => x"de",
          5769 => x"2e",
          5770 => x"63",
          5771 => x"80",
          5772 => x"cb",
          5773 => x"02",
          5774 => x"33",
          5775 => x"dd",
          5776 => x"c0",
          5777 => x"06",
          5778 => x"38",
          5779 => x"51",
          5780 => x"3f",
          5781 => x"ab",
          5782 => x"b0",
          5783 => x"39",
          5784 => x"f4",
          5785 => x"f8",
          5786 => x"81",
          5787 => x"de",
          5788 => x"2e",
          5789 => x"80",
          5790 => x"02",
          5791 => x"33",
          5792 => x"e6",
          5793 => x"c0",
          5794 => x"d7",
          5795 => x"fc",
          5796 => x"fe",
          5797 => x"fe",
          5798 => x"ff",
          5799 => x"81",
          5800 => x"80",
          5801 => x"63",
          5802 => x"d7",
          5803 => x"fe",
          5804 => x"fe",
          5805 => x"ff",
          5806 => x"81",
          5807 => x"86",
          5808 => x"c0",
          5809 => x"53",
          5810 => x"52",
          5811 => x"fe",
          5812 => x"80",
          5813 => x"53",
          5814 => x"84",
          5815 => x"df",
          5816 => x"ff",
          5817 => x"81",
          5818 => x"81",
          5819 => x"d7",
          5820 => x"f8",
          5821 => x"5d",
          5822 => x"b7",
          5823 => x"05",
          5824 => x"d0",
          5825 => x"c0",
          5826 => x"fe",
          5827 => x"5b",
          5828 => x"3f",
          5829 => x"de",
          5830 => x"7a",
          5831 => x"3f",
          5832 => x"b7",
          5833 => x"05",
          5834 => x"a8",
          5835 => x"c0",
          5836 => x"fe",
          5837 => x"5b",
          5838 => x"3f",
          5839 => x"08",
          5840 => x"f8",
          5841 => x"fe",
          5842 => x"81",
          5843 => x"b8",
          5844 => x"05",
          5845 => x"e5",
          5846 => x"db",
          5847 => x"de",
          5848 => x"56",
          5849 => x"de",
          5850 => x"ff",
          5851 => x"53",
          5852 => x"51",
          5853 => x"81",
          5854 => x"80",
          5855 => x"38",
          5856 => x"08",
          5857 => x"3f",
          5858 => x"b7",
          5859 => x"11",
          5860 => x"05",
          5861 => x"83",
          5862 => x"c0",
          5863 => x"fa",
          5864 => x"3d",
          5865 => x"53",
          5866 => x"51",
          5867 => x"3f",
          5868 => x"08",
          5869 => x"cb",
          5870 => x"fe",
          5871 => x"fe",
          5872 => x"fe",
          5873 => x"81",
          5874 => x"86",
          5875 => x"c0",
          5876 => x"d7",
          5877 => x"f6",
          5878 => x"63",
          5879 => x"7b",
          5880 => x"38",
          5881 => x"7a",
          5882 => x"5c",
          5883 => x"26",
          5884 => x"d5",
          5885 => x"fe",
          5886 => x"fe",
          5887 => x"fe",
          5888 => x"81",
          5889 => x"80",
          5890 => x"db",
          5891 => x"78",
          5892 => x"38",
          5893 => x"08",
          5894 => x"39",
          5895 => x"33",
          5896 => x"2e",
          5897 => x"db",
          5898 => x"bc",
          5899 => x"d6",
          5900 => x"80",
          5901 => x"81",
          5902 => x"44",
          5903 => x"db",
          5904 => x"78",
          5905 => x"38",
          5906 => x"08",
          5907 => x"81",
          5908 => x"59",
          5909 => x"88",
          5910 => x"ac",
          5911 => x"39",
          5912 => x"08",
          5913 => x"44",
          5914 => x"f0",
          5915 => x"f8",
          5916 => x"fd",
          5917 => x"de",
          5918 => x"de",
          5919 => x"d4",
          5920 => x"80",
          5921 => x"81",
          5922 => x"43",
          5923 => x"81",
          5924 => x"59",
          5925 => x"88",
          5926 => x"98",
          5927 => x"39",
          5928 => x"33",
          5929 => x"2e",
          5930 => x"db",
          5931 => x"aa",
          5932 => x"d7",
          5933 => x"80",
          5934 => x"81",
          5935 => x"43",
          5936 => x"db",
          5937 => x"78",
          5938 => x"38",
          5939 => x"08",
          5940 => x"81",
          5941 => x"88",
          5942 => x"3d",
          5943 => x"53",
          5944 => x"51",
          5945 => x"3f",
          5946 => x"08",
          5947 => x"38",
          5948 => x"59",
          5949 => x"83",
          5950 => x"79",
          5951 => x"38",
          5952 => x"88",
          5953 => x"2e",
          5954 => x"42",
          5955 => x"51",
          5956 => x"3f",
          5957 => x"54",
          5958 => x"52",
          5959 => x"c5",
          5960 => x"f4",
          5961 => x"39",
          5962 => x"f4",
          5963 => x"f8",
          5964 => x"fb",
          5965 => x"de",
          5966 => x"2e",
          5967 => x"b7",
          5968 => x"11",
          5969 => x"05",
          5970 => x"cf",
          5971 => x"c0",
          5972 => x"a5",
          5973 => x"02",
          5974 => x"33",
          5975 => x"81",
          5976 => x"3d",
          5977 => x"53",
          5978 => x"51",
          5979 => x"3f",
          5980 => x"08",
          5981 => x"8b",
          5982 => x"33",
          5983 => x"d8",
          5984 => x"f9",
          5985 => x"f8",
          5986 => x"fe",
          5987 => x"79",
          5988 => x"59",
          5989 => x"f6",
          5990 => x"79",
          5991 => x"b7",
          5992 => x"11",
          5993 => x"05",
          5994 => x"ef",
          5995 => x"c0",
          5996 => x"91",
          5997 => x"02",
          5998 => x"33",
          5999 => x"81",
          6000 => x"b5",
          6001 => x"8c",
          6002 => x"f6",
          6003 => x"39",
          6004 => x"e8",
          6005 => x"f8",
          6006 => x"fc",
          6007 => x"de",
          6008 => x"2e",
          6009 => x"b7",
          6010 => x"11",
          6011 => x"05",
          6012 => x"99",
          6013 => x"c0",
          6014 => x"a6",
          6015 => x"02",
          6016 => x"79",
          6017 => x"5b",
          6018 => x"b7",
          6019 => x"11",
          6020 => x"05",
          6021 => x"f5",
          6022 => x"c0",
          6023 => x"f5",
          6024 => x"70",
          6025 => x"81",
          6026 => x"fe",
          6027 => x"80",
          6028 => x"51",
          6029 => x"3f",
          6030 => x"33",
          6031 => x"2e",
          6032 => x"78",
          6033 => x"38",
          6034 => x"41",
          6035 => x"3d",
          6036 => x"53",
          6037 => x"51",
          6038 => x"3f",
          6039 => x"08",
          6040 => x"38",
          6041 => x"be",
          6042 => x"70",
          6043 => x"23",
          6044 => x"ae",
          6045 => x"8c",
          6046 => x"c6",
          6047 => x"39",
          6048 => x"e8",
          6049 => x"f8",
          6050 => x"fb",
          6051 => x"de",
          6052 => x"2e",
          6053 => x"b7",
          6054 => x"11",
          6055 => x"05",
          6056 => x"e9",
          6057 => x"c0",
          6058 => x"a1",
          6059 => x"71",
          6060 => x"84",
          6061 => x"3d",
          6062 => x"53",
          6063 => x"51",
          6064 => x"3f",
          6065 => x"08",
          6066 => x"b7",
          6067 => x"08",
          6068 => x"d8",
          6069 => x"f6",
          6070 => x"f8",
          6071 => x"fe",
          6072 => x"79",
          6073 => x"59",
          6074 => x"f4",
          6075 => x"79",
          6076 => x"b7",
          6077 => x"11",
          6078 => x"05",
          6079 => x"8d",
          6080 => x"c0",
          6081 => x"8d",
          6082 => x"71",
          6083 => x"84",
          6084 => x"b9",
          6085 => x"8c",
          6086 => x"a6",
          6087 => x"39",
          6088 => x"f4",
          6089 => x"f8",
          6090 => x"f7",
          6091 => x"de",
          6092 => x"df",
          6093 => x"d4",
          6094 => x"80",
          6095 => x"81",
          6096 => x"44",
          6097 => x"81",
          6098 => x"59",
          6099 => x"88",
          6100 => x"94",
          6101 => x"39",
          6102 => x"33",
          6103 => x"2e",
          6104 => x"db",
          6105 => x"ab",
          6106 => x"d7",
          6107 => x"80",
          6108 => x"81",
          6109 => x"44",
          6110 => x"db",
          6111 => x"78",
          6112 => x"38",
          6113 => x"08",
          6114 => x"81",
          6115 => x"fc",
          6116 => x"b7",
          6117 => x"11",
          6118 => x"05",
          6119 => x"fb",
          6120 => x"c0",
          6121 => x"38",
          6122 => x"33",
          6123 => x"2e",
          6124 => x"db",
          6125 => x"80",
          6126 => x"db",
          6127 => x"78",
          6128 => x"38",
          6129 => x"08",
          6130 => x"81",
          6131 => x"59",
          6132 => x"88",
          6133 => x"a0",
          6134 => x"39",
          6135 => x"33",
          6136 => x"2e",
          6137 => x"db",
          6138 => x"99",
          6139 => x"d2",
          6140 => x"80",
          6141 => x"81",
          6142 => x"43",
          6143 => x"db",
          6144 => x"05",
          6145 => x"fe",
          6146 => x"fe",
          6147 => x"fe",
          6148 => x"81",
          6149 => x"86",
          6150 => x"c0",
          6151 => x"d8",
          6152 => x"ee",
          6153 => x"5a",
          6154 => x"9d",
          6155 => x"59",
          6156 => x"09",
          6157 => x"38",
          6158 => x"52",
          6159 => x"51",
          6160 => x"3f",
          6161 => x"e0",
          6162 => x"9c",
          6163 => x"81",
          6164 => x"fe",
          6165 => x"82",
          6166 => x"da",
          6167 => x"39",
          6168 => x"51",
          6169 => x"3f",
          6170 => x"ec",
          6171 => x"93",
          6172 => x"81",
          6173 => x"94",
          6174 => x"80",
          6175 => x"c0",
          6176 => x"81",
          6177 => x"fe",
          6178 => x"f0",
          6179 => x"d9",
          6180 => x"ed",
          6181 => x"80",
          6182 => x"c0",
          6183 => x"8c",
          6184 => x"87",
          6185 => x"0c",
          6186 => x"b7",
          6187 => x"11",
          6188 => x"05",
          6189 => x"e3",
          6190 => x"c0",
          6191 => x"f0",
          6192 => x"52",
          6193 => x"51",
          6194 => x"3f",
          6195 => x"04",
          6196 => x"f4",
          6197 => x"f8",
          6198 => x"f4",
          6199 => x"de",
          6200 => x"2e",
          6201 => x"63",
          6202 => x"c0",
          6203 => x"b6",
          6204 => x"78",
          6205 => x"c0",
          6206 => x"de",
          6207 => x"2e",
          6208 => x"81",
          6209 => x"52",
          6210 => x"51",
          6211 => x"3f",
          6212 => x"81",
          6213 => x"fe",
          6214 => x"fe",
          6215 => x"ef",
          6216 => x"da",
          6217 => x"ec",
          6218 => x"59",
          6219 => x"fe",
          6220 => x"ef",
          6221 => x"70",
          6222 => x"78",
          6223 => x"c3",
          6224 => x"2e",
          6225 => x"81",
          6226 => x"5a",
          6227 => x"2e",
          6228 => x"b7",
          6229 => x"05",
          6230 => x"f8",
          6231 => x"c0",
          6232 => x"5b",
          6233 => x"b2",
          6234 => x"24",
          6235 => x"81",
          6236 => x"80",
          6237 => x"83",
          6238 => x"80",
          6239 => x"da",
          6240 => x"55",
          6241 => x"54",
          6242 => x"da",
          6243 => x"3d",
          6244 => x"51",
          6245 => x"3f",
          6246 => x"da",
          6247 => x"3d",
          6248 => x"51",
          6249 => x"3f",
          6250 => x"55",
          6251 => x"54",
          6252 => x"da",
          6253 => x"3d",
          6254 => x"51",
          6255 => x"3f",
          6256 => x"54",
          6257 => x"da",
          6258 => x"3d",
          6259 => x"51",
          6260 => x"3f",
          6261 => x"58",
          6262 => x"57",
          6263 => x"81",
          6264 => x"05",
          6265 => x"82",
          6266 => x"82",
          6267 => x"b7",
          6268 => x"05",
          6269 => x"3f",
          6270 => x"08",
          6271 => x"08",
          6272 => x"70",
          6273 => x"25",
          6274 => x"5e",
          6275 => x"92",
          6276 => x"2e",
          6277 => x"1c",
          6278 => x"06",
          6279 => x"fe",
          6280 => x"81",
          6281 => x"32",
          6282 => x"8a",
          6283 => x"2e",
          6284 => x"ed",
          6285 => x"da",
          6286 => x"ef",
          6287 => x"c3",
          6288 => x"0d",
          6289 => x"de",
          6290 => x"c0",
          6291 => x"08",
          6292 => x"84",
          6293 => x"51",
          6294 => x"3f",
          6295 => x"08",
          6296 => x"08",
          6297 => x"84",
          6298 => x"51",
          6299 => x"3f",
          6300 => x"c0",
          6301 => x"0c",
          6302 => x"9c",
          6303 => x"55",
          6304 => x"52",
          6305 => x"cd",
          6306 => x"de",
          6307 => x"2b",
          6308 => x"53",
          6309 => x"52",
          6310 => x"cd",
          6311 => x"81",
          6312 => x"07",
          6313 => x"80",
          6314 => x"c0",
          6315 => x"8c",
          6316 => x"87",
          6317 => x"0c",
          6318 => x"81",
          6319 => x"a2",
          6320 => x"de",
          6321 => x"de",
          6322 => x"e7",
          6323 => x"da",
          6324 => x"db",
          6325 => x"da",
          6326 => x"e8",
          6327 => x"ac",
          6328 => x"e7",
          6329 => x"51",
          6330 => x"eb",
          6331 => x"04",
          6332 => x"00",
          6333 => x"ff",
          6334 => x"ff",
          6335 => x"ff",
          6336 => x"00",
          6337 => x"00",
          6338 => x"00",
          6339 => x"00",
          6340 => x"00",
          6341 => x"00",
          6342 => x"00",
          6343 => x"00",
          6344 => x"00",
          6345 => x"00",
          6346 => x"00",
          6347 => x"00",
          6348 => x"00",
          6349 => x"00",
          6350 => x"00",
          6351 => x"00",
          6352 => x"00",
          6353 => x"00",
          6354 => x"00",
          6355 => x"00",
          6356 => x"00",
          6357 => x"00",
          6358 => x"00",
          6359 => x"00",
          6360 => x"00",
          6361 => x"25",
          6362 => x"64",
          6363 => x"20",
          6364 => x"25",
          6365 => x"64",
          6366 => x"25",
          6367 => x"53",
          6368 => x"43",
          6369 => x"69",
          6370 => x"61",
          6371 => x"6e",
          6372 => x"20",
          6373 => x"6f",
          6374 => x"6f",
          6375 => x"6f",
          6376 => x"67",
          6377 => x"3a",
          6378 => x"76",
          6379 => x"73",
          6380 => x"70",
          6381 => x"65",
          6382 => x"64",
          6383 => x"20",
          6384 => x"57",
          6385 => x"44",
          6386 => x"20",
          6387 => x"30",
          6388 => x"25",
          6389 => x"29",
          6390 => x"20",
          6391 => x"53",
          6392 => x"4d",
          6393 => x"20",
          6394 => x"30",
          6395 => x"25",
          6396 => x"29",
          6397 => x"20",
          6398 => x"49",
          6399 => x"20",
          6400 => x"4d",
          6401 => x"30",
          6402 => x"25",
          6403 => x"29",
          6404 => x"20",
          6405 => x"42",
          6406 => x"20",
          6407 => x"20",
          6408 => x"30",
          6409 => x"25",
          6410 => x"29",
          6411 => x"20",
          6412 => x"52",
          6413 => x"20",
          6414 => x"20",
          6415 => x"30",
          6416 => x"25",
          6417 => x"29",
          6418 => x"20",
          6419 => x"53",
          6420 => x"41",
          6421 => x"20",
          6422 => x"65",
          6423 => x"65",
          6424 => x"25",
          6425 => x"29",
          6426 => x"20",
          6427 => x"54",
          6428 => x"52",
          6429 => x"20",
          6430 => x"69",
          6431 => x"73",
          6432 => x"25",
          6433 => x"29",
          6434 => x"20",
          6435 => x"49",
          6436 => x"20",
          6437 => x"4c",
          6438 => x"68",
          6439 => x"65",
          6440 => x"25",
          6441 => x"29",
          6442 => x"20",
          6443 => x"57",
          6444 => x"42",
          6445 => x"20",
          6446 => x"0a",
          6447 => x"20",
          6448 => x"57",
          6449 => x"32",
          6450 => x"20",
          6451 => x"49",
          6452 => x"4c",
          6453 => x"20",
          6454 => x"50",
          6455 => x"00",
          6456 => x"20",
          6457 => x"53",
          6458 => x"00",
          6459 => x"41",
          6460 => x"65",
          6461 => x"73",
          6462 => x"20",
          6463 => x"43",
          6464 => x"52",
          6465 => x"74",
          6466 => x"63",
          6467 => x"20",
          6468 => x"72",
          6469 => x"20",
          6470 => x"30",
          6471 => x"00",
          6472 => x"20",
          6473 => x"43",
          6474 => x"4d",
          6475 => x"72",
          6476 => x"74",
          6477 => x"20",
          6478 => x"72",
          6479 => x"20",
          6480 => x"30",
          6481 => x"00",
          6482 => x"20",
          6483 => x"53",
          6484 => x"6b",
          6485 => x"61",
          6486 => x"41",
          6487 => x"65",
          6488 => x"20",
          6489 => x"20",
          6490 => x"30",
          6491 => x"00",
          6492 => x"4d",
          6493 => x"3a",
          6494 => x"20",
          6495 => x"5a",
          6496 => x"49",
          6497 => x"20",
          6498 => x"20",
          6499 => x"20",
          6500 => x"20",
          6501 => x"20",
          6502 => x"30",
          6503 => x"00",
          6504 => x"20",
          6505 => x"53",
          6506 => x"65",
          6507 => x"6c",
          6508 => x"20",
          6509 => x"71",
          6510 => x"20",
          6511 => x"20",
          6512 => x"64",
          6513 => x"34",
          6514 => x"7a",
          6515 => x"20",
          6516 => x"53",
          6517 => x"4d",
          6518 => x"6f",
          6519 => x"46",
          6520 => x"20",
          6521 => x"20",
          6522 => x"20",
          6523 => x"64",
          6524 => x"34",
          6525 => x"7a",
          6526 => x"20",
          6527 => x"57",
          6528 => x"62",
          6529 => x"20",
          6530 => x"41",
          6531 => x"6c",
          6532 => x"20",
          6533 => x"71",
          6534 => x"64",
          6535 => x"34",
          6536 => x"7a",
          6537 => x"53",
          6538 => x"6c",
          6539 => x"4d",
          6540 => x"75",
          6541 => x"46",
          6542 => x"00",
          6543 => x"45",
          6544 => x"45",
          6545 => x"69",
          6546 => x"55",
          6547 => x"6f",
          6548 => x"53",
          6549 => x"22",
          6550 => x"3a",
          6551 => x"3e",
          6552 => x"7c",
          6553 => x"46",
          6554 => x"46",
          6555 => x"32",
          6556 => x"eb",
          6557 => x"53",
          6558 => x"35",
          6559 => x"4e",
          6560 => x"41",
          6561 => x"20",
          6562 => x"41",
          6563 => x"20",
          6564 => x"4e",
          6565 => x"41",
          6566 => x"20",
          6567 => x"41",
          6568 => x"20",
          6569 => x"00",
          6570 => x"00",
          6571 => x"00",
          6572 => x"00",
          6573 => x"80",
          6574 => x"8e",
          6575 => x"45",
          6576 => x"49",
          6577 => x"90",
          6578 => x"99",
          6579 => x"59",
          6580 => x"9c",
          6581 => x"41",
          6582 => x"a5",
          6583 => x"a8",
          6584 => x"ac",
          6585 => x"b0",
          6586 => x"b4",
          6587 => x"b8",
          6588 => x"bc",
          6589 => x"c0",
          6590 => x"c4",
          6591 => x"c8",
          6592 => x"cc",
          6593 => x"d0",
          6594 => x"d4",
          6595 => x"d8",
          6596 => x"dc",
          6597 => x"e0",
          6598 => x"e4",
          6599 => x"e8",
          6600 => x"ec",
          6601 => x"f0",
          6602 => x"f4",
          6603 => x"f8",
          6604 => x"fc",
          6605 => x"2b",
          6606 => x"3d",
          6607 => x"5c",
          6608 => x"3c",
          6609 => x"7f",
          6610 => x"00",
          6611 => x"00",
          6612 => x"01",
          6613 => x"00",
          6614 => x"00",
          6615 => x"00",
          6616 => x"00",
          6617 => x"00",
          6618 => x"64",
          6619 => x"74",
          6620 => x"64",
          6621 => x"74",
          6622 => x"66",
          6623 => x"74",
          6624 => x"66",
          6625 => x"64",
          6626 => x"66",
          6627 => x"63",
          6628 => x"6d",
          6629 => x"61",
          6630 => x"6d",
          6631 => x"70",
          6632 => x"6d",
          6633 => x"68",
          6634 => x"6d",
          6635 => x"6d",
          6636 => x"6d",
          6637 => x"68",
          6638 => x"68",
          6639 => x"68",
          6640 => x"68",
          6641 => x"63",
          6642 => x"00",
          6643 => x"6a",
          6644 => x"72",
          6645 => x"61",
          6646 => x"72",
          6647 => x"74",
          6648 => x"69",
          6649 => x"00",
          6650 => x"74",
          6651 => x"00",
          6652 => x"44",
          6653 => x"20",
          6654 => x"6f",
          6655 => x"49",
          6656 => x"72",
          6657 => x"20",
          6658 => x"6f",
          6659 => x"00",
          6660 => x"44",
          6661 => x"20",
          6662 => x"20",
          6663 => x"64",
          6664 => x"00",
          6665 => x"4e",
          6666 => x"69",
          6667 => x"66",
          6668 => x"64",
          6669 => x"4e",
          6670 => x"61",
          6671 => x"66",
          6672 => x"64",
          6673 => x"49",
          6674 => x"6c",
          6675 => x"66",
          6676 => x"6e",
          6677 => x"2e",
          6678 => x"41",
          6679 => x"73",
          6680 => x"65",
          6681 => x"64",
          6682 => x"46",
          6683 => x"20",
          6684 => x"65",
          6685 => x"20",
          6686 => x"73",
          6687 => x"0a",
          6688 => x"46",
          6689 => x"20",
          6690 => x"64",
          6691 => x"69",
          6692 => x"6c",
          6693 => x"0a",
          6694 => x"53",
          6695 => x"73",
          6696 => x"69",
          6697 => x"70",
          6698 => x"65",
          6699 => x"64",
          6700 => x"44",
          6701 => x"65",
          6702 => x"6d",
          6703 => x"20",
          6704 => x"69",
          6705 => x"6c",
          6706 => x"0a",
          6707 => x"44",
          6708 => x"20",
          6709 => x"20",
          6710 => x"62",
          6711 => x"2e",
          6712 => x"4e",
          6713 => x"6f",
          6714 => x"74",
          6715 => x"65",
          6716 => x"6c",
          6717 => x"73",
          6718 => x"20",
          6719 => x"6e",
          6720 => x"6e",
          6721 => x"73",
          6722 => x"00",
          6723 => x"46",
          6724 => x"61",
          6725 => x"62",
          6726 => x"65",
          6727 => x"00",
          6728 => x"54",
          6729 => x"6f",
          6730 => x"20",
          6731 => x"72",
          6732 => x"6f",
          6733 => x"61",
          6734 => x"6c",
          6735 => x"2e",
          6736 => x"46",
          6737 => x"20",
          6738 => x"6c",
          6739 => x"65",
          6740 => x"00",
          6741 => x"49",
          6742 => x"66",
          6743 => x"69",
          6744 => x"20",
          6745 => x"6f",
          6746 => x"0a",
          6747 => x"54",
          6748 => x"6d",
          6749 => x"20",
          6750 => x"6e",
          6751 => x"6c",
          6752 => x"0a",
          6753 => x"50",
          6754 => x"6d",
          6755 => x"72",
          6756 => x"6e",
          6757 => x"72",
          6758 => x"2e",
          6759 => x"53",
          6760 => x"65",
          6761 => x"0a",
          6762 => x"55",
          6763 => x"6f",
          6764 => x"65",
          6765 => x"72",
          6766 => x"0a",
          6767 => x"20",
          6768 => x"65",
          6769 => x"73",
          6770 => x"20",
          6771 => x"20",
          6772 => x"65",
          6773 => x"65",
          6774 => x"00",
          6775 => x"25",
          6776 => x"00",
          6777 => x"3a",
          6778 => x"25",
          6779 => x"00",
          6780 => x"20",
          6781 => x"20",
          6782 => x"00",
          6783 => x"25",
          6784 => x"00",
          6785 => x"20",
          6786 => x"20",
          6787 => x"7c",
          6788 => x"72",
          6789 => x"00",
          6790 => x"5a",
          6791 => x"41",
          6792 => x"0a",
          6793 => x"25",
          6794 => x"00",
          6795 => x"32",
          6796 => x"32",
          6797 => x"31",
          6798 => x"76",
          6799 => x"00",
          6800 => x"20",
          6801 => x"2c",
          6802 => x"76",
          6803 => x"32",
          6804 => x"25",
          6805 => x"73",
          6806 => x"0a",
          6807 => x"5a",
          6808 => x"41",
          6809 => x"74",
          6810 => x"75",
          6811 => x"48",
          6812 => x"6c",
          6813 => x"00",
          6814 => x"54",
          6815 => x"72",
          6816 => x"74",
          6817 => x"75",
          6818 => x"00",
          6819 => x"50",
          6820 => x"69",
          6821 => x"72",
          6822 => x"74",
          6823 => x"49",
          6824 => x"4c",
          6825 => x"20",
          6826 => x"65",
          6827 => x"70",
          6828 => x"49",
          6829 => x"4c",
          6830 => x"20",
          6831 => x"65",
          6832 => x"70",
          6833 => x"55",
          6834 => x"30",
          6835 => x"20",
          6836 => x"65",
          6837 => x"70",
          6838 => x"55",
          6839 => x"30",
          6840 => x"20",
          6841 => x"65",
          6842 => x"70",
          6843 => x"55",
          6844 => x"31",
          6845 => x"20",
          6846 => x"65",
          6847 => x"70",
          6848 => x"55",
          6849 => x"31",
          6850 => x"20",
          6851 => x"65",
          6852 => x"70",
          6853 => x"53",
          6854 => x"69",
          6855 => x"75",
          6856 => x"69",
          6857 => x"2e",
          6858 => x"00",
          6859 => x"45",
          6860 => x"6c",
          6861 => x"20",
          6862 => x"65",
          6863 => x"2e",
          6864 => x"61",
          6865 => x"65",
          6866 => x"2e",
          6867 => x"00",
          6868 => x"30",
          6869 => x"46",
          6870 => x"65",
          6871 => x"6f",
          6872 => x"69",
          6873 => x"6c",
          6874 => x"20",
          6875 => x"63",
          6876 => x"20",
          6877 => x"70",
          6878 => x"73",
          6879 => x"6e",
          6880 => x"6d",
          6881 => x"61",
          6882 => x"2e",
          6883 => x"2a",
          6884 => x"42",
          6885 => x"64",
          6886 => x"20",
          6887 => x"0a",
          6888 => x"49",
          6889 => x"69",
          6890 => x"73",
          6891 => x"0a",
          6892 => x"46",
          6893 => x"65",
          6894 => x"6f",
          6895 => x"69",
          6896 => x"6c",
          6897 => x"2e",
          6898 => x"72",
          6899 => x"64",
          6900 => x"25",
          6901 => x"43",
          6902 => x"72",
          6903 => x"2e",
          6904 => x"00",
          6905 => x"44",
          6906 => x"20",
          6907 => x"6f",
          6908 => x"00",
          6909 => x"0a",
          6910 => x"70",
          6911 => x"65",
          6912 => x"25",
          6913 => x"20",
          6914 => x"58",
          6915 => x"3f",
          6916 => x"00",
          6917 => x"25",
          6918 => x"20",
          6919 => x"58",
          6920 => x"25",
          6921 => x"20",
          6922 => x"58",
          6923 => x"53",
          6924 => x"63",
          6925 => x"67",
          6926 => x"00",
          6927 => x"25",
          6928 => x"78",
          6929 => x"30",
          6930 => x"0a",
          6931 => x"44",
          6932 => x"62",
          6933 => x"67",
          6934 => x"74",
          6935 => x"75",
          6936 => x"0a",
          6937 => x"45",
          6938 => x"6c",
          6939 => x"20",
          6940 => x"65",
          6941 => x"70",
          6942 => x"00",
          6943 => x"44",
          6944 => x"62",
          6945 => x"20",
          6946 => x"74",
          6947 => x"66",
          6948 => x"45",
          6949 => x"6c",
          6950 => x"20",
          6951 => x"74",
          6952 => x"66",
          6953 => x"45",
          6954 => x"75",
          6955 => x"67",
          6956 => x"64",
          6957 => x"20",
          6958 => x"78",
          6959 => x"2e",
          6960 => x"43",
          6961 => x"69",
          6962 => x"63",
          6963 => x"20",
          6964 => x"30",
          6965 => x"2e",
          6966 => x"00",
          6967 => x"43",
          6968 => x"20",
          6969 => x"75",
          6970 => x"64",
          6971 => x"64",
          6972 => x"25",
          6973 => x"0a",
          6974 => x"52",
          6975 => x"61",
          6976 => x"6e",
          6977 => x"70",
          6978 => x"63",
          6979 => x"6f",
          6980 => x"2e",
          6981 => x"43",
          6982 => x"20",
          6983 => x"6f",
          6984 => x"6e",
          6985 => x"2e",
          6986 => x"5a",
          6987 => x"62",
          6988 => x"25",
          6989 => x"25",
          6990 => x"73",
          6991 => x"00",
          6992 => x"25",
          6993 => x"25",
          6994 => x"73",
          6995 => x"25",
          6996 => x"25",
          6997 => x"42",
          6998 => x"63",
          6999 => x"61",
          7000 => x"0a",
          7001 => x"52",
          7002 => x"69",
          7003 => x"2e",
          7004 => x"45",
          7005 => x"6c",
          7006 => x"20",
          7007 => x"65",
          7008 => x"70",
          7009 => x"2e",
          7010 => x"00",
          7011 => x"00",
          7012 => x"00",
          7013 => x"00",
          7014 => x"00",
          7015 => x"00",
          7016 => x"00",
          7017 => x"00",
          7018 => x"00",
          7019 => x"01",
          7020 => x"01",
          7021 => x"00",
          7022 => x"00",
          7023 => x"00",
          7024 => x"00",
          7025 => x"05",
          7026 => x"05",
          7027 => x"05",
          7028 => x"00",
          7029 => x"01",
          7030 => x"01",
          7031 => x"01",
          7032 => x"01",
          7033 => x"00",
          7034 => x"01",
          7035 => x"00",
          7036 => x"00",
          7037 => x"01",
          7038 => x"00",
          7039 => x"00",
          7040 => x"00",
          7041 => x"01",
          7042 => x"00",
          7043 => x"00",
          7044 => x"00",
          7045 => x"01",
          7046 => x"00",
          7047 => x"00",
          7048 => x"00",
          7049 => x"01",
          7050 => x"00",
          7051 => x"00",
          7052 => x"00",
          7053 => x"01",
          7054 => x"00",
          7055 => x"00",
          7056 => x"00",
          7057 => x"01",
          7058 => x"00",
          7059 => x"00",
          7060 => x"00",
          7061 => x"01",
          7062 => x"00",
          7063 => x"00",
          7064 => x"00",
          7065 => x"01",
          7066 => x"00",
          7067 => x"00",
          7068 => x"00",
          7069 => x"01",
          7070 => x"00",
          7071 => x"00",
          7072 => x"00",
          7073 => x"01",
          7074 => x"00",
          7075 => x"00",
          7076 => x"00",
          7077 => x"01",
          7078 => x"00",
          7079 => x"00",
          7080 => x"00",
          7081 => x"01",
          7082 => x"00",
          7083 => x"00",
          7084 => x"00",
          7085 => x"01",
          7086 => x"00",
          7087 => x"00",
          7088 => x"00",
          7089 => x"01",
          7090 => x"00",
          7091 => x"00",
          7092 => x"00",
          7093 => x"01",
          7094 => x"00",
          7095 => x"00",
          7096 => x"00",
          7097 => x"01",
          7098 => x"00",
          7099 => x"00",
          7100 => x"00",
          7101 => x"01",
          7102 => x"00",
          7103 => x"00",
          7104 => x"00",
          7105 => x"01",
          7106 => x"00",
          7107 => x"00",
          7108 => x"00",
          7109 => x"01",
          7110 => x"00",
          7111 => x"00",
          7112 => x"00",
          7113 => x"01",
          7114 => x"00",
          7115 => x"00",
          7116 => x"00",
          7117 => x"01",
          7118 => x"00",
          7119 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
