-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.softZPU_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"b0",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"bd",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"ac",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"ab",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8f",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"90",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"91",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"92",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"d4",
           386 => x"87",
           387 => x"d4",
           388 => x"80",
           389 => x"b9",
           390 => x"ee",
           391 => x"d4",
           392 => x"80",
           393 => x"b9",
           394 => x"f3",
           395 => x"d4",
           396 => x"80",
           397 => x"b9",
           398 => x"e0",
           399 => x"d4",
           400 => x"80",
           401 => x"b9",
           402 => x"a3",
           403 => x"d4",
           404 => x"80",
           405 => x"b9",
           406 => x"f6",
           407 => x"d4",
           408 => x"80",
           409 => x"b9",
           410 => x"86",
           411 => x"d4",
           412 => x"80",
           413 => x"b9",
           414 => x"82",
           415 => x"d4",
           416 => x"80",
           417 => x"b9",
           418 => x"88",
           419 => x"d4",
           420 => x"80",
           421 => x"b9",
           422 => x"a8",
           423 => x"d4",
           424 => x"80",
           425 => x"b9",
           426 => x"d1",
           427 => x"d4",
           428 => x"80",
           429 => x"b9",
           430 => x"8a",
           431 => x"d4",
           432 => x"80",
           433 => x"b9",
           434 => x"d4",
           435 => x"b9",
           436 => x"c0",
           437 => x"84",
           438 => x"80",
           439 => x"84",
           440 => x"80",
           441 => x"04",
           442 => x"0c",
           443 => x"2d",
           444 => x"08",
           445 => x"90",
           446 => x"d4",
           447 => x"db",
           448 => x"d4",
           449 => x"80",
           450 => x"b9",
           451 => x"c9",
           452 => x"b9",
           453 => x"c0",
           454 => x"84",
           455 => x"82",
           456 => x"84",
           457 => x"80",
           458 => x"04",
           459 => x"0c",
           460 => x"2d",
           461 => x"08",
           462 => x"90",
           463 => x"d4",
           464 => x"c0",
           465 => x"d4",
           466 => x"80",
           467 => x"b9",
           468 => x"ed",
           469 => x"b9",
           470 => x"c0",
           471 => x"84",
           472 => x"82",
           473 => x"84",
           474 => x"80",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"90",
           480 => x"d4",
           481 => x"be",
           482 => x"d4",
           483 => x"80",
           484 => x"b9",
           485 => x"f3",
           486 => x"b9",
           487 => x"c0",
           488 => x"84",
           489 => x"82",
           490 => x"84",
           491 => x"80",
           492 => x"04",
           493 => x"0c",
           494 => x"2d",
           495 => x"08",
           496 => x"90",
           497 => x"d4",
           498 => x"e7",
           499 => x"d4",
           500 => x"80",
           501 => x"b9",
           502 => x"8b",
           503 => x"b9",
           504 => x"c0",
           505 => x"84",
           506 => x"82",
           507 => x"84",
           508 => x"80",
           509 => x"04",
           510 => x"0c",
           511 => x"2d",
           512 => x"08",
           513 => x"90",
           514 => x"d4",
           515 => x"88",
           516 => x"d4",
           517 => x"80",
           518 => x"b9",
           519 => x"e5",
           520 => x"b9",
           521 => x"c0",
           522 => x"84",
           523 => x"82",
           524 => x"84",
           525 => x"80",
           526 => x"04",
           527 => x"0c",
           528 => x"2d",
           529 => x"08",
           530 => x"90",
           531 => x"d4",
           532 => x"a7",
           533 => x"d4",
           534 => x"80",
           535 => x"b9",
           536 => x"96",
           537 => x"b9",
           538 => x"c0",
           539 => x"84",
           540 => x"83",
           541 => x"84",
           542 => x"80",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"90",
           548 => x"d4",
           549 => x"ff",
           550 => x"d4",
           551 => x"80",
           552 => x"b9",
           553 => x"a4",
           554 => x"b9",
           555 => x"c0",
           556 => x"84",
           557 => x"83",
           558 => x"84",
           559 => x"80",
           560 => x"04",
           561 => x"0c",
           562 => x"2d",
           563 => x"08",
           564 => x"90",
           565 => x"d4",
           566 => x"e3",
           567 => x"d4",
           568 => x"80",
           569 => x"b9",
           570 => x"f4",
           571 => x"b9",
           572 => x"c0",
           573 => x"84",
           574 => x"81",
           575 => x"84",
           576 => x"80",
           577 => x"04",
           578 => x"0c",
           579 => x"2d",
           580 => x"08",
           581 => x"90",
           582 => x"d4",
           583 => x"fa",
           584 => x"d4",
           585 => x"80",
           586 => x"b9",
           587 => x"d7",
           588 => x"b9",
           589 => x"c0",
           590 => x"84",
           591 => x"b1",
           592 => x"b9",
           593 => x"c0",
           594 => x"84",
           595 => x"81",
           596 => x"84",
           597 => x"80",
           598 => x"04",
           599 => x"0c",
           600 => x"2d",
           601 => x"08",
           602 => x"90",
           603 => x"d4",
           604 => x"bd",
           605 => x"d4",
           606 => x"80",
           607 => x"b9",
           608 => x"d5",
           609 => x"b9",
           610 => x"c0",
           611 => x"3c",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"00",
           621 => x"ff",
           622 => x"06",
           623 => x"83",
           624 => x"10",
           625 => x"fc",
           626 => x"51",
           627 => x"80",
           628 => x"ff",
           629 => x"06",
           630 => x"52",
           631 => x"0a",
           632 => x"38",
           633 => x"51",
           634 => x"c8",
           635 => x"b4",
           636 => x"80",
           637 => x"05",
           638 => x"0b",
           639 => x"04",
           640 => x"80",
           641 => x"00",
           642 => x"87",
           643 => x"84",
           644 => x"56",
           645 => x"84",
           646 => x"51",
           647 => x"86",
           648 => x"fa",
           649 => x"7a",
           650 => x"33",
           651 => x"06",
           652 => x"07",
           653 => x"57",
           654 => x"72",
           655 => x"06",
           656 => x"ff",
           657 => x"8a",
           658 => x"70",
           659 => x"2a",
           660 => x"56",
           661 => x"25",
           662 => x"80",
           663 => x"75",
           664 => x"3f",
           665 => x"08",
           666 => x"c8",
           667 => x"ae",
           668 => x"c8",
           669 => x"81",
           670 => x"ff",
           671 => x"32",
           672 => x"72",
           673 => x"51",
           674 => x"73",
           675 => x"38",
           676 => x"76",
           677 => x"b9",
           678 => x"3d",
           679 => x"0b",
           680 => x"0c",
           681 => x"04",
           682 => x"7d",
           683 => x"84",
           684 => x"34",
           685 => x"0a",
           686 => x"88",
           687 => x"52",
           688 => x"05",
           689 => x"73",
           690 => x"74",
           691 => x"0d",
           692 => x"0d",
           693 => x"05",
           694 => x"75",
           695 => x"85",
           696 => x"f1",
           697 => x"63",
           698 => x"5d",
           699 => x"1f",
           700 => x"33",
           701 => x"81",
           702 => x"55",
           703 => x"54",
           704 => x"09",
           705 => x"d2",
           706 => x"57",
           707 => x"80",
           708 => x"1c",
           709 => x"54",
           710 => x"2e",
           711 => x"d0",
           712 => x"89",
           713 => x"38",
           714 => x"70",
           715 => x"25",
           716 => x"78",
           717 => x"80",
           718 => x"7a",
           719 => x"81",
           720 => x"40",
           721 => x"2e",
           722 => x"82",
           723 => x"7b",
           724 => x"ff",
           725 => x"1d",
           726 => x"84",
           727 => x"91",
           728 => x"7a",
           729 => x"78",
           730 => x"79",
           731 => x"98",
           732 => x"2c",
           733 => x"80",
           734 => x"0a",
           735 => x"2c",
           736 => x"56",
           737 => x"24",
           738 => x"73",
           739 => x"72",
           740 => x"78",
           741 => x"58",
           742 => x"38",
           743 => x"76",
           744 => x"81",
           745 => x"81",
           746 => x"5a",
           747 => x"33",
           748 => x"fe",
           749 => x"9e",
           750 => x"76",
           751 => x"3f",
           752 => x"76",
           753 => x"ff",
           754 => x"83",
           755 => x"06",
           756 => x"8a",
           757 => x"74",
           758 => x"7e",
           759 => x"17",
           760 => x"d8",
           761 => x"72",
           762 => x"ca",
           763 => x"73",
           764 => x"e0",
           765 => x"80",
           766 => x"eb",
           767 => x"76",
           768 => x"3f",
           769 => x"58",
           770 => x"86",
           771 => x"39",
           772 => x"fe",
           773 => x"5a",
           774 => x"05",
           775 => x"83",
           776 => x"5e",
           777 => x"84",
           778 => x"79",
           779 => x"93",
           780 => x"b9",
           781 => x"ff",
           782 => x"c8",
           783 => x"05",
           784 => x"89",
           785 => x"84",
           786 => x"b0",
           787 => x"7e",
           788 => x"40",
           789 => x"75",
           790 => x"3f",
           791 => x"08",
           792 => x"c8",
           793 => x"7d",
           794 => x"31",
           795 => x"b2",
           796 => x"7e",
           797 => x"38",
           798 => x"80",
           799 => x"80",
           800 => x"2c",
           801 => x"86",
           802 => x"06",
           803 => x"80",
           804 => x"77",
           805 => x"29",
           806 => x"05",
           807 => x"2e",
           808 => x"84",
           809 => x"fc",
           810 => x"53",
           811 => x"58",
           812 => x"70",
           813 => x"55",
           814 => x"9e",
           815 => x"2c",
           816 => x"06",
           817 => x"73",
           818 => x"38",
           819 => x"f7",
           820 => x"2a",
           821 => x"41",
           822 => x"81",
           823 => x"80",
           824 => x"38",
           825 => x"90",
           826 => x"2c",
           827 => x"06",
           828 => x"73",
           829 => x"96",
           830 => x"2a",
           831 => x"73",
           832 => x"7a",
           833 => x"06",
           834 => x"98",
           835 => x"2a",
           836 => x"73",
           837 => x"7e",
           838 => x"73",
           839 => x"7a",
           840 => x"06",
           841 => x"2e",
           842 => x"78",
           843 => x"29",
           844 => x"05",
           845 => x"5a",
           846 => x"74",
           847 => x"7c",
           848 => x"88",
           849 => x"78",
           850 => x"29",
           851 => x"05",
           852 => x"5a",
           853 => x"80",
           854 => x"74",
           855 => x"72",
           856 => x"38",
           857 => x"80",
           858 => x"ff",
           859 => x"98",
           860 => x"55",
           861 => x"9d",
           862 => x"b0",
           863 => x"3f",
           864 => x"80",
           865 => x"ff",
           866 => x"98",
           867 => x"55",
           868 => x"e5",
           869 => x"2a",
           870 => x"5c",
           871 => x"2e",
           872 => x"76",
           873 => x"84",
           874 => x"80",
           875 => x"ca",
           876 => x"d3",
           877 => x"38",
           878 => x"d8",
           879 => x"7c",
           880 => x"70",
           881 => x"87",
           882 => x"84",
           883 => x"09",
           884 => x"38",
           885 => x"5b",
           886 => x"fc",
           887 => x"78",
           888 => x"29",
           889 => x"05",
           890 => x"5a",
           891 => x"75",
           892 => x"38",
           893 => x"51",
           894 => x"e2",
           895 => x"07",
           896 => x"07",
           897 => x"5b",
           898 => x"38",
           899 => x"7a",
           900 => x"5b",
           901 => x"90",
           902 => x"05",
           903 => x"83",
           904 => x"5f",
           905 => x"5a",
           906 => x"7f",
           907 => x"77",
           908 => x"06",
           909 => x"70",
           910 => x"07",
           911 => x"80",
           912 => x"80",
           913 => x"2c",
           914 => x"56",
           915 => x"7a",
           916 => x"81",
           917 => x"7a",
           918 => x"77",
           919 => x"80",
           920 => x"80",
           921 => x"2c",
           922 => x"80",
           923 => x"b3",
           924 => x"a0",
           925 => x"3f",
           926 => x"1a",
           927 => x"ff",
           928 => x"79",
           929 => x"2e",
           930 => x"7c",
           931 => x"81",
           932 => x"51",
           933 => x"e2",
           934 => x"70",
           935 => x"06",
           936 => x"83",
           937 => x"fe",
           938 => x"52",
           939 => x"05",
           940 => x"85",
           941 => x"39",
           942 => x"06",
           943 => x"07",
           944 => x"80",
           945 => x"80",
           946 => x"2c",
           947 => x"80",
           948 => x"2a",
           949 => x"5d",
           950 => x"fd",
           951 => x"fb",
           952 => x"84",
           953 => x"70",
           954 => x"56",
           955 => x"82",
           956 => x"83",
           957 => x"5b",
           958 => x"5e",
           959 => x"7a",
           960 => x"33",
           961 => x"f8",
           962 => x"ca",
           963 => x"07",
           964 => x"33",
           965 => x"f7",
           966 => x"ba",
           967 => x"84",
           968 => x"77",
           969 => x"58",
           970 => x"82",
           971 => x"51",
           972 => x"84",
           973 => x"83",
           974 => x"78",
           975 => x"2b",
           976 => x"90",
           977 => x"87",
           978 => x"c0",
           979 => x"58",
           980 => x"be",
           981 => x"39",
           982 => x"05",
           983 => x"81",
           984 => x"41",
           985 => x"cf",
           986 => x"87",
           987 => x"b9",
           988 => x"ff",
           989 => x"71",
           990 => x"54",
           991 => x"7a",
           992 => x"7c",
           993 => x"76",
           994 => x"f7",
           995 => x"78",
           996 => x"29",
           997 => x"05",
           998 => x"5a",
           999 => x"74",
          1000 => x"38",
          1001 => x"51",
          1002 => x"e2",
          1003 => x"b0",
          1004 => x"3f",
          1005 => x"09",
          1006 => x"e3",
          1007 => x"76",
          1008 => x"3f",
          1009 => x"81",
          1010 => x"80",
          1011 => x"38",
          1012 => x"75",
          1013 => x"71",
          1014 => x"70",
          1015 => x"83",
          1016 => x"5a",
          1017 => x"fa",
          1018 => x"a2",
          1019 => x"ad",
          1020 => x"3f",
          1021 => x"54",
          1022 => x"fa",
          1023 => x"ad",
          1024 => x"75",
          1025 => x"82",
          1026 => x"81",
          1027 => x"80",
          1028 => x"38",
          1029 => x"78",
          1030 => x"2b",
          1031 => x"5a",
          1032 => x"39",
          1033 => x"51",
          1034 => x"c8",
          1035 => x"a0",
          1036 => x"3f",
          1037 => x"78",
          1038 => x"88",
          1039 => x"b9",
          1040 => x"ff",
          1041 => x"71",
          1042 => x"54",
          1043 => x"39",
          1044 => x"7e",
          1045 => x"ff",
          1046 => x"57",
          1047 => x"39",
          1048 => x"84",
          1049 => x"53",
          1050 => x"51",
          1051 => x"84",
          1052 => x"fa",
          1053 => x"55",
          1054 => x"d5",
          1055 => x"11",
          1056 => x"2a",
          1057 => x"81",
          1058 => x"58",
          1059 => x"56",
          1060 => x"09",
          1061 => x"d5",
          1062 => x"81",
          1063 => x"53",
          1064 => x"b0",
          1065 => x"ac",
          1066 => x"51",
          1067 => x"53",
          1068 => x"b9",
          1069 => x"2e",
          1070 => x"57",
          1071 => x"05",
          1072 => x"72",
          1073 => x"38",
          1074 => x"08",
          1075 => x"84",
          1076 => x"54",
          1077 => x"08",
          1078 => x"90",
          1079 => x"74",
          1080 => x"c8",
          1081 => x"83",
          1082 => x"76",
          1083 => x"b9",
          1084 => x"3d",
          1085 => x"3d",
          1086 => x"56",
          1087 => x"85",
          1088 => x"81",
          1089 => x"70",
          1090 => x"55",
          1091 => x"56",
          1092 => x"09",
          1093 => x"38",
          1094 => x"05",
          1095 => x"72",
          1096 => x"81",
          1097 => x"76",
          1098 => x"b9",
          1099 => x"3d",
          1100 => x"70",
          1101 => x"33",
          1102 => x"2e",
          1103 => x"52",
          1104 => x"15",
          1105 => x"2d",
          1106 => x"08",
          1107 => x"38",
          1108 => x"81",
          1109 => x"54",
          1110 => x"38",
          1111 => x"3d",
          1112 => x"ac",
          1113 => x"51",
          1114 => x"3d",
          1115 => x"3d",
          1116 => x"85",
          1117 => x"81",
          1118 => x"81",
          1119 => x"56",
          1120 => x"72",
          1121 => x"82",
          1122 => x"54",
          1123 => x"ac",
          1124 => x"08",
          1125 => x"16",
          1126 => x"38",
          1127 => x"76",
          1128 => x"08",
          1129 => x"0c",
          1130 => x"53",
          1131 => x"16",
          1132 => x"75",
          1133 => x"0c",
          1134 => x"04",
          1135 => x"81",
          1136 => x"90",
          1137 => x"73",
          1138 => x"84",
          1139 => x"e3",
          1140 => x"08",
          1141 => x"16",
          1142 => x"d7",
          1143 => x"0d",
          1144 => x"33",
          1145 => x"06",
          1146 => x"81",
          1147 => x"56",
          1148 => x"71",
          1149 => x"86",
          1150 => x"52",
          1151 => x"72",
          1152 => x"06",
          1153 => x"2e",
          1154 => x"75",
          1155 => x"53",
          1156 => x"2e",
          1157 => x"81",
          1158 => x"8c",
          1159 => x"05",
          1160 => x"71",
          1161 => x"54",
          1162 => x"c8",
          1163 => x"0d",
          1164 => x"bf",
          1165 => x"85",
          1166 => x"16",
          1167 => x"8c",
          1168 => x"16",
          1169 => x"c8",
          1170 => x"0d",
          1171 => x"94",
          1172 => x"74",
          1173 => x"c8",
          1174 => x"b9",
          1175 => x"25",
          1176 => x"85",
          1177 => x"90",
          1178 => x"84",
          1179 => x"ff",
          1180 => x"71",
          1181 => x"72",
          1182 => x"ff",
          1183 => x"b9",
          1184 => x"3d",
          1185 => x"a0",
          1186 => x"85",
          1187 => x"54",
          1188 => x"3d",
          1189 => x"71",
          1190 => x"71",
          1191 => x"53",
          1192 => x"f7",
          1193 => x"52",
          1194 => x"05",
          1195 => x"70",
          1196 => x"05",
          1197 => x"f0",
          1198 => x"b9",
          1199 => x"3d",
          1200 => x"3d",
          1201 => x"71",
          1202 => x"52",
          1203 => x"2e",
          1204 => x"72",
          1205 => x"70",
          1206 => x"38",
          1207 => x"05",
          1208 => x"70",
          1209 => x"34",
          1210 => x"70",
          1211 => x"84",
          1212 => x"86",
          1213 => x"70",
          1214 => x"75",
          1215 => x"70",
          1216 => x"53",
          1217 => x"13",
          1218 => x"33",
          1219 => x"11",
          1220 => x"2e",
          1221 => x"13",
          1222 => x"53",
          1223 => x"34",
          1224 => x"70",
          1225 => x"39",
          1226 => x"74",
          1227 => x"71",
          1228 => x"53",
          1229 => x"f7",
          1230 => x"70",
          1231 => x"b9",
          1232 => x"84",
          1233 => x"fd",
          1234 => x"77",
          1235 => x"54",
          1236 => x"05",
          1237 => x"70",
          1238 => x"05",
          1239 => x"f0",
          1240 => x"b9",
          1241 => x"3d",
          1242 => x"3d",
          1243 => x"71",
          1244 => x"52",
          1245 => x"2e",
          1246 => x"70",
          1247 => x"33",
          1248 => x"05",
          1249 => x"11",
          1250 => x"38",
          1251 => x"c8",
          1252 => x"0d",
          1253 => x"0d",
          1254 => x"55",
          1255 => x"80",
          1256 => x"73",
          1257 => x"81",
          1258 => x"52",
          1259 => x"2e",
          1260 => x"9a",
          1261 => x"54",
          1262 => x"b7",
          1263 => x"53",
          1264 => x"80",
          1265 => x"b9",
          1266 => x"3d",
          1267 => x"80",
          1268 => x"73",
          1269 => x"51",
          1270 => x"e9",
          1271 => x"33",
          1272 => x"71",
          1273 => x"38",
          1274 => x"84",
          1275 => x"86",
          1276 => x"71",
          1277 => x"0c",
          1278 => x"04",
          1279 => x"77",
          1280 => x"52",
          1281 => x"3f",
          1282 => x"08",
          1283 => x"08",
          1284 => x"55",
          1285 => x"3f",
          1286 => x"08",
          1287 => x"c8",
          1288 => x"9b",
          1289 => x"c8",
          1290 => x"80",
          1291 => x"53",
          1292 => x"b9",
          1293 => x"fe",
          1294 => x"b9",
          1295 => x"73",
          1296 => x"0c",
          1297 => x"04",
          1298 => x"75",
          1299 => x"54",
          1300 => x"71",
          1301 => x"38",
          1302 => x"05",
          1303 => x"70",
          1304 => x"38",
          1305 => x"71",
          1306 => x"81",
          1307 => x"ff",
          1308 => x"31",
          1309 => x"84",
          1310 => x"85",
          1311 => x"fd",
          1312 => x"77",
          1313 => x"53",
          1314 => x"80",
          1315 => x"72",
          1316 => x"05",
          1317 => x"11",
          1318 => x"38",
          1319 => x"c8",
          1320 => x"0d",
          1321 => x"0d",
          1322 => x"54",
          1323 => x"80",
          1324 => x"76",
          1325 => x"3f",
          1326 => x"08",
          1327 => x"53",
          1328 => x"8d",
          1329 => x"80",
          1330 => x"84",
          1331 => x"31",
          1332 => x"72",
          1333 => x"cb",
          1334 => x"72",
          1335 => x"c3",
          1336 => x"74",
          1337 => x"72",
          1338 => x"2b",
          1339 => x"55",
          1340 => x"76",
          1341 => x"72",
          1342 => x"2a",
          1343 => x"77",
          1344 => x"31",
          1345 => x"2c",
          1346 => x"7b",
          1347 => x"71",
          1348 => x"5c",
          1349 => x"55",
          1350 => x"74",
          1351 => x"10",
          1352 => x"71",
          1353 => x"0c",
          1354 => x"04",
          1355 => x"76",
          1356 => x"80",
          1357 => x"70",
          1358 => x"25",
          1359 => x"90",
          1360 => x"71",
          1361 => x"fe",
          1362 => x"30",
          1363 => x"83",
          1364 => x"31",
          1365 => x"70",
          1366 => x"70",
          1367 => x"25",
          1368 => x"71",
          1369 => x"2a",
          1370 => x"1b",
          1371 => x"06",
          1372 => x"80",
          1373 => x"71",
          1374 => x"2a",
          1375 => x"81",
          1376 => x"06",
          1377 => x"74",
          1378 => x"19",
          1379 => x"c8",
          1380 => x"54",
          1381 => x"56",
          1382 => x"55",
          1383 => x"56",
          1384 => x"58",
          1385 => x"86",
          1386 => x"fd",
          1387 => x"77",
          1388 => x"53",
          1389 => x"94",
          1390 => x"c8",
          1391 => x"74",
          1392 => x"b9",
          1393 => x"85",
          1394 => x"fa",
          1395 => x"7a",
          1396 => x"53",
          1397 => x"8b",
          1398 => x"fe",
          1399 => x"b9",
          1400 => x"e0",
          1401 => x"80",
          1402 => x"73",
          1403 => x"3f",
          1404 => x"c8",
          1405 => x"73",
          1406 => x"26",
          1407 => x"80",
          1408 => x"2e",
          1409 => x"12",
          1410 => x"a0",
          1411 => x"71",
          1412 => x"54",
          1413 => x"74",
          1414 => x"38",
          1415 => x"9f",
          1416 => x"10",
          1417 => x"72",
          1418 => x"9f",
          1419 => x"06",
          1420 => x"75",
          1421 => x"1c",
          1422 => x"52",
          1423 => x"53",
          1424 => x"72",
          1425 => x"0c",
          1426 => x"04",
          1427 => x"78",
          1428 => x"9f",
          1429 => x"2c",
          1430 => x"9f",
          1431 => x"73",
          1432 => x"74",
          1433 => x"75",
          1434 => x"56",
          1435 => x"fc",
          1436 => x"b9",
          1437 => x"32",
          1438 => x"b9",
          1439 => x"3d",
          1440 => x"3d",
          1441 => x"5b",
          1442 => x"7b",
          1443 => x"70",
          1444 => x"59",
          1445 => x"09",
          1446 => x"38",
          1447 => x"78",
          1448 => x"55",
          1449 => x"2e",
          1450 => x"ad",
          1451 => x"38",
          1452 => x"81",
          1453 => x"14",
          1454 => x"77",
          1455 => x"db",
          1456 => x"80",
          1457 => x"27",
          1458 => x"80",
          1459 => x"89",
          1460 => x"70",
          1461 => x"55",
          1462 => x"70",
          1463 => x"51",
          1464 => x"27",
          1465 => x"13",
          1466 => x"06",
          1467 => x"73",
          1468 => x"38",
          1469 => x"81",
          1470 => x"76",
          1471 => x"16",
          1472 => x"70",
          1473 => x"56",
          1474 => x"ff",
          1475 => x"80",
          1476 => x"75",
          1477 => x"7a",
          1478 => x"75",
          1479 => x"0c",
          1480 => x"04",
          1481 => x"70",
          1482 => x"33",
          1483 => x"73",
          1484 => x"81",
          1485 => x"38",
          1486 => x"78",
          1487 => x"55",
          1488 => x"e2",
          1489 => x"90",
          1490 => x"f8",
          1491 => x"81",
          1492 => x"27",
          1493 => x"14",
          1494 => x"88",
          1495 => x"27",
          1496 => x"75",
          1497 => x"0c",
          1498 => x"04",
          1499 => x"15",
          1500 => x"70",
          1501 => x"80",
          1502 => x"39",
          1503 => x"b9",
          1504 => x"3d",
          1505 => x"3d",
          1506 => x"5b",
          1507 => x"7b",
          1508 => x"70",
          1509 => x"59",
          1510 => x"09",
          1511 => x"38",
          1512 => x"78",
          1513 => x"55",
          1514 => x"2e",
          1515 => x"ad",
          1516 => x"38",
          1517 => x"81",
          1518 => x"14",
          1519 => x"77",
          1520 => x"db",
          1521 => x"80",
          1522 => x"27",
          1523 => x"80",
          1524 => x"89",
          1525 => x"70",
          1526 => x"55",
          1527 => x"70",
          1528 => x"51",
          1529 => x"27",
          1530 => x"13",
          1531 => x"06",
          1532 => x"73",
          1533 => x"38",
          1534 => x"81",
          1535 => x"76",
          1536 => x"16",
          1537 => x"70",
          1538 => x"56",
          1539 => x"ff",
          1540 => x"80",
          1541 => x"75",
          1542 => x"7a",
          1543 => x"75",
          1544 => x"0c",
          1545 => x"04",
          1546 => x"70",
          1547 => x"33",
          1548 => x"73",
          1549 => x"81",
          1550 => x"38",
          1551 => x"78",
          1552 => x"55",
          1553 => x"e2",
          1554 => x"90",
          1555 => x"f8",
          1556 => x"81",
          1557 => x"27",
          1558 => x"14",
          1559 => x"88",
          1560 => x"27",
          1561 => x"75",
          1562 => x"0c",
          1563 => x"04",
          1564 => x"15",
          1565 => x"70",
          1566 => x"80",
          1567 => x"39",
          1568 => x"b9",
          1569 => x"3d",
          1570 => x"d6",
          1571 => x"b9",
          1572 => x"ff",
          1573 => x"c8",
          1574 => x"3d",
          1575 => x"71",
          1576 => x"38",
          1577 => x"83",
          1578 => x"52",
          1579 => x"83",
          1580 => x"ef",
          1581 => x"3d",
          1582 => x"ce",
          1583 => x"b3",
          1584 => x"0d",
          1585 => x"c4",
          1586 => x"3f",
          1587 => x"04",
          1588 => x"51",
          1589 => x"83",
          1590 => x"83",
          1591 => x"ef",
          1592 => x"3d",
          1593 => x"cf",
          1594 => x"87",
          1595 => x"0d",
          1596 => x"a4",
          1597 => x"3f",
          1598 => x"04",
          1599 => x"51",
          1600 => x"83",
          1601 => x"83",
          1602 => x"ee",
          1603 => x"3d",
          1604 => x"cf",
          1605 => x"db",
          1606 => x"0d",
          1607 => x"8c",
          1608 => x"3f",
          1609 => x"04",
          1610 => x"51",
          1611 => x"83",
          1612 => x"83",
          1613 => x"ee",
          1614 => x"3d",
          1615 => x"d0",
          1616 => x"af",
          1617 => x"0d",
          1618 => x"e4",
          1619 => x"3f",
          1620 => x"04",
          1621 => x"51",
          1622 => x"83",
          1623 => x"83",
          1624 => x"ee",
          1625 => x"3d",
          1626 => x"d1",
          1627 => x"83",
          1628 => x"0d",
          1629 => x"a8",
          1630 => x"3f",
          1631 => x"04",
          1632 => x"51",
          1633 => x"83",
          1634 => x"83",
          1635 => x"ed",
          1636 => x"3d",
          1637 => x"3d",
          1638 => x"84",
          1639 => x"05",
          1640 => x"80",
          1641 => x"70",
          1642 => x"25",
          1643 => x"59",
          1644 => x"87",
          1645 => x"38",
          1646 => x"77",
          1647 => x"ff",
          1648 => x"93",
          1649 => x"e2",
          1650 => x"77",
          1651 => x"70",
          1652 => x"95",
          1653 => x"b9",
          1654 => x"84",
          1655 => x"80",
          1656 => x"38",
          1657 => x"af",
          1658 => x"30",
          1659 => x"80",
          1660 => x"70",
          1661 => x"06",
          1662 => x"58",
          1663 => x"aa",
          1664 => x"98",
          1665 => x"74",
          1666 => x"80",
          1667 => x"52",
          1668 => x"29",
          1669 => x"3f",
          1670 => x"08",
          1671 => x"f4",
          1672 => x"83",
          1673 => x"df",
          1674 => x"84",
          1675 => x"96",
          1676 => x"84",
          1677 => x"87",
          1678 => x"0c",
          1679 => x"08",
          1680 => x"d4",
          1681 => x"80",
          1682 => x"77",
          1683 => x"ce",
          1684 => x"c8",
          1685 => x"b9",
          1686 => x"88",
          1687 => x"74",
          1688 => x"80",
          1689 => x"75",
          1690 => x"d5",
          1691 => x"52",
          1692 => x"b1",
          1693 => x"c8",
          1694 => x"51",
          1695 => x"84",
          1696 => x"54",
          1697 => x"53",
          1698 => x"d1",
          1699 => x"f8",
          1700 => x"39",
          1701 => x"7c",
          1702 => x"b7",
          1703 => x"59",
          1704 => x"53",
          1705 => x"51",
          1706 => x"84",
          1707 => x"8b",
          1708 => x"2e",
          1709 => x"81",
          1710 => x"77",
          1711 => x"0c",
          1712 => x"04",
          1713 => x"d5",
          1714 => x"55",
          1715 => x"b9",
          1716 => x"52",
          1717 => x"2d",
          1718 => x"08",
          1719 => x"0c",
          1720 => x"04",
          1721 => x"7f",
          1722 => x"8c",
          1723 => x"05",
          1724 => x"15",
          1725 => x"5c",
          1726 => x"5e",
          1727 => x"83",
          1728 => x"52",
          1729 => x"51",
          1730 => x"83",
          1731 => x"dd",
          1732 => x"54",
          1733 => x"b2",
          1734 => x"2e",
          1735 => x"7c",
          1736 => x"a8",
          1737 => x"53",
          1738 => x"81",
          1739 => x"33",
          1740 => x"88",
          1741 => x"3f",
          1742 => x"d5",
          1743 => x"54",
          1744 => x"aa",
          1745 => x"26",
          1746 => x"d2",
          1747 => x"b8",
          1748 => x"75",
          1749 => x"c0",
          1750 => x"70",
          1751 => x"80",
          1752 => x"27",
          1753 => x"55",
          1754 => x"74",
          1755 => x"81",
          1756 => x"06",
          1757 => x"06",
          1758 => x"80",
          1759 => x"80",
          1760 => x"81",
          1761 => x"d5",
          1762 => x"a0",
          1763 => x"3f",
          1764 => x"78",
          1765 => x"38",
          1766 => x"51",
          1767 => x"78",
          1768 => x"5c",
          1769 => x"9d",
          1770 => x"b9",
          1771 => x"2b",
          1772 => x"58",
          1773 => x"2e",
          1774 => x"76",
          1775 => x"c3",
          1776 => x"57",
          1777 => x"fe",
          1778 => x"0b",
          1779 => x"0c",
          1780 => x"04",
          1781 => x"51",
          1782 => x"81",
          1783 => x"ac",
          1784 => x"a0",
          1785 => x"3f",
          1786 => x"fe",
          1787 => x"da",
          1788 => x"a8",
          1789 => x"3f",
          1790 => x"d5",
          1791 => x"54",
          1792 => x"ea",
          1793 => x"27",
          1794 => x"73",
          1795 => x"7a",
          1796 => x"72",
          1797 => x"d2",
          1798 => x"ec",
          1799 => x"84",
          1800 => x"53",
          1801 => x"ea",
          1802 => x"74",
          1803 => x"fe",
          1804 => x"d2",
          1805 => x"d0",
          1806 => x"84",
          1807 => x"53",
          1808 => x"ea",
          1809 => x"79",
          1810 => x"38",
          1811 => x"72",
          1812 => x"38",
          1813 => x"83",
          1814 => x"db",
          1815 => x"14",
          1816 => x"08",
          1817 => x"51",
          1818 => x"78",
          1819 => x"38",
          1820 => x"84",
          1821 => x"52",
          1822 => x"f2",
          1823 => x"56",
          1824 => x"80",
          1825 => x"84",
          1826 => x"81",
          1827 => x"88",
          1828 => x"2e",
          1829 => x"a0",
          1830 => x"d0",
          1831 => x"06",
          1832 => x"90",
          1833 => x"39",
          1834 => x"c0",
          1835 => x"c8",
          1836 => x"70",
          1837 => x"a0",
          1838 => x"72",
          1839 => x"30",
          1840 => x"73",
          1841 => x"51",
          1842 => x"57",
          1843 => x"80",
          1844 => x"38",
          1845 => x"94",
          1846 => x"c8",
          1847 => x"70",
          1848 => x"a0",
          1849 => x"72",
          1850 => x"30",
          1851 => x"73",
          1852 => x"51",
          1853 => x"57",
          1854 => x"73",
          1855 => x"38",
          1856 => x"80",
          1857 => x"c8",
          1858 => x"0d",
          1859 => x"0d",
          1860 => x"80",
          1861 => x"d7",
          1862 => x"9d",
          1863 => x"d3",
          1864 => x"99",
          1865 => x"9c",
          1866 => x"81",
          1867 => x"06",
          1868 => x"82",
          1869 => x"82",
          1870 => x"06",
          1871 => x"82",
          1872 => x"83",
          1873 => x"06",
          1874 => x"81",
          1875 => x"84",
          1876 => x"06",
          1877 => x"81",
          1878 => x"85",
          1879 => x"06",
          1880 => x"80",
          1881 => x"86",
          1882 => x"06",
          1883 => x"80",
          1884 => x"87",
          1885 => x"06",
          1886 => x"a9",
          1887 => x"2a",
          1888 => x"72",
          1889 => x"ef",
          1890 => x"0d",
          1891 => x"9c",
          1892 => x"d3",
          1893 => x"a5",
          1894 => x"9c",
          1895 => x"d7",
          1896 => x"0d",
          1897 => x"9b",
          1898 => x"d3",
          1899 => x"8d",
          1900 => x"9b",
          1901 => x"88",
          1902 => x"53",
          1903 => x"c6",
          1904 => x"81",
          1905 => x"3f",
          1906 => x"51",
          1907 => x"80",
          1908 => x"3f",
          1909 => x"70",
          1910 => x"52",
          1911 => x"ff",
          1912 => x"39",
          1913 => x"bd",
          1914 => x"94",
          1915 => x"3f",
          1916 => x"b1",
          1917 => x"2a",
          1918 => x"51",
          1919 => x"2e",
          1920 => x"ff",
          1921 => x"51",
          1922 => x"83",
          1923 => x"9b",
          1924 => x"51",
          1925 => x"72",
          1926 => x"81",
          1927 => x"71",
          1928 => x"c2",
          1929 => x"39",
          1930 => x"f9",
          1931 => x"bc",
          1932 => x"3f",
          1933 => x"ed",
          1934 => x"2a",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"ff",
          1938 => x"51",
          1939 => x"83",
          1940 => x"9a",
          1941 => x"51",
          1942 => x"72",
          1943 => x"81",
          1944 => x"71",
          1945 => x"e6",
          1946 => x"39",
          1947 => x"b5",
          1948 => x"e0",
          1949 => x"3f",
          1950 => x"a9",
          1951 => x"2a",
          1952 => x"51",
          1953 => x"2e",
          1954 => x"ff",
          1955 => x"3d",
          1956 => x"41",
          1957 => x"84",
          1958 => x"42",
          1959 => x"51",
          1960 => x"3f",
          1961 => x"08",
          1962 => x"9b",
          1963 => x"78",
          1964 => x"b1",
          1965 => x"b4",
          1966 => x"3f",
          1967 => x"83",
          1968 => x"d6",
          1969 => x"48",
          1970 => x"80",
          1971 => x"eb",
          1972 => x"0b",
          1973 => x"33",
          1974 => x"06",
          1975 => x"80",
          1976 => x"38",
          1977 => x"83",
          1978 => x"81",
          1979 => x"7d",
          1980 => x"c1",
          1981 => x"5a",
          1982 => x"2e",
          1983 => x"79",
          1984 => x"a0",
          1985 => x"06",
          1986 => x"1a",
          1987 => x"5a",
          1988 => x"f6",
          1989 => x"7b",
          1990 => x"38",
          1991 => x"83",
          1992 => x"70",
          1993 => x"e7",
          1994 => x"b9",
          1995 => x"b9",
          1996 => x"7a",
          1997 => x"52",
          1998 => x"3f",
          1999 => x"08",
          2000 => x"1b",
          2001 => x"81",
          2002 => x"38",
          2003 => x"81",
          2004 => x"5b",
          2005 => x"c4",
          2006 => x"33",
          2007 => x"2e",
          2008 => x"80",
          2009 => x"51",
          2010 => x"84",
          2011 => x"5e",
          2012 => x"08",
          2013 => x"c9",
          2014 => x"c8",
          2015 => x"3d",
          2016 => x"51",
          2017 => x"84",
          2018 => x"60",
          2019 => x"5c",
          2020 => x"81",
          2021 => x"b9",
          2022 => x"e7",
          2023 => x"b9",
          2024 => x"26",
          2025 => x"81",
          2026 => x"5e",
          2027 => x"2e",
          2028 => x"7a",
          2029 => x"e2",
          2030 => x"2e",
          2031 => x"7b",
          2032 => x"83",
          2033 => x"7c",
          2034 => x"3f",
          2035 => x"58",
          2036 => x"57",
          2037 => x"55",
          2038 => x"80",
          2039 => x"80",
          2040 => x"51",
          2041 => x"84",
          2042 => x"84",
          2043 => x"09",
          2044 => x"72",
          2045 => x"51",
          2046 => x"80",
          2047 => x"26",
          2048 => x"5a",
          2049 => x"59",
          2050 => x"8d",
          2051 => x"70",
          2052 => x"5c",
          2053 => x"95",
          2054 => x"32",
          2055 => x"07",
          2056 => x"ee",
          2057 => x"2e",
          2058 => x"7d",
          2059 => x"e1",
          2060 => x"ec",
          2061 => x"3f",
          2062 => x"f8",
          2063 => x"7e",
          2064 => x"3f",
          2065 => x"ee",
          2066 => x"81",
          2067 => x"59",
          2068 => x"38",
          2069 => x"d5",
          2070 => x"d0",
          2071 => x"88",
          2072 => x"b9",
          2073 => x"c5",
          2074 => x"0b",
          2075 => x"bc",
          2076 => x"d8",
          2077 => x"52",
          2078 => x"f6",
          2079 => x"b9",
          2080 => x"2e",
          2081 => x"b9",
          2082 => x"df",
          2083 => x"0b",
          2084 => x"33",
          2085 => x"06",
          2086 => x"82",
          2087 => x"06",
          2088 => x"91",
          2089 => x"d8",
          2090 => x"d4",
          2091 => x"0b",
          2092 => x"bc",
          2093 => x"a8",
          2094 => x"52",
          2095 => x"d4",
          2096 => x"5a",
          2097 => x"b7",
          2098 => x"7c",
          2099 => x"85",
          2100 => x"78",
          2101 => x"fd",
          2102 => x"10",
          2103 => x"d4",
          2104 => x"08",
          2105 => x"83",
          2106 => x"7e",
          2107 => x"3f",
          2108 => x"52",
          2109 => x"51",
          2110 => x"3f",
          2111 => x"08",
          2112 => x"81",
          2113 => x"38",
          2114 => x"3d",
          2115 => x"fb",
          2116 => x"d5",
          2117 => x"db",
          2118 => x"81",
          2119 => x"fe",
          2120 => x"d6",
          2121 => x"55",
          2122 => x"54",
          2123 => x"d6",
          2124 => x"51",
          2125 => x"fd",
          2126 => x"8c",
          2127 => x"ff",
          2128 => x"3f",
          2129 => x"81",
          2130 => x"bf",
          2131 => x"ef",
          2132 => x"d6",
          2133 => x"39",
          2134 => x"51",
          2135 => x"80",
          2136 => x"83",
          2137 => x"de",
          2138 => x"fd",
          2139 => x"39",
          2140 => x"84",
          2141 => x"80",
          2142 => x"8a",
          2143 => x"c8",
          2144 => x"fa",
          2145 => x"52",
          2146 => x"51",
          2147 => x"68",
          2148 => x"84",
          2149 => x"80",
          2150 => x"38",
          2151 => x"08",
          2152 => x"f0",
          2153 => x"3f",
          2154 => x"b8",
          2155 => x"11",
          2156 => x"05",
          2157 => x"3f",
          2158 => x"08",
          2159 => x"ff",
          2160 => x"83",
          2161 => x"d0",
          2162 => x"59",
          2163 => x"3d",
          2164 => x"53",
          2165 => x"51",
          2166 => x"84",
          2167 => x"80",
          2168 => x"38",
          2169 => x"f0",
          2170 => x"80",
          2171 => x"92",
          2172 => x"c8",
          2173 => x"38",
          2174 => x"08",
          2175 => x"83",
          2176 => x"d0",
          2177 => x"d5",
          2178 => x"80",
          2179 => x"51",
          2180 => x"7e",
          2181 => x"59",
          2182 => x"f9",
          2183 => x"9f",
          2184 => x"38",
          2185 => x"70",
          2186 => x"39",
          2187 => x"f4",
          2188 => x"80",
          2189 => x"ca",
          2190 => x"c8",
          2191 => x"f8",
          2192 => x"3d",
          2193 => x"53",
          2194 => x"51",
          2195 => x"84",
          2196 => x"86",
          2197 => x"59",
          2198 => x"78",
          2199 => x"b8",
          2200 => x"3f",
          2201 => x"08",
          2202 => x"52",
          2203 => x"b3",
          2204 => x"7e",
          2205 => x"ae",
          2206 => x"38",
          2207 => x"87",
          2208 => x"82",
          2209 => x"59",
          2210 => x"3d",
          2211 => x"53",
          2212 => x"51",
          2213 => x"84",
          2214 => x"80",
          2215 => x"38",
          2216 => x"fc",
          2217 => x"80",
          2218 => x"da",
          2219 => x"c8",
          2220 => x"f8",
          2221 => x"3d",
          2222 => x"53",
          2223 => x"51",
          2224 => x"84",
          2225 => x"80",
          2226 => x"38",
          2227 => x"51",
          2228 => x"68",
          2229 => x"78",
          2230 => x"8d",
          2231 => x"33",
          2232 => x"5c",
          2233 => x"2e",
          2234 => x"55",
          2235 => x"33",
          2236 => x"83",
          2237 => x"ce",
          2238 => x"66",
          2239 => x"19",
          2240 => x"59",
          2241 => x"3d",
          2242 => x"53",
          2243 => x"51",
          2244 => x"84",
          2245 => x"80",
          2246 => x"38",
          2247 => x"fc",
          2248 => x"80",
          2249 => x"de",
          2250 => x"c8",
          2251 => x"f7",
          2252 => x"3d",
          2253 => x"53",
          2254 => x"51",
          2255 => x"84",
          2256 => x"80",
          2257 => x"38",
          2258 => x"51",
          2259 => x"68",
          2260 => x"27",
          2261 => x"65",
          2262 => x"81",
          2263 => x"7c",
          2264 => x"05",
          2265 => x"b8",
          2266 => x"11",
          2267 => x"05",
          2268 => x"3f",
          2269 => x"08",
          2270 => x"c3",
          2271 => x"fe",
          2272 => x"ff",
          2273 => x"e7",
          2274 => x"b9",
          2275 => x"38",
          2276 => x"54",
          2277 => x"fc",
          2278 => x"3f",
          2279 => x"08",
          2280 => x"52",
          2281 => x"fb",
          2282 => x"7e",
          2283 => x"ae",
          2284 => x"38",
          2285 => x"84",
          2286 => x"81",
          2287 => x"39",
          2288 => x"80",
          2289 => x"79",
          2290 => x"05",
          2291 => x"fe",
          2292 => x"ff",
          2293 => x"e7",
          2294 => x"b9",
          2295 => x"2e",
          2296 => x"68",
          2297 => x"db",
          2298 => x"34",
          2299 => x"49",
          2300 => x"fc",
          2301 => x"80",
          2302 => x"8a",
          2303 => x"c8",
          2304 => x"38",
          2305 => x"b8",
          2306 => x"11",
          2307 => x"05",
          2308 => x"3f",
          2309 => x"08",
          2310 => x"a3",
          2311 => x"fe",
          2312 => x"ff",
          2313 => x"e6",
          2314 => x"b9",
          2315 => x"2e",
          2316 => x"b8",
          2317 => x"11",
          2318 => x"05",
          2319 => x"3f",
          2320 => x"08",
          2321 => x"b9",
          2322 => x"83",
          2323 => x"cb",
          2324 => x"67",
          2325 => x"7a",
          2326 => x"65",
          2327 => x"70",
          2328 => x"0c",
          2329 => x"f5",
          2330 => x"d9",
          2331 => x"cf",
          2332 => x"ff",
          2333 => x"87",
          2334 => x"b9",
          2335 => x"3d",
          2336 => x"52",
          2337 => x"3f",
          2338 => x"b9",
          2339 => x"78",
          2340 => x"3f",
          2341 => x"08",
          2342 => x"a3",
          2343 => x"c8",
          2344 => x"f6",
          2345 => x"39",
          2346 => x"84",
          2347 => x"80",
          2348 => x"d2",
          2349 => x"c8",
          2350 => x"83",
          2351 => x"5a",
          2352 => x"83",
          2353 => x"f2",
          2354 => x"b8",
          2355 => x"11",
          2356 => x"05",
          2357 => x"3f",
          2358 => x"08",
          2359 => x"f2",
          2360 => x"79",
          2361 => x"8a",
          2362 => x"88",
          2363 => x"3d",
          2364 => x"53",
          2365 => x"51",
          2366 => x"84",
          2367 => x"80",
          2368 => x"80",
          2369 => x"7a",
          2370 => x"38",
          2371 => x"90",
          2372 => x"70",
          2373 => x"2a",
          2374 => x"5f",
          2375 => x"2e",
          2376 => x"a0",
          2377 => x"88",
          2378 => x"98",
          2379 => x"3f",
          2380 => x"54",
          2381 => x"52",
          2382 => x"a8",
          2383 => x"a4",
          2384 => x"3f",
          2385 => x"64",
          2386 => x"59",
          2387 => x"45",
          2388 => x"f0",
          2389 => x"80",
          2390 => x"a6",
          2391 => x"c8",
          2392 => x"f2",
          2393 => x"64",
          2394 => x"64",
          2395 => x"b8",
          2396 => x"11",
          2397 => x"05",
          2398 => x"3f",
          2399 => x"08",
          2400 => x"bb",
          2401 => x"02",
          2402 => x"22",
          2403 => x"05",
          2404 => x"45",
          2405 => x"f0",
          2406 => x"80",
          2407 => x"e2",
          2408 => x"c8",
          2409 => x"f2",
          2410 => x"5e",
          2411 => x"05",
          2412 => x"82",
          2413 => x"7d",
          2414 => x"fe",
          2415 => x"ff",
          2416 => x"e1",
          2417 => x"b9",
          2418 => x"b9",
          2419 => x"39",
          2420 => x"fc",
          2421 => x"80",
          2422 => x"aa",
          2423 => x"c8",
          2424 => x"81",
          2425 => x"5c",
          2426 => x"05",
          2427 => x"68",
          2428 => x"fb",
          2429 => x"3d",
          2430 => x"53",
          2431 => x"51",
          2432 => x"84",
          2433 => x"80",
          2434 => x"38",
          2435 => x"0c",
          2436 => x"05",
          2437 => x"f7",
          2438 => x"83",
          2439 => x"06",
          2440 => x"7b",
          2441 => x"90",
          2442 => x"83",
          2443 => x"7c",
          2444 => x"3f",
          2445 => x"7b",
          2446 => x"da",
          2447 => x"8c",
          2448 => x"bc",
          2449 => x"3f",
          2450 => x"b8",
          2451 => x"11",
          2452 => x"05",
          2453 => x"3f",
          2454 => x"08",
          2455 => x"38",
          2456 => x"80",
          2457 => x"79",
          2458 => x"5b",
          2459 => x"f7",
          2460 => x"f2",
          2461 => x"7b",
          2462 => x"cf",
          2463 => x"90",
          2464 => x"ea",
          2465 => x"cd",
          2466 => x"80",
          2467 => x"83",
          2468 => x"49",
          2469 => x"83",
          2470 => x"d3",
          2471 => x"59",
          2472 => x"83",
          2473 => x"d3",
          2474 => x"59",
          2475 => x"83",
          2476 => x"59",
          2477 => x"a5",
          2478 => x"94",
          2479 => x"8b",
          2480 => x"e8",
          2481 => x"3f",
          2482 => x"83",
          2483 => x"59",
          2484 => x"9b",
          2485 => x"98",
          2486 => x"92",
          2487 => x"cf",
          2488 => x"80",
          2489 => x"83",
          2490 => x"49",
          2491 => x"83",
          2492 => x"5e",
          2493 => x"9b",
          2494 => x"a0",
          2495 => x"ee",
          2496 => x"ca",
          2497 => x"80",
          2498 => x"83",
          2499 => x"49",
          2500 => x"83",
          2501 => x"5d",
          2502 => x"94",
          2503 => x"a8",
          2504 => x"ca",
          2505 => x"b4",
          2506 => x"05",
          2507 => x"39",
          2508 => x"08",
          2509 => x"fb",
          2510 => x"3d",
          2511 => x"84",
          2512 => x"87",
          2513 => x"70",
          2514 => x"87",
          2515 => x"74",
          2516 => x"3f",
          2517 => x"08",
          2518 => x"08",
          2519 => x"84",
          2520 => x"51",
          2521 => x"74",
          2522 => x"08",
          2523 => x"87",
          2524 => x"70",
          2525 => x"87",
          2526 => x"74",
          2527 => x"3f",
          2528 => x"08",
          2529 => x"08",
          2530 => x"84",
          2531 => x"51",
          2532 => x"74",
          2533 => x"08",
          2534 => x"8c",
          2535 => x"87",
          2536 => x"0c",
          2537 => x"0b",
          2538 => x"94",
          2539 => x"f2",
          2540 => x"f1",
          2541 => x"84",
          2542 => x"34",
          2543 => x"d5",
          2544 => x"3d",
          2545 => x"0c",
          2546 => x"84",
          2547 => x"56",
          2548 => x"89",
          2549 => x"97",
          2550 => x"51",
          2551 => x"83",
          2552 => x"83",
          2553 => x"c4",
          2554 => x"f2",
          2555 => x"52",
          2556 => x"3f",
          2557 => x"54",
          2558 => x"53",
          2559 => x"52",
          2560 => x"51",
          2561 => x"8d",
          2562 => x"d2",
          2563 => x"e3",
          2564 => x"83",
          2565 => x"c3",
          2566 => x"80",
          2567 => x"d3",
          2568 => x"e4",
          2569 => x"3f",
          2570 => x"3d",
          2571 => x"08",
          2572 => x"75",
          2573 => x"73",
          2574 => x"38",
          2575 => x"81",
          2576 => x"52",
          2577 => x"09",
          2578 => x"38",
          2579 => x"33",
          2580 => x"06",
          2581 => x"70",
          2582 => x"38",
          2583 => x"06",
          2584 => x"2e",
          2585 => x"74",
          2586 => x"2e",
          2587 => x"80",
          2588 => x"81",
          2589 => x"54",
          2590 => x"2e",
          2591 => x"54",
          2592 => x"8b",
          2593 => x"2e",
          2594 => x"12",
          2595 => x"80",
          2596 => x"06",
          2597 => x"a0",
          2598 => x"06",
          2599 => x"54",
          2600 => x"70",
          2601 => x"25",
          2602 => x"52",
          2603 => x"2e",
          2604 => x"72",
          2605 => x"54",
          2606 => x"0c",
          2607 => x"84",
          2608 => x"87",
          2609 => x"70",
          2610 => x"38",
          2611 => x"ff",
          2612 => x"12",
          2613 => x"33",
          2614 => x"06",
          2615 => x"70",
          2616 => x"38",
          2617 => x"39",
          2618 => x"81",
          2619 => x"72",
          2620 => x"81",
          2621 => x"38",
          2622 => x"3d",
          2623 => x"72",
          2624 => x"80",
          2625 => x"c8",
          2626 => x"0d",
          2627 => x"fc",
          2628 => x"51",
          2629 => x"84",
          2630 => x"80",
          2631 => x"74",
          2632 => x"0c",
          2633 => x"04",
          2634 => x"76",
          2635 => x"ff",
          2636 => x"81",
          2637 => x"26",
          2638 => x"83",
          2639 => x"05",
          2640 => x"73",
          2641 => x"8a",
          2642 => x"33",
          2643 => x"70",
          2644 => x"fe",
          2645 => x"33",
          2646 => x"73",
          2647 => x"f2",
          2648 => x"33",
          2649 => x"74",
          2650 => x"e6",
          2651 => x"22",
          2652 => x"74",
          2653 => x"80",
          2654 => x"13",
          2655 => x"52",
          2656 => x"26",
          2657 => x"81",
          2658 => x"98",
          2659 => x"22",
          2660 => x"bc",
          2661 => x"33",
          2662 => x"b8",
          2663 => x"33",
          2664 => x"b4",
          2665 => x"33",
          2666 => x"b0",
          2667 => x"33",
          2668 => x"ac",
          2669 => x"33",
          2670 => x"a8",
          2671 => x"c0",
          2672 => x"73",
          2673 => x"a0",
          2674 => x"87",
          2675 => x"0c",
          2676 => x"84",
          2677 => x"86",
          2678 => x"f3",
          2679 => x"5b",
          2680 => x"9c",
          2681 => x"0c",
          2682 => x"bc",
          2683 => x"7b",
          2684 => x"98",
          2685 => x"7b",
          2686 => x"87",
          2687 => x"08",
          2688 => x"1c",
          2689 => x"98",
          2690 => x"7b",
          2691 => x"87",
          2692 => x"08",
          2693 => x"1c",
          2694 => x"98",
          2695 => x"7b",
          2696 => x"87",
          2697 => x"08",
          2698 => x"1c",
          2699 => x"98",
          2700 => x"79",
          2701 => x"80",
          2702 => x"83",
          2703 => x"59",
          2704 => x"ff",
          2705 => x"1b",
          2706 => x"1b",
          2707 => x"1b",
          2708 => x"1b",
          2709 => x"1b",
          2710 => x"83",
          2711 => x"52",
          2712 => x"51",
          2713 => x"3f",
          2714 => x"04",
          2715 => x"02",
          2716 => x"53",
          2717 => x"a8",
          2718 => x"80",
          2719 => x"84",
          2720 => x"98",
          2721 => x"2c",
          2722 => x"ff",
          2723 => x"06",
          2724 => x"83",
          2725 => x"71",
          2726 => x"0c",
          2727 => x"04",
          2728 => x"e7",
          2729 => x"b9",
          2730 => x"2b",
          2731 => x"51",
          2732 => x"2e",
          2733 => x"df",
          2734 => x"80",
          2735 => x"84",
          2736 => x"98",
          2737 => x"2c",
          2738 => x"ff",
          2739 => x"c7",
          2740 => x"0d",
          2741 => x"52",
          2742 => x"54",
          2743 => x"e7",
          2744 => x"b9",
          2745 => x"2b",
          2746 => x"51",
          2747 => x"2e",
          2748 => x"72",
          2749 => x"54",
          2750 => x"25",
          2751 => x"84",
          2752 => x"85",
          2753 => x"fc",
          2754 => x"9b",
          2755 => x"f2",
          2756 => x"81",
          2757 => x"55",
          2758 => x"2e",
          2759 => x"87",
          2760 => x"08",
          2761 => x"70",
          2762 => x"54",
          2763 => x"2e",
          2764 => x"91",
          2765 => x"06",
          2766 => x"e3",
          2767 => x"32",
          2768 => x"72",
          2769 => x"38",
          2770 => x"81",
          2771 => x"cf",
          2772 => x"ff",
          2773 => x"c0",
          2774 => x"70",
          2775 => x"38",
          2776 => x"90",
          2777 => x"0c",
          2778 => x"c8",
          2779 => x"0d",
          2780 => x"2a",
          2781 => x"51",
          2782 => x"38",
          2783 => x"81",
          2784 => x"80",
          2785 => x"71",
          2786 => x"06",
          2787 => x"2e",
          2788 => x"c0",
          2789 => x"70",
          2790 => x"81",
          2791 => x"52",
          2792 => x"d8",
          2793 => x"0d",
          2794 => x"33",
          2795 => x"9f",
          2796 => x"52",
          2797 => x"80",
          2798 => x"0d",
          2799 => x"0d",
          2800 => x"75",
          2801 => x"52",
          2802 => x"2e",
          2803 => x"81",
          2804 => x"80",
          2805 => x"ff",
          2806 => x"55",
          2807 => x"80",
          2808 => x"c0",
          2809 => x"70",
          2810 => x"81",
          2811 => x"52",
          2812 => x"8c",
          2813 => x"2a",
          2814 => x"51",
          2815 => x"38",
          2816 => x"81",
          2817 => x"80",
          2818 => x"71",
          2819 => x"06",
          2820 => x"38",
          2821 => x"06",
          2822 => x"94",
          2823 => x"80",
          2824 => x"87",
          2825 => x"52",
          2826 => x"81",
          2827 => x"55",
          2828 => x"9b",
          2829 => x"b9",
          2830 => x"3d",
          2831 => x"91",
          2832 => x"06",
          2833 => x"98",
          2834 => x"32",
          2835 => x"72",
          2836 => x"38",
          2837 => x"81",
          2838 => x"80",
          2839 => x"38",
          2840 => x"84",
          2841 => x"2a",
          2842 => x"53",
          2843 => x"ce",
          2844 => x"ff",
          2845 => x"c0",
          2846 => x"70",
          2847 => x"06",
          2848 => x"80",
          2849 => x"38",
          2850 => x"a4",
          2851 => x"84",
          2852 => x"9e",
          2853 => x"f2",
          2854 => x"c0",
          2855 => x"83",
          2856 => x"87",
          2857 => x"08",
          2858 => x"0c",
          2859 => x"9c",
          2860 => x"94",
          2861 => x"9e",
          2862 => x"f2",
          2863 => x"c0",
          2864 => x"83",
          2865 => x"87",
          2866 => x"08",
          2867 => x"0c",
          2868 => x"b4",
          2869 => x"a4",
          2870 => x"9e",
          2871 => x"f2",
          2872 => x"c0",
          2873 => x"83",
          2874 => x"87",
          2875 => x"08",
          2876 => x"0c",
          2877 => x"c4",
          2878 => x"b4",
          2879 => x"9e",
          2880 => x"71",
          2881 => x"23",
          2882 => x"84",
          2883 => x"bc",
          2884 => x"9e",
          2885 => x"f2",
          2886 => x"c0",
          2887 => x"83",
          2888 => x"81",
          2889 => x"c8",
          2890 => x"87",
          2891 => x"08",
          2892 => x"0a",
          2893 => x"52",
          2894 => x"38",
          2895 => x"c9",
          2896 => x"87",
          2897 => x"08",
          2898 => x"0a",
          2899 => x"52",
          2900 => x"83",
          2901 => x"71",
          2902 => x"34",
          2903 => x"c0",
          2904 => x"70",
          2905 => x"06",
          2906 => x"70",
          2907 => x"38",
          2908 => x"83",
          2909 => x"80",
          2910 => x"9e",
          2911 => x"88",
          2912 => x"51",
          2913 => x"80",
          2914 => x"81",
          2915 => x"f2",
          2916 => x"0b",
          2917 => x"90",
          2918 => x"80",
          2919 => x"52",
          2920 => x"2e",
          2921 => x"52",
          2922 => x"cd",
          2923 => x"87",
          2924 => x"08",
          2925 => x"80",
          2926 => x"52",
          2927 => x"83",
          2928 => x"71",
          2929 => x"34",
          2930 => x"c0",
          2931 => x"70",
          2932 => x"06",
          2933 => x"70",
          2934 => x"38",
          2935 => x"83",
          2936 => x"80",
          2937 => x"9e",
          2938 => x"82",
          2939 => x"51",
          2940 => x"80",
          2941 => x"81",
          2942 => x"f2",
          2943 => x"0b",
          2944 => x"90",
          2945 => x"80",
          2946 => x"52",
          2947 => x"2e",
          2948 => x"52",
          2949 => x"d1",
          2950 => x"87",
          2951 => x"08",
          2952 => x"80",
          2953 => x"52",
          2954 => x"83",
          2955 => x"71",
          2956 => x"34",
          2957 => x"c0",
          2958 => x"70",
          2959 => x"51",
          2960 => x"80",
          2961 => x"81",
          2962 => x"f2",
          2963 => x"c0",
          2964 => x"98",
          2965 => x"8a",
          2966 => x"71",
          2967 => x"34",
          2968 => x"c0",
          2969 => x"70",
          2970 => x"51",
          2971 => x"80",
          2972 => x"81",
          2973 => x"f2",
          2974 => x"c0",
          2975 => x"83",
          2976 => x"84",
          2977 => x"71",
          2978 => x"34",
          2979 => x"c0",
          2980 => x"70",
          2981 => x"52",
          2982 => x"2e",
          2983 => x"52",
          2984 => x"d7",
          2985 => x"9e",
          2986 => x"06",
          2987 => x"f2",
          2988 => x"3d",
          2989 => x"52",
          2990 => x"fb",
          2991 => x"d9",
          2992 => x"b6",
          2993 => x"f2",
          2994 => x"73",
          2995 => x"83",
          2996 => x"c3",
          2997 => x"f2",
          2998 => x"74",
          2999 => x"83",
          3000 => x"54",
          3001 => x"38",
          3002 => x"33",
          3003 => x"9d",
          3004 => x"cd",
          3005 => x"84",
          3006 => x"f2",
          3007 => x"73",
          3008 => x"83",
          3009 => x"56",
          3010 => x"38",
          3011 => x"33",
          3012 => x"85",
          3013 => x"d5",
          3014 => x"83",
          3015 => x"f2",
          3016 => x"75",
          3017 => x"83",
          3018 => x"54",
          3019 => x"38",
          3020 => x"33",
          3021 => x"88",
          3022 => x"d1",
          3023 => x"82",
          3024 => x"f2",
          3025 => x"73",
          3026 => x"83",
          3027 => x"c2",
          3028 => x"f2",
          3029 => x"83",
          3030 => x"ff",
          3031 => x"83",
          3032 => x"52",
          3033 => x"51",
          3034 => x"3f",
          3035 => x"08",
          3036 => x"8c",
          3037 => x"90",
          3038 => x"b4",
          3039 => x"3f",
          3040 => x"22",
          3041 => x"bc",
          3042 => x"fc",
          3043 => x"bc",
          3044 => x"84",
          3045 => x"51",
          3046 => x"84",
          3047 => x"bd",
          3048 => x"76",
          3049 => x"54",
          3050 => x"08",
          3051 => x"e4",
          3052 => x"d4",
          3053 => x"cf",
          3054 => x"b9",
          3055 => x"ca",
          3056 => x"85",
          3057 => x"0d",
          3058 => x"c4",
          3059 => x"84",
          3060 => x"51",
          3061 => x"84",
          3062 => x"bd",
          3063 => x"76",
          3064 => x"54",
          3065 => x"08",
          3066 => x"90",
          3067 => x"98",
          3068 => x"0d",
          3069 => x"c0",
          3070 => x"84",
          3071 => x"51",
          3072 => x"84",
          3073 => x"bd",
          3074 => x"76",
          3075 => x"54",
          3076 => x"08",
          3077 => x"bc",
          3078 => x"ec",
          3079 => x"ca",
          3080 => x"80",
          3081 => x"38",
          3082 => x"83",
          3083 => x"c0",
          3084 => x"d9",
          3085 => x"bb",
          3086 => x"ac",
          3087 => x"d9",
          3088 => x"b3",
          3089 => x"f2",
          3090 => x"83",
          3091 => x"ff",
          3092 => x"83",
          3093 => x"52",
          3094 => x"51",
          3095 => x"3f",
          3096 => x"51",
          3097 => x"83",
          3098 => x"52",
          3099 => x"51",
          3100 => x"3f",
          3101 => x"08",
          3102 => x"c0",
          3103 => x"c8",
          3104 => x"b9",
          3105 => x"84",
          3106 => x"71",
          3107 => x"84",
          3108 => x"52",
          3109 => x"51",
          3110 => x"3f",
          3111 => x"33",
          3112 => x"2e",
          3113 => x"fe",
          3114 => x"db",
          3115 => x"bf",
          3116 => x"f2",
          3117 => x"73",
          3118 => x"8f",
          3119 => x"39",
          3120 => x"51",
          3121 => x"3f",
          3122 => x"33",
          3123 => x"2e",
          3124 => x"d6",
          3125 => x"84",
          3126 => x"97",
          3127 => x"d0",
          3128 => x"80",
          3129 => x"38",
          3130 => x"dc",
          3131 => x"bf",
          3132 => x"f2",
          3133 => x"73",
          3134 => x"b4",
          3135 => x"83",
          3136 => x"52",
          3137 => x"51",
          3138 => x"3f",
          3139 => x"33",
          3140 => x"2e",
          3141 => x"d2",
          3142 => x"d8",
          3143 => x"dc",
          3144 => x"b1",
          3145 => x"f2",
          3146 => x"74",
          3147 => x"ee",
          3148 => x"83",
          3149 => x"52",
          3150 => x"51",
          3151 => x"3f",
          3152 => x"33",
          3153 => x"2e",
          3154 => x"cd",
          3155 => x"94",
          3156 => x"98",
          3157 => x"52",
          3158 => x"51",
          3159 => x"3f",
          3160 => x"33",
          3161 => x"2e",
          3162 => x"c7",
          3163 => x"8c",
          3164 => x"90",
          3165 => x"52",
          3166 => x"51",
          3167 => x"3f",
          3168 => x"33",
          3169 => x"2e",
          3170 => x"c1",
          3171 => x"84",
          3172 => x"88",
          3173 => x"52",
          3174 => x"51",
          3175 => x"3f",
          3176 => x"33",
          3177 => x"2e",
          3178 => x"c1",
          3179 => x"9c",
          3180 => x"a0",
          3181 => x"52",
          3182 => x"51",
          3183 => x"3f",
          3184 => x"33",
          3185 => x"2e",
          3186 => x"c1",
          3187 => x"a4",
          3188 => x"a8",
          3189 => x"52",
          3190 => x"51",
          3191 => x"3f",
          3192 => x"33",
          3193 => x"2e",
          3194 => x"c1",
          3195 => x"90",
          3196 => x"94",
          3197 => x"98",
          3198 => x"f7",
          3199 => x"ca",
          3200 => x"80",
          3201 => x"38",
          3202 => x"3d",
          3203 => x"05",
          3204 => x"85",
          3205 => x"71",
          3206 => x"c2",
          3207 => x"71",
          3208 => x"de",
          3209 => x"af",
          3210 => x"3d",
          3211 => x"de",
          3212 => x"af",
          3213 => x"3d",
          3214 => x"de",
          3215 => x"af",
          3216 => x"3d",
          3217 => x"de",
          3218 => x"af",
          3219 => x"3d",
          3220 => x"de",
          3221 => x"af",
          3222 => x"3d",
          3223 => x"de",
          3224 => x"af",
          3225 => x"3d",
          3226 => x"88",
          3227 => x"80",
          3228 => x"96",
          3229 => x"83",
          3230 => x"87",
          3231 => x"0c",
          3232 => x"0d",
          3233 => x"ad",
          3234 => x"5a",
          3235 => x"58",
          3236 => x"f3",
          3237 => x"82",
          3238 => x"84",
          3239 => x"80",
          3240 => x"3d",
          3241 => x"83",
          3242 => x"54",
          3243 => x"52",
          3244 => x"d2",
          3245 => x"b9",
          3246 => x"2e",
          3247 => x"51",
          3248 => x"84",
          3249 => x"81",
          3250 => x"80",
          3251 => x"c8",
          3252 => x"38",
          3253 => x"08",
          3254 => x"18",
          3255 => x"74",
          3256 => x"70",
          3257 => x"07",
          3258 => x"55",
          3259 => x"2e",
          3260 => x"ff",
          3261 => x"f3",
          3262 => x"11",
          3263 => x"82",
          3264 => x"84",
          3265 => x"8f",
          3266 => x"2e",
          3267 => x"84",
          3268 => x"a9",
          3269 => x"83",
          3270 => x"ff",
          3271 => x"78",
          3272 => x"81",
          3273 => x"76",
          3274 => x"c0",
          3275 => x"51",
          3276 => x"3f",
          3277 => x"56",
          3278 => x"08",
          3279 => x"52",
          3280 => x"51",
          3281 => x"3f",
          3282 => x"b9",
          3283 => x"3d",
          3284 => x"3d",
          3285 => x"08",
          3286 => x"71",
          3287 => x"33",
          3288 => x"57",
          3289 => x"81",
          3290 => x"0b",
          3291 => x"56",
          3292 => x"10",
          3293 => x"05",
          3294 => x"54",
          3295 => x"3f",
          3296 => x"08",
          3297 => x"73",
          3298 => x"89",
          3299 => x"c8",
          3300 => x"84",
          3301 => x"73",
          3302 => x"88",
          3303 => x"2e",
          3304 => x"16",
          3305 => x"06",
          3306 => x"76",
          3307 => x"80",
          3308 => x"b9",
          3309 => x"3d",
          3310 => x"1a",
          3311 => x"ff",
          3312 => x"ff",
          3313 => x"c7",
          3314 => x"b9",
          3315 => x"2e",
          3316 => x"1b",
          3317 => x"76",
          3318 => x"3f",
          3319 => x"08",
          3320 => x"54",
          3321 => x"c9",
          3322 => x"70",
          3323 => x"57",
          3324 => x"27",
          3325 => x"ff",
          3326 => x"33",
          3327 => x"76",
          3328 => x"e6",
          3329 => x"70",
          3330 => x"55",
          3331 => x"2e",
          3332 => x"fe",
          3333 => x"75",
          3334 => x"80",
          3335 => x"59",
          3336 => x"39",
          3337 => x"c8",
          3338 => x"f3",
          3339 => x"56",
          3340 => x"3f",
          3341 => x"08",
          3342 => x"83",
          3343 => x"53",
          3344 => x"77",
          3345 => x"fd",
          3346 => x"c8",
          3347 => x"ba",
          3348 => x"ff",
          3349 => x"84",
          3350 => x"55",
          3351 => x"b9",
          3352 => x"9d",
          3353 => x"c8",
          3354 => x"70",
          3355 => x"80",
          3356 => x"53",
          3357 => x"16",
          3358 => x"52",
          3359 => x"88",
          3360 => x"2e",
          3361 => x"ff",
          3362 => x"0b",
          3363 => x"0c",
          3364 => x"04",
          3365 => x"b5",
          3366 => x"3d",
          3367 => x"08",
          3368 => x"80",
          3369 => x"34",
          3370 => x"33",
          3371 => x"08",
          3372 => x"9e",
          3373 => x"f3",
          3374 => x"56",
          3375 => x"82",
          3376 => x"80",
          3377 => x"38",
          3378 => x"06",
          3379 => x"90",
          3380 => x"80",
          3381 => x"38",
          3382 => x"3d",
          3383 => x"51",
          3384 => x"84",
          3385 => x"98",
          3386 => x"2c",
          3387 => x"ff",
          3388 => x"79",
          3389 => x"84",
          3390 => x"70",
          3391 => x"98",
          3392 => x"80",
          3393 => x"2b",
          3394 => x"71",
          3395 => x"70",
          3396 => x"de",
          3397 => x"08",
          3398 => x"52",
          3399 => x"46",
          3400 => x"5c",
          3401 => x"74",
          3402 => x"cd",
          3403 => x"27",
          3404 => x"75",
          3405 => x"29",
          3406 => x"05",
          3407 => x"57",
          3408 => x"24",
          3409 => x"75",
          3410 => x"82",
          3411 => x"80",
          3412 => x"d4",
          3413 => x"57",
          3414 => x"91",
          3415 => x"d0",
          3416 => x"70",
          3417 => x"78",
          3418 => x"95",
          3419 => x"2e",
          3420 => x"84",
          3421 => x"81",
          3422 => x"2e",
          3423 => x"81",
          3424 => x"2b",
          3425 => x"84",
          3426 => x"70",
          3427 => x"97",
          3428 => x"2c",
          3429 => x"2b",
          3430 => x"11",
          3431 => x"5f",
          3432 => x"57",
          3433 => x"2e",
          3434 => x"76",
          3435 => x"34",
          3436 => x"81",
          3437 => x"ba",
          3438 => x"80",
          3439 => x"80",
          3440 => x"98",
          3441 => x"ff",
          3442 => x"41",
          3443 => x"80",
          3444 => x"10",
          3445 => x"2b",
          3446 => x"0b",
          3447 => x"16",
          3448 => x"77",
          3449 => x"38",
          3450 => x"15",
          3451 => x"33",
          3452 => x"61",
          3453 => x"38",
          3454 => x"ff",
          3455 => x"f2",
          3456 => x"76",
          3457 => x"ab",
          3458 => x"39",
          3459 => x"b2",
          3460 => x"76",
          3461 => x"76",
          3462 => x"34",
          3463 => x"80",
          3464 => x"34",
          3465 => x"62",
          3466 => x"26",
          3467 => x"74",
          3468 => x"c3",
          3469 => x"76",
          3470 => x"de",
          3471 => x"7f",
          3472 => x"84",
          3473 => x"80",
          3474 => x"80",
          3475 => x"84",
          3476 => x"56",
          3477 => x"fd",
          3478 => x"d5",
          3479 => x"88",
          3480 => x"8a",
          3481 => x"8c",
          3482 => x"57",
          3483 => x"8c",
          3484 => x"39",
          3485 => x"33",
          3486 => x"06",
          3487 => x"33",
          3488 => x"75",
          3489 => x"d6",
          3490 => x"ac",
          3491 => x"15",
          3492 => x"d1",
          3493 => x"16",
          3494 => x"55",
          3495 => x"3f",
          3496 => x"7c",
          3497 => x"da",
          3498 => x"10",
          3499 => x"05",
          3500 => x"59",
          3501 => x"38",
          3502 => x"88",
          3503 => x"34",
          3504 => x"33",
          3505 => x"33",
          3506 => x"80",
          3507 => x"84",
          3508 => x"52",
          3509 => x"b5",
          3510 => x"d5",
          3511 => x"a0",
          3512 => x"8a",
          3513 => x"ac",
          3514 => x"51",
          3515 => x"3f",
          3516 => x"33",
          3517 => x"7a",
          3518 => x"34",
          3519 => x"06",
          3520 => x"38",
          3521 => x"a5",
          3522 => x"84",
          3523 => x"fb",
          3524 => x"8a",
          3525 => x"ac",
          3526 => x"8d",
          3527 => x"10",
          3528 => x"e0",
          3529 => x"08",
          3530 => x"8e",
          3531 => x"08",
          3532 => x"2e",
          3533 => x"75",
          3534 => x"ec",
          3535 => x"c8",
          3536 => x"88",
          3537 => x"c8",
          3538 => x"06",
          3539 => x"75",
          3540 => x"ff",
          3541 => x"84",
          3542 => x"84",
          3543 => x"56",
          3544 => x"2e",
          3545 => x"84",
          3546 => x"52",
          3547 => x"b3",
          3548 => x"d5",
          3549 => x"a0",
          3550 => x"f2",
          3551 => x"ac",
          3552 => x"51",
          3553 => x"3f",
          3554 => x"33",
          3555 => x"74",
          3556 => x"34",
          3557 => x"06",
          3558 => x"84",
          3559 => x"70",
          3560 => x"84",
          3561 => x"5b",
          3562 => x"79",
          3563 => x"38",
          3564 => x"08",
          3565 => x"57",
          3566 => x"8c",
          3567 => x"70",
          3568 => x"ff",
          3569 => x"84",
          3570 => x"70",
          3571 => x"84",
          3572 => x"5a",
          3573 => x"78",
          3574 => x"38",
          3575 => x"08",
          3576 => x"57",
          3577 => x"8c",
          3578 => x"70",
          3579 => x"ff",
          3580 => x"84",
          3581 => x"70",
          3582 => x"84",
          3583 => x"5a",
          3584 => x"76",
          3585 => x"38",
          3586 => x"84",
          3587 => x"84",
          3588 => x"56",
          3589 => x"2e",
          3590 => x"ff",
          3591 => x"84",
          3592 => x"75",
          3593 => x"98",
          3594 => x"ff",
          3595 => x"5a",
          3596 => x"80",
          3597 => x"d5",
          3598 => x"a0",
          3599 => x"ae",
          3600 => x"8c",
          3601 => x"2b",
          3602 => x"84",
          3603 => x"5a",
          3604 => x"74",
          3605 => x"86",
          3606 => x"ac",
          3607 => x"51",
          3608 => x"3f",
          3609 => x"0a",
          3610 => x"0a",
          3611 => x"2c",
          3612 => x"33",
          3613 => x"74",
          3614 => x"e2",
          3615 => x"ac",
          3616 => x"51",
          3617 => x"3f",
          3618 => x"0a",
          3619 => x"0a",
          3620 => x"2c",
          3621 => x"33",
          3622 => x"7a",
          3623 => x"b9",
          3624 => x"39",
          3625 => x"81",
          3626 => x"34",
          3627 => x"08",
          3628 => x"51",
          3629 => x"3f",
          3630 => x"0a",
          3631 => x"0a",
          3632 => x"2c",
          3633 => x"33",
          3634 => x"75",
          3635 => x"e6",
          3636 => x"58",
          3637 => x"78",
          3638 => x"ac",
          3639 => x"33",
          3640 => x"8a",
          3641 => x"80",
          3642 => x"80",
          3643 => x"98",
          3644 => x"88",
          3645 => x"55",
          3646 => x"ff",
          3647 => x"b6",
          3648 => x"8c",
          3649 => x"80",
          3650 => x"38",
          3651 => x"08",
          3652 => x"ff",
          3653 => x"84",
          3654 => x"ff",
          3655 => x"84",
          3656 => x"76",
          3657 => x"55",
          3658 => x"d1",
          3659 => x"05",
          3660 => x"34",
          3661 => x"08",
          3662 => x"ff",
          3663 => x"84",
          3664 => x"7b",
          3665 => x"3f",
          3666 => x"08",
          3667 => x"58",
          3668 => x"38",
          3669 => x"33",
          3670 => x"2e",
          3671 => x"83",
          3672 => x"70",
          3673 => x"f2",
          3674 => x"08",
          3675 => x"74",
          3676 => x"75",
          3677 => x"fc",
          3678 => x"e0",
          3679 => x"70",
          3680 => x"80",
          3681 => x"84",
          3682 => x"7b",
          3683 => x"b8",
          3684 => x"10",
          3685 => x"05",
          3686 => x"41",
          3687 => x"ad",
          3688 => x"b4",
          3689 => x"80",
          3690 => x"83",
          3691 => x"58",
          3692 => x"8b",
          3693 => x"0b",
          3694 => x"34",
          3695 => x"d1",
          3696 => x"84",
          3697 => x"b4",
          3698 => x"84",
          3699 => x"55",
          3700 => x"b6",
          3701 => x"ac",
          3702 => x"51",
          3703 => x"3f",
          3704 => x"08",
          3705 => x"ff",
          3706 => x"84",
          3707 => x"52",
          3708 => x"ae",
          3709 => x"d1",
          3710 => x"05",
          3711 => x"d1",
          3712 => x"81",
          3713 => x"74",
          3714 => x"d1",
          3715 => x"9f",
          3716 => x"0b",
          3717 => x"34",
          3718 => x"d1",
          3719 => x"be",
          3720 => x"34",
          3721 => x"1d",
          3722 => x"8c",
          3723 => x"80",
          3724 => x"84",
          3725 => x"52",
          3726 => x"ae",
          3727 => x"d5",
          3728 => x"a0",
          3729 => x"a6",
          3730 => x"ac",
          3731 => x"51",
          3732 => x"3f",
          3733 => x"33",
          3734 => x"7c",
          3735 => x"34",
          3736 => x"06",
          3737 => x"38",
          3738 => x"51",
          3739 => x"3f",
          3740 => x"d1",
          3741 => x"0b",
          3742 => x"34",
          3743 => x"c8",
          3744 => x"0d",
          3745 => x"8c",
          3746 => x"ff",
          3747 => x"7a",
          3748 => x"ca",
          3749 => x"88",
          3750 => x"59",
          3751 => x"88",
          3752 => x"58",
          3753 => x"8c",
          3754 => x"ac",
          3755 => x"51",
          3756 => x"3f",
          3757 => x"33",
          3758 => x"70",
          3759 => x"d1",
          3760 => x"52",
          3761 => x"76",
          3762 => x"38",
          3763 => x"08",
          3764 => x"ff",
          3765 => x"84",
          3766 => x"70",
          3767 => x"98",
          3768 => x"88",
          3769 => x"59",
          3770 => x"24",
          3771 => x"84",
          3772 => x"52",
          3773 => x"ac",
          3774 => x"81",
          3775 => x"81",
          3776 => x"70",
          3777 => x"d1",
          3778 => x"51",
          3779 => x"24",
          3780 => x"84",
          3781 => x"52",
          3782 => x"ac",
          3783 => x"81",
          3784 => x"81",
          3785 => x"70",
          3786 => x"d1",
          3787 => x"51",
          3788 => x"25",
          3789 => x"f3",
          3790 => x"16",
          3791 => x"33",
          3792 => x"d5",
          3793 => x"76",
          3794 => x"ac",
          3795 => x"81",
          3796 => x"81",
          3797 => x"70",
          3798 => x"d1",
          3799 => x"57",
          3800 => x"25",
          3801 => x"7b",
          3802 => x"17",
          3803 => x"84",
          3804 => x"52",
          3805 => x"ff",
          3806 => x"75",
          3807 => x"29",
          3808 => x"05",
          3809 => x"84",
          3810 => x"43",
          3811 => x"76",
          3812 => x"38",
          3813 => x"84",
          3814 => x"70",
          3815 => x"58",
          3816 => x"2e",
          3817 => x"84",
          3818 => x"55",
          3819 => x"ae",
          3820 => x"2b",
          3821 => x"57",
          3822 => x"24",
          3823 => x"16",
          3824 => x"81",
          3825 => x"81",
          3826 => x"81",
          3827 => x"70",
          3828 => x"d1",
          3829 => x"57",
          3830 => x"25",
          3831 => x"18",
          3832 => x"d1",
          3833 => x"81",
          3834 => x"05",
          3835 => x"33",
          3836 => x"d1",
          3837 => x"76",
          3838 => x"38",
          3839 => x"75",
          3840 => x"34",
          3841 => x"d1",
          3842 => x"81",
          3843 => x"81",
          3844 => x"70",
          3845 => x"81",
          3846 => x"58",
          3847 => x"76",
          3848 => x"38",
          3849 => x"70",
          3850 => x"81",
          3851 => x"57",
          3852 => x"25",
          3853 => x"84",
          3854 => x"52",
          3855 => x"aa",
          3856 => x"81",
          3857 => x"81",
          3858 => x"70",
          3859 => x"d1",
          3860 => x"57",
          3861 => x"25",
          3862 => x"84",
          3863 => x"52",
          3864 => x"aa",
          3865 => x"81",
          3866 => x"81",
          3867 => x"70",
          3868 => x"d1",
          3869 => x"57",
          3870 => x"24",
          3871 => x"f0",
          3872 => x"f2",
          3873 => x"75",
          3874 => x"9d",
          3875 => x"ff",
          3876 => x"84",
          3877 => x"84",
          3878 => x"84",
          3879 => x"81",
          3880 => x"05",
          3881 => x"7b",
          3882 => x"be",
          3883 => x"88",
          3884 => x"8c",
          3885 => x"74",
          3886 => x"c8",
          3887 => x"ac",
          3888 => x"51",
          3889 => x"3f",
          3890 => x"08",
          3891 => x"ff",
          3892 => x"84",
          3893 => x"52",
          3894 => x"a9",
          3895 => x"d1",
          3896 => x"05",
          3897 => x"d1",
          3898 => x"81",
          3899 => x"c7",
          3900 => x"80",
          3901 => x"84",
          3902 => x"83",
          3903 => x"84",
          3904 => x"85",
          3905 => x"83",
          3906 => x"77",
          3907 => x"80",
          3908 => x"d5",
          3909 => x"7b",
          3910 => x"52",
          3911 => x"ce",
          3912 => x"80",
          3913 => x"80",
          3914 => x"98",
          3915 => x"88",
          3916 => x"57",
          3917 => x"da",
          3918 => x"8c",
          3919 => x"2b",
          3920 => x"79",
          3921 => x"5d",
          3922 => x"75",
          3923 => x"8e",
          3924 => x"39",
          3925 => x"08",
          3926 => x"fc",
          3927 => x"e0",
          3928 => x"76",
          3929 => x"bb",
          3930 => x"84",
          3931 => x"75",
          3932 => x"38",
          3933 => x"f3",
          3934 => x"f3",
          3935 => x"74",
          3936 => x"d4",
          3937 => x"81",
          3938 => x"83",
          3939 => x"51",
          3940 => x"3f",
          3941 => x"f3",
          3942 => x"3d",
          3943 => x"5f",
          3944 => x"74",
          3945 => x"e9",
          3946 => x"0c",
          3947 => x"18",
          3948 => x"80",
          3949 => x"38",
          3950 => x"75",
          3951 => x"e8",
          3952 => x"c8",
          3953 => x"88",
          3954 => x"c8",
          3955 => x"06",
          3956 => x"75",
          3957 => x"ff",
          3958 => x"93",
          3959 => x"88",
          3960 => x"8c",
          3961 => x"5d",
          3962 => x"f2",
          3963 => x"d5",
          3964 => x"88",
          3965 => x"f6",
          3966 => x"ac",
          3967 => x"51",
          3968 => x"3f",
          3969 => x"08",
          3970 => x"ff",
          3971 => x"84",
          3972 => x"ff",
          3973 => x"84",
          3974 => x"79",
          3975 => x"55",
          3976 => x"7c",
          3977 => x"84",
          3978 => x"80",
          3979 => x"88",
          3980 => x"b9",
          3981 => x"3d",
          3982 => x"51",
          3983 => x"3f",
          3984 => x"08",
          3985 => x"34",
          3986 => x"08",
          3987 => x"81",
          3988 => x"52",
          3989 => x"aa",
          3990 => x"1d",
          3991 => x"06",
          3992 => x"33",
          3993 => x"33",
          3994 => x"56",
          3995 => x"f1",
          3996 => x"d5",
          3997 => x"88",
          3998 => x"f2",
          3999 => x"ac",
          4000 => x"51",
          4001 => x"3f",
          4002 => x"08",
          4003 => x"ff",
          4004 => x"84",
          4005 => x"ff",
          4006 => x"84",
          4007 => x"76",
          4008 => x"55",
          4009 => x"51",
          4010 => x"3f",
          4011 => x"08",
          4012 => x"34",
          4013 => x"08",
          4014 => x"81",
          4015 => x"52",
          4016 => x"a9",
          4017 => x"1d",
          4018 => x"06",
          4019 => x"33",
          4020 => x"33",
          4021 => x"58",
          4022 => x"f0",
          4023 => x"d5",
          4024 => x"88",
          4025 => x"86",
          4026 => x"ac",
          4027 => x"51",
          4028 => x"3f",
          4029 => x"08",
          4030 => x"ff",
          4031 => x"84",
          4032 => x"ff",
          4033 => x"84",
          4034 => x"60",
          4035 => x"55",
          4036 => x"51",
          4037 => x"3f",
          4038 => x"33",
          4039 => x"87",
          4040 => x"f2",
          4041 => x"19",
          4042 => x"5c",
          4043 => x"d1",
          4044 => x"c8",
          4045 => x"83",
          4046 => x"70",
          4047 => x"f2",
          4048 => x"08",
          4049 => x"74",
          4050 => x"d5",
          4051 => x"7b",
          4052 => x"ff",
          4053 => x"83",
          4054 => x"81",
          4055 => x"ff",
          4056 => x"93",
          4057 => x"f2",
          4058 => x"f3",
          4059 => x"b1",
          4060 => x"fe",
          4061 => x"76",
          4062 => x"75",
          4063 => x"c0",
          4064 => x"b4",
          4065 => x"51",
          4066 => x"3f",
          4067 => x"08",
          4068 => x"f3",
          4069 => x"84",
          4070 => x"80",
          4071 => x"88",
          4072 => x"b9",
          4073 => x"3d",
          4074 => x"53",
          4075 => x"b9",
          4076 => x"81",
          4077 => x"84",
          4078 => x"82",
          4079 => x"b9",
          4080 => x"3d",
          4081 => x"f3",
          4082 => x"80",
          4083 => x"51",
          4084 => x"3f",
          4085 => x"08",
          4086 => x"c8",
          4087 => x"09",
          4088 => x"ee",
          4089 => x"c8",
          4090 => x"a6",
          4091 => x"b9",
          4092 => x"80",
          4093 => x"c8",
          4094 => x"e3",
          4095 => x"c8",
          4096 => x"70",
          4097 => x"80",
          4098 => x"81",
          4099 => x"f3",
          4100 => x"10",
          4101 => x"e0",
          4102 => x"58",
          4103 => x"74",
          4104 => x"76",
          4105 => x"fc",
          4106 => x"e0",
          4107 => x"70",
          4108 => x"80",
          4109 => x"84",
          4110 => x"75",
          4111 => x"b8",
          4112 => x"10",
          4113 => x"05",
          4114 => x"40",
          4115 => x"38",
          4116 => x"81",
          4117 => x"57",
          4118 => x"83",
          4119 => x"75",
          4120 => x"81",
          4121 => x"38",
          4122 => x"38",
          4123 => x"76",
          4124 => x"74",
          4125 => x"f2",
          4126 => x"b8",
          4127 => x"70",
          4128 => x"5b",
          4129 => x"27",
          4130 => x"80",
          4131 => x"b8",
          4132 => x"39",
          4133 => x"d3",
          4134 => x"f3",
          4135 => x"82",
          4136 => x"06",
          4137 => x"05",
          4138 => x"54",
          4139 => x"80",
          4140 => x"84",
          4141 => x"75",
          4142 => x"b8",
          4143 => x"10",
          4144 => x"05",
          4145 => x"40",
          4146 => x"2e",
          4147 => x"ff",
          4148 => x"83",
          4149 => x"fe",
          4150 => x"83",
          4151 => x"f1",
          4152 => x"e1",
          4153 => x"9f",
          4154 => x"e7",
          4155 => x"e4",
          4156 => x"0d",
          4157 => x"05",
          4158 => x"05",
          4159 => x"33",
          4160 => x"83",
          4161 => x"38",
          4162 => x"81",
          4163 => x"73",
          4164 => x"38",
          4165 => x"82",
          4166 => x"a7",
          4167 => x"86",
          4168 => x"70",
          4169 => x"56",
          4170 => x"79",
          4171 => x"38",
          4172 => x"f8",
          4173 => x"f8",
          4174 => x"83",
          4175 => x"83",
          4176 => x"70",
          4177 => x"90",
          4178 => x"88",
          4179 => x"07",
          4180 => x"56",
          4181 => x"77",
          4182 => x"80",
          4183 => x"05",
          4184 => x"73",
          4185 => x"55",
          4186 => x"26",
          4187 => x"78",
          4188 => x"83",
          4189 => x"84",
          4190 => x"79",
          4191 => x"55",
          4192 => x"e0",
          4193 => x"74",
          4194 => x"05",
          4195 => x"13",
          4196 => x"38",
          4197 => x"04",
          4198 => x"80",
          4199 => x"f8",
          4200 => x"10",
          4201 => x"f9",
          4202 => x"29",
          4203 => x"5b",
          4204 => x"59",
          4205 => x"80",
          4206 => x"bc",
          4207 => x"ff",
          4208 => x"bb",
          4209 => x"ff",
          4210 => x"f6",
          4211 => x"ff",
          4212 => x"75",
          4213 => x"5d",
          4214 => x"5b",
          4215 => x"26",
          4216 => x"74",
          4217 => x"56",
          4218 => x"06",
          4219 => x"06",
          4220 => x"06",
          4221 => x"ff",
          4222 => x"ff",
          4223 => x"29",
          4224 => x"57",
          4225 => x"74",
          4226 => x"38",
          4227 => x"33",
          4228 => x"05",
          4229 => x"1b",
          4230 => x"83",
          4231 => x"80",
          4232 => x"38",
          4233 => x"53",
          4234 => x"fe",
          4235 => x"73",
          4236 => x"55",
          4237 => x"f4",
          4238 => x"81",
          4239 => x"e8",
          4240 => x"a0",
          4241 => x"a7",
          4242 => x"84",
          4243 => x"70",
          4244 => x"84",
          4245 => x"70",
          4246 => x"83",
          4247 => x"70",
          4248 => x"5b",
          4249 => x"56",
          4250 => x"78",
          4251 => x"38",
          4252 => x"06",
          4253 => x"06",
          4254 => x"18",
          4255 => x"79",
          4256 => x"bb",
          4257 => x"83",
          4258 => x"80",
          4259 => x"f9",
          4260 => x"f4",
          4261 => x"2b",
          4262 => x"07",
          4263 => x"07",
          4264 => x"7f",
          4265 => x"5b",
          4266 => x"fd",
          4267 => x"be",
          4268 => x"e6",
          4269 => x"f8",
          4270 => x"ff",
          4271 => x"10",
          4272 => x"f9",
          4273 => x"29",
          4274 => x"a0",
          4275 => x"57",
          4276 => x"5f",
          4277 => x"80",
          4278 => x"b7",
          4279 => x"81",
          4280 => x"b7",
          4281 => x"81",
          4282 => x"f8",
          4283 => x"83",
          4284 => x"7c",
          4285 => x"05",
          4286 => x"5f",
          4287 => x"5e",
          4288 => x"26",
          4289 => x"7a",
          4290 => x"7d",
          4291 => x"53",
          4292 => x"06",
          4293 => x"06",
          4294 => x"7d",
          4295 => x"06",
          4296 => x"06",
          4297 => x"58",
          4298 => x"5d",
          4299 => x"26",
          4300 => x"75",
          4301 => x"73",
          4302 => x"83",
          4303 => x"79",
          4304 => x"76",
          4305 => x"7b",
          4306 => x"fb",
          4307 => x"78",
          4308 => x"56",
          4309 => x"fb",
          4310 => x"8e",
          4311 => x"ff",
          4312 => x"87",
          4313 => x"73",
          4314 => x"34",
          4315 => x"9c",
          4316 => x"75",
          4317 => x"75",
          4318 => x"80",
          4319 => x"76",
          4320 => x"34",
          4321 => x"94",
          4322 => x"34",
          4323 => x"ff",
          4324 => x"81",
          4325 => x"fa",
          4326 => x"a0",
          4327 => x"08",
          4328 => x"f8",
          4329 => x"81",
          4330 => x"06",
          4331 => x"55",
          4332 => x"73",
          4333 => x"ff",
          4334 => x"07",
          4335 => x"75",
          4336 => x"87",
          4337 => x"77",
          4338 => x"51",
          4339 => x"a0",
          4340 => x"73",
          4341 => x"06",
          4342 => x"72",
          4343 => x"d0",
          4344 => x"bc",
          4345 => x"84",
          4346 => x"87",
          4347 => x"84",
          4348 => x"84",
          4349 => x"04",
          4350 => x"02",
          4351 => x"02",
          4352 => x"05",
          4353 => x"bb",
          4354 => x"56",
          4355 => x"79",
          4356 => x"38",
          4357 => x"33",
          4358 => x"33",
          4359 => x"33",
          4360 => x"12",
          4361 => x"80",
          4362 => x"f6",
          4363 => x"57",
          4364 => x"29",
          4365 => x"ff",
          4366 => x"f7",
          4367 => x"57",
          4368 => x"81",
          4369 => x"38",
          4370 => x"22",
          4371 => x"74",
          4372 => x"23",
          4373 => x"33",
          4374 => x"81",
          4375 => x"81",
          4376 => x"5b",
          4377 => x"26",
          4378 => x"ff",
          4379 => x"83",
          4380 => x"83",
          4381 => x"70",
          4382 => x"06",
          4383 => x"33",
          4384 => x"79",
          4385 => x"89",
          4386 => x"bc",
          4387 => x"29",
          4388 => x"54",
          4389 => x"26",
          4390 => x"98",
          4391 => x"54",
          4392 => x"13",
          4393 => x"16",
          4394 => x"81",
          4395 => x"75",
          4396 => x"57",
          4397 => x"54",
          4398 => x"73",
          4399 => x"73",
          4400 => x"a1",
          4401 => x"f4",
          4402 => x"9a",
          4403 => x"a0",
          4404 => x"14",
          4405 => x"70",
          4406 => x"34",
          4407 => x"9f",
          4408 => x"eb",
          4409 => x"ba",
          4410 => x"56",
          4411 => x"f6",
          4412 => x"78",
          4413 => x"77",
          4414 => x"06",
          4415 => x"73",
          4416 => x"38",
          4417 => x"81",
          4418 => x"bc",
          4419 => x"29",
          4420 => x"75",
          4421 => x"a0",
          4422 => x"a7",
          4423 => x"81",
          4424 => x"81",
          4425 => x"71",
          4426 => x"5c",
          4427 => x"79",
          4428 => x"84",
          4429 => x"54",
          4430 => x"33",
          4431 => x"c4",
          4432 => x"70",
          4433 => x"34",
          4434 => x"05",
          4435 => x"70",
          4436 => x"34",
          4437 => x"b7",
          4438 => x"b7",
          4439 => x"71",
          4440 => x"5c",
          4441 => x"75",
          4442 => x"80",
          4443 => x"b9",
          4444 => x"3d",
          4445 => x"83",
          4446 => x"83",
          4447 => x"70",
          4448 => x"06",
          4449 => x"33",
          4450 => x"73",
          4451 => x"f9",
          4452 => x"2e",
          4453 => x"78",
          4454 => x"ff",
          4455 => x"f8",
          4456 => x"72",
          4457 => x"81",
          4458 => x"38",
          4459 => x"81",
          4460 => x"bc",
          4461 => x"29",
          4462 => x"11",
          4463 => x"54",
          4464 => x"fe",
          4465 => x"f8",
          4466 => x"98",
          4467 => x"76",
          4468 => x"56",
          4469 => x"e0",
          4470 => x"75",
          4471 => x"57",
          4472 => x"53",
          4473 => x"fe",
          4474 => x"0b",
          4475 => x"34",
          4476 => x"81",
          4477 => x"ff",
          4478 => x"d8",
          4479 => x"39",
          4480 => x"b7",
          4481 => x"56",
          4482 => x"83",
          4483 => x"33",
          4484 => x"c4",
          4485 => x"34",
          4486 => x"33",
          4487 => x"39",
          4488 => x"76",
          4489 => x"9f",
          4490 => x"51",
          4491 => x"9b",
          4492 => x"10",
          4493 => x"05",
          4494 => x"04",
          4495 => x"33",
          4496 => x"27",
          4497 => x"83",
          4498 => x"80",
          4499 => x"c8",
          4500 => x"0d",
          4501 => x"83",
          4502 => x"83",
          4503 => x"70",
          4504 => x"54",
          4505 => x"2e",
          4506 => x"12",
          4507 => x"f8",
          4508 => x"0b",
          4509 => x"0c",
          4510 => x"04",
          4511 => x"33",
          4512 => x"70",
          4513 => x"2c",
          4514 => x"55",
          4515 => x"83",
          4516 => x"de",
          4517 => x"f8",
          4518 => x"84",
          4519 => x"ff",
          4520 => x"51",
          4521 => x"83",
          4522 => x"72",
          4523 => x"34",
          4524 => x"b9",
          4525 => x"3d",
          4526 => x"f8",
          4527 => x"73",
          4528 => x"70",
          4529 => x"06",
          4530 => x"55",
          4531 => x"f9",
          4532 => x"84",
          4533 => x"86",
          4534 => x"83",
          4535 => x"72",
          4536 => x"bc",
          4537 => x"55",
          4538 => x"74",
          4539 => x"70",
          4540 => x"f8",
          4541 => x"0b",
          4542 => x"0c",
          4543 => x"04",
          4544 => x"f8",
          4545 => x"f8",
          4546 => x"b7",
          4547 => x"05",
          4548 => x"75",
          4549 => x"38",
          4550 => x"70",
          4551 => x"34",
          4552 => x"ff",
          4553 => x"8f",
          4554 => x"70",
          4555 => x"38",
          4556 => x"83",
          4557 => x"51",
          4558 => x"83",
          4559 => x"70",
          4560 => x"71",
          4561 => x"f0",
          4562 => x"84",
          4563 => x"52",
          4564 => x"80",
          4565 => x"81",
          4566 => x"80",
          4567 => x"f8",
          4568 => x"0b",
          4569 => x"0c",
          4570 => x"04",
          4571 => x"33",
          4572 => x"90",
          4573 => x"83",
          4574 => x"80",
          4575 => x"c8",
          4576 => x"0d",
          4577 => x"f4",
          4578 => x"07",
          4579 => x"f8",
          4580 => x"39",
          4581 => x"33",
          4582 => x"86",
          4583 => x"83",
          4584 => x"d7",
          4585 => x"0b",
          4586 => x"34",
          4587 => x"b9",
          4588 => x"3d",
          4589 => x"f8",
          4590 => x"fc",
          4591 => x"51",
          4592 => x"f4",
          4593 => x"39",
          4594 => x"33",
          4595 => x"70",
          4596 => x"34",
          4597 => x"83",
          4598 => x"81",
          4599 => x"07",
          4600 => x"f8",
          4601 => x"93",
          4602 => x"f4",
          4603 => x"06",
          4604 => x"70",
          4605 => x"34",
          4606 => x"83",
          4607 => x"81",
          4608 => x"07",
          4609 => x"f8",
          4610 => x"ef",
          4611 => x"f4",
          4612 => x"06",
          4613 => x"f8",
          4614 => x"df",
          4615 => x"f4",
          4616 => x"06",
          4617 => x"51",
          4618 => x"f4",
          4619 => x"39",
          4620 => x"33",
          4621 => x"b0",
          4622 => x"83",
          4623 => x"fe",
          4624 => x"f8",
          4625 => x"ef",
          4626 => x"07",
          4627 => x"f8",
          4628 => x"a7",
          4629 => x"f4",
          4630 => x"06",
          4631 => x"51",
          4632 => x"f4",
          4633 => x"39",
          4634 => x"33",
          4635 => x"a0",
          4636 => x"83",
          4637 => x"fe",
          4638 => x"f8",
          4639 => x"8f",
          4640 => x"83",
          4641 => x"fd",
          4642 => x"f8",
          4643 => x"fa",
          4644 => x"51",
          4645 => x"f4",
          4646 => x"39",
          4647 => x"02",
          4648 => x"02",
          4649 => x"c3",
          4650 => x"f8",
          4651 => x"f8",
          4652 => x"f8",
          4653 => x"b7",
          4654 => x"41",
          4655 => x"59",
          4656 => x"82",
          4657 => x"82",
          4658 => x"78",
          4659 => x"82",
          4660 => x"b7",
          4661 => x"0b",
          4662 => x"34",
          4663 => x"f8",
          4664 => x"f8",
          4665 => x"83",
          4666 => x"8f",
          4667 => x"78",
          4668 => x"81",
          4669 => x"80",
          4670 => x"be",
          4671 => x"84",
          4672 => x"82",
          4673 => x"f8",
          4674 => x"83",
          4675 => x"82",
          4676 => x"f6",
          4677 => x"84",
          4678 => x"57",
          4679 => x"33",
          4680 => x"ba",
          4681 => x"54",
          4682 => x"52",
          4683 => x"51",
          4684 => x"3f",
          4685 => x"be",
          4686 => x"84",
          4687 => x"7a",
          4688 => x"34",
          4689 => x"f6",
          4690 => x"f8",
          4691 => x"3d",
          4692 => x"0b",
          4693 => x"34",
          4694 => x"b7",
          4695 => x"0b",
          4696 => x"34",
          4697 => x"f8",
          4698 => x"0b",
          4699 => x"23",
          4700 => x"33",
          4701 => x"ca",
          4702 => x"b8",
          4703 => x"79",
          4704 => x"7c",
          4705 => x"83",
          4706 => x"ff",
          4707 => x"80",
          4708 => x"c9",
          4709 => x"79",
          4710 => x"38",
          4711 => x"b9",
          4712 => x"22",
          4713 => x"e3",
          4714 => x"80",
          4715 => x"1a",
          4716 => x"06",
          4717 => x"33",
          4718 => x"78",
          4719 => x"38",
          4720 => x"51",
          4721 => x"3f",
          4722 => x"be",
          4723 => x"84",
          4724 => x"7a",
          4725 => x"34",
          4726 => x"f6",
          4727 => x"f8",
          4728 => x"3d",
          4729 => x"0b",
          4730 => x"34",
          4731 => x"b7",
          4732 => x"0b",
          4733 => x"34",
          4734 => x"f8",
          4735 => x"0b",
          4736 => x"23",
          4737 => x"51",
          4738 => x"3f",
          4739 => x"08",
          4740 => x"f4",
          4741 => x"f0",
          4742 => x"83",
          4743 => x"ff",
          4744 => x"78",
          4745 => x"08",
          4746 => x"38",
          4747 => x"19",
          4748 => x"e3",
          4749 => x"ff",
          4750 => x"19",
          4751 => x"06",
          4752 => x"39",
          4753 => x"7a",
          4754 => x"a7",
          4755 => x"b7",
          4756 => x"f8",
          4757 => x"f8",
          4758 => x"71",
          4759 => x"a7",
          4760 => x"83",
          4761 => x"53",
          4762 => x"71",
          4763 => x"70",
          4764 => x"06",
          4765 => x"33",
          4766 => x"55",
          4767 => x"81",
          4768 => x"38",
          4769 => x"81",
          4770 => x"89",
          4771 => x"38",
          4772 => x"83",
          4773 => x"88",
          4774 => x"38",
          4775 => x"33",
          4776 => x"33",
          4777 => x"33",
          4778 => x"05",
          4779 => x"84",
          4780 => x"33",
          4781 => x"80",
          4782 => x"b7",
          4783 => x"f8",
          4784 => x"f8",
          4785 => x"71",
          4786 => x"5a",
          4787 => x"83",
          4788 => x"34",
          4789 => x"33",
          4790 => x"16",
          4791 => x"f8",
          4792 => x"a7",
          4793 => x"34",
          4794 => x"33",
          4795 => x"06",
          4796 => x"22",
          4797 => x"33",
          4798 => x"11",
          4799 => x"55",
          4800 => x"f4",
          4801 => x"9a",
          4802 => x"18",
          4803 => x"06",
          4804 => x"78",
          4805 => x"38",
          4806 => x"33",
          4807 => x"ea",
          4808 => x"53",
          4809 => x"f9",
          4810 => x"bf",
          4811 => x"80",
          4812 => x"84",
          4813 => x"57",
          4814 => x"80",
          4815 => x"0b",
          4816 => x"0c",
          4817 => x"04",
          4818 => x"97",
          4819 => x"24",
          4820 => x"75",
          4821 => x"81",
          4822 => x"38",
          4823 => x"51",
          4824 => x"80",
          4825 => x"f9",
          4826 => x"39",
          4827 => x"15",
          4828 => x"b7",
          4829 => x"74",
          4830 => x"2e",
          4831 => x"fe",
          4832 => x"53",
          4833 => x"51",
          4834 => x"81",
          4835 => x"ff",
          4836 => x"72",
          4837 => x"91",
          4838 => x"a0",
          4839 => x"3f",
          4840 => x"81",
          4841 => x"54",
          4842 => x"d8",
          4843 => x"39",
          4844 => x"f9",
          4845 => x"39",
          4846 => x"51",
          4847 => x"80",
          4848 => x"c8",
          4849 => x"0d",
          4850 => x"ff",
          4851 => x"06",
          4852 => x"83",
          4853 => x"70",
          4854 => x"55",
          4855 => x"73",
          4856 => x"53",
          4857 => x"f9",
          4858 => x"a0",
          4859 => x"3f",
          4860 => x"33",
          4861 => x"06",
          4862 => x"53",
          4863 => x"38",
          4864 => x"83",
          4865 => x"fe",
          4866 => x"0b",
          4867 => x"34",
          4868 => x"51",
          4869 => x"fe",
          4870 => x"52",
          4871 => x"d8",
          4872 => x"39",
          4873 => x"02",
          4874 => x"33",
          4875 => x"08",
          4876 => x"81",
          4877 => x"38",
          4878 => x"83",
          4879 => x"8a",
          4880 => x"38",
          4881 => x"82",
          4882 => x"88",
          4883 => x"38",
          4884 => x"88",
          4885 => x"b7",
          4886 => x"f8",
          4887 => x"f8",
          4888 => x"72",
          4889 => x"5e",
          4890 => x"c4",
          4891 => x"a7",
          4892 => x"34",
          4893 => x"33",
          4894 => x"33",
          4895 => x"22",
          4896 => x"12",
          4897 => x"40",
          4898 => x"fa",
          4899 => x"f8",
          4900 => x"71",
          4901 => x"40",
          4902 => x"f4",
          4903 => x"a7",
          4904 => x"34",
          4905 => x"33",
          4906 => x"06",
          4907 => x"22",
          4908 => x"33",
          4909 => x"11",
          4910 => x"58",
          4911 => x"f4",
          4912 => x"9a",
          4913 => x"1d",
          4914 => x"06",
          4915 => x"61",
          4916 => x"38",
          4917 => x"33",
          4918 => x"f1",
          4919 => x"56",
          4920 => x"f9",
          4921 => x"84",
          4922 => x"9c",
          4923 => x"78",
          4924 => x"8a",
          4925 => x"25",
          4926 => x"78",
          4927 => x"b3",
          4928 => x"db",
          4929 => x"38",
          4930 => x"b8",
          4931 => x"b7",
          4932 => x"f8",
          4933 => x"f8",
          4934 => x"72",
          4935 => x"40",
          4936 => x"c4",
          4937 => x"a7",
          4938 => x"34",
          4939 => x"33",
          4940 => x"33",
          4941 => x"22",
          4942 => x"12",
          4943 => x"56",
          4944 => x"fa",
          4945 => x"f8",
          4946 => x"71",
          4947 => x"57",
          4948 => x"33",
          4949 => x"80",
          4950 => x"b7",
          4951 => x"81",
          4952 => x"f8",
          4953 => x"f8",
          4954 => x"72",
          4955 => x"42",
          4956 => x"83",
          4957 => x"60",
          4958 => x"05",
          4959 => x"58",
          4960 => x"06",
          4961 => x"27",
          4962 => x"77",
          4963 => x"34",
          4964 => x"b9",
          4965 => x"3d",
          4966 => x"9b",
          4967 => x"38",
          4968 => x"83",
          4969 => x"8d",
          4970 => x"06",
          4971 => x"80",
          4972 => x"f9",
          4973 => x"84",
          4974 => x"9c",
          4975 => x"78",
          4976 => x"aa",
          4977 => x"56",
          4978 => x"84",
          4979 => x"b8",
          4980 => x"11",
          4981 => x"84",
          4982 => x"78",
          4983 => x"18",
          4984 => x"ff",
          4985 => x"0b",
          4986 => x"1a",
          4987 => x"84",
          4988 => x"9c",
          4989 => x"78",
          4990 => x"e9",
          4991 => x"84",
          4992 => x"84",
          4993 => x"83",
          4994 => x"83",
          4995 => x"72",
          4996 => x"5e",
          4997 => x"b7",
          4998 => x"86",
          4999 => x"1d",
          5000 => x"bc",
          5001 => x"f9",
          5002 => x"f6",
          5003 => x"29",
          5004 => x"59",
          5005 => x"f8",
          5006 => x"83",
          5007 => x"76",
          5008 => x"5b",
          5009 => x"f4",
          5010 => x"b0",
          5011 => x"84",
          5012 => x"70",
          5013 => x"83",
          5014 => x"83",
          5015 => x"72",
          5016 => x"44",
          5017 => x"59",
          5018 => x"33",
          5019 => x"9a",
          5020 => x"1f",
          5021 => x"39",
          5022 => x"51",
          5023 => x"80",
          5024 => x"f9",
          5025 => x"39",
          5026 => x"33",
          5027 => x"33",
          5028 => x"06",
          5029 => x"33",
          5030 => x"12",
          5031 => x"80",
          5032 => x"f6",
          5033 => x"5d",
          5034 => x"05",
          5035 => x"ff",
          5036 => x"ce",
          5037 => x"59",
          5038 => x"81",
          5039 => x"38",
          5040 => x"06",
          5041 => x"57",
          5042 => x"38",
          5043 => x"83",
          5044 => x"fc",
          5045 => x"0b",
          5046 => x"34",
          5047 => x"b8",
          5048 => x"0b",
          5049 => x"34",
          5050 => x"b8",
          5051 => x"0b",
          5052 => x"0c",
          5053 => x"b9",
          5054 => x"3d",
          5055 => x"f8",
          5056 => x"b9",
          5057 => x"f8",
          5058 => x"b9",
          5059 => x"f8",
          5060 => x"b9",
          5061 => x"0b",
          5062 => x"0c",
          5063 => x"b9",
          5064 => x"3d",
          5065 => x"80",
          5066 => x"81",
          5067 => x"38",
          5068 => x"33",
          5069 => x"33",
          5070 => x"06",
          5071 => x"33",
          5072 => x"06",
          5073 => x"11",
          5074 => x"80",
          5075 => x"f6",
          5076 => x"72",
          5077 => x"70",
          5078 => x"06",
          5079 => x"33",
          5080 => x"5c",
          5081 => x"7d",
          5082 => x"fe",
          5083 => x"ff",
          5084 => x"58",
          5085 => x"38",
          5086 => x"83",
          5087 => x"7b",
          5088 => x"7a",
          5089 => x"78",
          5090 => x"72",
          5091 => x"5f",
          5092 => x"b7",
          5093 => x"a7",
          5094 => x"34",
          5095 => x"33",
          5096 => x"33",
          5097 => x"22",
          5098 => x"12",
          5099 => x"40",
          5100 => x"f8",
          5101 => x"83",
          5102 => x"60",
          5103 => x"05",
          5104 => x"f8",
          5105 => x"a7",
          5106 => x"34",
          5107 => x"33",
          5108 => x"06",
          5109 => x"22",
          5110 => x"33",
          5111 => x"11",
          5112 => x"5e",
          5113 => x"f4",
          5114 => x"98",
          5115 => x"81",
          5116 => x"ff",
          5117 => x"7c",
          5118 => x"ea",
          5119 => x"bd",
          5120 => x"96",
          5121 => x"19",
          5122 => x"f8",
          5123 => x"f8",
          5124 => x"81",
          5125 => x"ff",
          5126 => x"ac",
          5127 => x"2e",
          5128 => x"78",
          5129 => x"d7",
          5130 => x"2e",
          5131 => x"84",
          5132 => x"5f",
          5133 => x"38",
          5134 => x"56",
          5135 => x"84",
          5136 => x"10",
          5137 => x"d0",
          5138 => x"08",
          5139 => x"83",
          5140 => x"80",
          5141 => x"e7",
          5142 => x"0b",
          5143 => x"0c",
          5144 => x"04",
          5145 => x"33",
          5146 => x"33",
          5147 => x"06",
          5148 => x"33",
          5149 => x"06",
          5150 => x"11",
          5151 => x"80",
          5152 => x"f6",
          5153 => x"72",
          5154 => x"70",
          5155 => x"06",
          5156 => x"33",
          5157 => x"5c",
          5158 => x"7f",
          5159 => x"ef",
          5160 => x"7a",
          5161 => x"7a",
          5162 => x"7a",
          5163 => x"72",
          5164 => x"5c",
          5165 => x"b7",
          5166 => x"a7",
          5167 => x"34",
          5168 => x"33",
          5169 => x"33",
          5170 => x"22",
          5171 => x"12",
          5172 => x"56",
          5173 => x"f8",
          5174 => x"83",
          5175 => x"76",
          5176 => x"5a",
          5177 => x"f4",
          5178 => x"b0",
          5179 => x"84",
          5180 => x"70",
          5181 => x"83",
          5182 => x"83",
          5183 => x"72",
          5184 => x"5b",
          5185 => x"59",
          5186 => x"33",
          5187 => x"18",
          5188 => x"05",
          5189 => x"06",
          5190 => x"7a",
          5191 => x"38",
          5192 => x"33",
          5193 => x"fb",
          5194 => x"56",
          5195 => x"f9",
          5196 => x"70",
          5197 => x"5d",
          5198 => x"26",
          5199 => x"83",
          5200 => x"84",
          5201 => x"83",
          5202 => x"72",
          5203 => x"72",
          5204 => x"72",
          5205 => x"72",
          5206 => x"54",
          5207 => x"5b",
          5208 => x"e4",
          5209 => x"a0",
          5210 => x"84",
          5211 => x"83",
          5212 => x"83",
          5213 => x"72",
          5214 => x"5e",
          5215 => x"a0",
          5216 => x"fa",
          5217 => x"f8",
          5218 => x"71",
          5219 => x"5e",
          5220 => x"33",
          5221 => x"80",
          5222 => x"b7",
          5223 => x"81",
          5224 => x"f8",
          5225 => x"f8",
          5226 => x"72",
          5227 => x"44",
          5228 => x"83",
          5229 => x"84",
          5230 => x"34",
          5231 => x"70",
          5232 => x"5b",
          5233 => x"27",
          5234 => x"77",
          5235 => x"34",
          5236 => x"82",
          5237 => x"c4",
          5238 => x"84",
          5239 => x"9c",
          5240 => x"83",
          5241 => x"33",
          5242 => x"c4",
          5243 => x"34",
          5244 => x"33",
          5245 => x"06",
          5246 => x"56",
          5247 => x"81",
          5248 => x"ca",
          5249 => x"84",
          5250 => x"9c",
          5251 => x"83",
          5252 => x"33",
          5253 => x"c4",
          5254 => x"34",
          5255 => x"33",
          5256 => x"33",
          5257 => x"33",
          5258 => x"80",
          5259 => x"39",
          5260 => x"42",
          5261 => x"11",
          5262 => x"51",
          5263 => x"3f",
          5264 => x"08",
          5265 => x"f0",
          5266 => x"c9",
          5267 => x"57",
          5268 => x"b8",
          5269 => x"10",
          5270 => x"41",
          5271 => x"05",
          5272 => x"b9",
          5273 => x"fb",
          5274 => x"f8",
          5275 => x"5c",
          5276 => x"1c",
          5277 => x"83",
          5278 => x"84",
          5279 => x"83",
          5280 => x"5b",
          5281 => x"e5",
          5282 => x"bc",
          5283 => x"f8",
          5284 => x"f9",
          5285 => x"29",
          5286 => x"5b",
          5287 => x"19",
          5288 => x"a7",
          5289 => x"34",
          5290 => x"33",
          5291 => x"33",
          5292 => x"22",
          5293 => x"12",
          5294 => x"56",
          5295 => x"fa",
          5296 => x"f8",
          5297 => x"71",
          5298 => x"5e",
          5299 => x"33",
          5300 => x"b0",
          5301 => x"84",
          5302 => x"70",
          5303 => x"83",
          5304 => x"83",
          5305 => x"72",
          5306 => x"41",
          5307 => x"5a",
          5308 => x"33",
          5309 => x"1e",
          5310 => x"70",
          5311 => x"5c",
          5312 => x"26",
          5313 => x"84",
          5314 => x"58",
          5315 => x"38",
          5316 => x"75",
          5317 => x"34",
          5318 => x"b8",
          5319 => x"b7",
          5320 => x"7f",
          5321 => x"bd",
          5322 => x"c0",
          5323 => x"f3",
          5324 => x"52",
          5325 => x"e4",
          5326 => x"84",
          5327 => x"9c",
          5328 => x"84",
          5329 => x"83",
          5330 => x"84",
          5331 => x"83",
          5332 => x"84",
          5333 => x"57",
          5334 => x"f6",
          5335 => x"39",
          5336 => x"33",
          5337 => x"34",
          5338 => x"33",
          5339 => x"34",
          5340 => x"33",
          5341 => x"34",
          5342 => x"84",
          5343 => x"5b",
          5344 => x"ff",
          5345 => x"b9",
          5346 => x"7c",
          5347 => x"81",
          5348 => x"38",
          5349 => x"33",
          5350 => x"83",
          5351 => x"81",
          5352 => x"53",
          5353 => x"52",
          5354 => x"52",
          5355 => x"f8",
          5356 => x"fe",
          5357 => x"84",
          5358 => x"81",
          5359 => x"f7",
          5360 => x"76",
          5361 => x"a0",
          5362 => x"38",
          5363 => x"f7",
          5364 => x"fd",
          5365 => x"c0",
          5366 => x"84",
          5367 => x"5b",
          5368 => x"ff",
          5369 => x"7b",
          5370 => x"38",
          5371 => x"b9",
          5372 => x"11",
          5373 => x"75",
          5374 => x"a5",
          5375 => x"10",
          5376 => x"05",
          5377 => x"04",
          5378 => x"33",
          5379 => x"2e",
          5380 => x"83",
          5381 => x"84",
          5382 => x"71",
          5383 => x"09",
          5384 => x"72",
          5385 => x"59",
          5386 => x"83",
          5387 => x"fd",
          5388 => x"b8",
          5389 => x"75",
          5390 => x"e7",
          5391 => x"9d",
          5392 => x"70",
          5393 => x"84",
          5394 => x"5d",
          5395 => x"7b",
          5396 => x"38",
          5397 => x"f9",
          5398 => x"39",
          5399 => x"f8",
          5400 => x"f8",
          5401 => x"81",
          5402 => x"57",
          5403 => x"fd",
          5404 => x"17",
          5405 => x"f8",
          5406 => x"9c",
          5407 => x"83",
          5408 => x"83",
          5409 => x"84",
          5410 => x"ff",
          5411 => x"76",
          5412 => x"84",
          5413 => x"56",
          5414 => x"f8",
          5415 => x"39",
          5416 => x"33",
          5417 => x"2e",
          5418 => x"83",
          5419 => x"84",
          5420 => x"71",
          5421 => x"09",
          5422 => x"72",
          5423 => x"59",
          5424 => x"83",
          5425 => x"fc",
          5426 => x"b8",
          5427 => x"7a",
          5428 => x"c4",
          5429 => x"9c",
          5430 => x"99",
          5431 => x"06",
          5432 => x"84",
          5433 => x"83",
          5434 => x"83",
          5435 => x"72",
          5436 => x"86",
          5437 => x"11",
          5438 => x"22",
          5439 => x"58",
          5440 => x"05",
          5441 => x"ff",
          5442 => x"cc",
          5443 => x"fe",
          5444 => x"5a",
          5445 => x"84",
          5446 => x"92",
          5447 => x"0b",
          5448 => x"34",
          5449 => x"84",
          5450 => x"5a",
          5451 => x"fb",
          5452 => x"b9",
          5453 => x"77",
          5454 => x"81",
          5455 => x"38",
          5456 => x"f7",
          5457 => x"d0",
          5458 => x"c9",
          5459 => x"80",
          5460 => x"38",
          5461 => x"33",
          5462 => x"33",
          5463 => x"84",
          5464 => x"ff",
          5465 => x"56",
          5466 => x"83",
          5467 => x"76",
          5468 => x"34",
          5469 => x"84",
          5470 => x"57",
          5471 => x"8c",
          5472 => x"b9",
          5473 => x"f8",
          5474 => x"61",
          5475 => x"bb",
          5476 => x"59",
          5477 => x"60",
          5478 => x"75",
          5479 => x"f8",
          5480 => x"f4",
          5481 => x"90",
          5482 => x"dc",
          5483 => x"84",
          5484 => x"57",
          5485 => x"27",
          5486 => x"76",
          5487 => x"9c",
          5488 => x"53",
          5489 => x"f0",
          5490 => x"bc",
          5491 => x"70",
          5492 => x"84",
          5493 => x"58",
          5494 => x"39",
          5495 => x"b8",
          5496 => x"57",
          5497 => x"8d",
          5498 => x"9c",
          5499 => x"83",
          5500 => x"75",
          5501 => x"76",
          5502 => x"51",
          5503 => x"fa",
          5504 => x"b8",
          5505 => x"81",
          5506 => x"b7",
          5507 => x"9f",
          5508 => x"70",
          5509 => x"84",
          5510 => x"ff",
          5511 => x"ff",
          5512 => x"bb",
          5513 => x"ff",
          5514 => x"40",
          5515 => x"59",
          5516 => x"7e",
          5517 => x"77",
          5518 => x"f8",
          5519 => x"81",
          5520 => x"18",
          5521 => x"7f",
          5522 => x"77",
          5523 => x"f8",
          5524 => x"b7",
          5525 => x"11",
          5526 => x"60",
          5527 => x"38",
          5528 => x"83",
          5529 => x"f9",
          5530 => x"b8",
          5531 => x"7e",
          5532 => x"ef",
          5533 => x"9d",
          5534 => x"bb",
          5535 => x"7a",
          5536 => x"94",
          5537 => x"f8",
          5538 => x"bc",
          5539 => x"ff",
          5540 => x"f9",
          5541 => x"29",
          5542 => x"a0",
          5543 => x"f8",
          5544 => x"40",
          5545 => x"05",
          5546 => x"ff",
          5547 => x"ce",
          5548 => x"59",
          5549 => x"60",
          5550 => x"f0",
          5551 => x"ff",
          5552 => x"7c",
          5553 => x"80",
          5554 => x"fe",
          5555 => x"bb",
          5556 => x"76",
          5557 => x"38",
          5558 => x"75",
          5559 => x"23",
          5560 => x"06",
          5561 => x"41",
          5562 => x"24",
          5563 => x"84",
          5564 => x"56",
          5565 => x"8d",
          5566 => x"16",
          5567 => x"f8",
          5568 => x"81",
          5569 => x"f8",
          5570 => x"57",
          5571 => x"76",
          5572 => x"75",
          5573 => x"05",
          5574 => x"06",
          5575 => x"5c",
          5576 => x"58",
          5577 => x"80",
          5578 => x"b0",
          5579 => x"ff",
          5580 => x"ff",
          5581 => x"29",
          5582 => x"42",
          5583 => x"27",
          5584 => x"84",
          5585 => x"57",
          5586 => x"33",
          5587 => x"c4",
          5588 => x"70",
          5589 => x"34",
          5590 => x"05",
          5591 => x"70",
          5592 => x"34",
          5593 => x"b7",
          5594 => x"b7",
          5595 => x"71",
          5596 => x"40",
          5597 => x"60",
          5598 => x"38",
          5599 => x"33",
          5600 => x"c4",
          5601 => x"70",
          5602 => x"34",
          5603 => x"05",
          5604 => x"70",
          5605 => x"34",
          5606 => x"b7",
          5607 => x"b7",
          5608 => x"71",
          5609 => x"40",
          5610 => x"78",
          5611 => x"38",
          5612 => x"84",
          5613 => x"56",
          5614 => x"87",
          5615 => x"52",
          5616 => x"33",
          5617 => x"3f",
          5618 => x"80",
          5619 => x"bc",
          5620 => x"84",
          5621 => x"5d",
          5622 => x"79",
          5623 => x"38",
          5624 => x"22",
          5625 => x"2e",
          5626 => x"8b",
          5627 => x"f8",
          5628 => x"76",
          5629 => x"83",
          5630 => x"79",
          5631 => x"76",
          5632 => x"ed",
          5633 => x"bb",
          5634 => x"60",
          5635 => x"38",
          5636 => x"06",
          5637 => x"26",
          5638 => x"7b",
          5639 => x"7d",
          5640 => x"76",
          5641 => x"7a",
          5642 => x"70",
          5643 => x"05",
          5644 => x"80",
          5645 => x"5d",
          5646 => x"b0",
          5647 => x"83",
          5648 => x"5d",
          5649 => x"38",
          5650 => x"57",
          5651 => x"38",
          5652 => x"33",
          5653 => x"71",
          5654 => x"71",
          5655 => x"71",
          5656 => x"59",
          5657 => x"77",
          5658 => x"38",
          5659 => x"84",
          5660 => x"7d",
          5661 => x"05",
          5662 => x"77",
          5663 => x"84",
          5664 => x"84",
          5665 => x"41",
          5666 => x"ff",
          5667 => x"ff",
          5668 => x"f6",
          5669 => x"29",
          5670 => x"59",
          5671 => x"77",
          5672 => x"76",
          5673 => x"70",
          5674 => x"05",
          5675 => x"76",
          5676 => x"76",
          5677 => x"e0",
          5678 => x"f4",
          5679 => x"9a",
          5680 => x"a0",
          5681 => x"19",
          5682 => x"70",
          5683 => x"34",
          5684 => x"76",
          5685 => x"c0",
          5686 => x"e0",
          5687 => x"79",
          5688 => x"05",
          5689 => x"17",
          5690 => x"27",
          5691 => x"a8",
          5692 => x"70",
          5693 => x"5d",
          5694 => x"39",
          5695 => x"33",
          5696 => x"06",
          5697 => x"80",
          5698 => x"84",
          5699 => x"5d",
          5700 => x"f0",
          5701 => x"06",
          5702 => x"f2",
          5703 => x"f4",
          5704 => x"70",
          5705 => x"59",
          5706 => x"39",
          5707 => x"17",
          5708 => x"b7",
          5709 => x"7c",
          5710 => x"f8",
          5711 => x"bc",
          5712 => x"f6",
          5713 => x"bb",
          5714 => x"5f",
          5715 => x"39",
          5716 => x"33",
          5717 => x"75",
          5718 => x"34",
          5719 => x"81",
          5720 => x"56",
          5721 => x"83",
          5722 => x"81",
          5723 => x"07",
          5724 => x"f8",
          5725 => x"39",
          5726 => x"33",
          5727 => x"83",
          5728 => x"83",
          5729 => x"d4",
          5730 => x"f4",
          5731 => x"06",
          5732 => x"75",
          5733 => x"34",
          5734 => x"f8",
          5735 => x"9f",
          5736 => x"56",
          5737 => x"f4",
          5738 => x"39",
          5739 => x"83",
          5740 => x"81",
          5741 => x"ff",
          5742 => x"f4",
          5743 => x"f8",
          5744 => x"8f",
          5745 => x"83",
          5746 => x"ff",
          5747 => x"f8",
          5748 => x"9f",
          5749 => x"56",
          5750 => x"f4",
          5751 => x"39",
          5752 => x"33",
          5753 => x"80",
          5754 => x"75",
          5755 => x"34",
          5756 => x"83",
          5757 => x"81",
          5758 => x"c0",
          5759 => x"83",
          5760 => x"fe",
          5761 => x"f8",
          5762 => x"af",
          5763 => x"56",
          5764 => x"f4",
          5765 => x"39",
          5766 => x"33",
          5767 => x"86",
          5768 => x"83",
          5769 => x"fe",
          5770 => x"f8",
          5771 => x"fc",
          5772 => x"56",
          5773 => x"f4",
          5774 => x"39",
          5775 => x"33",
          5776 => x"82",
          5777 => x"83",
          5778 => x"fe",
          5779 => x"f8",
          5780 => x"f8",
          5781 => x"83",
          5782 => x"fd",
          5783 => x"f8",
          5784 => x"f0",
          5785 => x"83",
          5786 => x"fd",
          5787 => x"f8",
          5788 => x"f0",
          5789 => x"83",
          5790 => x"fd",
          5791 => x"f8",
          5792 => x"df",
          5793 => x"07",
          5794 => x"f8",
          5795 => x"cc",
          5796 => x"f4",
          5797 => x"06",
          5798 => x"75",
          5799 => x"34",
          5800 => x"80",
          5801 => x"f9",
          5802 => x"81",
          5803 => x"3f",
          5804 => x"84",
          5805 => x"83",
          5806 => x"84",
          5807 => x"83",
          5808 => x"84",
          5809 => x"59",
          5810 => x"f6",
          5811 => x"84",
          5812 => x"e8",
          5813 => x"0b",
          5814 => x"34",
          5815 => x"b9",
          5816 => x"3d",
          5817 => x"83",
          5818 => x"83",
          5819 => x"70",
          5820 => x"58",
          5821 => x"e7",
          5822 => x"b8",
          5823 => x"3d",
          5824 => x"d8",
          5825 => x"f8",
          5826 => x"b9",
          5827 => x"38",
          5828 => x"08",
          5829 => x"0c",
          5830 => x"b8",
          5831 => x"0b",
          5832 => x"0c",
          5833 => x"04",
          5834 => x"f9",
          5835 => x"39",
          5836 => x"33",
          5837 => x"5c",
          5838 => x"c9",
          5839 => x"83",
          5840 => x"02",
          5841 => x"22",
          5842 => x"1e",
          5843 => x"84",
          5844 => x"ca",
          5845 => x"83",
          5846 => x"80",
          5847 => x"d1",
          5848 => x"f8",
          5849 => x"81",
          5850 => x"ff",
          5851 => x"d8",
          5852 => x"83",
          5853 => x"80",
          5854 => x"d0",
          5855 => x"98",
          5856 => x"fe",
          5857 => x"ef",
          5858 => x"f8",
          5859 => x"05",
          5860 => x"9f",
          5861 => x"58",
          5862 => x"a6",
          5863 => x"81",
          5864 => x"84",
          5865 => x"40",
          5866 => x"ee",
          5867 => x"83",
          5868 => x"ee",
          5869 => x"f8",
          5870 => x"05",
          5871 => x"9f",
          5872 => x"58",
          5873 => x"e2",
          5874 => x"f8",
          5875 => x"84",
          5876 => x"ff",
          5877 => x"56",
          5878 => x"f3",
          5879 => x"57",
          5880 => x"84",
          5881 => x"70",
          5882 => x"58",
          5883 => x"26",
          5884 => x"83",
          5885 => x"84",
          5886 => x"70",
          5887 => x"83",
          5888 => x"71",
          5889 => x"86",
          5890 => x"05",
          5891 => x"22",
          5892 => x"7e",
          5893 => x"83",
          5894 => x"83",
          5895 => x"5d",
          5896 => x"5f",
          5897 => x"2e",
          5898 => x"79",
          5899 => x"06",
          5900 => x"57",
          5901 => x"84",
          5902 => x"b7",
          5903 => x"76",
          5904 => x"98",
          5905 => x"56",
          5906 => x"f6",
          5907 => x"ff",
          5908 => x"57",
          5909 => x"24",
          5910 => x"84",
          5911 => x"56",
          5912 => x"82",
          5913 => x"16",
          5914 => x"f8",
          5915 => x"81",
          5916 => x"f8",
          5917 => x"57",
          5918 => x"76",
          5919 => x"75",
          5920 => x"05",
          5921 => x"06",
          5922 => x"5c",
          5923 => x"58",
          5924 => x"80",
          5925 => x"b0",
          5926 => x"ff",
          5927 => x"ff",
          5928 => x"29",
          5929 => x"42",
          5930 => x"27",
          5931 => x"84",
          5932 => x"57",
          5933 => x"33",
          5934 => x"c4",
          5935 => x"70",
          5936 => x"34",
          5937 => x"05",
          5938 => x"70",
          5939 => x"34",
          5940 => x"b7",
          5941 => x"b7",
          5942 => x"71",
          5943 => x"41",
          5944 => x"76",
          5945 => x"38",
          5946 => x"33",
          5947 => x"c4",
          5948 => x"70",
          5949 => x"34",
          5950 => x"05",
          5951 => x"70",
          5952 => x"34",
          5953 => x"b7",
          5954 => x"b7",
          5955 => x"71",
          5956 => x"41",
          5957 => x"78",
          5958 => x"38",
          5959 => x"83",
          5960 => x"33",
          5961 => x"c4",
          5962 => x"34",
          5963 => x"33",
          5964 => x"33",
          5965 => x"22",
          5966 => x"33",
          5967 => x"5d",
          5968 => x"76",
          5969 => x"84",
          5970 => x"70",
          5971 => x"ff",
          5972 => x"58",
          5973 => x"83",
          5974 => x"79",
          5975 => x"23",
          5976 => x"06",
          5977 => x"5a",
          5978 => x"83",
          5979 => x"76",
          5980 => x"34",
          5981 => x"33",
          5982 => x"06",
          5983 => x"59",
          5984 => x"27",
          5985 => x"80",
          5986 => x"f8",
          5987 => x"88",
          5988 => x"f9",
          5989 => x"84",
          5990 => x"ff",
          5991 => x"56",
          5992 => x"ef",
          5993 => x"57",
          5994 => x"75",
          5995 => x"81",
          5996 => x"38",
          5997 => x"33",
          5998 => x"06",
          5999 => x"33",
          6000 => x"5d",
          6001 => x"2e",
          6002 => x"f4",
          6003 => x"a1",
          6004 => x"56",
          6005 => x"f8",
          6006 => x"39",
          6007 => x"75",
          6008 => x"23",
          6009 => x"7c",
          6010 => x"75",
          6011 => x"34",
          6012 => x"77",
          6013 => x"77",
          6014 => x"8d",
          6015 => x"70",
          6016 => x"34",
          6017 => x"33",
          6018 => x"05",
          6019 => x"7a",
          6020 => x"38",
          6021 => x"81",
          6022 => x"83",
          6023 => x"77",
          6024 => x"59",
          6025 => x"27",
          6026 => x"d3",
          6027 => x"31",
          6028 => x"f8",
          6029 => x"a8",
          6030 => x"83",
          6031 => x"fc",
          6032 => x"83",
          6033 => x"fc",
          6034 => x"0b",
          6035 => x"23",
          6036 => x"80",
          6037 => x"f8",
          6038 => x"39",
          6039 => x"18",
          6040 => x"b7",
          6041 => x"77",
          6042 => x"83",
          6043 => x"e9",
          6044 => x"3d",
          6045 => x"05",
          6046 => x"be",
          6047 => x"72",
          6048 => x"38",
          6049 => x"9c",
          6050 => x"84",
          6051 => x"85",
          6052 => x"76",
          6053 => x"d7",
          6054 => x"0b",
          6055 => x"0c",
          6056 => x"04",
          6057 => x"02",
          6058 => x"5c",
          6059 => x"f7",
          6060 => x"81",
          6061 => x"f7",
          6062 => x"58",
          6063 => x"74",
          6064 => x"d6",
          6065 => x"56",
          6066 => x"cc",
          6067 => x"78",
          6068 => x"0c",
          6069 => x"04",
          6070 => x"08",
          6071 => x"73",
          6072 => x"38",
          6073 => x"70",
          6074 => x"70",
          6075 => x"2a",
          6076 => x"58",
          6077 => x"a8",
          6078 => x"80",
          6079 => x"2e",
          6080 => x"83",
          6081 => x"7b",
          6082 => x"30",
          6083 => x"76",
          6084 => x"5d",
          6085 => x"85",
          6086 => x"b7",
          6087 => x"f8",
          6088 => x"f8",
          6089 => x"71",
          6090 => x"a7",
          6091 => x"83",
          6092 => x"5b",
          6093 => x"79",
          6094 => x"83",
          6095 => x"83",
          6096 => x"58",
          6097 => x"74",
          6098 => x"8c",
          6099 => x"54",
          6100 => x"80",
          6101 => x"0b",
          6102 => x"88",
          6103 => x"98",
          6104 => x"75",
          6105 => x"38",
          6106 => x"84",
          6107 => x"83",
          6108 => x"34",
          6109 => x"81",
          6110 => x"55",
          6111 => x"27",
          6112 => x"54",
          6113 => x"14",
          6114 => x"ff",
          6115 => x"f2",
          6116 => x"54",
          6117 => x"2e",
          6118 => x"72",
          6119 => x"86",
          6120 => x"83",
          6121 => x"34",
          6122 => x"06",
          6123 => x"ff",
          6124 => x"38",
          6125 => x"86",
          6126 => x"f6",
          6127 => x"83",
          6128 => x"34",
          6129 => x"81",
          6130 => x"5e",
          6131 => x"ff",
          6132 => x"f6",
          6133 => x"98",
          6134 => x"25",
          6135 => x"75",
          6136 => x"34",
          6137 => x"06",
          6138 => x"81",
          6139 => x"06",
          6140 => x"72",
          6141 => x"e7",
          6142 => x"83",
          6143 => x"73",
          6144 => x"53",
          6145 => x"85",
          6146 => x"0b",
          6147 => x"34",
          6148 => x"f7",
          6149 => x"f7",
          6150 => x"f7",
          6151 => x"83",
          6152 => x"83",
          6153 => x"5d",
          6154 => x"5c",
          6155 => x"f6",
          6156 => x"55",
          6157 => x"2e",
          6158 => x"f7",
          6159 => x"54",
          6160 => x"82",
          6161 => x"f7",
          6162 => x"53",
          6163 => x"2e",
          6164 => x"f7",
          6165 => x"54",
          6166 => x"38",
          6167 => x"06",
          6168 => x"ff",
          6169 => x"83",
          6170 => x"33",
          6171 => x"2e",
          6172 => x"74",
          6173 => x"53",
          6174 => x"2e",
          6175 => x"83",
          6176 => x"33",
          6177 => x"27",
          6178 => x"83",
          6179 => x"87",
          6180 => x"c0",
          6181 => x"54",
          6182 => x"27",
          6183 => x"81",
          6184 => x"98",
          6185 => x"f7",
          6186 => x"81",
          6187 => x"ff",
          6188 => x"89",
          6189 => x"f6",
          6190 => x"f7",
          6191 => x"83",
          6192 => x"fe",
          6193 => x"72",
          6194 => x"8b",
          6195 => x"10",
          6196 => x"05",
          6197 => x"04",
          6198 => x"08",
          6199 => x"2e",
          6200 => x"f4",
          6201 => x"98",
          6202 => x"5e",
          6203 => x"fc",
          6204 => x"0b",
          6205 => x"33",
          6206 => x"81",
          6207 => x"74",
          6208 => x"f7",
          6209 => x"c0",
          6210 => x"83",
          6211 => x"73",
          6212 => x"58",
          6213 => x"94",
          6214 => x"fa",
          6215 => x"84",
          6216 => x"33",
          6217 => x"f0",
          6218 => x"39",
          6219 => x"08",
          6220 => x"2e",
          6221 => x"72",
          6222 => x"f4",
          6223 => x"76",
          6224 => x"54",
          6225 => x"80",
          6226 => x"39",
          6227 => x"57",
          6228 => x"81",
          6229 => x"79",
          6230 => x"81",
          6231 => x"38",
          6232 => x"80",
          6233 => x"81",
          6234 => x"38",
          6235 => x"06",
          6236 => x"27",
          6237 => x"54",
          6238 => x"25",
          6239 => x"80",
          6240 => x"81",
          6241 => x"ff",
          6242 => x"81",
          6243 => x"72",
          6244 => x"2b",
          6245 => x"58",
          6246 => x"24",
          6247 => x"10",
          6248 => x"10",
          6249 => x"83",
          6250 => x"83",
          6251 => x"70",
          6252 => x"54",
          6253 => x"98",
          6254 => x"f7",
          6255 => x"fd",
          6256 => x"59",
          6257 => x"ff",
          6258 => x"81",
          6259 => x"ff",
          6260 => x"59",
          6261 => x"78",
          6262 => x"9f",
          6263 => x"84",
          6264 => x"54",
          6265 => x"2e",
          6266 => x"7b",
          6267 => x"30",
          6268 => x"76",
          6269 => x"56",
          6270 => x"7b",
          6271 => x"81",
          6272 => x"38",
          6273 => x"f9",
          6274 => x"53",
          6275 => x"10",
          6276 => x"05",
          6277 => x"54",
          6278 => x"83",
          6279 => x"13",
          6280 => x"06",
          6281 => x"73",
          6282 => x"84",
          6283 => x"53",
          6284 => x"f9",
          6285 => x"b7",
          6286 => x"74",
          6287 => x"78",
          6288 => x"52",
          6289 => x"d4",
          6290 => x"b9",
          6291 => x"3d",
          6292 => x"76",
          6293 => x"54",
          6294 => x"72",
          6295 => x"92",
          6296 => x"90",
          6297 => x"05",
          6298 => x"f7",
          6299 => x"fa",
          6300 => x"0b",
          6301 => x"15",
          6302 => x"83",
          6303 => x"34",
          6304 => x"f7",
          6305 => x"fa",
          6306 => x"81",
          6307 => x"72",
          6308 => x"fc",
          6309 => x"f7",
          6310 => x"55",
          6311 => x"fc",
          6312 => x"81",
          6313 => x"73",
          6314 => x"81",
          6315 => x"38",
          6316 => x"08",
          6317 => x"87",
          6318 => x"08",
          6319 => x"73",
          6320 => x"38",
          6321 => x"9c",
          6322 => x"9c",
          6323 => x"ff",
          6324 => x"d7",
          6325 => x"83",
          6326 => x"34",
          6327 => x"72",
          6328 => x"34",
          6329 => x"06",
          6330 => x"9e",
          6331 => x"f7",
          6332 => x"0b",
          6333 => x"33",
          6334 => x"08",
          6335 => x"33",
          6336 => x"a4",
          6337 => x"a3",
          6338 => x"42",
          6339 => x"56",
          6340 => x"79",
          6341 => x"81",
          6342 => x"38",
          6343 => x"81",
          6344 => x"38",
          6345 => x"09",
          6346 => x"c0",
          6347 => x"39",
          6348 => x"81",
          6349 => x"98",
          6350 => x"84",
          6351 => x"57",
          6352 => x"38",
          6353 => x"84",
          6354 => x"ff",
          6355 => x"39",
          6356 => x"b7",
          6357 => x"54",
          6358 => x"81",
          6359 => x"b7",
          6360 => x"59",
          6361 => x"81",
          6362 => x"a8",
          6363 => x"f7",
          6364 => x"0b",
          6365 => x"0c",
          6366 => x"84",
          6367 => x"70",
          6368 => x"ff",
          6369 => x"54",
          6370 => x"83",
          6371 => x"74",
          6372 => x"23",
          6373 => x"06",
          6374 => x"53",
          6375 => x"83",
          6376 => x"73",
          6377 => x"34",
          6378 => x"33",
          6379 => x"06",
          6380 => x"53",
          6381 => x"83",
          6382 => x"72",
          6383 => x"34",
          6384 => x"b7",
          6385 => x"83",
          6386 => x"a5",
          6387 => x"f6",
          6388 => x"54",
          6389 => x"84",
          6390 => x"83",
          6391 => x"fe",
          6392 => x"81",
          6393 => x"cc",
          6394 => x"ac",
          6395 => x"bb",
          6396 => x"0d",
          6397 => x"ac",
          6398 => x"0d",
          6399 => x"0d",
          6400 => x"f3",
          6401 => x"57",
          6402 => x"33",
          6403 => x"83",
          6404 => x"51",
          6405 => x"34",
          6406 => x"f3",
          6407 => x"56",
          6408 => x"15",
          6409 => x"87",
          6410 => x"34",
          6411 => x"9c",
          6412 => x"d4",
          6413 => x"ce",
          6414 => x"87",
          6415 => x"08",
          6416 => x"98",
          6417 => x"70",
          6418 => x"38",
          6419 => x"87",
          6420 => x"08",
          6421 => x"73",
          6422 => x"71",
          6423 => x"db",
          6424 => x"98",
          6425 => x"ff",
          6426 => x"27",
          6427 => x"71",
          6428 => x"2e",
          6429 => x"87",
          6430 => x"08",
          6431 => x"05",
          6432 => x"98",
          6433 => x"87",
          6434 => x"08",
          6435 => x"2e",
          6436 => x"14",
          6437 => x"98",
          6438 => x"52",
          6439 => x"87",
          6440 => x"ff",
          6441 => x"87",
          6442 => x"08",
          6443 => x"26",
          6444 => x"52",
          6445 => x"16",
          6446 => x"06",
          6447 => x"80",
          6448 => x"74",
          6449 => x"52",
          6450 => x"38",
          6451 => x"8a",
          6452 => x"b9",
          6453 => x"3d",
          6454 => x"0b",
          6455 => x"0c",
          6456 => x"04",
          6457 => x"79",
          6458 => x"a3",
          6459 => x"52",
          6460 => x"f3",
          6461 => x"88",
          6462 => x"80",
          6463 => x"75",
          6464 => x"51",
          6465 => x"71",
          6466 => x"72",
          6467 => x"70",
          6468 => x"71",
          6469 => x"75",
          6470 => x"72",
          6471 => x"83",
          6472 => x"52",
          6473 => x"34",
          6474 => x"08",
          6475 => x"71",
          6476 => x"83",
          6477 => x"55",
          6478 => x"81",
          6479 => x"0b",
          6480 => x"e8",
          6481 => x"98",
          6482 => x"f3",
          6483 => x"80",
          6484 => x"53",
          6485 => x"9c",
          6486 => x"c0",
          6487 => x"51",
          6488 => x"f6",
          6489 => x"33",
          6490 => x"9c",
          6491 => x"74",
          6492 => x"38",
          6493 => x"2e",
          6494 => x"c0",
          6495 => x"51",
          6496 => x"73",
          6497 => x"38",
          6498 => x"ff",
          6499 => x"38",
          6500 => x"9c",
          6501 => x"90",
          6502 => x"c0",
          6503 => x"52",
          6504 => x"9c",
          6505 => x"72",
          6506 => x"81",
          6507 => x"c0",
          6508 => x"52",
          6509 => x"27",
          6510 => x"81",
          6511 => x"38",
          6512 => x"a4",
          6513 => x"75",
          6514 => x"ff",
          6515 => x"ff",
          6516 => x"ff",
          6517 => x"75",
          6518 => x"c7",
          6519 => x"ff",
          6520 => x"fe",
          6521 => x"51",
          6522 => x"06",
          6523 => x"38",
          6524 => x"7b",
          6525 => x"55",
          6526 => x"73",
          6527 => x"71",
          6528 => x"53",
          6529 => x"81",
          6530 => x"72",
          6531 => x"38",
          6532 => x"c8",
          6533 => x"0d",
          6534 => x"84",
          6535 => x"88",
          6536 => x"ff",
          6537 => x"fa",
          6538 => x"02",
          6539 => x"05",
          6540 => x"80",
          6541 => x"d4",
          6542 => x"2b",
          6543 => x"80",
          6544 => x"98",
          6545 => x"55",
          6546 => x"83",
          6547 => x"90",
          6548 => x"84",
          6549 => x"90",
          6550 => x"85",
          6551 => x"86",
          6552 => x"83",
          6553 => x"80",
          6554 => x"80",
          6555 => x"55",
          6556 => x"27",
          6557 => x"70",
          6558 => x"33",
          6559 => x"05",
          6560 => x"71",
          6561 => x"83",
          6562 => x"54",
          6563 => x"34",
          6564 => x"08",
          6565 => x"75",
          6566 => x"83",
          6567 => x"55",
          6568 => x"81",
          6569 => x"0b",
          6570 => x"e8",
          6571 => x"98",
          6572 => x"f3",
          6573 => x"80",
          6574 => x"53",
          6575 => x"9c",
          6576 => x"c0",
          6577 => x"51",
          6578 => x"f6",
          6579 => x"33",
          6580 => x"9c",
          6581 => x"74",
          6582 => x"38",
          6583 => x"2e",
          6584 => x"c0",
          6585 => x"51",
          6586 => x"73",
          6587 => x"38",
          6588 => x"ff",
          6589 => x"38",
          6590 => x"9c",
          6591 => x"90",
          6592 => x"c0",
          6593 => x"52",
          6594 => x"9c",
          6595 => x"72",
          6596 => x"81",
          6597 => x"c0",
          6598 => x"52",
          6599 => x"27",
          6600 => x"81",
          6601 => x"38",
          6602 => x"a4",
          6603 => x"75",
          6604 => x"ff",
          6605 => x"ff",
          6606 => x"ff",
          6607 => x"75",
          6608 => x"38",
          6609 => x"06",
          6610 => x"d5",
          6611 => x"70",
          6612 => x"54",
          6613 => x"83",
          6614 => x"76",
          6615 => x"0c",
          6616 => x"04",
          6617 => x"39",
          6618 => x"83",
          6619 => x"51",
          6620 => x"34",
          6621 => x"f3",
          6622 => x"56",
          6623 => x"16",
          6624 => x"87",
          6625 => x"34",
          6626 => x"9c",
          6627 => x"d4",
          6628 => x"ce",
          6629 => x"87",
          6630 => x"08",
          6631 => x"98",
          6632 => x"72",
          6633 => x"38",
          6634 => x"87",
          6635 => x"08",
          6636 => x"74",
          6637 => x"71",
          6638 => x"db",
          6639 => x"98",
          6640 => x"ff",
          6641 => x"27",
          6642 => x"71",
          6643 => x"2e",
          6644 => x"87",
          6645 => x"08",
          6646 => x"05",
          6647 => x"98",
          6648 => x"87",
          6649 => x"08",
          6650 => x"2e",
          6651 => x"15",
          6652 => x"98",
          6653 => x"52",
          6654 => x"87",
          6655 => x"ff",
          6656 => x"87",
          6657 => x"08",
          6658 => x"26",
          6659 => x"52",
          6660 => x"16",
          6661 => x"06",
          6662 => x"80",
          6663 => x"72",
          6664 => x"54",
          6665 => x"38",
          6666 => x"3d",
          6667 => x"cc",
          6668 => x"bf",
          6669 => x"0d",
          6670 => x"0d",
          6671 => x"08",
          6672 => x"83",
          6673 => x"ff",
          6674 => x"83",
          6675 => x"70",
          6676 => x"33",
          6677 => x"71",
          6678 => x"77",
          6679 => x"81",
          6680 => x"98",
          6681 => x"2b",
          6682 => x"41",
          6683 => x"57",
          6684 => x"57",
          6685 => x"24",
          6686 => x"72",
          6687 => x"33",
          6688 => x"71",
          6689 => x"83",
          6690 => x"05",
          6691 => x"12",
          6692 => x"2b",
          6693 => x"07",
          6694 => x"52",
          6695 => x"80",
          6696 => x"9e",
          6697 => x"33",
          6698 => x"71",
          6699 => x"83",
          6700 => x"05",
          6701 => x"52",
          6702 => x"74",
          6703 => x"73",
          6704 => x"54",
          6705 => x"34",
          6706 => x"08",
          6707 => x"12",
          6708 => x"33",
          6709 => x"07",
          6710 => x"5c",
          6711 => x"51",
          6712 => x"34",
          6713 => x"34",
          6714 => x"08",
          6715 => x"0b",
          6716 => x"80",
          6717 => x"34",
          6718 => x"08",
          6719 => x"14",
          6720 => x"14",
          6721 => x"b8",
          6722 => x"33",
          6723 => x"71",
          6724 => x"82",
          6725 => x"70",
          6726 => x"58",
          6727 => x"72",
          6728 => x"13",
          6729 => x"0d",
          6730 => x"33",
          6731 => x"71",
          6732 => x"83",
          6733 => x"11",
          6734 => x"85",
          6735 => x"88",
          6736 => x"88",
          6737 => x"54",
          6738 => x"58",
          6739 => x"34",
          6740 => x"34",
          6741 => x"08",
          6742 => x"11",
          6743 => x"33",
          6744 => x"71",
          6745 => x"56",
          6746 => x"72",
          6747 => x"33",
          6748 => x"71",
          6749 => x"70",
          6750 => x"55",
          6751 => x"86",
          6752 => x"87",
          6753 => x"b9",
          6754 => x"70",
          6755 => x"33",
          6756 => x"07",
          6757 => x"06",
          6758 => x"5a",
          6759 => x"76",
          6760 => x"81",
          6761 => x"b9",
          6762 => x"17",
          6763 => x"12",
          6764 => x"2b",
          6765 => x"07",
          6766 => x"33",
          6767 => x"71",
          6768 => x"70",
          6769 => x"ff",
          6770 => x"05",
          6771 => x"54",
          6772 => x"5c",
          6773 => x"52",
          6774 => x"34",
          6775 => x"34",
          6776 => x"08",
          6777 => x"33",
          6778 => x"71",
          6779 => x"83",
          6780 => x"05",
          6781 => x"12",
          6782 => x"2b",
          6783 => x"ff",
          6784 => x"2a",
          6785 => x"55",
          6786 => x"52",
          6787 => x"70",
          6788 => x"84",
          6789 => x"70",
          6790 => x"33",
          6791 => x"71",
          6792 => x"83",
          6793 => x"05",
          6794 => x"12",
          6795 => x"2b",
          6796 => x"07",
          6797 => x"52",
          6798 => x"53",
          6799 => x"fc",
          6800 => x"33",
          6801 => x"71",
          6802 => x"82",
          6803 => x"70",
          6804 => x"59",
          6805 => x"34",
          6806 => x"34",
          6807 => x"08",
          6808 => x"33",
          6809 => x"71",
          6810 => x"83",
          6811 => x"05",
          6812 => x"83",
          6813 => x"88",
          6814 => x"88",
          6815 => x"5c",
          6816 => x"52",
          6817 => x"15",
          6818 => x"15",
          6819 => x"0d",
          6820 => x"0d",
          6821 => x"b8",
          6822 => x"76",
          6823 => x"38",
          6824 => x"86",
          6825 => x"fb",
          6826 => x"3d",
          6827 => x"ff",
          6828 => x"b9",
          6829 => x"80",
          6830 => x"b4",
          6831 => x"80",
          6832 => x"84",
          6833 => x"fe",
          6834 => x"84",
          6835 => x"55",
          6836 => x"81",
          6837 => x"34",
          6838 => x"08",
          6839 => x"15",
          6840 => x"85",
          6841 => x"b9",
          6842 => x"76",
          6843 => x"81",
          6844 => x"34",
          6845 => x"08",
          6846 => x"22",
          6847 => x"80",
          6848 => x"83",
          6849 => x"70",
          6850 => x"51",
          6851 => x"88",
          6852 => x"89",
          6853 => x"b9",
          6854 => x"10",
          6855 => x"b9",
          6856 => x"f8",
          6857 => x"76",
          6858 => x"81",
          6859 => x"34",
          6860 => x"f7",
          6861 => x"52",
          6862 => x"51",
          6863 => x"8e",
          6864 => x"83",
          6865 => x"70",
          6866 => x"06",
          6867 => x"83",
          6868 => x"84",
          6869 => x"84",
          6870 => x"12",
          6871 => x"2b",
          6872 => x"59",
          6873 => x"81",
          6874 => x"75",
          6875 => x"cc",
          6876 => x"10",
          6877 => x"33",
          6878 => x"71",
          6879 => x"70",
          6880 => x"06",
          6881 => x"83",
          6882 => x"70",
          6883 => x"53",
          6884 => x"52",
          6885 => x"8a",
          6886 => x"2e",
          6887 => x"73",
          6888 => x"12",
          6889 => x"33",
          6890 => x"07",
          6891 => x"c1",
          6892 => x"ff",
          6893 => x"38",
          6894 => x"56",
          6895 => x"2b",
          6896 => x"33",
          6897 => x"71",
          6898 => x"70",
          6899 => x"06",
          6900 => x"56",
          6901 => x"79",
          6902 => x"81",
          6903 => x"74",
          6904 => x"8d",
          6905 => x"78",
          6906 => x"85",
          6907 => x"2e",
          6908 => x"74",
          6909 => x"2b",
          6910 => x"82",
          6911 => x"70",
          6912 => x"5c",
          6913 => x"76",
          6914 => x"81",
          6915 => x"b9",
          6916 => x"76",
          6917 => x"53",
          6918 => x"34",
          6919 => x"34",
          6920 => x"08",
          6921 => x"33",
          6922 => x"71",
          6923 => x"70",
          6924 => x"ff",
          6925 => x"05",
          6926 => x"ff",
          6927 => x"2a",
          6928 => x"57",
          6929 => x"75",
          6930 => x"72",
          6931 => x"53",
          6932 => x"34",
          6933 => x"08",
          6934 => x"74",
          6935 => x"15",
          6936 => x"b8",
          6937 => x"86",
          6938 => x"12",
          6939 => x"2b",
          6940 => x"07",
          6941 => x"5c",
          6942 => x"75",
          6943 => x"72",
          6944 => x"84",
          6945 => x"70",
          6946 => x"05",
          6947 => x"87",
          6948 => x"88",
          6949 => x"88",
          6950 => x"58",
          6951 => x"15",
          6952 => x"15",
          6953 => x"b8",
          6954 => x"84",
          6955 => x"12",
          6956 => x"2b",
          6957 => x"07",
          6958 => x"5a",
          6959 => x"75",
          6960 => x"72",
          6961 => x"84",
          6962 => x"70",
          6963 => x"05",
          6964 => x"85",
          6965 => x"88",
          6966 => x"88",
          6967 => x"57",
          6968 => x"15",
          6969 => x"15",
          6970 => x"b8",
          6971 => x"05",
          6972 => x"b9",
          6973 => x"3d",
          6974 => x"14",
          6975 => x"33",
          6976 => x"71",
          6977 => x"79",
          6978 => x"33",
          6979 => x"71",
          6980 => x"70",
          6981 => x"5b",
          6982 => x"52",
          6983 => x"34",
          6984 => x"34",
          6985 => x"08",
          6986 => x"11",
          6987 => x"33",
          6988 => x"71",
          6989 => x"74",
          6990 => x"33",
          6991 => x"71",
          6992 => x"70",
          6993 => x"5d",
          6994 => x"5b",
          6995 => x"86",
          6996 => x"87",
          6997 => x"b9",
          6998 => x"70",
          6999 => x"33",
          7000 => x"07",
          7001 => x"06",
          7002 => x"59",
          7003 => x"75",
          7004 => x"81",
          7005 => x"b9",
          7006 => x"84",
          7007 => x"f1",
          7008 => x"0d",
          7009 => x"b8",
          7010 => x"76",
          7011 => x"38",
          7012 => x"8a",
          7013 => x"b9",
          7014 => x"3d",
          7015 => x"51",
          7016 => x"84",
          7017 => x"84",
          7018 => x"89",
          7019 => x"84",
          7020 => x"84",
          7021 => x"a0",
          7022 => x"b9",
          7023 => x"80",
          7024 => x"52",
          7025 => x"51",
          7026 => x"3f",
          7027 => x"08",
          7028 => x"34",
          7029 => x"16",
          7030 => x"b8",
          7031 => x"84",
          7032 => x"0b",
          7033 => x"84",
          7034 => x"56",
          7035 => x"34",
          7036 => x"17",
          7037 => x"b8",
          7038 => x"b4",
          7039 => x"fe",
          7040 => x"70",
          7041 => x"06",
          7042 => x"58",
          7043 => x"74",
          7044 => x"73",
          7045 => x"84",
          7046 => x"70",
          7047 => x"84",
          7048 => x"05",
          7049 => x"55",
          7050 => x"34",
          7051 => x"15",
          7052 => x"77",
          7053 => x"dd",
          7054 => x"39",
          7055 => x"65",
          7056 => x"80",
          7057 => x"b8",
          7058 => x"41",
          7059 => x"84",
          7060 => x"80",
          7061 => x"38",
          7062 => x"88",
          7063 => x"54",
          7064 => x"8f",
          7065 => x"05",
          7066 => x"05",
          7067 => x"ff",
          7068 => x"73",
          7069 => x"06",
          7070 => x"83",
          7071 => x"ff",
          7072 => x"83",
          7073 => x"70",
          7074 => x"33",
          7075 => x"07",
          7076 => x"70",
          7077 => x"06",
          7078 => x"10",
          7079 => x"83",
          7080 => x"70",
          7081 => x"33",
          7082 => x"07",
          7083 => x"70",
          7084 => x"42",
          7085 => x"53",
          7086 => x"5c",
          7087 => x"5e",
          7088 => x"7a",
          7089 => x"38",
          7090 => x"83",
          7091 => x"88",
          7092 => x"10",
          7093 => x"70",
          7094 => x"33",
          7095 => x"71",
          7096 => x"53",
          7097 => x"56",
          7098 => x"24",
          7099 => x"7a",
          7100 => x"f6",
          7101 => x"58",
          7102 => x"87",
          7103 => x"80",
          7104 => x"38",
          7105 => x"77",
          7106 => x"be",
          7107 => x"59",
          7108 => x"92",
          7109 => x"1e",
          7110 => x"12",
          7111 => x"2b",
          7112 => x"07",
          7113 => x"33",
          7114 => x"71",
          7115 => x"90",
          7116 => x"43",
          7117 => x"57",
          7118 => x"60",
          7119 => x"38",
          7120 => x"11",
          7121 => x"33",
          7122 => x"71",
          7123 => x"7a",
          7124 => x"33",
          7125 => x"71",
          7126 => x"83",
          7127 => x"05",
          7128 => x"85",
          7129 => x"88",
          7130 => x"88",
          7131 => x"48",
          7132 => x"58",
          7133 => x"56",
          7134 => x"34",
          7135 => x"34",
          7136 => x"08",
          7137 => x"11",
          7138 => x"33",
          7139 => x"71",
          7140 => x"74",
          7141 => x"33",
          7142 => x"71",
          7143 => x"70",
          7144 => x"42",
          7145 => x"57",
          7146 => x"86",
          7147 => x"87",
          7148 => x"b9",
          7149 => x"70",
          7150 => x"33",
          7151 => x"07",
          7152 => x"06",
          7153 => x"5a",
          7154 => x"76",
          7155 => x"81",
          7156 => x"b9",
          7157 => x"1f",
          7158 => x"83",
          7159 => x"8b",
          7160 => x"2b",
          7161 => x"73",
          7162 => x"33",
          7163 => x"07",
          7164 => x"41",
          7165 => x"5f",
          7166 => x"79",
          7167 => x"81",
          7168 => x"b9",
          7169 => x"1f",
          7170 => x"12",
          7171 => x"2b",
          7172 => x"07",
          7173 => x"14",
          7174 => x"33",
          7175 => x"07",
          7176 => x"41",
          7177 => x"5f",
          7178 => x"79",
          7179 => x"75",
          7180 => x"84",
          7181 => x"70",
          7182 => x"33",
          7183 => x"71",
          7184 => x"66",
          7185 => x"70",
          7186 => x"52",
          7187 => x"05",
          7188 => x"fe",
          7189 => x"84",
          7190 => x"1e",
          7191 => x"65",
          7192 => x"83",
          7193 => x"5d",
          7194 => x"62",
          7195 => x"38",
          7196 => x"84",
          7197 => x"95",
          7198 => x"84",
          7199 => x"84",
          7200 => x"a0",
          7201 => x"b9",
          7202 => x"80",
          7203 => x"52",
          7204 => x"51",
          7205 => x"3f",
          7206 => x"08",
          7207 => x"34",
          7208 => x"1f",
          7209 => x"b8",
          7210 => x"84",
          7211 => x"0b",
          7212 => x"84",
          7213 => x"5c",
          7214 => x"34",
          7215 => x"1d",
          7216 => x"b8",
          7217 => x"b4",
          7218 => x"fe",
          7219 => x"70",
          7220 => x"06",
          7221 => x"5c",
          7222 => x"78",
          7223 => x"77",
          7224 => x"84",
          7225 => x"70",
          7226 => x"84",
          7227 => x"05",
          7228 => x"56",
          7229 => x"34",
          7230 => x"15",
          7231 => x"b8",
          7232 => x"fa",
          7233 => x"80",
          7234 => x"38",
          7235 => x"80",
          7236 => x"38",
          7237 => x"9b",
          7238 => x"c8",
          7239 => x"c8",
          7240 => x"0d",
          7241 => x"84",
          7242 => x"71",
          7243 => x"11",
          7244 => x"05",
          7245 => x"12",
          7246 => x"2b",
          7247 => x"ff",
          7248 => x"2a",
          7249 => x"5e",
          7250 => x"34",
          7251 => x"34",
          7252 => x"b8",
          7253 => x"88",
          7254 => x"75",
          7255 => x"7b",
          7256 => x"84",
          7257 => x"70",
          7258 => x"81",
          7259 => x"88",
          7260 => x"83",
          7261 => x"f8",
          7262 => x"64",
          7263 => x"06",
          7264 => x"4a",
          7265 => x"5e",
          7266 => x"63",
          7267 => x"76",
          7268 => x"41",
          7269 => x"05",
          7270 => x"b8",
          7271 => x"63",
          7272 => x"81",
          7273 => x"84",
          7274 => x"05",
          7275 => x"ed",
          7276 => x"54",
          7277 => x"7b",
          7278 => x"83",
          7279 => x"42",
          7280 => x"39",
          7281 => x"ff",
          7282 => x"70",
          7283 => x"06",
          7284 => x"83",
          7285 => x"88",
          7286 => x"10",
          7287 => x"70",
          7288 => x"33",
          7289 => x"71",
          7290 => x"53",
          7291 => x"58",
          7292 => x"73",
          7293 => x"f7",
          7294 => x"39",
          7295 => x"fa",
          7296 => x"7a",
          7297 => x"38",
          7298 => x"ff",
          7299 => x"7b",
          7300 => x"38",
          7301 => x"84",
          7302 => x"84",
          7303 => x"a0",
          7304 => x"b9",
          7305 => x"80",
          7306 => x"52",
          7307 => x"51",
          7308 => x"3f",
          7309 => x"08",
          7310 => x"34",
          7311 => x"1b",
          7312 => x"b8",
          7313 => x"84",
          7314 => x"0b",
          7315 => x"84",
          7316 => x"58",
          7317 => x"34",
          7318 => x"19",
          7319 => x"b8",
          7320 => x"b4",
          7321 => x"fe",
          7322 => x"70",
          7323 => x"06",
          7324 => x"58",
          7325 => x"74",
          7326 => x"34",
          7327 => x"05",
          7328 => x"b4",
          7329 => x"10",
          7330 => x"b8",
          7331 => x"05",
          7332 => x"61",
          7333 => x"81",
          7334 => x"34",
          7335 => x"80",
          7336 => x"de",
          7337 => x"ff",
          7338 => x"61",
          7339 => x"c0",
          7340 => x"39",
          7341 => x"82",
          7342 => x"51",
          7343 => x"7f",
          7344 => x"b9",
          7345 => x"3d",
          7346 => x"1e",
          7347 => x"83",
          7348 => x"8b",
          7349 => x"2b",
          7350 => x"86",
          7351 => x"12",
          7352 => x"2b",
          7353 => x"07",
          7354 => x"14",
          7355 => x"33",
          7356 => x"07",
          7357 => x"43",
          7358 => x"5b",
          7359 => x"5c",
          7360 => x"64",
          7361 => x"7a",
          7362 => x"34",
          7363 => x"08",
          7364 => x"11",
          7365 => x"33",
          7366 => x"71",
          7367 => x"74",
          7368 => x"33",
          7369 => x"71",
          7370 => x"70",
          7371 => x"41",
          7372 => x"59",
          7373 => x"64",
          7374 => x"7a",
          7375 => x"34",
          7376 => x"08",
          7377 => x"81",
          7378 => x"88",
          7379 => x"ff",
          7380 => x"88",
          7381 => x"5a",
          7382 => x"34",
          7383 => x"34",
          7384 => x"08",
          7385 => x"11",
          7386 => x"33",
          7387 => x"71",
          7388 => x"74",
          7389 => x"81",
          7390 => x"88",
          7391 => x"88",
          7392 => x"5e",
          7393 => x"45",
          7394 => x"34",
          7395 => x"34",
          7396 => x"08",
          7397 => x"33",
          7398 => x"71",
          7399 => x"83",
          7400 => x"05",
          7401 => x"83",
          7402 => x"88",
          7403 => x"88",
          7404 => x"40",
          7405 => x"55",
          7406 => x"18",
          7407 => x"18",
          7408 => x"b8",
          7409 => x"82",
          7410 => x"12",
          7411 => x"2b",
          7412 => x"62",
          7413 => x"2b",
          7414 => x"5d",
          7415 => x"05",
          7416 => x"de",
          7417 => x"b8",
          7418 => x"05",
          7419 => x"ff",
          7420 => x"fc",
          7421 => x"ff",
          7422 => x"b9",
          7423 => x"80",
          7424 => x"b4",
          7425 => x"80",
          7426 => x"84",
          7427 => x"fe",
          7428 => x"84",
          7429 => x"56",
          7430 => x"81",
          7431 => x"34",
          7432 => x"08",
          7433 => x"16",
          7434 => x"85",
          7435 => x"b9",
          7436 => x"7f",
          7437 => x"81",
          7438 => x"34",
          7439 => x"08",
          7440 => x"22",
          7441 => x"80",
          7442 => x"83",
          7443 => x"70",
          7444 => x"43",
          7445 => x"88",
          7446 => x"89",
          7447 => x"b9",
          7448 => x"10",
          7449 => x"b9",
          7450 => x"f8",
          7451 => x"7f",
          7452 => x"81",
          7453 => x"34",
          7454 => x"bd",
          7455 => x"fc",
          7456 => x"19",
          7457 => x"33",
          7458 => x"71",
          7459 => x"79",
          7460 => x"33",
          7461 => x"71",
          7462 => x"70",
          7463 => x"48",
          7464 => x"55",
          7465 => x"05",
          7466 => x"85",
          7467 => x"b9",
          7468 => x"1e",
          7469 => x"85",
          7470 => x"8b",
          7471 => x"2b",
          7472 => x"86",
          7473 => x"15",
          7474 => x"2b",
          7475 => x"2a",
          7476 => x"48",
          7477 => x"40",
          7478 => x"05",
          7479 => x"87",
          7480 => x"b9",
          7481 => x"70",
          7482 => x"33",
          7483 => x"07",
          7484 => x"06",
          7485 => x"59",
          7486 => x"75",
          7487 => x"81",
          7488 => x"b9",
          7489 => x"1f",
          7490 => x"12",
          7491 => x"2b",
          7492 => x"07",
          7493 => x"33",
          7494 => x"71",
          7495 => x"70",
          7496 => x"ff",
          7497 => x"05",
          7498 => x"48",
          7499 => x"5d",
          7500 => x"41",
          7501 => x"34",
          7502 => x"34",
          7503 => x"08",
          7504 => x"33",
          7505 => x"71",
          7506 => x"83",
          7507 => x"05",
          7508 => x"12",
          7509 => x"2b",
          7510 => x"ff",
          7511 => x"2a",
          7512 => x"5e",
          7513 => x"5b",
          7514 => x"76",
          7515 => x"34",
          7516 => x"ff",
          7517 => x"b3",
          7518 => x"33",
          7519 => x"71",
          7520 => x"83",
          7521 => x"05",
          7522 => x"85",
          7523 => x"88",
          7524 => x"88",
          7525 => x"5a",
          7526 => x"78",
          7527 => x"79",
          7528 => x"84",
          7529 => x"70",
          7530 => x"33",
          7531 => x"71",
          7532 => x"83",
          7533 => x"05",
          7534 => x"87",
          7535 => x"88",
          7536 => x"88",
          7537 => x"5e",
          7538 => x"55",
          7539 => x"86",
          7540 => x"60",
          7541 => x"84",
          7542 => x"18",
          7543 => x"12",
          7544 => x"2b",
          7545 => x"ff",
          7546 => x"2a",
          7547 => x"55",
          7548 => x"78",
          7549 => x"84",
          7550 => x"70",
          7551 => x"81",
          7552 => x"8b",
          7553 => x"2b",
          7554 => x"70",
          7555 => x"33",
          7556 => x"07",
          7557 => x"8f",
          7558 => x"77",
          7559 => x"2a",
          7560 => x"5f",
          7561 => x"5e",
          7562 => x"17",
          7563 => x"17",
          7564 => x"b8",
          7565 => x"70",
          7566 => x"33",
          7567 => x"71",
          7568 => x"74",
          7569 => x"81",
          7570 => x"88",
          7571 => x"ff",
          7572 => x"88",
          7573 => x"5e",
          7574 => x"5d",
          7575 => x"34",
          7576 => x"34",
          7577 => x"08",
          7578 => x"11",
          7579 => x"33",
          7580 => x"71",
          7581 => x"74",
          7582 => x"33",
          7583 => x"71",
          7584 => x"83",
          7585 => x"05",
          7586 => x"85",
          7587 => x"88",
          7588 => x"88",
          7589 => x"49",
          7590 => x"59",
          7591 => x"57",
          7592 => x"1d",
          7593 => x"1d",
          7594 => x"b8",
          7595 => x"84",
          7596 => x"12",
          7597 => x"2b",
          7598 => x"07",
          7599 => x"14",
          7600 => x"33",
          7601 => x"07",
          7602 => x"5f",
          7603 => x"40",
          7604 => x"77",
          7605 => x"7b",
          7606 => x"84",
          7607 => x"16",
          7608 => x"12",
          7609 => x"2b",
          7610 => x"ff",
          7611 => x"2a",
          7612 => x"59",
          7613 => x"79",
          7614 => x"84",
          7615 => x"70",
          7616 => x"33",
          7617 => x"71",
          7618 => x"83",
          7619 => x"05",
          7620 => x"15",
          7621 => x"2b",
          7622 => x"2a",
          7623 => x"5d",
          7624 => x"55",
          7625 => x"75",
          7626 => x"84",
          7627 => x"70",
          7628 => x"81",
          7629 => x"8b",
          7630 => x"2b",
          7631 => x"82",
          7632 => x"15",
          7633 => x"2b",
          7634 => x"2a",
          7635 => x"5d",
          7636 => x"55",
          7637 => x"34",
          7638 => x"34",
          7639 => x"08",
          7640 => x"11",
          7641 => x"33",
          7642 => x"07",
          7643 => x"56",
          7644 => x"42",
          7645 => x"7e",
          7646 => x"51",
          7647 => x"3f",
          7648 => x"08",
          7649 => x"61",
          7650 => x"70",
          7651 => x"06",
          7652 => x"f1",
          7653 => x"19",
          7654 => x"33",
          7655 => x"71",
          7656 => x"79",
          7657 => x"33",
          7658 => x"71",
          7659 => x"70",
          7660 => x"48",
          7661 => x"55",
          7662 => x"05",
          7663 => x"85",
          7664 => x"b9",
          7665 => x"1e",
          7666 => x"85",
          7667 => x"8b",
          7668 => x"2b",
          7669 => x"86",
          7670 => x"15",
          7671 => x"2b",
          7672 => x"2a",
          7673 => x"48",
          7674 => x"56",
          7675 => x"05",
          7676 => x"87",
          7677 => x"b9",
          7678 => x"70",
          7679 => x"33",
          7680 => x"07",
          7681 => x"06",
          7682 => x"5c",
          7683 => x"78",
          7684 => x"81",
          7685 => x"b9",
          7686 => x"1f",
          7687 => x"12",
          7688 => x"2b",
          7689 => x"07",
          7690 => x"33",
          7691 => x"71",
          7692 => x"70",
          7693 => x"ff",
          7694 => x"05",
          7695 => x"5d",
          7696 => x"58",
          7697 => x"40",
          7698 => x"34",
          7699 => x"34",
          7700 => x"08",
          7701 => x"33",
          7702 => x"71",
          7703 => x"83",
          7704 => x"05",
          7705 => x"12",
          7706 => x"2b",
          7707 => x"ff",
          7708 => x"2a",
          7709 => x"58",
          7710 => x"5b",
          7711 => x"78",
          7712 => x"77",
          7713 => x"06",
          7714 => x"39",
          7715 => x"54",
          7716 => x"84",
          7717 => x"5f",
          7718 => x"08",
          7719 => x"38",
          7720 => x"52",
          7721 => x"08",
          7722 => x"be",
          7723 => x"df",
          7724 => x"5b",
          7725 => x"ef",
          7726 => x"e9",
          7727 => x"0d",
          7728 => x"84",
          7729 => x"58",
          7730 => x"2e",
          7731 => x"54",
          7732 => x"73",
          7733 => x"0c",
          7734 => x"04",
          7735 => x"d3",
          7736 => x"c8",
          7737 => x"b9",
          7738 => x"2e",
          7739 => x"53",
          7740 => x"b9",
          7741 => x"fe",
          7742 => x"73",
          7743 => x"0c",
          7744 => x"04",
          7745 => x"0b",
          7746 => x"0c",
          7747 => x"84",
          7748 => x"82",
          7749 => x"76",
          7750 => x"f4",
          7751 => x"df",
          7752 => x"b8",
          7753 => x"75",
          7754 => x"81",
          7755 => x"b9",
          7756 => x"76",
          7757 => x"81",
          7758 => x"34",
          7759 => x"08",
          7760 => x"17",
          7761 => x"87",
          7762 => x"b9",
          7763 => x"b9",
          7764 => x"05",
          7765 => x"07",
          7766 => x"ff",
          7767 => x"2a",
          7768 => x"56",
          7769 => x"34",
          7770 => x"34",
          7771 => x"22",
          7772 => x"10",
          7773 => x"08",
          7774 => x"55",
          7775 => x"15",
          7776 => x"83",
          7777 => x"54",
          7778 => x"fe",
          7779 => x"cc",
          7780 => x"0d",
          7781 => x"33",
          7782 => x"70",
          7783 => x"38",
          7784 => x"11",
          7785 => x"84",
          7786 => x"83",
          7787 => x"fe",
          7788 => x"93",
          7789 => x"83",
          7790 => x"26",
          7791 => x"51",
          7792 => x"84",
          7793 => x"81",
          7794 => x"72",
          7795 => x"84",
          7796 => x"34",
          7797 => x"12",
          7798 => x"84",
          7799 => x"84",
          7800 => x"f7",
          7801 => x"7e",
          7802 => x"05",
          7803 => x"5a",
          7804 => x"81",
          7805 => x"26",
          7806 => x"b9",
          7807 => x"54",
          7808 => x"54",
          7809 => x"bd",
          7810 => x"85",
          7811 => x"98",
          7812 => x"53",
          7813 => x"51",
          7814 => x"84",
          7815 => x"81",
          7816 => x"74",
          7817 => x"38",
          7818 => x"8c",
          7819 => x"e2",
          7820 => x"26",
          7821 => x"fc",
          7822 => x"54",
          7823 => x"83",
          7824 => x"73",
          7825 => x"b9",
          7826 => x"3d",
          7827 => x"80",
          7828 => x"70",
          7829 => x"5a",
          7830 => x"78",
          7831 => x"38",
          7832 => x"3d",
          7833 => x"60",
          7834 => x"af",
          7835 => x"5c",
          7836 => x"54",
          7837 => x"87",
          7838 => x"c4",
          7839 => x"73",
          7840 => x"83",
          7841 => x"38",
          7842 => x"0b",
          7843 => x"8c",
          7844 => x"75",
          7845 => x"d7",
          7846 => x"b9",
          7847 => x"ff",
          7848 => x"80",
          7849 => x"87",
          7850 => x"08",
          7851 => x"38",
          7852 => x"d6",
          7853 => x"80",
          7854 => x"73",
          7855 => x"38",
          7856 => x"55",
          7857 => x"c8",
          7858 => x"0d",
          7859 => x"16",
          7860 => x"81",
          7861 => x"55",
          7862 => x"26",
          7863 => x"d5",
          7864 => x"0d",
          7865 => x"05",
          7866 => x"02",
          7867 => x"05",
          7868 => x"55",
          7869 => x"73",
          7870 => x"84",
          7871 => x"33",
          7872 => x"06",
          7873 => x"73",
          7874 => x"0b",
          7875 => x"8c",
          7876 => x"70",
          7877 => x"38",
          7878 => x"ad",
          7879 => x"2e",
          7880 => x"53",
          7881 => x"c8",
          7882 => x"0d",
          7883 => x"0a",
          7884 => x"84",
          7885 => x"86",
          7886 => x"81",
          7887 => x"80",
          7888 => x"c8",
          7889 => x"0d",
          7890 => x"2b",
          7891 => x"8c",
          7892 => x"70",
          7893 => x"08",
          7894 => x"81",
          7895 => x"70",
          7896 => x"38",
          7897 => x"8c",
          7898 => x"ea",
          7899 => x"98",
          7900 => x"70",
          7901 => x"72",
          7902 => x"92",
          7903 => x"71",
          7904 => x"54",
          7905 => x"ff",
          7906 => x"08",
          7907 => x"73",
          7908 => x"90",
          7909 => x"0d",
          7910 => x"0b",
          7911 => x"71",
          7912 => x"74",
          7913 => x"81",
          7914 => x"77",
          7915 => x"83",
          7916 => x"38",
          7917 => x"52",
          7918 => x"51",
          7919 => x"84",
          7920 => x"80",
          7921 => x"81",
          7922 => x"b9",
          7923 => x"3d",
          7924 => x"54",
          7925 => x"53",
          7926 => x"53",
          7927 => x"52",
          7928 => x"3f",
          7929 => x"b9",
          7930 => x"2e",
          7931 => x"d9",
          7932 => x"c8",
          7933 => x"34",
          7934 => x"70",
          7935 => x"31",
          7936 => x"84",
          7937 => x"5c",
          7938 => x"74",
          7939 => x"9b",
          7940 => x"33",
          7941 => x"2e",
          7942 => x"ff",
          7943 => x"54",
          7944 => x"79",
          7945 => x"33",
          7946 => x"3f",
          7947 => x"57",
          7948 => x"2e",
          7949 => x"fe",
          7950 => x"18",
          7951 => x"81",
          7952 => x"06",
          7953 => x"b8",
          7954 => x"80",
          7955 => x"80",
          7956 => x"05",
          7957 => x"17",
          7958 => x"38",
          7959 => x"84",
          7960 => x"ff",
          7961 => x"b7",
          7962 => x"d2",
          7963 => x"d2",
          7964 => x"34",
          7965 => x"ba",
          7966 => x"c1",
          7967 => x"34",
          7968 => x"84",
          7969 => x"80",
          7970 => x"9d",
          7971 => x"c1",
          7972 => x"19",
          7973 => x"0b",
          7974 => x"34",
          7975 => x"55",
          7976 => x"19",
          7977 => x"2a",
          7978 => x"a1",
          7979 => x"90",
          7980 => x"84",
          7981 => x"74",
          7982 => x"7a",
          7983 => x"34",
          7984 => x"5b",
          7985 => x"19",
          7986 => x"2a",
          7987 => x"a5",
          7988 => x"90",
          7989 => x"84",
          7990 => x"7a",
          7991 => x"74",
          7992 => x"34",
          7993 => x"81",
          7994 => x"1a",
          7995 => x"54",
          7996 => x"52",
          7997 => x"51",
          7998 => x"76",
          7999 => x"80",
          8000 => x"81",
          8001 => x"fb",
          8002 => x"b9",
          8003 => x"2e",
          8004 => x"fd",
          8005 => x"3d",
          8006 => x"70",
          8007 => x"56",
          8008 => x"88",
          8009 => x"08",
          8010 => x"38",
          8011 => x"84",
          8012 => x"8f",
          8013 => x"ff",
          8014 => x"58",
          8015 => x"81",
          8016 => x"82",
          8017 => x"38",
          8018 => x"09",
          8019 => x"38",
          8020 => x"16",
          8021 => x"a8",
          8022 => x"5a",
          8023 => x"b4",
          8024 => x"2e",
          8025 => x"17",
          8026 => x"7b",
          8027 => x"06",
          8028 => x"81",
          8029 => x"b8",
          8030 => x"17",
          8031 => x"e3",
          8032 => x"c8",
          8033 => x"85",
          8034 => x"81",
          8035 => x"18",
          8036 => x"9a",
          8037 => x"ff",
          8038 => x"11",
          8039 => x"70",
          8040 => x"1b",
          8041 => x"5d",
          8042 => x"17",
          8043 => x"b5",
          8044 => x"83",
          8045 => x"5c",
          8046 => x"7d",
          8047 => x"06",
          8048 => x"81",
          8049 => x"b8",
          8050 => x"17",
          8051 => x"93",
          8052 => x"c8",
          8053 => x"85",
          8054 => x"81",
          8055 => x"18",
          8056 => x"ca",
          8057 => x"ff",
          8058 => x"11",
          8059 => x"2b",
          8060 => x"81",
          8061 => x"2a",
          8062 => x"59",
          8063 => x"ae",
          8064 => x"ff",
          8065 => x"c8",
          8066 => x"0d",
          8067 => x"2a",
          8068 => x"05",
          8069 => x"08",
          8070 => x"38",
          8071 => x"18",
          8072 => x"5d",
          8073 => x"2e",
          8074 => x"81",
          8075 => x"54",
          8076 => x"17",
          8077 => x"33",
          8078 => x"3f",
          8079 => x"08",
          8080 => x"38",
          8081 => x"5a",
          8082 => x"0c",
          8083 => x"38",
          8084 => x"fe",
          8085 => x"b8",
          8086 => x"33",
          8087 => x"88",
          8088 => x"b9",
          8089 => x"5b",
          8090 => x"04",
          8091 => x"09",
          8092 => x"b8",
          8093 => x"2a",
          8094 => x"05",
          8095 => x"08",
          8096 => x"38",
          8097 => x"18",
          8098 => x"5e",
          8099 => x"2e",
          8100 => x"82",
          8101 => x"54",
          8102 => x"17",
          8103 => x"33",
          8104 => x"3f",
          8105 => x"08",
          8106 => x"38",
          8107 => x"5a",
          8108 => x"0c",
          8109 => x"38",
          8110 => x"83",
          8111 => x"05",
          8112 => x"11",
          8113 => x"33",
          8114 => x"71",
          8115 => x"81",
          8116 => x"72",
          8117 => x"75",
          8118 => x"ff",
          8119 => x"06",
          8120 => x"c8",
          8121 => x"5e",
          8122 => x"8f",
          8123 => x"81",
          8124 => x"08",
          8125 => x"70",
          8126 => x"33",
          8127 => x"e2",
          8128 => x"84",
          8129 => x"7b",
          8130 => x"06",
          8131 => x"84",
          8132 => x"83",
          8133 => x"17",
          8134 => x"08",
          8135 => x"c8",
          8136 => x"7d",
          8137 => x"27",
          8138 => x"82",
          8139 => x"74",
          8140 => x"81",
          8141 => x"38",
          8142 => x"17",
          8143 => x"08",
          8144 => x"52",
          8145 => x"51",
          8146 => x"7a",
          8147 => x"39",
          8148 => x"17",
          8149 => x"17",
          8150 => x"18",
          8151 => x"f6",
          8152 => x"b9",
          8153 => x"2e",
          8154 => x"82",
          8155 => x"b9",
          8156 => x"18",
          8157 => x"08",
          8158 => x"31",
          8159 => x"18",
          8160 => x"38",
          8161 => x"5e",
          8162 => x"81",
          8163 => x"b9",
          8164 => x"fb",
          8165 => x"54",
          8166 => x"53",
          8167 => x"53",
          8168 => x"52",
          8169 => x"3f",
          8170 => x"b9",
          8171 => x"2e",
          8172 => x"fd",
          8173 => x"b9",
          8174 => x"18",
          8175 => x"08",
          8176 => x"31",
          8177 => x"08",
          8178 => x"a0",
          8179 => x"fd",
          8180 => x"17",
          8181 => x"82",
          8182 => x"06",
          8183 => x"81",
          8184 => x"08",
          8185 => x"05",
          8186 => x"81",
          8187 => x"f4",
          8188 => x"5a",
          8189 => x"81",
          8190 => x"08",
          8191 => x"70",
          8192 => x"33",
          8193 => x"da",
          8194 => x"84",
          8195 => x"7d",
          8196 => x"06",
          8197 => x"84",
          8198 => x"83",
          8199 => x"17",
          8200 => x"08",
          8201 => x"c8",
          8202 => x"74",
          8203 => x"27",
          8204 => x"82",
          8205 => x"74",
          8206 => x"81",
          8207 => x"38",
          8208 => x"17",
          8209 => x"08",
          8210 => x"52",
          8211 => x"51",
          8212 => x"7c",
          8213 => x"39",
          8214 => x"17",
          8215 => x"08",
          8216 => x"52",
          8217 => x"51",
          8218 => x"fa",
          8219 => x"5b",
          8220 => x"38",
          8221 => x"f2",
          8222 => x"62",
          8223 => x"59",
          8224 => x"76",
          8225 => x"75",
          8226 => x"27",
          8227 => x"33",
          8228 => x"2e",
          8229 => x"78",
          8230 => x"38",
          8231 => x"82",
          8232 => x"84",
          8233 => x"90",
          8234 => x"75",
          8235 => x"1a",
          8236 => x"80",
          8237 => x"08",
          8238 => x"78",
          8239 => x"38",
          8240 => x"7c",
          8241 => x"7c",
          8242 => x"06",
          8243 => x"81",
          8244 => x"b8",
          8245 => x"19",
          8246 => x"87",
          8247 => x"c8",
          8248 => x"85",
          8249 => x"81",
          8250 => x"1a",
          8251 => x"79",
          8252 => x"75",
          8253 => x"06",
          8254 => x"83",
          8255 => x"58",
          8256 => x"1f",
          8257 => x"2a",
          8258 => x"1f",
          8259 => x"83",
          8260 => x"84",
          8261 => x"90",
          8262 => x"74",
          8263 => x"81",
          8264 => x"38",
          8265 => x"a8",
          8266 => x"58",
          8267 => x"1a",
          8268 => x"76",
          8269 => x"e1",
          8270 => x"33",
          8271 => x"7c",
          8272 => x"81",
          8273 => x"38",
          8274 => x"53",
          8275 => x"81",
          8276 => x"f1",
          8277 => x"b9",
          8278 => x"2e",
          8279 => x"58",
          8280 => x"b4",
          8281 => x"58",
          8282 => x"38",
          8283 => x"83",
          8284 => x"05",
          8285 => x"11",
          8286 => x"2b",
          8287 => x"7e",
          8288 => x"07",
          8289 => x"5c",
          8290 => x"7d",
          8291 => x"75",
          8292 => x"7d",
          8293 => x"79",
          8294 => x"7d",
          8295 => x"7a",
          8296 => x"81",
          8297 => x"34",
          8298 => x"75",
          8299 => x"70",
          8300 => x"1b",
          8301 => x"1b",
          8302 => x"5a",
          8303 => x"b7",
          8304 => x"83",
          8305 => x"5e",
          8306 => x"7d",
          8307 => x"06",
          8308 => x"81",
          8309 => x"b8",
          8310 => x"19",
          8311 => x"83",
          8312 => x"c8",
          8313 => x"85",
          8314 => x"81",
          8315 => x"1a",
          8316 => x"7b",
          8317 => x"79",
          8318 => x"19",
          8319 => x"1b",
          8320 => x"5f",
          8321 => x"55",
          8322 => x"8f",
          8323 => x"2b",
          8324 => x"77",
          8325 => x"71",
          8326 => x"74",
          8327 => x"0b",
          8328 => x"7d",
          8329 => x"1a",
          8330 => x"80",
          8331 => x"08",
          8332 => x"76",
          8333 => x"38",
          8334 => x"53",
          8335 => x"53",
          8336 => x"52",
          8337 => x"3f",
          8338 => x"b9",
          8339 => x"2e",
          8340 => x"80",
          8341 => x"b9",
          8342 => x"1a",
          8343 => x"08",
          8344 => x"08",
          8345 => x"08",
          8346 => x"08",
          8347 => x"5c",
          8348 => x"8b",
          8349 => x"33",
          8350 => x"2e",
          8351 => x"81",
          8352 => x"76",
          8353 => x"33",
          8354 => x"3f",
          8355 => x"08",
          8356 => x"38",
          8357 => x"58",
          8358 => x"0c",
          8359 => x"38",
          8360 => x"06",
          8361 => x"7b",
          8362 => x"56",
          8363 => x"7a",
          8364 => x"33",
          8365 => x"71",
          8366 => x"56",
          8367 => x"34",
          8368 => x"1a",
          8369 => x"39",
          8370 => x"53",
          8371 => x"53",
          8372 => x"52",
          8373 => x"3f",
          8374 => x"b9",
          8375 => x"2e",
          8376 => x"fc",
          8377 => x"b9",
          8378 => x"1a",
          8379 => x"08",
          8380 => x"08",
          8381 => x"08",
          8382 => x"08",
          8383 => x"5e",
          8384 => x"fb",
          8385 => x"19",
          8386 => x"82",
          8387 => x"06",
          8388 => x"81",
          8389 => x"53",
          8390 => x"19",
          8391 => x"c2",
          8392 => x"fb",
          8393 => x"54",
          8394 => x"19",
          8395 => x"1a",
          8396 => x"ee",
          8397 => x"5c",
          8398 => x"08",
          8399 => x"81",
          8400 => x"38",
          8401 => x"08",
          8402 => x"b4",
          8403 => x"a8",
          8404 => x"a0",
          8405 => x"b9",
          8406 => x"40",
          8407 => x"7e",
          8408 => x"38",
          8409 => x"55",
          8410 => x"09",
          8411 => x"e3",
          8412 => x"7d",
          8413 => x"52",
          8414 => x"51",
          8415 => x"7c",
          8416 => x"39",
          8417 => x"53",
          8418 => x"53",
          8419 => x"52",
          8420 => x"3f",
          8421 => x"b9",
          8422 => x"2e",
          8423 => x"fb",
          8424 => x"b9",
          8425 => x"1a",
          8426 => x"08",
          8427 => x"08",
          8428 => x"08",
          8429 => x"08",
          8430 => x"5e",
          8431 => x"fb",
          8432 => x"19",
          8433 => x"82",
          8434 => x"06",
          8435 => x"81",
          8436 => x"53",
          8437 => x"19",
          8438 => x"86",
          8439 => x"fa",
          8440 => x"54",
          8441 => x"76",
          8442 => x"33",
          8443 => x"3f",
          8444 => x"8b",
          8445 => x"10",
          8446 => x"7a",
          8447 => x"ff",
          8448 => x"5f",
          8449 => x"1f",
          8450 => x"2a",
          8451 => x"1f",
          8452 => x"39",
          8453 => x"88",
          8454 => x"82",
          8455 => x"06",
          8456 => x"11",
          8457 => x"70",
          8458 => x"0a",
          8459 => x"0a",
          8460 => x"58",
          8461 => x"7d",
          8462 => x"88",
          8463 => x"b9",
          8464 => x"90",
          8465 => x"ba",
          8466 => x"98",
          8467 => x"bb",
          8468 => x"cf",
          8469 => x"0d",
          8470 => x"08",
          8471 => x"7a",
          8472 => x"90",
          8473 => x"76",
          8474 => x"f4",
          8475 => x"1a",
          8476 => x"ec",
          8477 => x"08",
          8478 => x"73",
          8479 => x"d7",
          8480 => x"2e",
          8481 => x"76",
          8482 => x"56",
          8483 => x"76",
          8484 => x"82",
          8485 => x"26",
          8486 => x"75",
          8487 => x"f0",
          8488 => x"b9",
          8489 => x"2e",
          8490 => x"80",
          8491 => x"c8",
          8492 => x"b1",
          8493 => x"c8",
          8494 => x"30",
          8495 => x"80",
          8496 => x"07",
          8497 => x"55",
          8498 => x"38",
          8499 => x"09",
          8500 => x"b5",
          8501 => x"74",
          8502 => x"0c",
          8503 => x"04",
          8504 => x"91",
          8505 => x"c8",
          8506 => x"39",
          8507 => x"51",
          8508 => x"81",
          8509 => x"b9",
          8510 => x"db",
          8511 => x"c8",
          8512 => x"b9",
          8513 => x"2e",
          8514 => x"19",
          8515 => x"c8",
          8516 => x"38",
          8517 => x"dd",
          8518 => x"56",
          8519 => x"76",
          8520 => x"82",
          8521 => x"79",
          8522 => x"3f",
          8523 => x"b9",
          8524 => x"2e",
          8525 => x"84",
          8526 => x"09",
          8527 => x"72",
          8528 => x"70",
          8529 => x"b9",
          8530 => x"51",
          8531 => x"73",
          8532 => x"84",
          8533 => x"80",
          8534 => x"90",
          8535 => x"81",
          8536 => x"a3",
          8537 => x"1a",
          8538 => x"9b",
          8539 => x"57",
          8540 => x"39",
          8541 => x"fe",
          8542 => x"53",
          8543 => x"51",
          8544 => x"84",
          8545 => x"84",
          8546 => x"30",
          8547 => x"c8",
          8548 => x"25",
          8549 => x"7a",
          8550 => x"74",
          8551 => x"75",
          8552 => x"9c",
          8553 => x"05",
          8554 => x"56",
          8555 => x"26",
          8556 => x"15",
          8557 => x"84",
          8558 => x"07",
          8559 => x"1a",
          8560 => x"74",
          8561 => x"0c",
          8562 => x"04",
          8563 => x"b9",
          8564 => x"3d",
          8565 => x"b9",
          8566 => x"fe",
          8567 => x"80",
          8568 => x"38",
          8569 => x"52",
          8570 => x"8b",
          8571 => x"c8",
          8572 => x"a7",
          8573 => x"c8",
          8574 => x"c8",
          8575 => x"0d",
          8576 => x"74",
          8577 => x"b9",
          8578 => x"ff",
          8579 => x"3d",
          8580 => x"71",
          8581 => x"58",
          8582 => x"0a",
          8583 => x"38",
          8584 => x"53",
          8585 => x"38",
          8586 => x"0c",
          8587 => x"55",
          8588 => x"38",
          8589 => x"75",
          8590 => x"cc",
          8591 => x"2a",
          8592 => x"88",
          8593 => x"56",
          8594 => x"a9",
          8595 => x"08",
          8596 => x"74",
          8597 => x"98",
          8598 => x"82",
          8599 => x"2e",
          8600 => x"89",
          8601 => x"19",
          8602 => x"ff",
          8603 => x"05",
          8604 => x"80",
          8605 => x"b9",
          8606 => x"3d",
          8607 => x"0b",
          8608 => x"0c",
          8609 => x"04",
          8610 => x"55",
          8611 => x"ff",
          8612 => x"17",
          8613 => x"2b",
          8614 => x"76",
          8615 => x"9c",
          8616 => x"fe",
          8617 => x"54",
          8618 => x"75",
          8619 => x"38",
          8620 => x"76",
          8621 => x"19",
          8622 => x"53",
          8623 => x"0c",
          8624 => x"74",
          8625 => x"ec",
          8626 => x"b9",
          8627 => x"84",
          8628 => x"ff",
          8629 => x"81",
          8630 => x"c8",
          8631 => x"9e",
          8632 => x"08",
          8633 => x"c8",
          8634 => x"ff",
          8635 => x"76",
          8636 => x"76",
          8637 => x"ff",
          8638 => x"0b",
          8639 => x"0c",
          8640 => x"04",
          8641 => x"7f",
          8642 => x"12",
          8643 => x"5c",
          8644 => x"80",
          8645 => x"86",
          8646 => x"98",
          8647 => x"17",
          8648 => x"56",
          8649 => x"b2",
          8650 => x"ff",
          8651 => x"9d",
          8652 => x"94",
          8653 => x"58",
          8654 => x"79",
          8655 => x"1a",
          8656 => x"74",
          8657 => x"f5",
          8658 => x"18",
          8659 => x"18",
          8660 => x"b8",
          8661 => x"0c",
          8662 => x"84",
          8663 => x"8f",
          8664 => x"77",
          8665 => x"8a",
          8666 => x"05",
          8667 => x"06",
          8668 => x"38",
          8669 => x"51",
          8670 => x"84",
          8671 => x"5d",
          8672 => x"0b",
          8673 => x"08",
          8674 => x"81",
          8675 => x"c8",
          8676 => x"c6",
          8677 => x"08",
          8678 => x"08",
          8679 => x"38",
          8680 => x"81",
          8681 => x"17",
          8682 => x"51",
          8683 => x"84",
          8684 => x"5d",
          8685 => x"b9",
          8686 => x"2e",
          8687 => x"82",
          8688 => x"c8",
          8689 => x"ff",
          8690 => x"56",
          8691 => x"08",
          8692 => x"86",
          8693 => x"c8",
          8694 => x"33",
          8695 => x"80",
          8696 => x"18",
          8697 => x"fe",
          8698 => x"80",
          8699 => x"27",
          8700 => x"19",
          8701 => x"29",
          8702 => x"05",
          8703 => x"b4",
          8704 => x"19",
          8705 => x"78",
          8706 => x"76",
          8707 => x"58",
          8708 => x"55",
          8709 => x"74",
          8710 => x"22",
          8711 => x"27",
          8712 => x"81",
          8713 => x"53",
          8714 => x"19",
          8715 => x"b2",
          8716 => x"c8",
          8717 => x"38",
          8718 => x"dd",
          8719 => x"18",
          8720 => x"84",
          8721 => x"8f",
          8722 => x"75",
          8723 => x"08",
          8724 => x"70",
          8725 => x"33",
          8726 => x"86",
          8727 => x"c8",
          8728 => x"38",
          8729 => x"08",
          8730 => x"b4",
          8731 => x"1a",
          8732 => x"74",
          8733 => x"27",
          8734 => x"82",
          8735 => x"7b",
          8736 => x"81",
          8737 => x"38",
          8738 => x"19",
          8739 => x"08",
          8740 => x"52",
          8741 => x"51",
          8742 => x"fe",
          8743 => x"19",
          8744 => x"83",
          8745 => x"55",
          8746 => x"09",
          8747 => x"38",
          8748 => x"0c",
          8749 => x"1a",
          8750 => x"5e",
          8751 => x"75",
          8752 => x"85",
          8753 => x"22",
          8754 => x"b0",
          8755 => x"98",
          8756 => x"fc",
          8757 => x"0b",
          8758 => x"0c",
          8759 => x"04",
          8760 => x"64",
          8761 => x"84",
          8762 => x"5b",
          8763 => x"98",
          8764 => x"5e",
          8765 => x"2e",
          8766 => x"b8",
          8767 => x"5a",
          8768 => x"19",
          8769 => x"82",
          8770 => x"19",
          8771 => x"55",
          8772 => x"09",
          8773 => x"94",
          8774 => x"75",
          8775 => x"52",
          8776 => x"51",
          8777 => x"84",
          8778 => x"80",
          8779 => x"ff",
          8780 => x"79",
          8781 => x"76",
          8782 => x"90",
          8783 => x"08",
          8784 => x"58",
          8785 => x"82",
          8786 => x"18",
          8787 => x"70",
          8788 => x"5b",
          8789 => x"1d",
          8790 => x"e5",
          8791 => x"78",
          8792 => x"30",
          8793 => x"71",
          8794 => x"54",
          8795 => x"55",
          8796 => x"74",
          8797 => x"43",
          8798 => x"2e",
          8799 => x"75",
          8800 => x"86",
          8801 => x"5d",
          8802 => x"51",
          8803 => x"84",
          8804 => x"5b",
          8805 => x"08",
          8806 => x"98",
          8807 => x"75",
          8808 => x"7a",
          8809 => x"0c",
          8810 => x"04",
          8811 => x"19",
          8812 => x"52",
          8813 => x"51",
          8814 => x"81",
          8815 => x"c8",
          8816 => x"09",
          8817 => x"ef",
          8818 => x"c8",
          8819 => x"34",
          8820 => x"a8",
          8821 => x"84",
          8822 => x"58",
          8823 => x"1a",
          8824 => x"b5",
          8825 => x"33",
          8826 => x"2e",
          8827 => x"fe",
          8828 => x"54",
          8829 => x"a0",
          8830 => x"53",
          8831 => x"19",
          8832 => x"de",
          8833 => x"fe",
          8834 => x"8f",
          8835 => x"06",
          8836 => x"76",
          8837 => x"06",
          8838 => x"2e",
          8839 => x"18",
          8840 => x"bf",
          8841 => x"1f",
          8842 => x"05",
          8843 => x"5e",
          8844 => x"ab",
          8845 => x"55",
          8846 => x"cc",
          8847 => x"75",
          8848 => x"81",
          8849 => x"38",
          8850 => x"5b",
          8851 => x"1d",
          8852 => x"b9",
          8853 => x"3d",
          8854 => x"5b",
          8855 => x"8d",
          8856 => x"7d",
          8857 => x"81",
          8858 => x"8c",
          8859 => x"19",
          8860 => x"33",
          8861 => x"07",
          8862 => x"75",
          8863 => x"77",
          8864 => x"bf",
          8865 => x"f3",
          8866 => x"81",
          8867 => x"83",
          8868 => x"33",
          8869 => x"11",
          8870 => x"71",
          8871 => x"52",
          8872 => x"80",
          8873 => x"38",
          8874 => x"26",
          8875 => x"79",
          8876 => x"76",
          8877 => x"62",
          8878 => x"5a",
          8879 => x"8c",
          8880 => x"38",
          8881 => x"86",
          8882 => x"59",
          8883 => x"2e",
          8884 => x"81",
          8885 => x"dd",
          8886 => x"61",
          8887 => x"63",
          8888 => x"70",
          8889 => x"5e",
          8890 => x"39",
          8891 => x"ff",
          8892 => x"81",
          8893 => x"c0",
          8894 => x"38",
          8895 => x"57",
          8896 => x"75",
          8897 => x"05",
          8898 => x"05",
          8899 => x"7f",
          8900 => x"ff",
          8901 => x"59",
          8902 => x"e4",
          8903 => x"2e",
          8904 => x"ff",
          8905 => x"0c",
          8906 => x"c8",
          8907 => x"0d",
          8908 => x"0d",
          8909 => x"5c",
          8910 => x"7b",
          8911 => x"3f",
          8912 => x"08",
          8913 => x"c8",
          8914 => x"38",
          8915 => x"40",
          8916 => x"ac",
          8917 => x"1b",
          8918 => x"08",
          8919 => x"b4",
          8920 => x"2e",
          8921 => x"83",
          8922 => x"58",
          8923 => x"2e",
          8924 => x"81",
          8925 => x"54",
          8926 => x"1b",
          8927 => x"33",
          8928 => x"3f",
          8929 => x"08",
          8930 => x"38",
          8931 => x"57",
          8932 => x"0c",
          8933 => x"81",
          8934 => x"1c",
          8935 => x"58",
          8936 => x"2e",
          8937 => x"8b",
          8938 => x"06",
          8939 => x"06",
          8940 => x"86",
          8941 => x"81",
          8942 => x"f2",
          8943 => x"2a",
          8944 => x"75",
          8945 => x"ef",
          8946 => x"e2",
          8947 => x"2e",
          8948 => x"7c",
          8949 => x"7d",
          8950 => x"57",
          8951 => x"75",
          8952 => x"05",
          8953 => x"05",
          8954 => x"76",
          8955 => x"ff",
          8956 => x"59",
          8957 => x"e4",
          8958 => x"2e",
          8959 => x"ab",
          8960 => x"06",
          8961 => x"38",
          8962 => x"1d",
          8963 => x"70",
          8964 => x"33",
          8965 => x"05",
          8966 => x"71",
          8967 => x"5a",
          8968 => x"76",
          8969 => x"dc",
          8970 => x"2e",
          8971 => x"ff",
          8972 => x"ac",
          8973 => x"52",
          8974 => x"c8",
          8975 => x"c8",
          8976 => x"b9",
          8977 => x"2e",
          8978 => x"79",
          8979 => x"0c",
          8980 => x"04",
          8981 => x"1b",
          8982 => x"52",
          8983 => x"51",
          8984 => x"81",
          8985 => x"c8",
          8986 => x"09",
          8987 => x"a4",
          8988 => x"c8",
          8989 => x"34",
          8990 => x"a8",
          8991 => x"84",
          8992 => x"58",
          8993 => x"1c",
          8994 => x"ea",
          8995 => x"33",
          8996 => x"2e",
          8997 => x"fd",
          8998 => x"54",
          8999 => x"a0",
          9000 => x"53",
          9001 => x"1b",
          9002 => x"b6",
          9003 => x"fd",
          9004 => x"5a",
          9005 => x"ab",
          9006 => x"86",
          9007 => x"42",
          9008 => x"f2",
          9009 => x"2a",
          9010 => x"79",
          9011 => x"38",
          9012 => x"77",
          9013 => x"70",
          9014 => x"7f",
          9015 => x"59",
          9016 => x"7d",
          9017 => x"81",
          9018 => x"5d",
          9019 => x"51",
          9020 => x"84",
          9021 => x"5a",
          9022 => x"08",
          9023 => x"d9",
          9024 => x"39",
          9025 => x"fe",
          9026 => x"ff",
          9027 => x"ac",
          9028 => x"a2",
          9029 => x"33",
          9030 => x"2e",
          9031 => x"c7",
          9032 => x"08",
          9033 => x"9a",
          9034 => x"88",
          9035 => x"42",
          9036 => x"b3",
          9037 => x"70",
          9038 => x"29",
          9039 => x"55",
          9040 => x"56",
          9041 => x"18",
          9042 => x"81",
          9043 => x"33",
          9044 => x"07",
          9045 => x"75",
          9046 => x"ed",
          9047 => x"fe",
          9048 => x"38",
          9049 => x"a1",
          9050 => x"b9",
          9051 => x"10",
          9052 => x"22",
          9053 => x"1b",
          9054 => x"a0",
          9055 => x"84",
          9056 => x"2e",
          9057 => x"fe",
          9058 => x"56",
          9059 => x"8c",
          9060 => x"b0",
          9061 => x"70",
          9062 => x"06",
          9063 => x"80",
          9064 => x"74",
          9065 => x"38",
          9066 => x"05",
          9067 => x"41",
          9068 => x"38",
          9069 => x"81",
          9070 => x"5a",
          9071 => x"84",
          9072 => x"c8",
          9073 => x"0d",
          9074 => x"ff",
          9075 => x"bc",
          9076 => x"55",
          9077 => x"ea",
          9078 => x"70",
          9079 => x"13",
          9080 => x"06",
          9081 => x"5e",
          9082 => x"85",
          9083 => x"8c",
          9084 => x"22",
          9085 => x"74",
          9086 => x"38",
          9087 => x"10",
          9088 => x"51",
          9089 => x"f4",
          9090 => x"a0",
          9091 => x"8c",
          9092 => x"58",
          9093 => x"81",
          9094 => x"77",
          9095 => x"59",
          9096 => x"55",
          9097 => x"02",
          9098 => x"33",
          9099 => x"58",
          9100 => x"2e",
          9101 => x"80",
          9102 => x"1f",
          9103 => x"94",
          9104 => x"8c",
          9105 => x"58",
          9106 => x"61",
          9107 => x"77",
          9108 => x"59",
          9109 => x"81",
          9110 => x"ff",
          9111 => x"ef",
          9112 => x"27",
          9113 => x"7a",
          9114 => x"57",
          9115 => x"b8",
          9116 => x"1a",
          9117 => x"58",
          9118 => x"77",
          9119 => x"81",
          9120 => x"ff",
          9121 => x"90",
          9122 => x"44",
          9123 => x"60",
          9124 => x"38",
          9125 => x"a1",
          9126 => x"18",
          9127 => x"25",
          9128 => x"22",
          9129 => x"38",
          9130 => x"05",
          9131 => x"57",
          9132 => x"07",
          9133 => x"b9",
          9134 => x"38",
          9135 => x"74",
          9136 => x"16",
          9137 => x"84",
          9138 => x"56",
          9139 => x"77",
          9140 => x"fe",
          9141 => x"7a",
          9142 => x"78",
          9143 => x"79",
          9144 => x"a0",
          9145 => x"81",
          9146 => x"78",
          9147 => x"38",
          9148 => x"33",
          9149 => x"a0",
          9150 => x"06",
          9151 => x"16",
          9152 => x"77",
          9153 => x"38",
          9154 => x"05",
          9155 => x"19",
          9156 => x"59",
          9157 => x"34",
          9158 => x"87",
          9159 => x"51",
          9160 => x"84",
          9161 => x"8b",
          9162 => x"5b",
          9163 => x"27",
          9164 => x"87",
          9165 => x"e4",
          9166 => x"38",
          9167 => x"08",
          9168 => x"c8",
          9169 => x"09",
          9170 => x"d6",
          9171 => x"db",
          9172 => x"1f",
          9173 => x"02",
          9174 => x"db",
          9175 => x"58",
          9176 => x"81",
          9177 => x"5b",
          9178 => x"90",
          9179 => x"8c",
          9180 => x"8a",
          9181 => x"b9",
          9182 => x"5b",
          9183 => x"51",
          9184 => x"84",
          9185 => x"56",
          9186 => x"08",
          9187 => x"84",
          9188 => x"b8",
          9189 => x"98",
          9190 => x"80",
          9191 => x"08",
          9192 => x"f3",
          9193 => x"33",
          9194 => x"2e",
          9195 => x"82",
          9196 => x"54",
          9197 => x"18",
          9198 => x"33",
          9199 => x"3f",
          9200 => x"08",
          9201 => x"38",
          9202 => x"57",
          9203 => x"0c",
          9204 => x"bc",
          9205 => x"08",
          9206 => x"42",
          9207 => x"2e",
          9208 => x"74",
          9209 => x"25",
          9210 => x"5f",
          9211 => x"81",
          9212 => x"19",
          9213 => x"2e",
          9214 => x"81",
          9215 => x"ee",
          9216 => x"b9",
          9217 => x"84",
          9218 => x"80",
          9219 => x"38",
          9220 => x"84",
          9221 => x"38",
          9222 => x"81",
          9223 => x"1b",
          9224 => x"f3",
          9225 => x"08",
          9226 => x"08",
          9227 => x"38",
          9228 => x"78",
          9229 => x"84",
          9230 => x"54",
          9231 => x"1c",
          9232 => x"33",
          9233 => x"3f",
          9234 => x"08",
          9235 => x"38",
          9236 => x"56",
          9237 => x"0c",
          9238 => x"80",
          9239 => x"0b",
          9240 => x"57",
          9241 => x"70",
          9242 => x"34",
          9243 => x"74",
          9244 => x"0b",
          9245 => x"7b",
          9246 => x"75",
          9247 => x"57",
          9248 => x"81",
          9249 => x"ff",
          9250 => x"ef",
          9251 => x"08",
          9252 => x"98",
          9253 => x"7c",
          9254 => x"81",
          9255 => x"34",
          9256 => x"84",
          9257 => x"98",
          9258 => x"81",
          9259 => x"80",
          9260 => x"57",
          9261 => x"fe",
          9262 => x"59",
          9263 => x"51",
          9264 => x"84",
          9265 => x"56",
          9266 => x"08",
          9267 => x"c7",
          9268 => x"39",
          9269 => x"18",
          9270 => x"52",
          9271 => x"51",
          9272 => x"84",
          9273 => x"77",
          9274 => x"06",
          9275 => x"84",
          9276 => x"83",
          9277 => x"18",
          9278 => x"08",
          9279 => x"a0",
          9280 => x"8b",
          9281 => x"33",
          9282 => x"2e",
          9283 => x"84",
          9284 => x"57",
          9285 => x"7f",
          9286 => x"1f",
          9287 => x"53",
          9288 => x"e9",
          9289 => x"b9",
          9290 => x"84",
          9291 => x"fe",
          9292 => x"84",
          9293 => x"56",
          9294 => x"74",
          9295 => x"81",
          9296 => x"78",
          9297 => x"5a",
          9298 => x"05",
          9299 => x"06",
          9300 => x"56",
          9301 => x"38",
          9302 => x"06",
          9303 => x"41",
          9304 => x"57",
          9305 => x"1c",
          9306 => x"b2",
          9307 => x"33",
          9308 => x"2e",
          9309 => x"82",
          9310 => x"54",
          9311 => x"1c",
          9312 => x"33",
          9313 => x"3f",
          9314 => x"08",
          9315 => x"38",
          9316 => x"56",
          9317 => x"0c",
          9318 => x"fe",
          9319 => x"1c",
          9320 => x"08",
          9321 => x"06",
          9322 => x"60",
          9323 => x"8f",
          9324 => x"34",
          9325 => x"34",
          9326 => x"34",
          9327 => x"34",
          9328 => x"f3",
          9329 => x"5a",
          9330 => x"83",
          9331 => x"8b",
          9332 => x"1f",
          9333 => x"1b",
          9334 => x"83",
          9335 => x"33",
          9336 => x"76",
          9337 => x"05",
          9338 => x"88",
          9339 => x"75",
          9340 => x"38",
          9341 => x"57",
          9342 => x"8c",
          9343 => x"38",
          9344 => x"ff",
          9345 => x"38",
          9346 => x"70",
          9347 => x"76",
          9348 => x"a6",
          9349 => x"34",
          9350 => x"1d",
          9351 => x"7d",
          9352 => x"3f",
          9353 => x"08",
          9354 => x"c8",
          9355 => x"38",
          9356 => x"40",
          9357 => x"38",
          9358 => x"81",
          9359 => x"08",
          9360 => x"70",
          9361 => x"33",
          9362 => x"96",
          9363 => x"84",
          9364 => x"fc",
          9365 => x"b9",
          9366 => x"1d",
          9367 => x"08",
          9368 => x"31",
          9369 => x"08",
          9370 => x"a0",
          9371 => x"fb",
          9372 => x"1c",
          9373 => x"82",
          9374 => x"06",
          9375 => x"81",
          9376 => x"08",
          9377 => x"05",
          9378 => x"81",
          9379 => x"cf",
          9380 => x"56",
          9381 => x"76",
          9382 => x"70",
          9383 => x"56",
          9384 => x"2e",
          9385 => x"fa",
          9386 => x"ff",
          9387 => x"57",
          9388 => x"2e",
          9389 => x"fa",
          9390 => x"80",
          9391 => x"fe",
          9392 => x"54",
          9393 => x"53",
          9394 => x"1c",
          9395 => x"92",
          9396 => x"c8",
          9397 => x"09",
          9398 => x"38",
          9399 => x"08",
          9400 => x"b4",
          9401 => x"1d",
          9402 => x"74",
          9403 => x"27",
          9404 => x"1c",
          9405 => x"82",
          9406 => x"84",
          9407 => x"56",
          9408 => x"75",
          9409 => x"58",
          9410 => x"fa",
          9411 => x"87",
          9412 => x"57",
          9413 => x"81",
          9414 => x"75",
          9415 => x"fe",
          9416 => x"39",
          9417 => x"1c",
          9418 => x"08",
          9419 => x"52",
          9420 => x"51",
          9421 => x"fc",
          9422 => x"54",
          9423 => x"a0",
          9424 => x"53",
          9425 => x"18",
          9426 => x"96",
          9427 => x"39",
          9428 => x"7f",
          9429 => x"40",
          9430 => x"0b",
          9431 => x"98",
          9432 => x"2e",
          9433 => x"ac",
          9434 => x"2e",
          9435 => x"80",
          9436 => x"8c",
          9437 => x"22",
          9438 => x"5c",
          9439 => x"2e",
          9440 => x"54",
          9441 => x"22",
          9442 => x"55",
          9443 => x"95",
          9444 => x"80",
          9445 => x"ff",
          9446 => x"5a",
          9447 => x"26",
          9448 => x"73",
          9449 => x"11",
          9450 => x"58",
          9451 => x"d4",
          9452 => x"70",
          9453 => x"30",
          9454 => x"5c",
          9455 => x"94",
          9456 => x"0b",
          9457 => x"80",
          9458 => x"59",
          9459 => x"1c",
          9460 => x"33",
          9461 => x"56",
          9462 => x"2e",
          9463 => x"85",
          9464 => x"38",
          9465 => x"70",
          9466 => x"07",
          9467 => x"5b",
          9468 => x"26",
          9469 => x"80",
          9470 => x"ae",
          9471 => x"05",
          9472 => x"18",
          9473 => x"70",
          9474 => x"34",
          9475 => x"8a",
          9476 => x"ba",
          9477 => x"88",
          9478 => x"0b",
          9479 => x"96",
          9480 => x"72",
          9481 => x"81",
          9482 => x"0b",
          9483 => x"81",
          9484 => x"94",
          9485 => x"0b",
          9486 => x"9c",
          9487 => x"11",
          9488 => x"73",
          9489 => x"89",
          9490 => x"1c",
          9491 => x"13",
          9492 => x"34",
          9493 => x"9c",
          9494 => x"33",
          9495 => x"71",
          9496 => x"88",
          9497 => x"14",
          9498 => x"07",
          9499 => x"33",
          9500 => x"0c",
          9501 => x"33",
          9502 => x"71",
          9503 => x"5f",
          9504 => x"5a",
          9505 => x"77",
          9506 => x"99",
          9507 => x"16",
          9508 => x"2b",
          9509 => x"7b",
          9510 => x"8f",
          9511 => x"81",
          9512 => x"c0",
          9513 => x"96",
          9514 => x"7a",
          9515 => x"57",
          9516 => x"7a",
          9517 => x"07",
          9518 => x"89",
          9519 => x"c8",
          9520 => x"ff",
          9521 => x"ff",
          9522 => x"38",
          9523 => x"81",
          9524 => x"88",
          9525 => x"7a",
          9526 => x"18",
          9527 => x"05",
          9528 => x"8c",
          9529 => x"5b",
          9530 => x"11",
          9531 => x"57",
          9532 => x"90",
          9533 => x"39",
          9534 => x"30",
          9535 => x"80",
          9536 => x"25",
          9537 => x"57",
          9538 => x"38",
          9539 => x"81",
          9540 => x"80",
          9541 => x"08",
          9542 => x"39",
          9543 => x"1f",
          9544 => x"57",
          9545 => x"fe",
          9546 => x"96",
          9547 => x"59",
          9548 => x"33",
          9549 => x"5a",
          9550 => x"26",
          9551 => x"1c",
          9552 => x"33",
          9553 => x"76",
          9554 => x"72",
          9555 => x"72",
          9556 => x"7d",
          9557 => x"38",
          9558 => x"83",
          9559 => x"55",
          9560 => x"70",
          9561 => x"34",
          9562 => x"16",
          9563 => x"89",
          9564 => x"57",
          9565 => x"79",
          9566 => x"fd",
          9567 => x"83",
          9568 => x"39",
          9569 => x"70",
          9570 => x"30",
          9571 => x"5d",
          9572 => x"a9",
          9573 => x"0d",
          9574 => x"70",
          9575 => x"80",
          9576 => x"57",
          9577 => x"af",
          9578 => x"81",
          9579 => x"dc",
          9580 => x"38",
          9581 => x"81",
          9582 => x"16",
          9583 => x"0c",
          9584 => x"3d",
          9585 => x"42",
          9586 => x"27",
          9587 => x"73",
          9588 => x"08",
          9589 => x"61",
          9590 => x"05",
          9591 => x"53",
          9592 => x"38",
          9593 => x"73",
          9594 => x"ec",
          9595 => x"ff",
          9596 => x"38",
          9597 => x"56",
          9598 => x"81",
          9599 => x"83",
          9600 => x"70",
          9601 => x"30",
          9602 => x"71",
          9603 => x"57",
          9604 => x"73",
          9605 => x"74",
          9606 => x"82",
          9607 => x"80",
          9608 => x"38",
          9609 => x"0b",
          9610 => x"33",
          9611 => x"06",
          9612 => x"73",
          9613 => x"ab",
          9614 => x"2e",
          9615 => x"16",
          9616 => x"81",
          9617 => x"54",
          9618 => x"38",
          9619 => x"06",
          9620 => x"84",
          9621 => x"fe",
          9622 => x"38",
          9623 => x"5d",
          9624 => x"81",
          9625 => x"70",
          9626 => x"33",
          9627 => x"73",
          9628 => x"f0",
          9629 => x"39",
          9630 => x"dc",
          9631 => x"70",
          9632 => x"07",
          9633 => x"55",
          9634 => x"a1",
          9635 => x"70",
          9636 => x"74",
          9637 => x"72",
          9638 => x"38",
          9639 => x"32",
          9640 => x"80",
          9641 => x"51",
          9642 => x"e1",
          9643 => x"1d",
          9644 => x"96",
          9645 => x"41",
          9646 => x"9f",
          9647 => x"38",
          9648 => x"b5",
          9649 => x"81",
          9650 => x"84",
          9651 => x"83",
          9652 => x"54",
          9653 => x"38",
          9654 => x"84",
          9655 => x"93",
          9656 => x"83",
          9657 => x"70",
          9658 => x"5c",
          9659 => x"2e",
          9660 => x"e4",
          9661 => x"0b",
          9662 => x"80",
          9663 => x"de",
          9664 => x"b9",
          9665 => x"b9",
          9666 => x"3d",
          9667 => x"73",
          9668 => x"70",
          9669 => x"25",
          9670 => x"55",
          9671 => x"80",
          9672 => x"81",
          9673 => x"62",
          9674 => x"55",
          9675 => x"2e",
          9676 => x"80",
          9677 => x"30",
          9678 => x"78",
          9679 => x"59",
          9680 => x"73",
          9681 => x"75",
          9682 => x"5a",
          9683 => x"84",
          9684 => x"82",
          9685 => x"38",
          9686 => x"76",
          9687 => x"38",
          9688 => x"11",
          9689 => x"22",
          9690 => x"70",
          9691 => x"2a",
          9692 => x"5f",
          9693 => x"ae",
          9694 => x"72",
          9695 => x"17",
          9696 => x"38",
          9697 => x"19",
          9698 => x"23",
          9699 => x"fe",
          9700 => x"78",
          9701 => x"ff",
          9702 => x"58",
          9703 => x"7a",
          9704 => x"e6",
          9705 => x"ff",
          9706 => x"72",
          9707 => x"f1",
          9708 => x"2e",
          9709 => x"19",
          9710 => x"22",
          9711 => x"ae",
          9712 => x"76",
          9713 => x"05",
          9714 => x"57",
          9715 => x"8f",
          9716 => x"70",
          9717 => x"7c",
          9718 => x"81",
          9719 => x"8b",
          9720 => x"55",
          9721 => x"70",
          9722 => x"34",
          9723 => x"72",
          9724 => x"73",
          9725 => x"78",
          9726 => x"81",
          9727 => x"54",
          9728 => x"2e",
          9729 => x"74",
          9730 => x"d0",
          9731 => x"32",
          9732 => x"80",
          9733 => x"54",
          9734 => x"85",
          9735 => x"83",
          9736 => x"59",
          9737 => x"83",
          9738 => x"75",
          9739 => x"30",
          9740 => x"80",
          9741 => x"07",
          9742 => x"54",
          9743 => x"83",
          9744 => x"8b",
          9745 => x"38",
          9746 => x"8a",
          9747 => x"07",
          9748 => x"26",
          9749 => x"56",
          9750 => x"7e",
          9751 => x"fc",
          9752 => x"57",
          9753 => x"15",
          9754 => x"18",
          9755 => x"74",
          9756 => x"a0",
          9757 => x"76",
          9758 => x"83",
          9759 => x"88",
          9760 => x"38",
          9761 => x"58",
          9762 => x"82",
          9763 => x"83",
          9764 => x"83",
          9765 => x"38",
          9766 => x"81",
          9767 => x"9d",
          9768 => x"06",
          9769 => x"2e",
          9770 => x"90",
          9771 => x"82",
          9772 => x"5e",
          9773 => x"85",
          9774 => x"07",
          9775 => x"1d",
          9776 => x"e4",
          9777 => x"b9",
          9778 => x"1d",
          9779 => x"84",
          9780 => x"80",
          9781 => x"38",
          9782 => x"08",
          9783 => x"81",
          9784 => x"38",
          9785 => x"81",
          9786 => x"80",
          9787 => x"38",
          9788 => x"81",
          9789 => x"82",
          9790 => x"08",
          9791 => x"73",
          9792 => x"08",
          9793 => x"f9",
          9794 => x"16",
          9795 => x"11",
          9796 => x"40",
          9797 => x"a0",
          9798 => x"75",
          9799 => x"85",
          9800 => x"07",
          9801 => x"39",
          9802 => x"56",
          9803 => x"09",
          9804 => x"ac",
          9805 => x"54",
          9806 => x"09",
          9807 => x"a0",
          9808 => x"18",
          9809 => x"23",
          9810 => x"1d",
          9811 => x"54",
          9812 => x"83",
          9813 => x"73",
          9814 => x"05",
          9815 => x"13",
          9816 => x"27",
          9817 => x"a0",
          9818 => x"ab",
          9819 => x"51",
          9820 => x"84",
          9821 => x"ab",
          9822 => x"54",
          9823 => x"08",
          9824 => x"74",
          9825 => x"06",
          9826 => x"ce",
          9827 => x"33",
          9828 => x"81",
          9829 => x"74",
          9830 => x"cd",
          9831 => x"08",
          9832 => x"60",
          9833 => x"11",
          9834 => x"12",
          9835 => x"2b",
          9836 => x"41",
          9837 => x"7d",
          9838 => x"d8",
          9839 => x"1d",
          9840 => x"65",
          9841 => x"b7",
          9842 => x"55",
          9843 => x"fe",
          9844 => x"17",
          9845 => x"88",
          9846 => x"39",
          9847 => x"76",
          9848 => x"fd",
          9849 => x"82",
          9850 => x"06",
          9851 => x"59",
          9852 => x"2e",
          9853 => x"fd",
          9854 => x"82",
          9855 => x"98",
          9856 => x"a0",
          9857 => x"88",
          9858 => x"06",
          9859 => x"d6",
          9860 => x"0b",
          9861 => x"80",
          9862 => x"c8",
          9863 => x"0d",
          9864 => x"ff",
          9865 => x"81",
          9866 => x"80",
          9867 => x"1d",
          9868 => x"26",
          9869 => x"79",
          9870 => x"77",
          9871 => x"5a",
          9872 => x"79",
          9873 => x"83",
          9874 => x"51",
          9875 => x"3f",
          9876 => x"08",
          9877 => x"06",
          9878 => x"81",
          9879 => x"78",
          9880 => x"38",
          9881 => x"06",
          9882 => x"11",
          9883 => x"74",
          9884 => x"ff",
          9885 => x"80",
          9886 => x"38",
          9887 => x"0b",
          9888 => x"33",
          9889 => x"06",
          9890 => x"73",
          9891 => x"e0",
          9892 => x"2e",
          9893 => x"19",
          9894 => x"81",
          9895 => x"54",
          9896 => x"38",
          9897 => x"06",
          9898 => x"d4",
          9899 => x"15",
          9900 => x"26",
          9901 => x"82",
          9902 => x"ff",
          9903 => x"ff",
          9904 => x"78",
          9905 => x"38",
          9906 => x"70",
          9907 => x"e0",
          9908 => x"ff",
          9909 => x"56",
          9910 => x"1b",
          9911 => x"74",
          9912 => x"1b",
          9913 => x"55",
          9914 => x"80",
          9915 => x"39",
          9916 => x"33",
          9917 => x"06",
          9918 => x"80",
          9919 => x"38",
          9920 => x"83",
          9921 => x"a0",
          9922 => x"55",
          9923 => x"81",
          9924 => x"39",
          9925 => x"33",
          9926 => x"33",
          9927 => x"71",
          9928 => x"77",
          9929 => x"0c",
          9930 => x"95",
          9931 => x"a0",
          9932 => x"2a",
          9933 => x"74",
          9934 => x"7c",
          9935 => x"5a",
          9936 => x"34",
          9937 => x"ff",
          9938 => x"83",
          9939 => x"33",
          9940 => x"81",
          9941 => x"81",
          9942 => x"38",
          9943 => x"74",
          9944 => x"06",
          9945 => x"f2",
          9946 => x"84",
          9947 => x"93",
          9948 => x"eb",
          9949 => x"69",
          9950 => x"80",
          9951 => x"42",
          9952 => x"61",
          9953 => x"08",
          9954 => x"42",
          9955 => x"85",
          9956 => x"70",
          9957 => x"33",
          9958 => x"56",
          9959 => x"2e",
          9960 => x"74",
          9961 => x"ba",
          9962 => x"38",
          9963 => x"33",
          9964 => x"24",
          9965 => x"75",
          9966 => x"d1",
          9967 => x"08",
          9968 => x"58",
          9969 => x"85",
          9970 => x"61",
          9971 => x"fe",
          9972 => x"5d",
          9973 => x"2e",
          9974 => x"17",
          9975 => x"bb",
          9976 => x"b9",
          9977 => x"ff",
          9978 => x"06",
          9979 => x"80",
          9980 => x"38",
          9981 => x"75",
          9982 => x"b9",
          9983 => x"81",
          9984 => x"52",
          9985 => x"51",
          9986 => x"3f",
          9987 => x"08",
          9988 => x"70",
          9989 => x"56",
          9990 => x"84",
          9991 => x"80",
          9992 => x"75",
          9993 => x"06",
          9994 => x"60",
          9995 => x"80",
          9996 => x"18",
          9997 => x"b4",
          9998 => x"7b",
          9999 => x"54",
         10000 => x"17",
         10001 => x"18",
         10002 => x"ff",
         10003 => x"84",
         10004 => x"7b",
         10005 => x"ff",
         10006 => x"74",
         10007 => x"84",
         10008 => x"38",
         10009 => x"33",
         10010 => x"33",
         10011 => x"07",
         10012 => x"56",
         10013 => x"d5",
         10014 => x"38",
         10015 => x"8b",
         10016 => x"bd",
         10017 => x"61",
         10018 => x"81",
         10019 => x"2e",
         10020 => x"8d",
         10021 => x"26",
         10022 => x"80",
         10023 => x"80",
         10024 => x"71",
         10025 => x"5e",
         10026 => x"80",
         10027 => x"06",
         10028 => x"80",
         10029 => x"80",
         10030 => x"71",
         10031 => x"57",
         10032 => x"38",
         10033 => x"83",
         10034 => x"12",
         10035 => x"2b",
         10036 => x"07",
         10037 => x"70",
         10038 => x"2b",
         10039 => x"07",
         10040 => x"43",
         10041 => x"75",
         10042 => x"80",
         10043 => x"82",
         10044 => x"c8",
         10045 => x"11",
         10046 => x"06",
         10047 => x"8d",
         10048 => x"26",
         10049 => x"78",
         10050 => x"76",
         10051 => x"c5",
         10052 => x"5f",
         10053 => x"18",
         10054 => x"77",
         10055 => x"c4",
         10056 => x"78",
         10057 => x"87",
         10058 => x"ca",
         10059 => x"c9",
         10060 => x"88",
         10061 => x"40",
         10062 => x"23",
         10063 => x"06",
         10064 => x"58",
         10065 => x"38",
         10066 => x"33",
         10067 => x"33",
         10068 => x"07",
         10069 => x"a4",
         10070 => x"17",
         10071 => x"82",
         10072 => x"90",
         10073 => x"2b",
         10074 => x"33",
         10075 => x"88",
         10076 => x"71",
         10077 => x"5a",
         10078 => x"42",
         10079 => x"33",
         10080 => x"33",
         10081 => x"07",
         10082 => x"58",
         10083 => x"81",
         10084 => x"1c",
         10085 => x"05",
         10086 => x"26",
         10087 => x"78",
         10088 => x"31",
         10089 => x"fd",
         10090 => x"c8",
         10091 => x"b9",
         10092 => x"2e",
         10093 => x"84",
         10094 => x"80",
         10095 => x"f5",
         10096 => x"83",
         10097 => x"ff",
         10098 => x"38",
         10099 => x"9f",
         10100 => x"eb",
         10101 => x"82",
         10102 => x"19",
         10103 => x"19",
         10104 => x"70",
         10105 => x"7b",
         10106 => x"0c",
         10107 => x"83",
         10108 => x"38",
         10109 => x"5c",
         10110 => x"80",
         10111 => x"38",
         10112 => x"18",
         10113 => x"55",
         10114 => x"8d",
         10115 => x"19",
         10116 => x"7a",
         10117 => x"56",
         10118 => x"15",
         10119 => x"8d",
         10120 => x"18",
         10121 => x"38",
         10122 => x"18",
         10123 => x"90",
         10124 => x"80",
         10125 => x"34",
         10126 => x"86",
         10127 => x"77",
         10128 => x"a0",
         10129 => x"5d",
         10130 => x"a0",
         10131 => x"18",
         10132 => x"a8",
         10133 => x"0c",
         10134 => x"18",
         10135 => x"77",
         10136 => x"0c",
         10137 => x"04",
         10138 => x"b9",
         10139 => x"3d",
         10140 => x"33",
         10141 => x"81",
         10142 => x"57",
         10143 => x"26",
         10144 => x"17",
         10145 => x"06",
         10146 => x"59",
         10147 => x"87",
         10148 => x"7e",
         10149 => x"b8",
         10150 => x"7c",
         10151 => x"5b",
         10152 => x"05",
         10153 => x"70",
         10154 => x"33",
         10155 => x"5a",
         10156 => x"99",
         10157 => x"e0",
         10158 => x"ff",
         10159 => x"ff",
         10160 => x"77",
         10161 => x"38",
         10162 => x"81",
         10163 => x"55",
         10164 => x"9f",
         10165 => x"75",
         10166 => x"81",
         10167 => x"77",
         10168 => x"78",
         10169 => x"30",
         10170 => x"9f",
         10171 => x"5d",
         10172 => x"80",
         10173 => x"38",
         10174 => x"1e",
         10175 => x"7c",
         10176 => x"38",
         10177 => x"a9",
         10178 => x"2e",
         10179 => x"77",
         10180 => x"06",
         10181 => x"7d",
         10182 => x"80",
         10183 => x"39",
         10184 => x"57",
         10185 => x"e9",
         10186 => x"06",
         10187 => x"59",
         10188 => x"32",
         10189 => x"80",
         10190 => x"5a",
         10191 => x"83",
         10192 => x"81",
         10193 => x"a6",
         10194 => x"77",
         10195 => x"59",
         10196 => x"33",
         10197 => x"7a",
         10198 => x"38",
         10199 => x"33",
         10200 => x"33",
         10201 => x"71",
         10202 => x"83",
         10203 => x"70",
         10204 => x"2b",
         10205 => x"33",
         10206 => x"59",
         10207 => x"40",
         10208 => x"84",
         10209 => x"ff",
         10210 => x"57",
         10211 => x"25",
         10212 => x"84",
         10213 => x"33",
         10214 => x"9f",
         10215 => x"31",
         10216 => x"10",
         10217 => x"05",
         10218 => x"44",
         10219 => x"5b",
         10220 => x"5b",
         10221 => x"80",
         10222 => x"38",
         10223 => x"18",
         10224 => x"b4",
         10225 => x"55",
         10226 => x"ff",
         10227 => x"81",
         10228 => x"b8",
         10229 => x"17",
         10230 => x"b4",
         10231 => x"b9",
         10232 => x"2e",
         10233 => x"55",
         10234 => x"b4",
         10235 => x"58",
         10236 => x"81",
         10237 => x"33",
         10238 => x"07",
         10239 => x"58",
         10240 => x"d5",
         10241 => x"06",
         10242 => x"0b",
         10243 => x"57",
         10244 => x"e9",
         10245 => x"38",
         10246 => x"32",
         10247 => x"80",
         10248 => x"42",
         10249 => x"bc",
         10250 => x"e8",
         10251 => x"82",
         10252 => x"ff",
         10253 => x"0b",
         10254 => x"1e",
         10255 => x"7b",
         10256 => x"81",
         10257 => x"81",
         10258 => x"27",
         10259 => x"77",
         10260 => x"b7",
         10261 => x"84",
         10262 => x"83",
         10263 => x"d1",
         10264 => x"39",
         10265 => x"ee",
         10266 => x"f8",
         10267 => x"7b",
         10268 => x"5d",
         10269 => x"81",
         10270 => x"71",
         10271 => x"1b",
         10272 => x"56",
         10273 => x"80",
         10274 => x"80",
         10275 => x"85",
         10276 => x"18",
         10277 => x"40",
         10278 => x"70",
         10279 => x"33",
         10280 => x"05",
         10281 => x"71",
         10282 => x"5b",
         10283 => x"77",
         10284 => x"8e",
         10285 => x"2e",
         10286 => x"58",
         10287 => x"8d",
         10288 => x"93",
         10289 => x"b9",
         10290 => x"3d",
         10291 => x"58",
         10292 => x"fe",
         10293 => x"0b",
         10294 => x"83",
         10295 => x"5d",
         10296 => x"39",
         10297 => x"b9",
         10298 => x"3d",
         10299 => x"0b",
         10300 => x"83",
         10301 => x"5a",
         10302 => x"81",
         10303 => x"7a",
         10304 => x"5c",
         10305 => x"31",
         10306 => x"57",
         10307 => x"80",
         10308 => x"38",
         10309 => x"e1",
         10310 => x"81",
         10311 => x"e4",
         10312 => x"58",
         10313 => x"05",
         10314 => x"70",
         10315 => x"33",
         10316 => x"ff",
         10317 => x"42",
         10318 => x"2e",
         10319 => x"75",
         10320 => x"38",
         10321 => x"57",
         10322 => x"fc",
         10323 => x"58",
         10324 => x"80",
         10325 => x"80",
         10326 => x"71",
         10327 => x"57",
         10328 => x"2e",
         10329 => x"f9",
         10330 => x"1b",
         10331 => x"b4",
         10332 => x"2e",
         10333 => x"17",
         10334 => x"7a",
         10335 => x"06",
         10336 => x"81",
         10337 => x"b8",
         10338 => x"17",
         10339 => x"b0",
         10340 => x"b9",
         10341 => x"2e",
         10342 => x"58",
         10343 => x"b4",
         10344 => x"f9",
         10345 => x"84",
         10346 => x"b7",
         10347 => x"b6",
         10348 => x"88",
         10349 => x"5e",
         10350 => x"d5",
         10351 => x"06",
         10352 => x"b8",
         10353 => x"33",
         10354 => x"71",
         10355 => x"88",
         10356 => x"14",
         10357 => x"07",
         10358 => x"33",
         10359 => x"41",
         10360 => x"5c",
         10361 => x"8b",
         10362 => x"2e",
         10363 => x"f8",
         10364 => x"9c",
         10365 => x"33",
         10366 => x"71",
         10367 => x"88",
         10368 => x"14",
         10369 => x"07",
         10370 => x"33",
         10371 => x"44",
         10372 => x"5a",
         10373 => x"8a",
         10374 => x"2e",
         10375 => x"f8",
         10376 => x"a0",
         10377 => x"33",
         10378 => x"71",
         10379 => x"88",
         10380 => x"14",
         10381 => x"07",
         10382 => x"33",
         10383 => x"1e",
         10384 => x"a4",
         10385 => x"33",
         10386 => x"71",
         10387 => x"88",
         10388 => x"14",
         10389 => x"07",
         10390 => x"33",
         10391 => x"90",
         10392 => x"44",
         10393 => x"45",
         10394 => x"56",
         10395 => x"34",
         10396 => x"22",
         10397 => x"7c",
         10398 => x"23",
         10399 => x"23",
         10400 => x"0b",
         10401 => x"80",
         10402 => x"0c",
         10403 => x"7b",
         10404 => x"f0",
         10405 => x"7f",
         10406 => x"95",
         10407 => x"b4",
         10408 => x"b8",
         10409 => x"81",
         10410 => x"59",
         10411 => x"3f",
         10412 => x"08",
         10413 => x"81",
         10414 => x"38",
         10415 => x"08",
         10416 => x"b4",
         10417 => x"18",
         10418 => x"7f",
         10419 => x"27",
         10420 => x"17",
         10421 => x"82",
         10422 => x"38",
         10423 => x"08",
         10424 => x"39",
         10425 => x"80",
         10426 => x"38",
         10427 => x"8a",
         10428 => x"fc",
         10429 => x"fc",
         10430 => x"e3",
         10431 => x"e2",
         10432 => x"88",
         10433 => x"5a",
         10434 => x"f6",
         10435 => x"17",
         10436 => x"f6",
         10437 => x"e4",
         10438 => x"33",
         10439 => x"71",
         10440 => x"88",
         10441 => x"14",
         10442 => x"07",
         10443 => x"33",
         10444 => x"1e",
         10445 => x"82",
         10446 => x"44",
         10447 => x"f5",
         10448 => x"58",
         10449 => x"f9",
         10450 => x"58",
         10451 => x"75",
         10452 => x"a8",
         10453 => x"77",
         10454 => x"59",
         10455 => x"75",
         10456 => x"da",
         10457 => x"39",
         10458 => x"17",
         10459 => x"08",
         10460 => x"52",
         10461 => x"51",
         10462 => x"3f",
         10463 => x"f0",
         10464 => x"80",
         10465 => x"64",
         10466 => x"3d",
         10467 => x"ff",
         10468 => x"75",
         10469 => x"e9",
         10470 => x"81",
         10471 => x"70",
         10472 => x"55",
         10473 => x"80",
         10474 => x"ed",
         10475 => x"2e",
         10476 => x"84",
         10477 => x"54",
         10478 => x"80",
         10479 => x"10",
         10480 => x"90",
         10481 => x"55",
         10482 => x"2e",
         10483 => x"74",
         10484 => x"73",
         10485 => x"38",
         10486 => x"62",
         10487 => x"0c",
         10488 => x"80",
         10489 => x"80",
         10490 => x"70",
         10491 => x"51",
         10492 => x"84",
         10493 => x"54",
         10494 => x"c8",
         10495 => x"0d",
         10496 => x"84",
         10497 => x"92",
         10498 => x"75",
         10499 => x"70",
         10500 => x"56",
         10501 => x"89",
         10502 => x"82",
         10503 => x"ff",
         10504 => x"5c",
         10505 => x"2e",
         10506 => x"80",
         10507 => x"e5",
         10508 => x"5b",
         10509 => x"59",
         10510 => x"81",
         10511 => x"78",
         10512 => x"5a",
         10513 => x"12",
         10514 => x"76",
         10515 => x"38",
         10516 => x"81",
         10517 => x"54",
         10518 => x"57",
         10519 => x"89",
         10520 => x"70",
         10521 => x"57",
         10522 => x"70",
         10523 => x"54",
         10524 => x"09",
         10525 => x"38",
         10526 => x"38",
         10527 => x"70",
         10528 => x"07",
         10529 => x"07",
         10530 => x"79",
         10531 => x"38",
         10532 => x"1d",
         10533 => x"7b",
         10534 => x"38",
         10535 => x"98",
         10536 => x"24",
         10537 => x"79",
         10538 => x"fe",
         10539 => x"3d",
         10540 => x"84",
         10541 => x"05",
         10542 => x"89",
         10543 => x"2e",
         10544 => x"bf",
         10545 => x"9d",
         10546 => x"53",
         10547 => x"05",
         10548 => x"9f",
         10549 => x"c8",
         10550 => x"b9",
         10551 => x"2e",
         10552 => x"79",
         10553 => x"75",
         10554 => x"0c",
         10555 => x"04",
         10556 => x"52",
         10557 => x"52",
         10558 => x"3f",
         10559 => x"08",
         10560 => x"c8",
         10561 => x"81",
         10562 => x"9c",
         10563 => x"80",
         10564 => x"38",
         10565 => x"83",
         10566 => x"84",
         10567 => x"38",
         10568 => x"58",
         10569 => x"38",
         10570 => x"81",
         10571 => x"80",
         10572 => x"38",
         10573 => x"33",
         10574 => x"71",
         10575 => x"61",
         10576 => x"58",
         10577 => x"7d",
         10578 => x"e9",
         10579 => x"8e",
         10580 => x"0b",
         10581 => x"a1",
         10582 => x"34",
         10583 => x"91",
         10584 => x"56",
         10585 => x"17",
         10586 => x"57",
         10587 => x"9a",
         10588 => x"0b",
         10589 => x"7d",
         10590 => x"83",
         10591 => x"38",
         10592 => x"0b",
         10593 => x"80",
         10594 => x"34",
         10595 => x"1c",
         10596 => x"9f",
         10597 => x"55",
         10598 => x"16",
         10599 => x"2e",
         10600 => x"7e",
         10601 => x"7d",
         10602 => x"57",
         10603 => x"7c",
         10604 => x"9c",
         10605 => x"26",
         10606 => x"82",
         10607 => x"0c",
         10608 => x"02",
         10609 => x"33",
         10610 => x"5d",
         10611 => x"25",
         10612 => x"86",
         10613 => x"5e",
         10614 => x"b8",
         10615 => x"82",
         10616 => x"c2",
         10617 => x"84",
         10618 => x"5d",
         10619 => x"91",
         10620 => x"2a",
         10621 => x"7d",
         10622 => x"38",
         10623 => x"5a",
         10624 => x"38",
         10625 => x"81",
         10626 => x"80",
         10627 => x"77",
         10628 => x"58",
         10629 => x"08",
         10630 => x"67",
         10631 => x"67",
         10632 => x"9a",
         10633 => x"88",
         10634 => x"33",
         10635 => x"57",
         10636 => x"2e",
         10637 => x"7a",
         10638 => x"9c",
         10639 => x"33",
         10640 => x"71",
         10641 => x"88",
         10642 => x"14",
         10643 => x"07",
         10644 => x"33",
         10645 => x"60",
         10646 => x"60",
         10647 => x"52",
         10648 => x"5d",
         10649 => x"22",
         10650 => x"77",
         10651 => x"80",
         10652 => x"34",
         10653 => x"1a",
         10654 => x"2a",
         10655 => x"74",
         10656 => x"ac",
         10657 => x"2e",
         10658 => x"75",
         10659 => x"8a",
         10660 => x"89",
         10661 => x"5b",
         10662 => x"70",
         10663 => x"25",
         10664 => x"76",
         10665 => x"38",
         10666 => x"06",
         10667 => x"80",
         10668 => x"38",
         10669 => x"51",
         10670 => x"3f",
         10671 => x"08",
         10672 => x"c8",
         10673 => x"83",
         10674 => x"84",
         10675 => x"ff",
         10676 => x"38",
         10677 => x"56",
         10678 => x"80",
         10679 => x"91",
         10680 => x"95",
         10681 => x"2a",
         10682 => x"74",
         10683 => x"b8",
         10684 => x"80",
         10685 => x"ed",
         10686 => x"80",
         10687 => x"e5",
         10688 => x"80",
         10689 => x"dd",
         10690 => x"cd",
         10691 => x"b9",
         10692 => x"88",
         10693 => x"76",
         10694 => x"fc",
         10695 => x"76",
         10696 => x"57",
         10697 => x"95",
         10698 => x"17",
         10699 => x"2b",
         10700 => x"07",
         10701 => x"5e",
         10702 => x"39",
         10703 => x"7b",
         10704 => x"38",
         10705 => x"51",
         10706 => x"3f",
         10707 => x"08",
         10708 => x"c8",
         10709 => x"81",
         10710 => x"b9",
         10711 => x"2e",
         10712 => x"84",
         10713 => x"ff",
         10714 => x"38",
         10715 => x"52",
         10716 => x"b2",
         10717 => x"b9",
         10718 => x"90",
         10719 => x"08",
         10720 => x"19",
         10721 => x"5b",
         10722 => x"ff",
         10723 => x"16",
         10724 => x"84",
         10725 => x"07",
         10726 => x"18",
         10727 => x"7a",
         10728 => x"a0",
         10729 => x"39",
         10730 => x"17",
         10731 => x"95",
         10732 => x"cc",
         10733 => x"33",
         10734 => x"71",
         10735 => x"90",
         10736 => x"07",
         10737 => x"80",
         10738 => x"34",
         10739 => x"17",
         10740 => x"90",
         10741 => x"cc",
         10742 => x"34",
         10743 => x"0b",
         10744 => x"7e",
         10745 => x"80",
         10746 => x"34",
         10747 => x"17",
         10748 => x"5d",
         10749 => x"09",
         10750 => x"84",
         10751 => x"39",
         10752 => x"72",
         10753 => x"5d",
         10754 => x"7e",
         10755 => x"83",
         10756 => x"79",
         10757 => x"81",
         10758 => x"81",
         10759 => x"b8",
         10760 => x"16",
         10761 => x"a3",
         10762 => x"b9",
         10763 => x"2e",
         10764 => x"57",
         10765 => x"b4",
         10766 => x"56",
         10767 => x"90",
         10768 => x"7a",
         10769 => x"bc",
         10770 => x"0c",
         10771 => x"81",
         10772 => x"08",
         10773 => x"70",
         10774 => x"33",
         10775 => x"a4",
         10776 => x"b9",
         10777 => x"2e",
         10778 => x"81",
         10779 => x"b9",
         10780 => x"17",
         10781 => x"08",
         10782 => x"31",
         10783 => x"08",
         10784 => x"a0",
         10785 => x"ff",
         10786 => x"16",
         10787 => x"82",
         10788 => x"06",
         10789 => x"81",
         10790 => x"08",
         10791 => x"05",
         10792 => x"81",
         10793 => x"ff",
         10794 => x"7c",
         10795 => x"39",
         10796 => x"0c",
         10797 => x"af",
         10798 => x"1a",
         10799 => x"a2",
         10800 => x"ff",
         10801 => x"80",
         10802 => x"38",
         10803 => x"9c",
         10804 => x"05",
         10805 => x"77",
         10806 => x"df",
         10807 => x"22",
         10808 => x"b0",
         10809 => x"56",
         10810 => x"2e",
         10811 => x"75",
         10812 => x"9c",
         10813 => x"56",
         10814 => x"75",
         10815 => x"76",
         10816 => x"39",
         10817 => x"79",
         10818 => x"39",
         10819 => x"08",
         10820 => x"0c",
         10821 => x"81",
         10822 => x"fe",
         10823 => x"3d",
         10824 => x"67",
         10825 => x"5d",
         10826 => x"0c",
         10827 => x"80",
         10828 => x"79",
         10829 => x"80",
         10830 => x"75",
         10831 => x"80",
         10832 => x"86",
         10833 => x"1b",
         10834 => x"78",
         10835 => x"b7",
         10836 => x"74",
         10837 => x"76",
         10838 => x"91",
         10839 => x"74",
         10840 => x"90",
         10841 => x"06",
         10842 => x"76",
         10843 => x"ed",
         10844 => x"08",
         10845 => x"71",
         10846 => x"7b",
         10847 => x"ef",
         10848 => x"2e",
         10849 => x"60",
         10850 => x"ff",
         10851 => x"81",
         10852 => x"19",
         10853 => x"76",
         10854 => x"5b",
         10855 => x"75",
         10856 => x"88",
         10857 => x"81",
         10858 => x"85",
         10859 => x"2e",
         10860 => x"74",
         10861 => x"60",
         10862 => x"08",
         10863 => x"1a",
         10864 => x"41",
         10865 => x"27",
         10866 => x"8a",
         10867 => x"78",
         10868 => x"08",
         10869 => x"74",
         10870 => x"d5",
         10871 => x"7c",
         10872 => x"57",
         10873 => x"83",
         10874 => x"1b",
         10875 => x"27",
         10876 => x"7b",
         10877 => x"54",
         10878 => x"52",
         10879 => x"51",
         10880 => x"3f",
         10881 => x"08",
         10882 => x"60",
         10883 => x"57",
         10884 => x"2e",
         10885 => x"19",
         10886 => x"56",
         10887 => x"9e",
         10888 => x"76",
         10889 => x"b8",
         10890 => x"55",
         10891 => x"05",
         10892 => x"70",
         10893 => x"34",
         10894 => x"74",
         10895 => x"89",
         10896 => x"78",
         10897 => x"19",
         10898 => x"1e",
         10899 => x"1a",
         10900 => x"1d",
         10901 => x"7b",
         10902 => x"80",
         10903 => x"b9",
         10904 => x"3d",
         10905 => x"84",
         10906 => x"92",
         10907 => x"74",
         10908 => x"39",
         10909 => x"57",
         10910 => x"06",
         10911 => x"31",
         10912 => x"78",
         10913 => x"7b",
         10914 => x"b4",
         10915 => x"2e",
         10916 => x"0b",
         10917 => x"71",
         10918 => x"7f",
         10919 => x"81",
         10920 => x"38",
         10921 => x"53",
         10922 => x"81",
         10923 => x"ff",
         10924 => x"84",
         10925 => x"80",
         10926 => x"ff",
         10927 => x"75",
         10928 => x"7a",
         10929 => x"60",
         10930 => x"83",
         10931 => x"79",
         10932 => x"b8",
         10933 => x"77",
         10934 => x"e6",
         10935 => x"81",
         10936 => x"77",
         10937 => x"59",
         10938 => x"56",
         10939 => x"fe",
         10940 => x"70",
         10941 => x"33",
         10942 => x"05",
         10943 => x"16",
         10944 => x"38",
         10945 => x"81",
         10946 => x"08",
         10947 => x"70",
         10948 => x"33",
         10949 => x"9e",
         10950 => x"5b",
         10951 => x"08",
         10952 => x"81",
         10953 => x"38",
         10954 => x"08",
         10955 => x"b4",
         10956 => x"1a",
         10957 => x"b9",
         10958 => x"55",
         10959 => x"08",
         10960 => x"38",
         10961 => x"55",
         10962 => x"09",
         10963 => x"d4",
         10964 => x"b4",
         10965 => x"1a",
         10966 => x"7f",
         10967 => x"33",
         10968 => x"fe",
         10969 => x"fe",
         10970 => x"9c",
         10971 => x"1a",
         10972 => x"84",
         10973 => x"08",
         10974 => x"ff",
         10975 => x"84",
         10976 => x"55",
         10977 => x"81",
         10978 => x"ff",
         10979 => x"84",
         10980 => x"81",
         10981 => x"fb",
         10982 => x"7a",
         10983 => x"fb",
         10984 => x"0b",
         10985 => x"81",
         10986 => x"c8",
         10987 => x"0d",
         10988 => x"91",
         10989 => x"0b",
         10990 => x"0c",
         10991 => x"04",
         10992 => x"62",
         10993 => x"40",
         10994 => x"80",
         10995 => x"57",
         10996 => x"9f",
         10997 => x"56",
         10998 => x"97",
         10999 => x"55",
         11000 => x"8f",
         11001 => x"22",
         11002 => x"59",
         11003 => x"2e",
         11004 => x"80",
         11005 => x"76",
         11006 => x"c4",
         11007 => x"33",
         11008 => x"bc",
         11009 => x"33",
         11010 => x"81",
         11011 => x"87",
         11012 => x"2e",
         11013 => x"94",
         11014 => x"11",
         11015 => x"77",
         11016 => x"76",
         11017 => x"80",
         11018 => x"38",
         11019 => x"06",
         11020 => x"a2",
         11021 => x"11",
         11022 => x"78",
         11023 => x"5a",
         11024 => x"38",
         11025 => x"38",
         11026 => x"55",
         11027 => x"84",
         11028 => x"81",
         11029 => x"38",
         11030 => x"86",
         11031 => x"98",
         11032 => x"1a",
         11033 => x"74",
         11034 => x"60",
         11035 => x"08",
         11036 => x"2e",
         11037 => x"98",
         11038 => x"05",
         11039 => x"fe",
         11040 => x"77",
         11041 => x"f0",
         11042 => x"22",
         11043 => x"b0",
         11044 => x"56",
         11045 => x"2e",
         11046 => x"78",
         11047 => x"2a",
         11048 => x"80",
         11049 => x"38",
         11050 => x"76",
         11051 => x"38",
         11052 => x"58",
         11053 => x"53",
         11054 => x"16",
         11055 => x"9b",
         11056 => x"b9",
         11057 => x"a1",
         11058 => x"11",
         11059 => x"56",
         11060 => x"27",
         11061 => x"80",
         11062 => x"76",
         11063 => x"57",
         11064 => x"70",
         11065 => x"33",
         11066 => x"05",
         11067 => x"16",
         11068 => x"38",
         11069 => x"83",
         11070 => x"89",
         11071 => x"79",
         11072 => x"1a",
         11073 => x"1e",
         11074 => x"1b",
         11075 => x"1f",
         11076 => x"08",
         11077 => x"5e",
         11078 => x"27",
         11079 => x"56",
         11080 => x"0c",
         11081 => x"38",
         11082 => x"58",
         11083 => x"07",
         11084 => x"1b",
         11085 => x"75",
         11086 => x"0c",
         11087 => x"04",
         11088 => x"c8",
         11089 => x"0d",
         11090 => x"33",
         11091 => x"c8",
         11092 => x"fe",
         11093 => x"9c",
         11094 => x"56",
         11095 => x"06",
         11096 => x"31",
         11097 => x"79",
         11098 => x"7a",
         11099 => x"b4",
         11100 => x"2e",
         11101 => x"0b",
         11102 => x"71",
         11103 => x"7f",
         11104 => x"81",
         11105 => x"38",
         11106 => x"53",
         11107 => x"81",
         11108 => x"ff",
         11109 => x"84",
         11110 => x"80",
         11111 => x"ff",
         11112 => x"76",
         11113 => x"7b",
         11114 => x"60",
         11115 => x"83",
         11116 => x"7a",
         11117 => x"7e",
         11118 => x"78",
         11119 => x"38",
         11120 => x"05",
         11121 => x"70",
         11122 => x"34",
         11123 => x"75",
         11124 => x"58",
         11125 => x"19",
         11126 => x"39",
         11127 => x"16",
         11128 => x"16",
         11129 => x"17",
         11130 => x"ff",
         11131 => x"81",
         11132 => x"c8",
         11133 => x"09",
         11134 => x"ab",
         11135 => x"c8",
         11136 => x"34",
         11137 => x"a8",
         11138 => x"84",
         11139 => x"5d",
         11140 => x"17",
         11141 => x"f0",
         11142 => x"33",
         11143 => x"2e",
         11144 => x"fe",
         11145 => x"54",
         11146 => x"a0",
         11147 => x"53",
         11148 => x"16",
         11149 => x"98",
         11150 => x"5c",
         11151 => x"94",
         11152 => x"8c",
         11153 => x"26",
         11154 => x"16",
         11155 => x"81",
         11156 => x"7c",
         11157 => x"94",
         11158 => x"56",
         11159 => x"1c",
         11160 => x"f8",
         11161 => x"08",
         11162 => x"ff",
         11163 => x"84",
         11164 => x"55",
         11165 => x"08",
         11166 => x"90",
         11167 => x"fd",
         11168 => x"52",
         11169 => x"ab",
         11170 => x"b9",
         11171 => x"84",
         11172 => x"fb",
         11173 => x"39",
         11174 => x"16",
         11175 => x"16",
         11176 => x"17",
         11177 => x"ff",
         11178 => x"84",
         11179 => x"81",
         11180 => x"b9",
         11181 => x"17",
         11182 => x"08",
         11183 => x"31",
         11184 => x"17",
         11185 => x"89",
         11186 => x"33",
         11187 => x"2e",
         11188 => x"fc",
         11189 => x"54",
         11190 => x"a0",
         11191 => x"53",
         11192 => x"16",
         11193 => x"96",
         11194 => x"56",
         11195 => x"81",
         11196 => x"ff",
         11197 => x"84",
         11198 => x"81",
         11199 => x"f9",
         11200 => x"7a",
         11201 => x"f9",
         11202 => x"54",
         11203 => x"53",
         11204 => x"53",
         11205 => x"52",
         11206 => x"c6",
         11207 => x"c8",
         11208 => x"38",
         11209 => x"08",
         11210 => x"b4",
         11211 => x"17",
         11212 => x"74",
         11213 => x"27",
         11214 => x"82",
         11215 => x"77",
         11216 => x"81",
         11217 => x"38",
         11218 => x"16",
         11219 => x"08",
         11220 => x"52",
         11221 => x"51",
         11222 => x"3f",
         11223 => x"12",
         11224 => x"08",
         11225 => x"f4",
         11226 => x"91",
         11227 => x"0b",
         11228 => x"0c",
         11229 => x"04",
         11230 => x"1b",
         11231 => x"84",
         11232 => x"92",
         11233 => x"f5",
         11234 => x"58",
         11235 => x"80",
         11236 => x"77",
         11237 => x"80",
         11238 => x"75",
         11239 => x"80",
         11240 => x"86",
         11241 => x"19",
         11242 => x"78",
         11243 => x"b5",
         11244 => x"74",
         11245 => x"79",
         11246 => x"90",
         11247 => x"86",
         11248 => x"5c",
         11249 => x"2e",
         11250 => x"7b",
         11251 => x"5a",
         11252 => x"08",
         11253 => x"38",
         11254 => x"5b",
         11255 => x"38",
         11256 => x"53",
         11257 => x"81",
         11258 => x"ff",
         11259 => x"84",
         11260 => x"80",
         11261 => x"ff",
         11262 => x"78",
         11263 => x"75",
         11264 => x"a4",
         11265 => x"11",
         11266 => x"5a",
         11267 => x"18",
         11268 => x"88",
         11269 => x"83",
         11270 => x"5d",
         11271 => x"9a",
         11272 => x"88",
         11273 => x"9b",
         11274 => x"17",
         11275 => x"19",
         11276 => x"74",
         11277 => x"c1",
         11278 => x"08",
         11279 => x"34",
         11280 => x"5b",
         11281 => x"34",
         11282 => x"56",
         11283 => x"34",
         11284 => x"59",
         11285 => x"34",
         11286 => x"80",
         11287 => x"34",
         11288 => x"18",
         11289 => x"0b",
         11290 => x"80",
         11291 => x"34",
         11292 => x"18",
         11293 => x"81",
         11294 => x"34",
         11295 => x"96",
         11296 => x"b9",
         11297 => x"19",
         11298 => x"06",
         11299 => x"90",
         11300 => x"84",
         11301 => x"8d",
         11302 => x"81",
         11303 => x"08",
         11304 => x"70",
         11305 => x"33",
         11306 => x"93",
         11307 => x"56",
         11308 => x"08",
         11309 => x"84",
         11310 => x"83",
         11311 => x"17",
         11312 => x"08",
         11313 => x"c8",
         11314 => x"74",
         11315 => x"27",
         11316 => x"82",
         11317 => x"74",
         11318 => x"81",
         11319 => x"38",
         11320 => x"17",
         11321 => x"08",
         11322 => x"52",
         11323 => x"51",
         11324 => x"3f",
         11325 => x"e8",
         11326 => x"2a",
         11327 => x"18",
         11328 => x"2a",
         11329 => x"18",
         11330 => x"08",
         11331 => x"34",
         11332 => x"5b",
         11333 => x"34",
         11334 => x"56",
         11335 => x"34",
         11336 => x"59",
         11337 => x"34",
         11338 => x"80",
         11339 => x"34",
         11340 => x"18",
         11341 => x"0b",
         11342 => x"80",
         11343 => x"34",
         11344 => x"18",
         11345 => x"81",
         11346 => x"34",
         11347 => x"94",
         11348 => x"b9",
         11349 => x"19",
         11350 => x"06",
         11351 => x"90",
         11352 => x"ae",
         11353 => x"33",
         11354 => x"a5",
         11355 => x"c8",
         11356 => x"55",
         11357 => x"38",
         11358 => x"56",
         11359 => x"39",
         11360 => x"79",
         11361 => x"fb",
         11362 => x"b9",
         11363 => x"84",
         11364 => x"b1",
         11365 => x"74",
         11366 => x"38",
         11367 => x"72",
         11368 => x"38",
         11369 => x"71",
         11370 => x"38",
         11371 => x"84",
         11372 => x"52",
         11373 => x"96",
         11374 => x"71",
         11375 => x"75",
         11376 => x"75",
         11377 => x"b9",
         11378 => x"3d",
         11379 => x"13",
         11380 => x"8f",
         11381 => x"b9",
         11382 => x"06",
         11383 => x"38",
         11384 => x"53",
         11385 => x"f6",
         11386 => x"7d",
         11387 => x"5b",
         11388 => x"b2",
         11389 => x"81",
         11390 => x"70",
         11391 => x"52",
         11392 => x"ac",
         11393 => x"38",
         11394 => x"a4",
         11395 => x"a4",
         11396 => x"71",
         11397 => x"70",
         11398 => x"34",
         11399 => x"b9",
         11400 => x"3d",
         11401 => x"0b",
         11402 => x"0c",
         11403 => x"04",
         11404 => x"11",
         11405 => x"06",
         11406 => x"70",
         11407 => x"38",
         11408 => x"81",
         11409 => x"05",
         11410 => x"76",
         11411 => x"38",
         11412 => x"e5",
         11413 => x"79",
         11414 => x"57",
         11415 => x"05",
         11416 => x"70",
         11417 => x"33",
         11418 => x"53",
         11419 => x"99",
         11420 => x"e0",
         11421 => x"ff",
         11422 => x"ff",
         11423 => x"70",
         11424 => x"38",
         11425 => x"81",
         11426 => x"54",
         11427 => x"9f",
         11428 => x"71",
         11429 => x"81",
         11430 => x"73",
         11431 => x"74",
         11432 => x"30",
         11433 => x"9f",
         11434 => x"59",
         11435 => x"80",
         11436 => x"81",
         11437 => x"5b",
         11438 => x"25",
         11439 => x"7a",
         11440 => x"39",
         11441 => x"f7",
         11442 => x"5e",
         11443 => x"39",
         11444 => x"80",
         11445 => x"cc",
         11446 => x"3d",
         11447 => x"3f",
         11448 => x"08",
         11449 => x"c8",
         11450 => x"8a",
         11451 => x"b9",
         11452 => x"3d",
         11453 => x"5c",
         11454 => x"3d",
         11455 => x"c5",
         11456 => x"b9",
         11457 => x"84",
         11458 => x"80",
         11459 => x"80",
         11460 => x"70",
         11461 => x"5a",
         11462 => x"80",
         11463 => x"b2",
         11464 => x"84",
         11465 => x"57",
         11466 => x"2e",
         11467 => x"63",
         11468 => x"9a",
         11469 => x"88",
         11470 => x"33",
         11471 => x"57",
         11472 => x"2e",
         11473 => x"98",
         11474 => x"84",
         11475 => x"98",
         11476 => x"84",
         11477 => x"84",
         11478 => x"06",
         11479 => x"85",
         11480 => x"c8",
         11481 => x"0d",
         11482 => x"33",
         11483 => x"71",
         11484 => x"90",
         11485 => x"07",
         11486 => x"5b",
         11487 => x"7a",
         11488 => x"0c",
         11489 => x"b9",
         11490 => x"3d",
         11491 => x"9e",
         11492 => x"e6",
         11493 => x"e6",
         11494 => x"40",
         11495 => x"80",
         11496 => x"3d",
         11497 => x"52",
         11498 => x"51",
         11499 => x"84",
         11500 => x"59",
         11501 => x"08",
         11502 => x"60",
         11503 => x"0c",
         11504 => x"11",
         11505 => x"3d",
         11506 => x"db",
         11507 => x"58",
         11508 => x"82",
         11509 => x"d8",
         11510 => x"40",
         11511 => x"7a",
         11512 => x"aa",
         11513 => x"c8",
         11514 => x"b9",
         11515 => x"92",
         11516 => x"df",
         11517 => x"56",
         11518 => x"77",
         11519 => x"84",
         11520 => x"83",
         11521 => x"5d",
         11522 => x"38",
         11523 => x"53",
         11524 => x"81",
         11525 => x"ff",
         11526 => x"84",
         11527 => x"80",
         11528 => x"ff",
         11529 => x"76",
         11530 => x"78",
         11531 => x"80",
         11532 => x"9b",
         11533 => x"12",
         11534 => x"2b",
         11535 => x"33",
         11536 => x"56",
         11537 => x"2e",
         11538 => x"76",
         11539 => x"0c",
         11540 => x"51",
         11541 => x"3f",
         11542 => x"08",
         11543 => x"c8",
         11544 => x"38",
         11545 => x"51",
         11546 => x"3f",
         11547 => x"08",
         11548 => x"c8",
         11549 => x"80",
         11550 => x"9b",
         11551 => x"12",
         11552 => x"2b",
         11553 => x"33",
         11554 => x"5e",
         11555 => x"2e",
         11556 => x"76",
         11557 => x"38",
         11558 => x"08",
         11559 => x"ff",
         11560 => x"84",
         11561 => x"59",
         11562 => x"08",
         11563 => x"b4",
         11564 => x"2e",
         11565 => x"78",
         11566 => x"80",
         11567 => x"b8",
         11568 => x"51",
         11569 => x"3f",
         11570 => x"05",
         11571 => x"79",
         11572 => x"38",
         11573 => x"81",
         11574 => x"70",
         11575 => x"57",
         11576 => x"81",
         11577 => x"78",
         11578 => x"38",
         11579 => x"9c",
         11580 => x"82",
         11581 => x"18",
         11582 => x"08",
         11583 => x"ff",
         11584 => x"56",
         11585 => x"75",
         11586 => x"38",
         11587 => x"e6",
         11588 => x"5f",
         11589 => x"34",
         11590 => x"08",
         11591 => x"bd",
         11592 => x"2e",
         11593 => x"80",
         11594 => x"a4",
         11595 => x"10",
         11596 => x"05",
         11597 => x"33",
         11598 => x"5e",
         11599 => x"2e",
         11600 => x"1a",
         11601 => x"33",
         11602 => x"74",
         11603 => x"1a",
         11604 => x"26",
         11605 => x"57",
         11606 => x"94",
         11607 => x"5f",
         11608 => x"70",
         11609 => x"34",
         11610 => x"79",
         11611 => x"38",
         11612 => x"81",
         11613 => x"76",
         11614 => x"81",
         11615 => x"38",
         11616 => x"7c",
         11617 => x"b9",
         11618 => x"e4",
         11619 => x"95",
         11620 => x"17",
         11621 => x"2b",
         11622 => x"07",
         11623 => x"56",
         11624 => x"39",
         11625 => x"94",
         11626 => x"98",
         11627 => x"2b",
         11628 => x"80",
         11629 => x"5a",
         11630 => x"7a",
         11631 => x"ce",
         11632 => x"c8",
         11633 => x"b9",
         11634 => x"2e",
         11635 => x"ff",
         11636 => x"54",
         11637 => x"53",
         11638 => x"53",
         11639 => x"52",
         11640 => x"fe",
         11641 => x"84",
         11642 => x"fc",
         11643 => x"b9",
         11644 => x"17",
         11645 => x"08",
         11646 => x"31",
         11647 => x"08",
         11648 => x"a0",
         11649 => x"fc",
         11650 => x"16",
         11651 => x"82",
         11652 => x"06",
         11653 => x"81",
         11654 => x"08",
         11655 => x"05",
         11656 => x"81",
         11657 => x"ff",
         11658 => x"7c",
         11659 => x"39",
         11660 => x"e6",
         11661 => x"5c",
         11662 => x"34",
         11663 => x"d1",
         11664 => x"10",
         11665 => x"b8",
         11666 => x"70",
         11667 => x"59",
         11668 => x"7a",
         11669 => x"06",
         11670 => x"fd",
         11671 => x"e5",
         11672 => x"81",
         11673 => x"79",
         11674 => x"81",
         11675 => x"77",
         11676 => x"8e",
         11677 => x"3d",
         11678 => x"19",
         11679 => x"33",
         11680 => x"05",
         11681 => x"78",
         11682 => x"fd",
         11683 => x"59",
         11684 => x"78",
         11685 => x"0c",
         11686 => x"0d",
         11687 => x"0d",
         11688 => x"55",
         11689 => x"80",
         11690 => x"74",
         11691 => x"80",
         11692 => x"73",
         11693 => x"80",
         11694 => x"86",
         11695 => x"16",
         11696 => x"78",
         11697 => x"a0",
         11698 => x"72",
         11699 => x"75",
         11700 => x"91",
         11701 => x"72",
         11702 => x"8c",
         11703 => x"76",
         11704 => x"b9",
         11705 => x"08",
         11706 => x"76",
         11707 => x"cc",
         11708 => x"11",
         11709 => x"2b",
         11710 => x"73",
         11711 => x"f7",
         11712 => x"ff",
         11713 => x"bb",
         11714 => x"b9",
         11715 => x"15",
         11716 => x"53",
         11717 => x"bb",
         11718 => x"b9",
         11719 => x"26",
         11720 => x"75",
         11721 => x"70",
         11722 => x"77",
         11723 => x"17",
         11724 => x"59",
         11725 => x"82",
         11726 => x"77",
         11727 => x"38",
         11728 => x"94",
         11729 => x"94",
         11730 => x"16",
         11731 => x"2a",
         11732 => x"5a",
         11733 => x"2e",
         11734 => x"73",
         11735 => x"ff",
         11736 => x"84",
         11737 => x"54",
         11738 => x"08",
         11739 => x"a3",
         11740 => x"2e",
         11741 => x"74",
         11742 => x"38",
         11743 => x"9c",
         11744 => x"82",
         11745 => x"98",
         11746 => x"ae",
         11747 => x"91",
         11748 => x"53",
         11749 => x"c8",
         11750 => x"0d",
         11751 => x"33",
         11752 => x"81",
         11753 => x"73",
         11754 => x"75",
         11755 => x"55",
         11756 => x"76",
         11757 => x"81",
         11758 => x"38",
         11759 => x"0c",
         11760 => x"54",
         11761 => x"90",
         11762 => x"16",
         11763 => x"33",
         11764 => x"57",
         11765 => x"34",
         11766 => x"06",
         11767 => x"2e",
         11768 => x"15",
         11769 => x"85",
         11770 => x"16",
         11771 => x"84",
         11772 => x"8b",
         11773 => x"80",
         11774 => x"0c",
         11775 => x"54",
         11776 => x"80",
         11777 => x"98",
         11778 => x"80",
         11779 => x"38",
         11780 => x"84",
         11781 => x"57",
         11782 => x"17",
         11783 => x"76",
         11784 => x"56",
         11785 => x"a9",
         11786 => x"15",
         11787 => x"fe",
         11788 => x"56",
         11789 => x"80",
         11790 => x"16",
         11791 => x"29",
         11792 => x"05",
         11793 => x"11",
         11794 => x"78",
         11795 => x"df",
         11796 => x"08",
         11797 => x"39",
         11798 => x"51",
         11799 => x"3f",
         11800 => x"08",
         11801 => x"39",
         11802 => x"51",
         11803 => x"3f",
         11804 => x"08",
         11805 => x"72",
         11806 => x"72",
         11807 => x"56",
         11808 => x"73",
         11809 => x"ff",
         11810 => x"84",
         11811 => x"54",
         11812 => x"08",
         11813 => x"38",
         11814 => x"08",
         11815 => x"ed",
         11816 => x"c8",
         11817 => x"0c",
         11818 => x"0c",
         11819 => x"82",
         11820 => x"34",
         11821 => x"b9",
         11822 => x"3d",
         11823 => x"3d",
         11824 => x"89",
         11825 => x"2e",
         11826 => x"53",
         11827 => x"05",
         11828 => x"84",
         11829 => x"9b",
         11830 => x"c8",
         11831 => x"b9",
         11832 => x"2e",
         11833 => x"76",
         11834 => x"73",
         11835 => x"0c",
         11836 => x"04",
         11837 => x"7d",
         11838 => x"ff",
         11839 => x"84",
         11840 => x"55",
         11841 => x"08",
         11842 => x"ab",
         11843 => x"98",
         11844 => x"80",
         11845 => x"38",
         11846 => x"70",
         11847 => x"06",
         11848 => x"80",
         11849 => x"38",
         11850 => x"9b",
         11851 => x"12",
         11852 => x"2b",
         11853 => x"33",
         11854 => x"55",
         11855 => x"2e",
         11856 => x"88",
         11857 => x"58",
         11858 => x"84",
         11859 => x"52",
         11860 => x"99",
         11861 => x"b9",
         11862 => x"74",
         11863 => x"38",
         11864 => x"ff",
         11865 => x"76",
         11866 => x"39",
         11867 => x"76",
         11868 => x"39",
         11869 => x"94",
         11870 => x"98",
         11871 => x"2b",
         11872 => x"88",
         11873 => x"5a",
         11874 => x"fa",
         11875 => x"55",
         11876 => x"80",
         11877 => x"74",
         11878 => x"80",
         11879 => x"72",
         11880 => x"80",
         11881 => x"86",
         11882 => x"16",
         11883 => x"71",
         11884 => x"38",
         11885 => x"57",
         11886 => x"73",
         11887 => x"84",
         11888 => x"88",
         11889 => x"81",
         11890 => x"fe",
         11891 => x"84",
         11892 => x"81",
         11893 => x"dc",
         11894 => x"08",
         11895 => x"39",
         11896 => x"7a",
         11897 => x"89",
         11898 => x"2e",
         11899 => x"08",
         11900 => x"2e",
         11901 => x"33",
         11902 => x"2e",
         11903 => x"14",
         11904 => x"22",
         11905 => x"78",
         11906 => x"38",
         11907 => x"59",
         11908 => x"80",
         11909 => x"80",
         11910 => x"38",
         11911 => x"51",
         11912 => x"3f",
         11913 => x"08",
         11914 => x"c8",
         11915 => x"b5",
         11916 => x"c8",
         11917 => x"76",
         11918 => x"ff",
         11919 => x"72",
         11920 => x"ff",
         11921 => x"84",
         11922 => x"84",
         11923 => x"70",
         11924 => x"2c",
         11925 => x"08",
         11926 => x"54",
         11927 => x"c8",
         11928 => x"0d",
         11929 => x"53",
         11930 => x"ff",
         11931 => x"72",
         11932 => x"ff",
         11933 => x"84",
         11934 => x"84",
         11935 => x"70",
         11936 => x"2c",
         11937 => x"08",
         11938 => x"54",
         11939 => x"52",
         11940 => x"96",
         11941 => x"b9",
         11942 => x"b9",
         11943 => x"3d",
         11944 => x"14",
         11945 => x"fd",
         11946 => x"b9",
         11947 => x"06",
         11948 => x"d8",
         11949 => x"08",
         11950 => x"d2",
         11951 => x"0d",
         11952 => x"53",
         11953 => x"53",
         11954 => x"56",
         11955 => x"84",
         11956 => x"55",
         11957 => x"08",
         11958 => x"38",
         11959 => x"c8",
         11960 => x"0d",
         11961 => x"75",
         11962 => x"a9",
         11963 => x"c8",
         11964 => x"b9",
         11965 => x"38",
         11966 => x"05",
         11967 => x"2b",
         11968 => x"74",
         11969 => x"76",
         11970 => x"38",
         11971 => x"51",
         11972 => x"3f",
         11973 => x"c8",
         11974 => x"0d",
         11975 => x"84",
         11976 => x"95",
         11977 => x"ed",
         11978 => x"68",
         11979 => x"53",
         11980 => x"05",
         11981 => x"51",
         11982 => x"84",
         11983 => x"5a",
         11984 => x"08",
         11985 => x"75",
         11986 => x"9c",
         11987 => x"11",
         11988 => x"59",
         11989 => x"75",
         11990 => x"38",
         11991 => x"79",
         11992 => x"0c",
         11993 => x"04",
         11994 => x"08",
         11995 => x"5b",
         11996 => x"82",
         11997 => x"a8",
         11998 => x"b9",
         11999 => x"5d",
         12000 => x"c1",
         12001 => x"1d",
         12002 => x"56",
         12003 => x"76",
         12004 => x"38",
         12005 => x"78",
         12006 => x"81",
         12007 => x"54",
         12008 => x"17",
         12009 => x"33",
         12010 => x"b7",
         12011 => x"c8",
         12012 => x"85",
         12013 => x"81",
         12014 => x"18",
         12015 => x"5b",
         12016 => x"cc",
         12017 => x"5e",
         12018 => x"82",
         12019 => x"17",
         12020 => x"11",
         12021 => x"33",
         12022 => x"71",
         12023 => x"81",
         12024 => x"72",
         12025 => x"75",
         12026 => x"ff",
         12027 => x"06",
         12028 => x"70",
         12029 => x"05",
         12030 => x"83",
         12031 => x"ff",
         12032 => x"43",
         12033 => x"53",
         12034 => x"56",
         12035 => x"38",
         12036 => x"7a",
         12037 => x"84",
         12038 => x"07",
         12039 => x"18",
         12040 => x"b9",
         12041 => x"3d",
         12042 => x"54",
         12043 => x"53",
         12044 => x"53",
         12045 => x"52",
         12046 => x"a6",
         12047 => x"84",
         12048 => x"fe",
         12049 => x"b9",
         12050 => x"18",
         12051 => x"08",
         12052 => x"31",
         12053 => x"08",
         12054 => x"a0",
         12055 => x"fe",
         12056 => x"17",
         12057 => x"82",
         12058 => x"06",
         12059 => x"81",
         12060 => x"08",
         12061 => x"05",
         12062 => x"81",
         12063 => x"fe",
         12064 => x"77",
         12065 => x"39",
         12066 => x"92",
         12067 => x"75",
         12068 => x"ff",
         12069 => x"84",
         12070 => x"ff",
         12071 => x"38",
         12072 => x"08",
         12073 => x"f7",
         12074 => x"c8",
         12075 => x"84",
         12076 => x"07",
         12077 => x"05",
         12078 => x"5a",
         12079 => x"9c",
         12080 => x"26",
         12081 => x"7f",
         12082 => x"18",
         12083 => x"33",
         12084 => x"77",
         12085 => x"fe",
         12086 => x"17",
         12087 => x"11",
         12088 => x"71",
         12089 => x"70",
         12090 => x"25",
         12091 => x"83",
         12092 => x"1f",
         12093 => x"59",
         12094 => x"78",
         12095 => x"fe",
         12096 => x"5a",
         12097 => x"81",
         12098 => x"7a",
         12099 => x"94",
         12100 => x"17",
         12101 => x"58",
         12102 => x"34",
         12103 => x"82",
         12104 => x"e7",
         12105 => x"0d",
         12106 => x"56",
         12107 => x"9f",
         12108 => x"55",
         12109 => x"97",
         12110 => x"54",
         12111 => x"8f",
         12112 => x"22",
         12113 => x"59",
         12114 => x"2e",
         12115 => x"80",
         12116 => x"75",
         12117 => x"91",
         12118 => x"75",
         12119 => x"90",
         12120 => x"81",
         12121 => x"55",
         12122 => x"73",
         12123 => x"c4",
         12124 => x"08",
         12125 => x"18",
         12126 => x"38",
         12127 => x"38",
         12128 => x"77",
         12129 => x"81",
         12130 => x"38",
         12131 => x"74",
         12132 => x"82",
         12133 => x"88",
         12134 => x"17",
         12135 => x"0c",
         12136 => x"07",
         12137 => x"18",
         12138 => x"2e",
         12139 => x"91",
         12140 => x"55",
         12141 => x"c8",
         12142 => x"0d",
         12143 => x"78",
         12144 => x"ff",
         12145 => x"76",
         12146 => x"ca",
         12147 => x"c8",
         12148 => x"b9",
         12149 => x"2e",
         12150 => x"84",
         12151 => x"81",
         12152 => x"38",
         12153 => x"08",
         12154 => x"e5",
         12155 => x"73",
         12156 => x"ff",
         12157 => x"84",
         12158 => x"82",
         12159 => x"16",
         12160 => x"94",
         12161 => x"55",
         12162 => x"27",
         12163 => x"81",
         12164 => x"0c",
         12165 => x"81",
         12166 => x"84",
         12167 => x"54",
         12168 => x"ff",
         12169 => x"39",
         12170 => x"51",
         12171 => x"3f",
         12172 => x"08",
         12173 => x"73",
         12174 => x"73",
         12175 => x"56",
         12176 => x"80",
         12177 => x"33",
         12178 => x"56",
         12179 => x"18",
         12180 => x"39",
         12181 => x"52",
         12182 => x"fd",
         12183 => x"b9",
         12184 => x"2e",
         12185 => x"84",
         12186 => x"81",
         12187 => x"38",
         12188 => x"38",
         12189 => x"b9",
         12190 => x"19",
         12191 => x"a1",
         12192 => x"c8",
         12193 => x"08",
         12194 => x"56",
         12195 => x"84",
         12196 => x"27",
         12197 => x"84",
         12198 => x"9c",
         12199 => x"81",
         12200 => x"80",
         12201 => x"ff",
         12202 => x"75",
         12203 => x"c7",
         12204 => x"c8",
         12205 => x"b9",
         12206 => x"e3",
         12207 => x"76",
         12208 => x"d2",
         12209 => x"c8",
         12210 => x"b9",
         12211 => x"2e",
         12212 => x"84",
         12213 => x"81",
         12214 => x"38",
         12215 => x"08",
         12216 => x"fe",
         12217 => x"73",
         12218 => x"ff",
         12219 => x"84",
         12220 => x"80",
         12221 => x"16",
         12222 => x"94",
         12223 => x"55",
         12224 => x"27",
         12225 => x"15",
         12226 => x"84",
         12227 => x"07",
         12228 => x"17",
         12229 => x"77",
         12230 => x"a1",
         12231 => x"74",
         12232 => x"33",
         12233 => x"39",
         12234 => x"bb",
         12235 => x"90",
         12236 => x"56",
         12237 => x"82",
         12238 => x"82",
         12239 => x"33",
         12240 => x"86",
         12241 => x"c8",
         12242 => x"33",
         12243 => x"fa",
         12244 => x"90",
         12245 => x"54",
         12246 => x"84",
         12247 => x"56",
         12248 => x"56",
         12249 => x"db",
         12250 => x"53",
         12251 => x"9c",
         12252 => x"3d",
         12253 => x"fb",
         12254 => x"c8",
         12255 => x"b9",
         12256 => x"2e",
         12257 => x"84",
         12258 => x"a7",
         12259 => x"7d",
         12260 => x"08",
         12261 => x"70",
         12262 => x"ab",
         12263 => x"b9",
         12264 => x"84",
         12265 => x"de",
         12266 => x"93",
         12267 => x"85",
         12268 => x"59",
         12269 => x"77",
         12270 => x"98",
         12271 => x"7b",
         12272 => x"02",
         12273 => x"33",
         12274 => x"5d",
         12275 => x"7b",
         12276 => x"7d",
         12277 => x"9b",
         12278 => x"12",
         12279 => x"2b",
         12280 => x"41",
         12281 => x"58",
         12282 => x"80",
         12283 => x"84",
         12284 => x"57",
         12285 => x"80",
         12286 => x"56",
         12287 => x"7b",
         12288 => x"38",
         12289 => x"41",
         12290 => x"08",
         12291 => x"70",
         12292 => x"8b",
         12293 => x"b9",
         12294 => x"84",
         12295 => x"fe",
         12296 => x"b9",
         12297 => x"74",
         12298 => x"b4",
         12299 => x"c8",
         12300 => x"b9",
         12301 => x"38",
         12302 => x"b9",
         12303 => x"3d",
         12304 => x"16",
         12305 => x"33",
         12306 => x"71",
         12307 => x"7d",
         12308 => x"5d",
         12309 => x"84",
         12310 => x"84",
         12311 => x"84",
         12312 => x"fe",
         12313 => x"08",
         12314 => x"08",
         12315 => x"74",
         12316 => x"d3",
         12317 => x"78",
         12318 => x"92",
         12319 => x"c8",
         12320 => x"b9",
         12321 => x"2e",
         12322 => x"30",
         12323 => x"80",
         12324 => x"7a",
         12325 => x"38",
         12326 => x"95",
         12327 => x"08",
         12328 => x"7b",
         12329 => x"9c",
         12330 => x"26",
         12331 => x"82",
         12332 => x"d2",
         12333 => x"fe",
         12334 => x"84",
         12335 => x"84",
         12336 => x"a7",
         12337 => x"b8",
         12338 => x"19",
         12339 => x"5a",
         12340 => x"76",
         12341 => x"38",
         12342 => x"7a",
         12343 => x"7a",
         12344 => x"06",
         12345 => x"81",
         12346 => x"b8",
         12347 => x"17",
         12348 => x"f1",
         12349 => x"b9",
         12350 => x"2e",
         12351 => x"56",
         12352 => x"b4",
         12353 => x"56",
         12354 => x"9c",
         12355 => x"e5",
         12356 => x"0b",
         12357 => x"90",
         12358 => x"27",
         12359 => x"80",
         12360 => x"ff",
         12361 => x"84",
         12362 => x"56",
         12363 => x"08",
         12364 => x"96",
         12365 => x"2e",
         12366 => x"fe",
         12367 => x"56",
         12368 => x"81",
         12369 => x"08",
         12370 => x"81",
         12371 => x"fe",
         12372 => x"81",
         12373 => x"c8",
         12374 => x"09",
         12375 => x"a6",
         12376 => x"c8",
         12377 => x"34",
         12378 => x"a8",
         12379 => x"84",
         12380 => x"59",
         12381 => x"18",
         12382 => x"eb",
         12383 => x"33",
         12384 => x"2e",
         12385 => x"fe",
         12386 => x"54",
         12387 => x"a0",
         12388 => x"53",
         12389 => x"17",
         12390 => x"f1",
         12391 => x"58",
         12392 => x"79",
         12393 => x"27",
         12394 => x"74",
         12395 => x"fe",
         12396 => x"84",
         12397 => x"5a",
         12398 => x"08",
         12399 => x"cb",
         12400 => x"c8",
         12401 => x"fd",
         12402 => x"b9",
         12403 => x"2e",
         12404 => x"80",
         12405 => x"76",
         12406 => x"9b",
         12407 => x"c8",
         12408 => x"9c",
         12409 => x"11",
         12410 => x"58",
         12411 => x"7b",
         12412 => x"38",
         12413 => x"18",
         12414 => x"33",
         12415 => x"7b",
         12416 => x"79",
         12417 => x"26",
         12418 => x"80",
         12419 => x"39",
         12420 => x"f7",
         12421 => x"c8",
         12422 => x"95",
         12423 => x"fd",
         12424 => x"3d",
         12425 => x"9f",
         12426 => x"05",
         12427 => x"51",
         12428 => x"3f",
         12429 => x"08",
         12430 => x"c8",
         12431 => x"8a",
         12432 => x"b9",
         12433 => x"3d",
         12434 => x"43",
         12435 => x"3d",
         12436 => x"ff",
         12437 => x"84",
         12438 => x"56",
         12439 => x"08",
         12440 => x"0b",
         12441 => x"0c",
         12442 => x"04",
         12443 => x"08",
         12444 => x"81",
         12445 => x"02",
         12446 => x"33",
         12447 => x"81",
         12448 => x"86",
         12449 => x"b9",
         12450 => x"74",
         12451 => x"70",
         12452 => x"83",
         12453 => x"b9",
         12454 => x"57",
         12455 => x"c8",
         12456 => x"87",
         12457 => x"c8",
         12458 => x"80",
         12459 => x"b9",
         12460 => x"2e",
         12461 => x"75",
         12462 => x"7d",
         12463 => x"08",
         12464 => x"5d",
         12465 => x"80",
         12466 => x"19",
         12467 => x"fe",
         12468 => x"80",
         12469 => x"27",
         12470 => x"17",
         12471 => x"29",
         12472 => x"05",
         12473 => x"b4",
         12474 => x"17",
         12475 => x"79",
         12476 => x"76",
         12477 => x"58",
         12478 => x"55",
         12479 => x"74",
         12480 => x"22",
         12481 => x"27",
         12482 => x"81",
         12483 => x"53",
         12484 => x"17",
         12485 => x"ee",
         12486 => x"b9",
         12487 => x"df",
         12488 => x"58",
         12489 => x"56",
         12490 => x"81",
         12491 => x"08",
         12492 => x"70",
         12493 => x"33",
         12494 => x"ee",
         12495 => x"56",
         12496 => x"08",
         12497 => x"b9",
         12498 => x"18",
         12499 => x"08",
         12500 => x"31",
         12501 => x"18",
         12502 => x"ee",
         12503 => x"33",
         12504 => x"2e",
         12505 => x"fe",
         12506 => x"54",
         12507 => x"a0",
         12508 => x"53",
         12509 => x"17",
         12510 => x"ed",
         12511 => x"ca",
         12512 => x"7b",
         12513 => x"55",
         12514 => x"fd",
         12515 => x"9c",
         12516 => x"fd",
         12517 => x"52",
         12518 => x"f2",
         12519 => x"b9",
         12520 => x"84",
         12521 => x"80",
         12522 => x"38",
         12523 => x"08",
         12524 => x"8d",
         12525 => x"c8",
         12526 => x"fd",
         12527 => x"53",
         12528 => x"51",
         12529 => x"3f",
         12530 => x"08",
         12531 => x"9c",
         12532 => x"11",
         12533 => x"5a",
         12534 => x"7b",
         12535 => x"81",
         12536 => x"0c",
         12537 => x"81",
         12538 => x"84",
         12539 => x"55",
         12540 => x"ff",
         12541 => x"84",
         12542 => x"9f",
         12543 => x"8a",
         12544 => x"74",
         12545 => x"06",
         12546 => x"76",
         12547 => x"81",
         12548 => x"38",
         12549 => x"1f",
         12550 => x"75",
         12551 => x"57",
         12552 => x"56",
         12553 => x"7d",
         12554 => x"b8",
         12555 => x"58",
         12556 => x"c3",
         12557 => x"59",
         12558 => x"1a",
         12559 => x"cf",
         12560 => x"0b",
         12561 => x"34",
         12562 => x"80",
         12563 => x"7d",
         12564 => x"ff",
         12565 => x"77",
         12566 => x"34",
         12567 => x"5b",
         12568 => x"17",
         12569 => x"55",
         12570 => x"81",
         12571 => x"59",
         12572 => x"d8",
         12573 => x"57",
         12574 => x"70",
         12575 => x"33",
         12576 => x"05",
         12577 => x"16",
         12578 => x"38",
         12579 => x"0b",
         12580 => x"34",
         12581 => x"83",
         12582 => x"5b",
         12583 => x"80",
         12584 => x"78",
         12585 => x"7a",
         12586 => x"34",
         12587 => x"74",
         12588 => x"f0",
         12589 => x"81",
         12590 => x"34",
         12591 => x"92",
         12592 => x"b9",
         12593 => x"84",
         12594 => x"fd",
         12595 => x"56",
         12596 => x"08",
         12597 => x"84",
         12598 => x"97",
         12599 => x"0b",
         12600 => x"80",
         12601 => x"17",
         12602 => x"58",
         12603 => x"18",
         12604 => x"2a",
         12605 => x"18",
         12606 => x"5a",
         12607 => x"80",
         12608 => x"55",
         12609 => x"16",
         12610 => x"81",
         12611 => x"34",
         12612 => x"ed",
         12613 => x"b9",
         12614 => x"75",
         12615 => x"0c",
         12616 => x"04",
         12617 => x"55",
         12618 => x"17",
         12619 => x"2a",
         12620 => x"ed",
         12621 => x"fd",
         12622 => x"2a",
         12623 => x"cc",
         12624 => x"88",
         12625 => x"80",
         12626 => x"7d",
         12627 => x"80",
         12628 => x"1b",
         12629 => x"fe",
         12630 => x"90",
         12631 => x"94",
         12632 => x"88",
         12633 => x"95",
         12634 => x"55",
         12635 => x"16",
         12636 => x"81",
         12637 => x"34",
         12638 => x"ec",
         12639 => x"b9",
         12640 => x"ff",
         12641 => x"3d",
         12642 => x"b4",
         12643 => x"59",
         12644 => x"80",
         12645 => x"79",
         12646 => x"5b",
         12647 => x"26",
         12648 => x"ba",
         12649 => x"38",
         12650 => x"75",
         12651 => x"af",
         12652 => x"b1",
         12653 => x"05",
         12654 => x"51",
         12655 => x"3f",
         12656 => x"08",
         12657 => x"c8",
         12658 => x"8a",
         12659 => x"b9",
         12660 => x"3d",
         12661 => x"a6",
         12662 => x"3d",
         12663 => x"3d",
         12664 => x"ff",
         12665 => x"84",
         12666 => x"56",
         12667 => x"08",
         12668 => x"81",
         12669 => x"81",
         12670 => x"86",
         12671 => x"38",
         12672 => x"3d",
         12673 => x"58",
         12674 => x"70",
         12675 => x"33",
         12676 => x"05",
         12677 => x"15",
         12678 => x"38",
         12679 => x"b0",
         12680 => x"58",
         12681 => x"81",
         12682 => x"77",
         12683 => x"59",
         12684 => x"55",
         12685 => x"b3",
         12686 => x"77",
         12687 => x"d5",
         12688 => x"c8",
         12689 => x"b9",
         12690 => x"d8",
         12691 => x"3d",
         12692 => x"cb",
         12693 => x"84",
         12694 => x"b1",
         12695 => x"76",
         12696 => x"70",
         12697 => x"57",
         12698 => x"89",
         12699 => x"82",
         12700 => x"ff",
         12701 => x"5d",
         12702 => x"2e",
         12703 => x"80",
         12704 => x"e5",
         12705 => x"72",
         12706 => x"5f",
         12707 => x"81",
         12708 => x"79",
         12709 => x"5b",
         12710 => x"12",
         12711 => x"77",
         12712 => x"38",
         12713 => x"81",
         12714 => x"55",
         12715 => x"58",
         12716 => x"89",
         12717 => x"70",
         12718 => x"58",
         12719 => x"70",
         12720 => x"55",
         12721 => x"09",
         12722 => x"38",
         12723 => x"38",
         12724 => x"70",
         12725 => x"07",
         12726 => x"07",
         12727 => x"7a",
         12728 => x"38",
         12729 => x"1e",
         12730 => x"83",
         12731 => x"38",
         12732 => x"5a",
         12733 => x"39",
         12734 => x"fd",
         12735 => x"7f",
         12736 => x"b1",
         12737 => x"05",
         12738 => x"51",
         12739 => x"3f",
         12740 => x"08",
         12741 => x"c8",
         12742 => x"38",
         12743 => x"6c",
         12744 => x"2e",
         12745 => x"fe",
         12746 => x"51",
         12747 => x"3f",
         12748 => x"08",
         12749 => x"c8",
         12750 => x"38",
         12751 => x"0b",
         12752 => x"88",
         12753 => x"05",
         12754 => x"75",
         12755 => x"57",
         12756 => x"81",
         12757 => x"ff",
         12758 => x"ef",
         12759 => x"cb",
         12760 => x"19",
         12761 => x"33",
         12762 => x"81",
         12763 => x"7e",
         12764 => x"a0",
         12765 => x"8b",
         12766 => x"5d",
         12767 => x"1e",
         12768 => x"33",
         12769 => x"81",
         12770 => x"75",
         12771 => x"c5",
         12772 => x"08",
         12773 => x"bd",
         12774 => x"19",
         12775 => x"33",
         12776 => x"07",
         12777 => x"58",
         12778 => x"83",
         12779 => x"38",
         12780 => x"18",
         12781 => x"5e",
         12782 => x"27",
         12783 => x"8a",
         12784 => x"71",
         12785 => x"08",
         12786 => x"75",
         12787 => x"b5",
         12788 => x"5d",
         12789 => x"08",
         12790 => x"38",
         12791 => x"5f",
         12792 => x"38",
         12793 => x"53",
         12794 => x"81",
         12795 => x"fe",
         12796 => x"84",
         12797 => x"80",
         12798 => x"ff",
         12799 => x"77",
         12800 => x"7f",
         12801 => x"d8",
         12802 => x"7b",
         12803 => x"81",
         12804 => x"79",
         12805 => x"81",
         12806 => x"6a",
         12807 => x"ff",
         12808 => x"7b",
         12809 => x"34",
         12810 => x"58",
         12811 => x"18",
         12812 => x"5b",
         12813 => x"09",
         12814 => x"38",
         12815 => x"5e",
         12816 => x"18",
         12817 => x"2a",
         12818 => x"ed",
         12819 => x"57",
         12820 => x"18",
         12821 => x"aa",
         12822 => x"3d",
         12823 => x"56",
         12824 => x"95",
         12825 => x"78",
         12826 => x"a2",
         12827 => x"c8",
         12828 => x"b9",
         12829 => x"f5",
         12830 => x"5c",
         12831 => x"57",
         12832 => x"16",
         12833 => x"b4",
         12834 => x"33",
         12835 => x"7e",
         12836 => x"81",
         12837 => x"38",
         12838 => x"53",
         12839 => x"81",
         12840 => x"fe",
         12841 => x"84",
         12842 => x"80",
         12843 => x"ff",
         12844 => x"76",
         12845 => x"77",
         12846 => x"38",
         12847 => x"5a",
         12848 => x"81",
         12849 => x"34",
         12850 => x"7b",
         12851 => x"80",
         12852 => x"fe",
         12853 => x"84",
         12854 => x"55",
         12855 => x"08",
         12856 => x"98",
         12857 => x"74",
         12858 => x"e1",
         12859 => x"74",
         12860 => x"7f",
         12861 => x"9d",
         12862 => x"c8",
         12863 => x"c8",
         12864 => x"0d",
         12865 => x"84",
         12866 => x"b1",
         12867 => x"95",
         12868 => x"19",
         12869 => x"2b",
         12870 => x"07",
         12871 => x"56",
         12872 => x"39",
         12873 => x"08",
         12874 => x"fe",
         12875 => x"c8",
         12876 => x"fe",
         12877 => x"84",
         12878 => x"b1",
         12879 => x"81",
         12880 => x"08",
         12881 => x"81",
         12882 => x"fe",
         12883 => x"81",
         12884 => x"c8",
         12885 => x"09",
         12886 => x"db",
         12887 => x"c8",
         12888 => x"34",
         12889 => x"a8",
         12890 => x"84",
         12891 => x"59",
         12892 => x"17",
         12893 => x"a0",
         12894 => x"33",
         12895 => x"2e",
         12896 => x"fe",
         12897 => x"54",
         12898 => x"a0",
         12899 => x"53",
         12900 => x"16",
         12901 => x"e1",
         12902 => x"58",
         12903 => x"81",
         12904 => x"08",
         12905 => x"70",
         12906 => x"33",
         12907 => x"e1",
         12908 => x"5c",
         12909 => x"08",
         12910 => x"84",
         12911 => x"83",
         12912 => x"17",
         12913 => x"08",
         12914 => x"c8",
         12915 => x"74",
         12916 => x"27",
         12917 => x"82",
         12918 => x"7c",
         12919 => x"81",
         12920 => x"38",
         12921 => x"17",
         12922 => x"08",
         12923 => x"52",
         12924 => x"51",
         12925 => x"3f",
         12926 => x"e8",
         12927 => x"0d",
         12928 => x"05",
         12929 => x"05",
         12930 => x"33",
         12931 => x"53",
         12932 => x"05",
         12933 => x"51",
         12934 => x"3f",
         12935 => x"08",
         12936 => x"c8",
         12937 => x"8a",
         12938 => x"b9",
         12939 => x"3d",
         12940 => x"5a",
         12941 => x"3d",
         12942 => x"ff",
         12943 => x"84",
         12944 => x"56",
         12945 => x"08",
         12946 => x"80",
         12947 => x"81",
         12948 => x"86",
         12949 => x"38",
         12950 => x"61",
         12951 => x"12",
         12952 => x"7a",
         12953 => x"51",
         12954 => x"73",
         12955 => x"78",
         12956 => x"83",
         12957 => x"51",
         12958 => x"3f",
         12959 => x"08",
         12960 => x"0c",
         12961 => x"04",
         12962 => x"67",
         12963 => x"96",
         12964 => x"52",
         12965 => x"ff",
         12966 => x"84",
         12967 => x"55",
         12968 => x"08",
         12969 => x"38",
         12970 => x"c8",
         12971 => x"0d",
         12972 => x"66",
         12973 => x"d0",
         12974 => x"95",
         12975 => x"b9",
         12976 => x"84",
         12977 => x"e0",
         12978 => x"cf",
         12979 => x"a0",
         12980 => x"55",
         12981 => x"60",
         12982 => x"86",
         12983 => x"90",
         12984 => x"59",
         12985 => x"17",
         12986 => x"2a",
         12987 => x"17",
         12988 => x"2a",
         12989 => x"17",
         12990 => x"2a",
         12991 => x"17",
         12992 => x"81",
         12993 => x"34",
         12994 => x"e1",
         12995 => x"b9",
         12996 => x"b9",
         12997 => x"3d",
         12998 => x"3d",
         12999 => x"5d",
         13000 => x"9a",
         13001 => x"52",
         13002 => x"ff",
         13003 => x"84",
         13004 => x"84",
         13005 => x"30",
         13006 => x"c8",
         13007 => x"25",
         13008 => x"7a",
         13009 => x"38",
         13010 => x"06",
         13011 => x"81",
         13012 => x"30",
         13013 => x"80",
         13014 => x"7b",
         13015 => x"8c",
         13016 => x"76",
         13017 => x"78",
         13018 => x"80",
         13019 => x"11",
         13020 => x"80",
         13021 => x"08",
         13022 => x"f6",
         13023 => x"33",
         13024 => x"74",
         13025 => x"81",
         13026 => x"38",
         13027 => x"53",
         13028 => x"81",
         13029 => x"fe",
         13030 => x"84",
         13031 => x"80",
         13032 => x"ff",
         13033 => x"76",
         13034 => x"78",
         13035 => x"38",
         13036 => x"56",
         13037 => x"56",
         13038 => x"8b",
         13039 => x"56",
         13040 => x"83",
         13041 => x"75",
         13042 => x"83",
         13043 => x"12",
         13044 => x"2b",
         13045 => x"07",
         13046 => x"70",
         13047 => x"2b",
         13048 => x"07",
         13049 => x"5d",
         13050 => x"56",
         13051 => x"c8",
         13052 => x"0d",
         13053 => x"80",
         13054 => x"8e",
         13055 => x"55",
         13056 => x"3f",
         13057 => x"08",
         13058 => x"c8",
         13059 => x"81",
         13060 => x"84",
         13061 => x"06",
         13062 => x"80",
         13063 => x"57",
         13064 => x"77",
         13065 => x"08",
         13066 => x"70",
         13067 => x"33",
         13068 => x"dc",
         13069 => x"59",
         13070 => x"08",
         13071 => x"81",
         13072 => x"38",
         13073 => x"08",
         13074 => x"b4",
         13075 => x"17",
         13076 => x"b9",
         13077 => x"55",
         13078 => x"08",
         13079 => x"38",
         13080 => x"55",
         13081 => x"09",
         13082 => x"a0",
         13083 => x"b4",
         13084 => x"17",
         13085 => x"7a",
         13086 => x"33",
         13087 => x"e2",
         13088 => x"81",
         13089 => x"b8",
         13090 => x"16",
         13091 => x"da",
         13092 => x"b9",
         13093 => x"2e",
         13094 => x"fe",
         13095 => x"52",
         13096 => x"f8",
         13097 => x"b9",
         13098 => x"84",
         13099 => x"fe",
         13100 => x"b9",
         13101 => x"b9",
         13102 => x"5c",
         13103 => x"18",
         13104 => x"1b",
         13105 => x"75",
         13106 => x"81",
         13107 => x"78",
         13108 => x"8b",
         13109 => x"58",
         13110 => x"77",
         13111 => x"f2",
         13112 => x"7b",
         13113 => x"5c",
         13114 => x"a0",
         13115 => x"fc",
         13116 => x"57",
         13117 => x"e1",
         13118 => x"53",
         13119 => x"b4",
         13120 => x"3d",
         13121 => x"eb",
         13122 => x"c8",
         13123 => x"b9",
         13124 => x"a6",
         13125 => x"5d",
         13126 => x"55",
         13127 => x"81",
         13128 => x"ff",
         13129 => x"f4",
         13130 => x"3d",
         13131 => x"70",
         13132 => x"5b",
         13133 => x"9f",
         13134 => x"b7",
         13135 => x"90",
         13136 => x"75",
         13137 => x"81",
         13138 => x"74",
         13139 => x"75",
         13140 => x"83",
         13141 => x"81",
         13142 => x"51",
         13143 => x"83",
         13144 => x"b9",
         13145 => x"9f",
         13146 => x"b9",
         13147 => x"ff",
         13148 => x"76",
         13149 => x"e0",
         13150 => x"d8",
         13151 => x"d8",
         13152 => x"ff",
         13153 => x"58",
         13154 => x"81",
         13155 => x"56",
         13156 => x"99",
         13157 => x"70",
         13158 => x"ff",
         13159 => x"58",
         13160 => x"89",
         13161 => x"2e",
         13162 => x"e9",
         13163 => x"ff",
         13164 => x"81",
         13165 => x"ff",
         13166 => x"f8",
         13167 => x"26",
         13168 => x"81",
         13169 => x"8f",
         13170 => x"2a",
         13171 => x"70",
         13172 => x"34",
         13173 => x"76",
         13174 => x"05",
         13175 => x"1a",
         13176 => x"70",
         13177 => x"ff",
         13178 => x"58",
         13179 => x"26",
         13180 => x"8f",
         13181 => x"86",
         13182 => x"e5",
         13183 => x"79",
         13184 => x"38",
         13185 => x"56",
         13186 => x"33",
         13187 => x"a0",
         13188 => x"06",
         13189 => x"1a",
         13190 => x"38",
         13191 => x"47",
         13192 => x"3d",
         13193 => x"fe",
         13194 => x"84",
         13195 => x"55",
         13196 => x"08",
         13197 => x"38",
         13198 => x"84",
         13199 => x"a1",
         13200 => x"83",
         13201 => x"51",
         13202 => x"84",
         13203 => x"83",
         13204 => x"55",
         13205 => x"38",
         13206 => x"84",
         13207 => x"a1",
         13208 => x"83",
         13209 => x"56",
         13210 => x"81",
         13211 => x"fe",
         13212 => x"84",
         13213 => x"55",
         13214 => x"08",
         13215 => x"79",
         13216 => x"c4",
         13217 => x"7e",
         13218 => x"76",
         13219 => x"58",
         13220 => x"81",
         13221 => x"ff",
         13222 => x"ef",
         13223 => x"81",
         13224 => x"34",
         13225 => x"d9",
         13226 => x"b9",
         13227 => x"74",
         13228 => x"39",
         13229 => x"fe",
         13230 => x"56",
         13231 => x"84",
         13232 => x"84",
         13233 => x"06",
         13234 => x"80",
         13235 => x"2e",
         13236 => x"75",
         13237 => x"76",
         13238 => x"ee",
         13239 => x"b9",
         13240 => x"84",
         13241 => x"75",
         13242 => x"06",
         13243 => x"84",
         13244 => x"b8",
         13245 => x"98",
         13246 => x"80",
         13247 => x"08",
         13248 => x"38",
         13249 => x"55",
         13250 => x"09",
         13251 => x"d7",
         13252 => x"76",
         13253 => x"52",
         13254 => x"51",
         13255 => x"3f",
         13256 => x"08",
         13257 => x"38",
         13258 => x"59",
         13259 => x"0c",
         13260 => x"be",
         13261 => x"17",
         13262 => x"57",
         13263 => x"81",
         13264 => x"9e",
         13265 => x"70",
         13266 => x"07",
         13267 => x"80",
         13268 => x"38",
         13269 => x"79",
         13270 => x"38",
         13271 => x"51",
         13272 => x"3f",
         13273 => x"08",
         13274 => x"c8",
         13275 => x"ff",
         13276 => x"55",
         13277 => x"fd",
         13278 => x"55",
         13279 => x"38",
         13280 => x"55",
         13281 => x"81",
         13282 => x"ff",
         13283 => x"f4",
         13284 => x"88",
         13285 => x"34",
         13286 => x"59",
         13287 => x"70",
         13288 => x"33",
         13289 => x"05",
         13290 => x"15",
         13291 => x"2e",
         13292 => x"76",
         13293 => x"58",
         13294 => x"81",
         13295 => x"ff",
         13296 => x"da",
         13297 => x"39",
         13298 => x"7a",
         13299 => x"81",
         13300 => x"34",
         13301 => x"d7",
         13302 => x"b9",
         13303 => x"fd",
         13304 => x"57",
         13305 => x"81",
         13306 => x"08",
         13307 => x"81",
         13308 => x"fe",
         13309 => x"84",
         13310 => x"79",
         13311 => x"06",
         13312 => x"84",
         13313 => x"83",
         13314 => x"18",
         13315 => x"08",
         13316 => x"a0",
         13317 => x"8a",
         13318 => x"33",
         13319 => x"2e",
         13320 => x"b9",
         13321 => x"fd",
         13322 => x"5a",
         13323 => x"51",
         13324 => x"3f",
         13325 => x"08",
         13326 => x"c8",
         13327 => x"fd",
         13328 => x"ae",
         13329 => x"58",
         13330 => x"2e",
         13331 => x"fe",
         13332 => x"54",
         13333 => x"a0",
         13334 => x"53",
         13335 => x"18",
         13336 => x"d3",
         13337 => x"a9",
         13338 => x"0d",
         13339 => x"88",
         13340 => x"05",
         13341 => x"57",
         13342 => x"80",
         13343 => x"76",
         13344 => x"80",
         13345 => x"74",
         13346 => x"80",
         13347 => x"86",
         13348 => x"18",
         13349 => x"78",
         13350 => x"c2",
         13351 => x"73",
         13352 => x"a5",
         13353 => x"33",
         13354 => x"9d",
         13355 => x"2e",
         13356 => x"8c",
         13357 => x"9c",
         13358 => x"33",
         13359 => x"81",
         13360 => x"74",
         13361 => x"8c",
         13362 => x"11",
         13363 => x"2b",
         13364 => x"54",
         13365 => x"fd",
         13366 => x"ff",
         13367 => x"70",
         13368 => x"07",
         13369 => x"b9",
         13370 => x"90",
         13371 => x"42",
         13372 => x"58",
         13373 => x"88",
         13374 => x"08",
         13375 => x"38",
         13376 => x"78",
         13377 => x"59",
         13378 => x"51",
         13379 => x"3f",
         13380 => x"55",
         13381 => x"08",
         13382 => x"38",
         13383 => x"b9",
         13384 => x"2e",
         13385 => x"84",
         13386 => x"ff",
         13387 => x"38",
         13388 => x"08",
         13389 => x"81",
         13390 => x"7d",
         13391 => x"74",
         13392 => x"81",
         13393 => x"87",
         13394 => x"73",
         13395 => x"0c",
         13396 => x"04",
         13397 => x"b9",
         13398 => x"3d",
         13399 => x"15",
         13400 => x"d0",
         13401 => x"b9",
         13402 => x"06",
         13403 => x"ad",
         13404 => x"08",
         13405 => x"a7",
         13406 => x"2e",
         13407 => x"7a",
         13408 => x"7c",
         13409 => x"38",
         13410 => x"74",
         13411 => x"e6",
         13412 => x"77",
         13413 => x"fe",
         13414 => x"84",
         13415 => x"56",
         13416 => x"08",
         13417 => x"77",
         13418 => x"17",
         13419 => x"74",
         13420 => x"7e",
         13421 => x"55",
         13422 => x"ff",
         13423 => x"88",
         13424 => x"8c",
         13425 => x"17",
         13426 => x"07",
         13427 => x"18",
         13428 => x"08",
         13429 => x"16",
         13430 => x"76",
         13431 => x"e9",
         13432 => x"31",
         13433 => x"84",
         13434 => x"07",
         13435 => x"16",
         13436 => x"fe",
         13437 => x"54",
         13438 => x"74",
         13439 => x"fe",
         13440 => x"54",
         13441 => x"81",
         13442 => x"39",
         13443 => x"ff",
         13444 => x"b9",
         13445 => x"3d",
         13446 => x"08",
         13447 => x"02",
         13448 => x"87",
         13449 => x"42",
         13450 => x"a2",
         13451 => x"5f",
         13452 => x"80",
         13453 => x"38",
         13454 => x"05",
         13455 => x"9f",
         13456 => x"75",
         13457 => x"9b",
         13458 => x"38",
         13459 => x"85",
         13460 => x"d1",
         13461 => x"80",
         13462 => x"e5",
         13463 => x"10",
         13464 => x"05",
         13465 => x"5a",
         13466 => x"84",
         13467 => x"34",
         13468 => x"b9",
         13469 => x"84",
         13470 => x"33",
         13471 => x"81",
         13472 => x"fe",
         13473 => x"84",
         13474 => x"81",
         13475 => x"81",
         13476 => x"83",
         13477 => x"ab",
         13478 => x"2a",
         13479 => x"8a",
         13480 => x"9f",
         13481 => x"fc",
         13482 => x"52",
         13483 => x"d0",
         13484 => x"b9",
         13485 => x"98",
         13486 => x"74",
         13487 => x"90",
         13488 => x"80",
         13489 => x"88",
         13490 => x"75",
         13491 => x"83",
         13492 => x"80",
         13493 => x"84",
         13494 => x"83",
         13495 => x"81",
         13496 => x"83",
         13497 => x"1f",
         13498 => x"74",
         13499 => x"7e",
         13500 => x"3d",
         13501 => x"70",
         13502 => x"59",
         13503 => x"60",
         13504 => x"ab",
         13505 => x"70",
         13506 => x"07",
         13507 => x"57",
         13508 => x"38",
         13509 => x"84",
         13510 => x"54",
         13511 => x"52",
         13512 => x"cd",
         13513 => x"57",
         13514 => x"08",
         13515 => x"60",
         13516 => x"33",
         13517 => x"05",
         13518 => x"2b",
         13519 => x"8e",
         13520 => x"d4",
         13521 => x"81",
         13522 => x"38",
         13523 => x"61",
         13524 => x"11",
         13525 => x"62",
         13526 => x"e7",
         13527 => x"18",
         13528 => x"82",
         13529 => x"90",
         13530 => x"2b",
         13531 => x"33",
         13532 => x"88",
         13533 => x"71",
         13534 => x"1f",
         13535 => x"82",
         13536 => x"90",
         13537 => x"2b",
         13538 => x"33",
         13539 => x"88",
         13540 => x"71",
         13541 => x"3d",
         13542 => x"3d",
         13543 => x"0c",
         13544 => x"45",
         13545 => x"5a",
         13546 => x"8e",
         13547 => x"79",
         13548 => x"38",
         13549 => x"81",
         13550 => x"87",
         13551 => x"2a",
         13552 => x"45",
         13553 => x"2e",
         13554 => x"61",
         13555 => x"64",
         13556 => x"38",
         13557 => x"47",
         13558 => x"38",
         13559 => x"30",
         13560 => x"7a",
         13561 => x"2e",
         13562 => x"7a",
         13563 => x"8c",
         13564 => x"0b",
         13565 => x"22",
         13566 => x"80",
         13567 => x"74",
         13568 => x"38",
         13569 => x"56",
         13570 => x"17",
         13571 => x"57",
         13572 => x"2e",
         13573 => x"75",
         13574 => x"77",
         13575 => x"fd",
         13576 => x"84",
         13577 => x"10",
         13578 => x"84",
         13579 => x"9f",
         13580 => x"38",
         13581 => x"b9",
         13582 => x"84",
         13583 => x"05",
         13584 => x"2a",
         13585 => x"4c",
         13586 => x"15",
         13587 => x"81",
         13588 => x"7b",
         13589 => x"68",
         13590 => x"ff",
         13591 => x"06",
         13592 => x"4e",
         13593 => x"83",
         13594 => x"38",
         13595 => x"77",
         13596 => x"70",
         13597 => x"57",
         13598 => x"82",
         13599 => x"7c",
         13600 => x"78",
         13601 => x"31",
         13602 => x"80",
         13603 => x"b9",
         13604 => x"62",
         13605 => x"f6",
         13606 => x"2e",
         13607 => x"82",
         13608 => x"ff",
         13609 => x"b9",
         13610 => x"82",
         13611 => x"89",
         13612 => x"18",
         13613 => x"c0",
         13614 => x"38",
         13615 => x"a3",
         13616 => x"76",
         13617 => x"0c",
         13618 => x"84",
         13619 => x"04",
         13620 => x"fe",
         13621 => x"84",
         13622 => x"9f",
         13623 => x"b9",
         13624 => x"7c",
         13625 => x"70",
         13626 => x"57",
         13627 => x"89",
         13628 => x"82",
         13629 => x"ff",
         13630 => x"5d",
         13631 => x"2e",
         13632 => x"80",
         13633 => x"b8",
         13634 => x"08",
         13635 => x"7a",
         13636 => x"5c",
         13637 => x"81",
         13638 => x"ff",
         13639 => x"59",
         13640 => x"26",
         13641 => x"17",
         13642 => x"06",
         13643 => x"9f",
         13644 => x"99",
         13645 => x"e0",
         13646 => x"ff",
         13647 => x"76",
         13648 => x"2a",
         13649 => x"78",
         13650 => x"06",
         13651 => x"ff",
         13652 => x"7a",
         13653 => x"70",
         13654 => x"2a",
         13655 => x"4a",
         13656 => x"2e",
         13657 => x"81",
         13658 => x"5f",
         13659 => x"25",
         13660 => x"7f",
         13661 => x"39",
         13662 => x"05",
         13663 => x"79",
         13664 => x"dd",
         13665 => x"84",
         13666 => x"fe",
         13667 => x"83",
         13668 => x"84",
         13669 => x"40",
         13670 => x"38",
         13671 => x"55",
         13672 => x"75",
         13673 => x"38",
         13674 => x"59",
         13675 => x"81",
         13676 => x"39",
         13677 => x"ff",
         13678 => x"7a",
         13679 => x"56",
         13680 => x"61",
         13681 => x"93",
         13682 => x"2e",
         13683 => x"82",
         13684 => x"4a",
         13685 => x"8b",
         13686 => x"c8",
         13687 => x"26",
         13688 => x"8b",
         13689 => x"5b",
         13690 => x"27",
         13691 => x"8e",
         13692 => x"b9",
         13693 => x"3d",
         13694 => x"d4",
         13695 => x"55",
         13696 => x"86",
         13697 => x"f5",
         13698 => x"38",
         13699 => x"5b",
         13700 => x"fd",
         13701 => x"80",
         13702 => x"80",
         13703 => x"05",
         13704 => x"15",
         13705 => x"38",
         13706 => x"e5",
         13707 => x"55",
         13708 => x"05",
         13709 => x"70",
         13710 => x"34",
         13711 => x"74",
         13712 => x"8b",
         13713 => x"65",
         13714 => x"8c",
         13715 => x"61",
         13716 => x"7b",
         13717 => x"06",
         13718 => x"8e",
         13719 => x"88",
         13720 => x"61",
         13721 => x"81",
         13722 => x"34",
         13723 => x"70",
         13724 => x"80",
         13725 => x"34",
         13726 => x"82",
         13727 => x"61",
         13728 => x"6c",
         13729 => x"ff",
         13730 => x"ad",
         13731 => x"ff",
         13732 => x"74",
         13733 => x"34",
         13734 => x"4c",
         13735 => x"05",
         13736 => x"95",
         13737 => x"61",
         13738 => x"80",
         13739 => x"34",
         13740 => x"05",
         13741 => x"9b",
         13742 => x"61",
         13743 => x"7e",
         13744 => x"67",
         13745 => x"34",
         13746 => x"4c",
         13747 => x"05",
         13748 => x"2a",
         13749 => x"0c",
         13750 => x"08",
         13751 => x"34",
         13752 => x"85",
         13753 => x"61",
         13754 => x"80",
         13755 => x"34",
         13756 => x"05",
         13757 => x"61",
         13758 => x"7c",
         13759 => x"06",
         13760 => x"96",
         13761 => x"88",
         13762 => x"61",
         13763 => x"ff",
         13764 => x"05",
         13765 => x"a6",
         13766 => x"61",
         13767 => x"e5",
         13768 => x"55",
         13769 => x"05",
         13770 => x"70",
         13771 => x"34",
         13772 => x"74",
         13773 => x"83",
         13774 => x"80",
         13775 => x"60",
         13776 => x"4b",
         13777 => x"34",
         13778 => x"53",
         13779 => x"51",
         13780 => x"3f",
         13781 => x"b9",
         13782 => x"e7",
         13783 => x"5c",
         13784 => x"87",
         13785 => x"61",
         13786 => x"76",
         13787 => x"58",
         13788 => x"55",
         13789 => x"63",
         13790 => x"62",
         13791 => x"c0",
         13792 => x"ff",
         13793 => x"81",
         13794 => x"f8",
         13795 => x"34",
         13796 => x"7c",
         13797 => x"64",
         13798 => x"46",
         13799 => x"2a",
         13800 => x"70",
         13801 => x"34",
         13802 => x"56",
         13803 => x"7c",
         13804 => x"76",
         13805 => x"38",
         13806 => x"54",
         13807 => x"52",
         13808 => x"c5",
         13809 => x"b9",
         13810 => x"e6",
         13811 => x"61",
         13812 => x"76",
         13813 => x"58",
         13814 => x"55",
         13815 => x"78",
         13816 => x"31",
         13817 => x"c9",
         13818 => x"05",
         13819 => x"2e",
         13820 => x"77",
         13821 => x"2e",
         13822 => x"56",
         13823 => x"66",
         13824 => x"75",
         13825 => x"7a",
         13826 => x"79",
         13827 => x"d2",
         13828 => x"c8",
         13829 => x"38",
         13830 => x"76",
         13831 => x"75",
         13832 => x"58",
         13833 => x"93",
         13834 => x"6c",
         13835 => x"26",
         13836 => x"58",
         13837 => x"83",
         13838 => x"7d",
         13839 => x"61",
         13840 => x"06",
         13841 => x"b3",
         13842 => x"61",
         13843 => x"75",
         13844 => x"57",
         13845 => x"59",
         13846 => x"80",
         13847 => x"ff",
         13848 => x"60",
         13849 => x"47",
         13850 => x"81",
         13851 => x"34",
         13852 => x"05",
         13853 => x"83",
         13854 => x"67",
         13855 => x"6c",
         13856 => x"c1",
         13857 => x"51",
         13858 => x"3f",
         13859 => x"05",
         13860 => x"c8",
         13861 => x"bf",
         13862 => x"67",
         13863 => x"84",
         13864 => x"67",
         13865 => x"7e",
         13866 => x"05",
         13867 => x"83",
         13868 => x"6b",
         13869 => x"05",
         13870 => x"d4",
         13871 => x"c9",
         13872 => x"61",
         13873 => x"34",
         13874 => x"45",
         13875 => x"cb",
         13876 => x"90",
         13877 => x"61",
         13878 => x"34",
         13879 => x"5f",
         13880 => x"cd",
         13881 => x"54",
         13882 => x"52",
         13883 => x"c2",
         13884 => x"57",
         13885 => x"08",
         13886 => x"80",
         13887 => x"79",
         13888 => x"dd",
         13889 => x"84",
         13890 => x"f7",
         13891 => x"b9",
         13892 => x"b9",
         13893 => x"3d",
         13894 => x"d4",
         13895 => x"55",
         13896 => x"74",
         13897 => x"45",
         13898 => x"39",
         13899 => x"78",
         13900 => x"81",
         13901 => x"fc",
         13902 => x"74",
         13903 => x"38",
         13904 => x"98",
         13905 => x"fc",
         13906 => x"82",
         13907 => x"57",
         13908 => x"80",
         13909 => x"76",
         13910 => x"38",
         13911 => x"51",
         13912 => x"3f",
         13913 => x"08",
         13914 => x"87",
         13915 => x"2a",
         13916 => x"5c",
         13917 => x"b9",
         13918 => x"80",
         13919 => x"47",
         13920 => x"0a",
         13921 => x"cb",
         13922 => x"f8",
         13923 => x"b9",
         13924 => x"ff",
         13925 => x"e6",
         13926 => x"d3",
         13927 => x"2a",
         13928 => x"bf",
         13929 => x"f8",
         13930 => x"81",
         13931 => x"80",
         13932 => x"38",
         13933 => x"ab",
         13934 => x"a0",
         13935 => x"88",
         13936 => x"61",
         13937 => x"75",
         13938 => x"7a",
         13939 => x"34",
         13940 => x"57",
         13941 => x"05",
         13942 => x"39",
         13943 => x"c3",
         13944 => x"61",
         13945 => x"34",
         13946 => x"c5",
         13947 => x"cc",
         13948 => x"05",
         13949 => x"a4",
         13950 => x"88",
         13951 => x"61",
         13952 => x"7c",
         13953 => x"78",
         13954 => x"34",
         13955 => x"56",
         13956 => x"05",
         13957 => x"ac",
         13958 => x"61",
         13959 => x"80",
         13960 => x"34",
         13961 => x"05",
         13962 => x"b0",
         13963 => x"61",
         13964 => x"86",
         13965 => x"34",
         13966 => x"05",
         13967 => x"61",
         13968 => x"34",
         13969 => x"c2",
         13970 => x"61",
         13971 => x"83",
         13972 => x"57",
         13973 => x"81",
         13974 => x"76",
         13975 => x"58",
         13976 => x"55",
         13977 => x"f9",
         13978 => x"70",
         13979 => x"33",
         13980 => x"05",
         13981 => x"15",
         13982 => x"38",
         13983 => x"81",
         13984 => x"60",
         13985 => x"fe",
         13986 => x"81",
         13987 => x"c8",
         13988 => x"38",
         13989 => x"61",
         13990 => x"62",
         13991 => x"34",
         13992 => x"b9",
         13993 => x"60",
         13994 => x"fe",
         13995 => x"fc",
         13996 => x"0b",
         13997 => x"0c",
         13998 => x"84",
         13999 => x"04",
         14000 => x"7b",
         14001 => x"70",
         14002 => x"34",
         14003 => x"81",
         14004 => x"ff",
         14005 => x"61",
         14006 => x"ff",
         14007 => x"34",
         14008 => x"05",
         14009 => x"87",
         14010 => x"61",
         14011 => x"ff",
         14012 => x"34",
         14013 => x"05",
         14014 => x"34",
         14015 => x"b1",
         14016 => x"86",
         14017 => x"52",
         14018 => x"be",
         14019 => x"80",
         14020 => x"80",
         14021 => x"05",
         14022 => x"17",
         14023 => x"38",
         14024 => x"d2",
         14025 => x"05",
         14026 => x"55",
         14027 => x"70",
         14028 => x"34",
         14029 => x"70",
         14030 => x"34",
         14031 => x"34",
         14032 => x"83",
         14033 => x"80",
         14034 => x"e5",
         14035 => x"c1",
         14036 => x"05",
         14037 => x"61",
         14038 => x"34",
         14039 => x"5b",
         14040 => x"e8",
         14041 => x"88",
         14042 => x"61",
         14043 => x"34",
         14044 => x"56",
         14045 => x"ea",
         14046 => x"98",
         14047 => x"61",
         14048 => x"34",
         14049 => x"ec",
         14050 => x"61",
         14051 => x"34",
         14052 => x"ee",
         14053 => x"61",
         14054 => x"34",
         14055 => x"34",
         14056 => x"34",
         14057 => x"1f",
         14058 => x"79",
         14059 => x"b2",
         14060 => x"81",
         14061 => x"52",
         14062 => x"bd",
         14063 => x"61",
         14064 => x"a6",
         14065 => x"0d",
         14066 => x"5b",
         14067 => x"ff",
         14068 => x"57",
         14069 => x"b8",
         14070 => x"59",
         14071 => x"05",
         14072 => x"78",
         14073 => x"ff",
         14074 => x"7b",
         14075 => x"81",
         14076 => x"8d",
         14077 => x"74",
         14078 => x"38",
         14079 => x"81",
         14080 => x"81",
         14081 => x"8a",
         14082 => x"77",
         14083 => x"38",
         14084 => x"7a",
         14085 => x"38",
         14086 => x"84",
         14087 => x"8e",
         14088 => x"f7",
         14089 => x"02",
         14090 => x"05",
         14091 => x"77",
         14092 => x"d5",
         14093 => x"08",
         14094 => x"24",
         14095 => x"17",
         14096 => x"8c",
         14097 => x"77",
         14098 => x"16",
         14099 => x"24",
         14100 => x"84",
         14101 => x"19",
         14102 => x"8b",
         14103 => x"8b",
         14104 => x"54",
         14105 => x"17",
         14106 => x"51",
         14107 => x"3f",
         14108 => x"70",
         14109 => x"07",
         14110 => x"30",
         14111 => x"81",
         14112 => x"0c",
         14113 => x"d3",
         14114 => x"76",
         14115 => x"3f",
         14116 => x"e3",
         14117 => x"80",
         14118 => x"8d",
         14119 => x"80",
         14120 => x"55",
         14121 => x"81",
         14122 => x"ff",
         14123 => x"f4",
         14124 => x"08",
         14125 => x"8a",
         14126 => x"38",
         14127 => x"76",
         14128 => x"38",
         14129 => x"8c",
         14130 => x"77",
         14131 => x"16",
         14132 => x"24",
         14133 => x"84",
         14134 => x"19",
         14135 => x"7c",
         14136 => x"24",
         14137 => x"3d",
         14138 => x"55",
         14139 => x"05",
         14140 => x"51",
         14141 => x"3f",
         14142 => x"08",
         14143 => x"7a",
         14144 => x"ff",
         14145 => x"c8",
         14146 => x"0d",
         14147 => x"ff",
         14148 => x"75",
         14149 => x"52",
         14150 => x"ff",
         14151 => x"74",
         14152 => x"30",
         14153 => x"9f",
         14154 => x"52",
         14155 => x"ff",
         14156 => x"52",
         14157 => x"eb",
         14158 => x"39",
         14159 => x"c8",
         14160 => x"0d",
         14161 => x"0d",
         14162 => x"05",
         14163 => x"52",
         14164 => x"72",
         14165 => x"90",
         14166 => x"ff",
         14167 => x"71",
         14168 => x"0c",
         14169 => x"04",
         14170 => x"73",
         14171 => x"83",
         14172 => x"81",
         14173 => x"73",
         14174 => x"38",
         14175 => x"22",
         14176 => x"2e",
         14177 => x"12",
         14178 => x"ff",
         14179 => x"71",
         14180 => x"8d",
         14181 => x"83",
         14182 => x"70",
         14183 => x"e1",
         14184 => x"12",
         14185 => x"06",
         14186 => x"0c",
         14187 => x"0d",
         14188 => x"0d",
         14189 => x"22",
         14190 => x"96",
         14191 => x"51",
         14192 => x"80",
         14193 => x"38",
         14194 => x"84",
         14195 => x"84",
         14196 => x"71",
         14197 => x"09",
         14198 => x"38",
         14199 => x"26",
         14200 => x"10",
         14201 => x"05",
         14202 => x"b9",
         14203 => x"84",
         14204 => x"fb",
         14205 => x"51",
         14206 => x"ff",
         14207 => x"38",
         14208 => x"ff",
         14209 => x"8c",
         14210 => x"9f",
         14211 => x"d9",
         14212 => x"82",
         14213 => x"75",
         14214 => x"80",
         14215 => x"26",
         14216 => x"53",
         14217 => x"38",
         14218 => x"05",
         14219 => x"71",
         14220 => x"56",
         14221 => x"70",
         14222 => x"70",
         14223 => x"38",
         14224 => x"73",
         14225 => x"70",
         14226 => x"22",
         14227 => x"70",
         14228 => x"79",
         14229 => x"55",
         14230 => x"2e",
         14231 => x"51",
         14232 => x"c8",
         14233 => x"0d",
         14234 => x"80",
         14235 => x"39",
         14236 => x"ea",
         14237 => x"10",
         14238 => x"05",
         14239 => x"04",
         14240 => x"70",
         14241 => x"06",
         14242 => x"51",
         14243 => x"b0",
         14244 => x"ff",
         14245 => x"51",
         14246 => x"16",
         14247 => x"ff",
         14248 => x"e6",
         14249 => x"70",
         14250 => x"06",
         14251 => x"39",
         14252 => x"83",
         14253 => x"57",
         14254 => x"e0",
         14255 => x"ff",
         14256 => x"51",
         14257 => x"16",
         14258 => x"ff",
         14259 => x"ff",
         14260 => x"73",
         14261 => x"76",
         14262 => x"83",
         14263 => x"58",
         14264 => x"a6",
         14265 => x"31",
         14266 => x"70",
         14267 => x"fe",
         14268 => x"00",
         14269 => x"ff",
         14270 => x"ff",
         14271 => x"ff",
         14272 => x"00",
         14273 => x"8b",
         14274 => x"80",
         14275 => x"75",
         14276 => x"6a",
         14277 => x"5f",
         14278 => x"54",
         14279 => x"49",
         14280 => x"3e",
         14281 => x"33",
         14282 => x"28",
         14283 => x"1d",
         14284 => x"12",
         14285 => x"07",
         14286 => x"fc",
         14287 => x"f1",
         14288 => x"e6",
         14289 => x"db",
         14290 => x"d0",
         14291 => x"c5",
         14292 => x"ba",
         14293 => x"bf",
         14294 => x"59",
         14295 => x"59",
         14296 => x"59",
         14297 => x"59",
         14298 => x"59",
         14299 => x"59",
         14300 => x"59",
         14301 => x"59",
         14302 => x"59",
         14303 => x"59",
         14304 => x"59",
         14305 => x"59",
         14306 => x"59",
         14307 => x"59",
         14308 => x"59",
         14309 => x"59",
         14310 => x"59",
         14311 => x"59",
         14312 => x"59",
         14313 => x"59",
         14314 => x"59",
         14315 => x"59",
         14316 => x"59",
         14317 => x"59",
         14318 => x"59",
         14319 => x"59",
         14320 => x"59",
         14321 => x"59",
         14322 => x"59",
         14323 => x"59",
         14324 => x"59",
         14325 => x"59",
         14326 => x"59",
         14327 => x"59",
         14328 => x"59",
         14329 => x"59",
         14330 => x"59",
         14331 => x"59",
         14332 => x"59",
         14333 => x"59",
         14334 => x"59",
         14335 => x"59",
         14336 => x"71",
         14337 => x"59",
         14338 => x"59",
         14339 => x"59",
         14340 => x"59",
         14341 => x"59",
         14342 => x"59",
         14343 => x"59",
         14344 => x"59",
         14345 => x"59",
         14346 => x"59",
         14347 => x"59",
         14348 => x"59",
         14349 => x"59",
         14350 => x"59",
         14351 => x"59",
         14352 => x"59",
         14353 => x"07",
         14354 => x"06",
         14355 => x"59",
         14356 => x"8a",
         14357 => x"a8",
         14358 => x"67",
         14359 => x"2c",
         14360 => x"ce",
         14361 => x"59",
         14362 => x"59",
         14363 => x"59",
         14364 => x"59",
         14365 => x"59",
         14366 => x"59",
         14367 => x"59",
         14368 => x"59",
         14369 => x"59",
         14370 => x"59",
         14371 => x"59",
         14372 => x"59",
         14373 => x"59",
         14374 => x"59",
         14375 => x"59",
         14376 => x"59",
         14377 => x"59",
         14378 => x"59",
         14379 => x"59",
         14380 => x"59",
         14381 => x"59",
         14382 => x"59",
         14383 => x"59",
         14384 => x"59",
         14385 => x"59",
         14386 => x"59",
         14387 => x"59",
         14388 => x"59",
         14389 => x"59",
         14390 => x"59",
         14391 => x"59",
         14392 => x"59",
         14393 => x"59",
         14394 => x"59",
         14395 => x"59",
         14396 => x"59",
         14397 => x"59",
         14398 => x"59",
         14399 => x"59",
         14400 => x"59",
         14401 => x"59",
         14402 => x"59",
         14403 => x"59",
         14404 => x"59",
         14405 => x"59",
         14406 => x"59",
         14407 => x"59",
         14408 => x"59",
         14409 => x"59",
         14410 => x"59",
         14411 => x"59",
         14412 => x"59",
         14413 => x"ab",
         14414 => x"70",
         14415 => x"59",
         14416 => x"59",
         14417 => x"59",
         14418 => x"59",
         14419 => x"59",
         14420 => x"59",
         14421 => x"59",
         14422 => x"59",
         14423 => x"63",
         14424 => x"58",
         14425 => x"59",
         14426 => x"41",
         14427 => x"59",
         14428 => x"51",
         14429 => x"47",
         14430 => x"3a",
         14431 => x"22",
         14432 => x"3a",
         14433 => x"46",
         14434 => x"52",
         14435 => x"5e",
         14436 => x"2e",
         14437 => x"97",
         14438 => x"85",
         14439 => x"01",
         14440 => x"4f",
         14441 => x"21",
         14442 => x"de",
         14443 => x"9b",
         14444 => x"74",
         14445 => x"cb",
         14446 => x"a3",
         14447 => x"12",
         14448 => x"2a",
         14449 => x"de",
         14450 => x"01",
         14451 => x"0b",
         14452 => x"9b",
         14453 => x"de",
         14454 => x"de",
         14455 => x"12",
         14456 => x"a3",
         14457 => x"74",
         14458 => x"4f",
         14459 => x"7c",
         14460 => x"95",
         14461 => x"ba",
         14462 => x"db",
         14463 => x"3c",
         14464 => x"00",
         14465 => x"55",
         14466 => x"a5",
         14467 => x"62",
         14468 => x"62",
         14469 => x"62",
         14470 => x"62",
         14471 => x"62",
         14472 => x"62",
         14473 => x"3b",
         14474 => x"62",
         14475 => x"62",
         14476 => x"62",
         14477 => x"62",
         14478 => x"62",
         14479 => x"62",
         14480 => x"62",
         14481 => x"62",
         14482 => x"62",
         14483 => x"62",
         14484 => x"62",
         14485 => x"62",
         14486 => x"62",
         14487 => x"62",
         14488 => x"62",
         14489 => x"62",
         14490 => x"62",
         14491 => x"62",
         14492 => x"62",
         14493 => x"62",
         14494 => x"62",
         14495 => x"62",
         14496 => x"7a",
         14497 => x"68",
         14498 => x"55",
         14499 => x"42",
         14500 => x"6c",
         14501 => x"30",
         14502 => x"1d",
         14503 => x"85",
         14504 => x"62",
         14505 => x"85",
         14506 => x"0d",
         14507 => x"8a",
         14508 => x"b6",
         14509 => x"94",
         14510 => x"fb",
         14511 => x"e9",
         14512 => x"d7",
         14513 => x"c8",
         14514 => x"62",
         14515 => x"6c",
         14516 => x"08",
         14517 => x"77",
         14518 => x"49",
         14519 => x"a0",
         14520 => x"7d",
         14521 => x"5c",
         14522 => x"32",
         14523 => x"02",
         14524 => x"89",
         14525 => x"dc",
         14526 => x"cb",
         14527 => x"89",
         14528 => x"89",
         14529 => x"89",
         14530 => x"89",
         14531 => x"89",
         14532 => x"89",
         14533 => x"a5",
         14534 => x"b3",
         14535 => x"6a",
         14536 => x"89",
         14537 => x"89",
         14538 => x"89",
         14539 => x"89",
         14540 => x"89",
         14541 => x"89",
         14542 => x"89",
         14543 => x"89",
         14544 => x"89",
         14545 => x"89",
         14546 => x"89",
         14547 => x"89",
         14548 => x"89",
         14549 => x"89",
         14550 => x"89",
         14551 => x"89",
         14552 => x"89",
         14553 => x"89",
         14554 => x"89",
         14555 => x"27",
         14556 => x"89",
         14557 => x"89",
         14558 => x"89",
         14559 => x"ca",
         14560 => x"d9",
         14561 => x"7b",
         14562 => x"89",
         14563 => x"89",
         14564 => x"89",
         14565 => x"89",
         14566 => x"60",
         14567 => x"89",
         14568 => x"43",
         14569 => x"ac",
         14570 => x"21",
         14571 => x"21",
         14572 => x"21",
         14573 => x"21",
         14574 => x"21",
         14575 => x"21",
         14576 => x"fc",
         14577 => x"21",
         14578 => x"21",
         14579 => x"21",
         14580 => x"21",
         14581 => x"21",
         14582 => x"21",
         14583 => x"21",
         14584 => x"21",
         14585 => x"21",
         14586 => x"21",
         14587 => x"21",
         14588 => x"21",
         14589 => x"21",
         14590 => x"21",
         14591 => x"21",
         14592 => x"21",
         14593 => x"21",
         14594 => x"21",
         14595 => x"21",
         14596 => x"21",
         14597 => x"21",
         14598 => x"21",
         14599 => x"be",
         14600 => x"06",
         14601 => x"f3",
         14602 => x"e0",
         14603 => x"ce",
         14604 => x"91",
         14605 => x"7e",
         14606 => x"6e",
         14607 => x"21",
         14608 => x"5e",
         14609 => x"4e",
         14610 => x"3c",
         14611 => x"2a",
         14612 => x"18",
         14613 => x"89",
         14614 => x"78",
         14615 => x"67",
         14616 => x"50",
         14617 => x"21",
         14618 => x"9a",
         14619 => x"7b",
         14620 => x"d7",
         14621 => x"d7",
         14622 => x"d7",
         14623 => x"d7",
         14624 => x"d7",
         14625 => x"d7",
         14626 => x"d7",
         14627 => x"d7",
         14628 => x"d7",
         14629 => x"d7",
         14630 => x"d7",
         14631 => x"d7",
         14632 => x"d7",
         14633 => x"f9",
         14634 => x"d7",
         14635 => x"d7",
         14636 => x"d7",
         14637 => x"d7",
         14638 => x"d7",
         14639 => x"d7",
         14640 => x"c5",
         14641 => x"d7",
         14642 => x"d7",
         14643 => x"50",
         14644 => x"d7",
         14645 => x"67",
         14646 => x"d8",
         14647 => x"39",
         14648 => x"e5",
         14649 => x"d2",
         14650 => x"c6",
         14651 => x"bb",
         14652 => x"b0",
         14653 => x"a5",
         14654 => x"9a",
         14655 => x"8e",
         14656 => x"80",
         14657 => x"01",
         14658 => x"fd",
         14659 => x"fd",
         14660 => x"49",
         14661 => x"fd",
         14662 => x"fd",
         14663 => x"fd",
         14664 => x"fd",
         14665 => x"fd",
         14666 => x"fd",
         14667 => x"fd",
         14668 => x"fd",
         14669 => x"fd",
         14670 => x"7f",
         14671 => x"0d",
         14672 => x"fd",
         14673 => x"fd",
         14674 => x"fd",
         14675 => x"fd",
         14676 => x"fd",
         14677 => x"fd",
         14678 => x"fd",
         14679 => x"fd",
         14680 => x"fd",
         14681 => x"fd",
         14682 => x"fd",
         14683 => x"fd",
         14684 => x"fd",
         14685 => x"fd",
         14686 => x"fd",
         14687 => x"fd",
         14688 => x"fd",
         14689 => x"fd",
         14690 => x"fd",
         14691 => x"fd",
         14692 => x"fd",
         14693 => x"fd",
         14694 => x"fd",
         14695 => x"fd",
         14696 => x"fd",
         14697 => x"fd",
         14698 => x"fd",
         14699 => x"fd",
         14700 => x"fd",
         14701 => x"fd",
         14702 => x"fd",
         14703 => x"fd",
         14704 => x"fd",
         14705 => x"fd",
         14706 => x"fd",
         14707 => x"fd",
         14708 => x"1d",
         14709 => x"fd",
         14710 => x"fd",
         14711 => x"fd",
         14712 => x"fd",
         14713 => x"17",
         14714 => x"fd",
         14715 => x"fd",
         14716 => x"fd",
         14717 => x"fd",
         14718 => x"fd",
         14719 => x"fd",
         14720 => x"fd",
         14721 => x"fd",
         14722 => x"fd",
         14723 => x"fd",
         14724 => x"2b",
         14725 => x"e1",
         14726 => x"b8",
         14727 => x"b8",
         14728 => x"b8",
         14729 => x"fd",
         14730 => x"e1",
         14731 => x"fd",
         14732 => x"fd",
         14733 => x"ff",
         14734 => x"fd",
         14735 => x"fd",
         14736 => x"16",
         14737 => x"0f",
         14738 => x"fd",
         14739 => x"fd",
         14740 => x"58",
         14741 => x"fd",
         14742 => x"18",
         14743 => x"fd",
         14744 => x"fd",
         14745 => x"17",
         14746 => x"69",
         14747 => x"00",
         14748 => x"63",
         14749 => x"00",
         14750 => x"69",
         14751 => x"00",
         14752 => x"61",
         14753 => x"00",
         14754 => x"65",
         14755 => x"00",
         14756 => x"65",
         14757 => x"00",
         14758 => x"70",
         14759 => x"00",
         14760 => x"66",
         14761 => x"00",
         14762 => x"6d",
         14763 => x"00",
         14764 => x"00",
         14765 => x"00",
         14766 => x"00",
         14767 => x"00",
         14768 => x"00",
         14769 => x"00",
         14770 => x"00",
         14771 => x"6c",
         14772 => x"00",
         14773 => x"00",
         14774 => x"74",
         14775 => x"00",
         14776 => x"65",
         14777 => x"00",
         14778 => x"6f",
         14779 => x"00",
         14780 => x"74",
         14781 => x"00",
         14782 => x"00",
         14783 => x"00",
         14784 => x"73",
         14785 => x"00",
         14786 => x"73",
         14787 => x"00",
         14788 => x"6f",
         14789 => x"00",
         14790 => x"00",
         14791 => x"6e",
         14792 => x"20",
         14793 => x"6f",
         14794 => x"00",
         14795 => x"61",
         14796 => x"65",
         14797 => x"69",
         14798 => x"72",
         14799 => x"74",
         14800 => x"00",
         14801 => x"20",
         14802 => x"79",
         14803 => x"65",
         14804 => x"69",
         14805 => x"2e",
         14806 => x"00",
         14807 => x"75",
         14808 => x"63",
         14809 => x"74",
         14810 => x"6d",
         14811 => x"2e",
         14812 => x"00",
         14813 => x"65",
         14814 => x"20",
         14815 => x"6b",
         14816 => x"00",
         14817 => x"65",
         14818 => x"2c",
         14819 => x"65",
         14820 => x"69",
         14821 => x"63",
         14822 => x"65",
         14823 => x"64",
         14824 => x"00",
         14825 => x"6d",
         14826 => x"61",
         14827 => x"74",
         14828 => x"00",
         14829 => x"63",
         14830 => x"61",
         14831 => x"6c",
         14832 => x"69",
         14833 => x"79",
         14834 => x"6d",
         14835 => x"75",
         14836 => x"6f",
         14837 => x"69",
         14838 => x"00",
         14839 => x"6b",
         14840 => x"74",
         14841 => x"61",
         14842 => x"64",
         14843 => x"00",
         14844 => x"76",
         14845 => x"75",
         14846 => x"72",
         14847 => x"20",
         14848 => x"61",
         14849 => x"2e",
         14850 => x"00",
         14851 => x"69",
         14852 => x"72",
         14853 => x"20",
         14854 => x"74",
         14855 => x"65",
         14856 => x"00",
         14857 => x"65",
         14858 => x"6e",
         14859 => x"20",
         14860 => x"61",
         14861 => x"2e",
         14862 => x"00",
         14863 => x"65",
         14864 => x"72",
         14865 => x"79",
         14866 => x"69",
         14867 => x"2e",
         14868 => x"00",
         14869 => x"65",
         14870 => x"64",
         14871 => x"65",
         14872 => x"00",
         14873 => x"61",
         14874 => x"20",
         14875 => x"65",
         14876 => x"65",
         14877 => x"00",
         14878 => x"70",
         14879 => x"20",
         14880 => x"6e",
         14881 => x"00",
         14882 => x"66",
         14883 => x"20",
         14884 => x"6e",
         14885 => x"00",
         14886 => x"6b",
         14887 => x"74",
         14888 => x"61",
         14889 => x"00",
         14890 => x"65",
         14891 => x"6c",
         14892 => x"72",
         14893 => x"00",
         14894 => x"6b",
         14895 => x"72",
         14896 => x"00",
         14897 => x"63",
         14898 => x"2e",
         14899 => x"00",
         14900 => x"75",
         14901 => x"74",
         14902 => x"25",
         14903 => x"74",
         14904 => x"75",
         14905 => x"74",
         14906 => x"73",
         14907 => x"0a",
         14908 => x"00",
         14909 => x"64",
         14910 => x"00",
         14911 => x"6c",
         14912 => x"00",
         14913 => x"00",
         14914 => x"58",
         14915 => x"00",
         14916 => x"00",
         14917 => x"00",
         14918 => x"00",
         14919 => x"58",
         14920 => x"00",
         14921 => x"20",
         14922 => x"20",
         14923 => x"00",
         14924 => x"00",
         14925 => x"25",
         14926 => x"00",
         14927 => x"30",
         14928 => x"30",
         14929 => x"00",
         14930 => x"32",
         14931 => x"00",
         14932 => x"55",
         14933 => x"65",
         14934 => x"30",
         14935 => x"20",
         14936 => x"25",
         14937 => x"2a",
         14938 => x"00",
         14939 => x"00",
         14940 => x"20",
         14941 => x"65",
         14942 => x"64",
         14943 => x"73",
         14944 => x"20",
         14945 => x"20",
         14946 => x"20",
         14947 => x"25",
         14948 => x"78",
         14949 => x"00",
         14950 => x"20",
         14951 => x"20",
         14952 => x"72",
         14953 => x"20",
         14954 => x"20",
         14955 => x"20",
         14956 => x"20",
         14957 => x"25",
         14958 => x"78",
         14959 => x"00",
         14960 => x"20",
         14961 => x"65",
         14962 => x"70",
         14963 => x"61",
         14964 => x"65",
         14965 => x"00",
         14966 => x"54",
         14967 => x"58",
         14968 => x"74",
         14969 => x"75",
         14970 => x"00",
         14971 => x"54",
         14972 => x"58",
         14973 => x"74",
         14974 => x"75",
         14975 => x"00",
         14976 => x"54",
         14977 => x"58",
         14978 => x"74",
         14979 => x"75",
         14980 => x"00",
         14981 => x"54",
         14982 => x"58",
         14983 => x"74",
         14984 => x"75",
         14985 => x"00",
         14986 => x"54",
         14987 => x"52",
         14988 => x"74",
         14989 => x"75",
         14990 => x"00",
         14991 => x"54",
         14992 => x"44",
         14993 => x"74",
         14994 => x"75",
         14995 => x"00",
         14996 => x"20",
         14997 => x"65",
         14998 => x"70",
         14999 => x"00",
         15000 => x"65",
         15001 => x"6e",
         15002 => x"72",
         15003 => x"00",
         15004 => x"74",
         15005 => x"20",
         15006 => x"74",
         15007 => x"72",
         15008 => x"00",
         15009 => x"62",
         15010 => x"67",
         15011 => x"6d",
         15012 => x"2e",
         15013 => x"00",
         15014 => x"6f",
         15015 => x"63",
         15016 => x"74",
         15017 => x"00",
         15018 => x"5f",
         15019 => x"2e",
         15020 => x"00",
         15021 => x"6c",
         15022 => x"74",
         15023 => x"6e",
         15024 => x"61",
         15025 => x"65",
         15026 => x"20",
         15027 => x"64",
         15028 => x"20",
         15029 => x"61",
         15030 => x"69",
         15031 => x"20",
         15032 => x"75",
         15033 => x"79",
         15034 => x"00",
         15035 => x"00",
         15036 => x"5c",
         15037 => x"00",
         15038 => x"00",
         15039 => x"20",
         15040 => x"6d",
         15041 => x"2e",
         15042 => x"00",
         15043 => x"00",
         15044 => x"00",
         15045 => x"5c",
         15046 => x"25",
         15047 => x"73",
         15048 => x"00",
         15049 => x"64",
         15050 => x"62",
         15051 => x"69",
         15052 => x"2e",
         15053 => x"00",
         15054 => x"74",
         15055 => x"69",
         15056 => x"61",
         15057 => x"69",
         15058 => x"69",
         15059 => x"2e",
         15060 => x"00",
         15061 => x"6c",
         15062 => x"20",
         15063 => x"65",
         15064 => x"25",
         15065 => x"78",
         15066 => x"2e",
         15067 => x"00",
         15068 => x"6c",
         15069 => x"74",
         15070 => x"65",
         15071 => x"6f",
         15072 => x"28",
         15073 => x"2e",
         15074 => x"00",
         15075 => x"63",
         15076 => x"6e",
         15077 => x"6f",
         15078 => x"40",
         15079 => x"38",
         15080 => x"2e",
         15081 => x"00",
         15082 => x"6c",
         15083 => x"30",
         15084 => x"2d",
         15085 => x"00",
         15086 => x"6c",
         15087 => x"30",
         15088 => x"00",
         15089 => x"70",
         15090 => x"6e",
         15091 => x"2e",
         15092 => x"00",
         15093 => x"6c",
         15094 => x"30",
         15095 => x"2d",
         15096 => x"38",
         15097 => x"25",
         15098 => x"29",
         15099 => x"00",
         15100 => x"79",
         15101 => x"2e",
         15102 => x"00",
         15103 => x"6c",
         15104 => x"30",
         15105 => x"00",
         15106 => x"61",
         15107 => x"67",
         15108 => x"2e",
         15109 => x"00",
         15110 => x"70",
         15111 => x"6d",
         15112 => x"00",
         15113 => x"6d",
         15114 => x"74",
         15115 => x"00",
         15116 => x"5c",
         15117 => x"25",
         15118 => x"00",
         15119 => x"6f",
         15120 => x"65",
         15121 => x"75",
         15122 => x"64",
         15123 => x"61",
         15124 => x"74",
         15125 => x"6f",
         15126 => x"73",
         15127 => x"6d",
         15128 => x"64",
         15129 => x"00",
         15130 => x"00",
         15131 => x"25",
         15132 => x"64",
         15133 => x"3a",
         15134 => x"25",
         15135 => x"64",
         15136 => x"00",
         15137 => x"20",
         15138 => x"66",
         15139 => x"72",
         15140 => x"6f",
         15141 => x"00",
         15142 => x"65",
         15143 => x"65",
         15144 => x"6d",
         15145 => x"6d",
         15146 => x"65",
         15147 => x"00",
         15148 => x"72",
         15149 => x"65",
         15150 => x"00",
         15151 => x"20",
         15152 => x"20",
         15153 => x"65",
         15154 => x"65",
         15155 => x"72",
         15156 => x"64",
         15157 => x"73",
         15158 => x"25",
         15159 => x"0a",
         15160 => x"00",
         15161 => x"20",
         15162 => x"20",
         15163 => x"6f",
         15164 => x"53",
         15165 => x"74",
         15166 => x"64",
         15167 => x"73",
         15168 => x"25",
         15169 => x"0a",
         15170 => x"00",
         15171 => x"20",
         15172 => x"63",
         15173 => x"74",
         15174 => x"20",
         15175 => x"72",
         15176 => x"20",
         15177 => x"20",
         15178 => x"25",
         15179 => x"0a",
         15180 => x"00",
         15181 => x"63",
         15182 => x"00",
         15183 => x"20",
         15184 => x"20",
         15185 => x"20",
         15186 => x"20",
         15187 => x"20",
         15188 => x"20",
         15189 => x"20",
         15190 => x"25",
         15191 => x"0a",
         15192 => x"00",
         15193 => x"20",
         15194 => x"74",
         15195 => x"43",
         15196 => x"6b",
         15197 => x"65",
         15198 => x"20",
         15199 => x"20",
         15200 => x"25",
         15201 => x"30",
         15202 => x"48",
         15203 => x"00",
         15204 => x"20",
         15205 => x"68",
         15206 => x"65",
         15207 => x"52",
         15208 => x"43",
         15209 => x"6b",
         15210 => x"65",
         15211 => x"25",
         15212 => x"30",
         15213 => x"48",
         15214 => x"00",
         15215 => x"20",
         15216 => x"41",
         15217 => x"6c",
         15218 => x"20",
         15219 => x"71",
         15220 => x"20",
         15221 => x"20",
         15222 => x"25",
         15223 => x"30",
         15224 => x"48",
         15225 => x"00",
         15226 => x"20",
         15227 => x"00",
         15228 => x"20",
         15229 => x"00",
         15230 => x"20",
         15231 => x"54",
         15232 => x"00",
         15233 => x"20",
         15234 => x"49",
         15235 => x"00",
         15236 => x"20",
         15237 => x"48",
         15238 => x"45",
         15239 => x"53",
         15240 => x"00",
         15241 => x"20",
         15242 => x"52",
         15243 => x"52",
         15244 => x"43",
         15245 => x"6e",
         15246 => x"3d",
         15247 => x"64",
         15248 => x"00",
         15249 => x"20",
         15250 => x"45",
         15251 => x"20",
         15252 => x"54",
         15253 => x"72",
         15254 => x"3d",
         15255 => x"64",
         15256 => x"00",
         15257 => x"20",
         15258 => x"43",
         15259 => x"20",
         15260 => x"44",
         15261 => x"63",
         15262 => x"3d",
         15263 => x"64",
         15264 => x"00",
         15265 => x"20",
         15266 => x"20",
         15267 => x"20",
         15268 => x"25",
         15269 => x"3a",
         15270 => x"58",
         15271 => x"00",
         15272 => x"20",
         15273 => x"4d",
         15274 => x"20",
         15275 => x"25",
         15276 => x"3a",
         15277 => x"58",
         15278 => x"00",
         15279 => x"20",
         15280 => x"4e",
         15281 => x"41",
         15282 => x"25",
         15283 => x"3a",
         15284 => x"58",
         15285 => x"00",
         15286 => x"20",
         15287 => x"41",
         15288 => x"20",
         15289 => x"25",
         15290 => x"3a",
         15291 => x"58",
         15292 => x"00",
         15293 => x"20",
         15294 => x"53",
         15295 => x"4d",
         15296 => x"25",
         15297 => x"3a",
         15298 => x"58",
         15299 => x"00",
         15300 => x"72",
         15301 => x"53",
         15302 => x"63",
         15303 => x"69",
         15304 => x"00",
         15305 => x"6e",
         15306 => x"00",
         15307 => x"6d",
         15308 => x"00",
         15309 => x"6c",
         15310 => x"00",
         15311 => x"69",
         15312 => x"00",
         15313 => x"78",
         15314 => x"00",
         15315 => x"00",
         15316 => x"ac",
         15317 => x"00",
         15318 => x"02",
         15319 => x"a8",
         15320 => x"00",
         15321 => x"03",
         15322 => x"a4",
         15323 => x"00",
         15324 => x"04",
         15325 => x"a0",
         15326 => x"00",
         15327 => x"05",
         15328 => x"9c",
         15329 => x"00",
         15330 => x"06",
         15331 => x"98",
         15332 => x"00",
         15333 => x"07",
         15334 => x"94",
         15335 => x"00",
         15336 => x"01",
         15337 => x"90",
         15338 => x"00",
         15339 => x"08",
         15340 => x"8c",
         15341 => x"00",
         15342 => x"0b",
         15343 => x"88",
         15344 => x"00",
         15345 => x"09",
         15346 => x"84",
         15347 => x"00",
         15348 => x"0a",
         15349 => x"80",
         15350 => x"00",
         15351 => x"0d",
         15352 => x"7c",
         15353 => x"00",
         15354 => x"0c",
         15355 => x"78",
         15356 => x"00",
         15357 => x"0e",
         15358 => x"74",
         15359 => x"00",
         15360 => x"0f",
         15361 => x"70",
         15362 => x"00",
         15363 => x"0f",
         15364 => x"6c",
         15365 => x"00",
         15366 => x"10",
         15367 => x"68",
         15368 => x"00",
         15369 => x"11",
         15370 => x"64",
         15371 => x"00",
         15372 => x"12",
         15373 => x"60",
         15374 => x"00",
         15375 => x"13",
         15376 => x"5c",
         15377 => x"00",
         15378 => x"14",
         15379 => x"58",
         15380 => x"00",
         15381 => x"15",
         15382 => x"00",
         15383 => x"00",
         15384 => x"00",
         15385 => x"00",
         15386 => x"7e",
         15387 => x"7e",
         15388 => x"7e",
         15389 => x"00",
         15390 => x"7e",
         15391 => x"7e",
         15392 => x"7e",
         15393 => x"00",
         15394 => x"00",
         15395 => x"00",
         15396 => x"00",
         15397 => x"00",
         15398 => x"00",
         15399 => x"00",
         15400 => x"00",
         15401 => x"00",
         15402 => x"00",
         15403 => x"00",
         15404 => x"6e",
         15405 => x"6f",
         15406 => x"2f",
         15407 => x"61",
         15408 => x"68",
         15409 => x"6f",
         15410 => x"66",
         15411 => x"2c",
         15412 => x"73",
         15413 => x"69",
         15414 => x"00",
         15415 => x"74",
         15416 => x"00",
         15417 => x"74",
         15418 => x"00",
         15419 => x"00",
         15420 => x"6c",
         15421 => x"25",
         15422 => x"00",
         15423 => x"6c",
         15424 => x"74",
         15425 => x"65",
         15426 => x"20",
         15427 => x"20",
         15428 => x"74",
         15429 => x"20",
         15430 => x"65",
         15431 => x"20",
         15432 => x"2e",
         15433 => x"00",
         15434 => x"0a",
         15435 => x"00",
         15436 => x"7e",
         15437 => x"00",
         15438 => x"00",
         15439 => x"00",
         15440 => x"00",
         15441 => x"00",
         15442 => x"30",
         15443 => x"00",
         15444 => x"31",
         15445 => x"00",
         15446 => x"32",
         15447 => x"00",
         15448 => x"33",
         15449 => x"00",
         15450 => x"34",
         15451 => x"00",
         15452 => x"35",
         15453 => x"00",
         15454 => x"37",
         15455 => x"00",
         15456 => x"38",
         15457 => x"00",
         15458 => x"39",
         15459 => x"00",
         15460 => x"30",
         15461 => x"00",
         15462 => x"7e",
         15463 => x"00",
         15464 => x"7e",
         15465 => x"00",
         15466 => x"00",
         15467 => x"7e",
         15468 => x"00",
         15469 => x"7e",
         15470 => x"00",
         15471 => x"64",
         15472 => x"2c",
         15473 => x"25",
         15474 => x"64",
         15475 => x"3a",
         15476 => x"78",
         15477 => x"00",
         15478 => x"64",
         15479 => x"2d",
         15480 => x"25",
         15481 => x"64",
         15482 => x"2c",
         15483 => x"00",
         15484 => x"00",
         15485 => x"64",
         15486 => x"00",
         15487 => x"78",
         15488 => x"00",
         15489 => x"25",
         15490 => x"64",
         15491 => x"00",
         15492 => x"6f",
         15493 => x"43",
         15494 => x"6f",
         15495 => x"00",
         15496 => x"25",
         15497 => x"20",
         15498 => x"78",
         15499 => x"00",
         15500 => x"25",
         15501 => x"20",
         15502 => x"78",
         15503 => x"00",
         15504 => x"25",
         15505 => x"20",
         15506 => x"00",
         15507 => x"74",
         15508 => x"20",
         15509 => x"69",
         15510 => x"2e",
         15511 => x"00",
         15512 => x"00",
         15513 => x"3c",
         15514 => x"7f",
         15515 => x"00",
         15516 => x"3d",
         15517 => x"00",
         15518 => x"00",
         15519 => x"33",
         15520 => x"00",
         15521 => x"4d",
         15522 => x"53",
         15523 => x"00",
         15524 => x"4e",
         15525 => x"20",
         15526 => x"46",
         15527 => x"20",
         15528 => x"00",
         15529 => x"4e",
         15530 => x"20",
         15531 => x"46",
         15532 => x"32",
         15533 => x"00",
         15534 => x"60",
         15535 => x"00",
         15536 => x"00",
         15537 => x"00",
         15538 => x"07",
         15539 => x"12",
         15540 => x"1c",
         15541 => x"00",
         15542 => x"41",
         15543 => x"80",
         15544 => x"49",
         15545 => x"8f",
         15546 => x"4f",
         15547 => x"55",
         15548 => x"9b",
         15549 => x"9f",
         15550 => x"55",
         15551 => x"a7",
         15552 => x"ab",
         15553 => x"af",
         15554 => x"b3",
         15555 => x"b7",
         15556 => x"bb",
         15557 => x"bf",
         15558 => x"c3",
         15559 => x"c7",
         15560 => x"cb",
         15561 => x"cf",
         15562 => x"d3",
         15563 => x"d7",
         15564 => x"db",
         15565 => x"df",
         15566 => x"e3",
         15567 => x"e7",
         15568 => x"eb",
         15569 => x"ef",
         15570 => x"f3",
         15571 => x"f7",
         15572 => x"fb",
         15573 => x"ff",
         15574 => x"3b",
         15575 => x"2f",
         15576 => x"3a",
         15577 => x"7c",
         15578 => x"00",
         15579 => x"04",
         15580 => x"40",
         15581 => x"00",
         15582 => x"00",
         15583 => x"02",
         15584 => x"08",
         15585 => x"20",
         15586 => x"00",
         15587 => x"fc",
         15588 => x"e2",
         15589 => x"e0",
         15590 => x"e7",
         15591 => x"eb",
         15592 => x"ef",
         15593 => x"ec",
         15594 => x"c5",
         15595 => x"e6",
         15596 => x"f4",
         15597 => x"f2",
         15598 => x"f9",
         15599 => x"d6",
         15600 => x"a2",
         15601 => x"a5",
         15602 => x"92",
         15603 => x"ed",
         15604 => x"fa",
         15605 => x"d1",
         15606 => x"ba",
         15607 => x"10",
         15608 => x"bd",
         15609 => x"a1",
         15610 => x"bb",
         15611 => x"92",
         15612 => x"02",
         15613 => x"61",
         15614 => x"56",
         15615 => x"63",
         15616 => x"57",
         15617 => x"5c",
         15618 => x"10",
         15619 => x"34",
         15620 => x"1c",
         15621 => x"3c",
         15622 => x"5f",
         15623 => x"54",
         15624 => x"66",
         15625 => x"50",
         15626 => x"67",
         15627 => x"64",
         15628 => x"59",
         15629 => x"52",
         15630 => x"6b",
         15631 => x"18",
         15632 => x"88",
         15633 => x"8c",
         15634 => x"80",
         15635 => x"df",
         15636 => x"c0",
         15637 => x"c3",
         15638 => x"c4",
         15639 => x"98",
         15640 => x"b4",
         15641 => x"c6",
         15642 => x"29",
         15643 => x"b1",
         15644 => x"64",
         15645 => x"21",
         15646 => x"48",
         15647 => x"19",
         15648 => x"1a",
         15649 => x"b2",
         15650 => x"a0",
         15651 => x"1a",
         15652 => x"17",
         15653 => x"07",
         15654 => x"01",
         15655 => x"00",
         15656 => x"32",
         15657 => x"39",
         15658 => x"4a",
         15659 => x"79",
         15660 => x"80",
         15661 => x"43",
         15662 => x"82",
         15663 => x"84",
         15664 => x"86",
         15665 => x"87",
         15666 => x"8a",
         15667 => x"8b",
         15668 => x"8e",
         15669 => x"90",
         15670 => x"91",
         15671 => x"94",
         15672 => x"96",
         15673 => x"98",
         15674 => x"3d",
         15675 => x"9c",
         15676 => x"20",
         15677 => x"a0",
         15678 => x"a2",
         15679 => x"a4",
         15680 => x"a6",
         15681 => x"a7",
         15682 => x"aa",
         15683 => x"ac",
         15684 => x"ae",
         15685 => x"af",
         15686 => x"b2",
         15687 => x"b3",
         15688 => x"b5",
         15689 => x"b8",
         15690 => x"ba",
         15691 => x"bc",
         15692 => x"be",
         15693 => x"c0",
         15694 => x"c2",
         15695 => x"c4",
         15696 => x"c4",
         15697 => x"c8",
         15698 => x"ca",
         15699 => x"ca",
         15700 => x"10",
         15701 => x"01",
         15702 => x"de",
         15703 => x"f3",
         15704 => x"f1",
         15705 => x"f4",
         15706 => x"28",
         15707 => x"12",
         15708 => x"09",
         15709 => x"3b",
         15710 => x"3d",
         15711 => x"3f",
         15712 => x"41",
         15713 => x"46",
         15714 => x"53",
         15715 => x"81",
         15716 => x"55",
         15717 => x"8a",
         15718 => x"8f",
         15719 => x"90",
         15720 => x"5d",
         15721 => x"5f",
         15722 => x"61",
         15723 => x"94",
         15724 => x"65",
         15725 => x"67",
         15726 => x"96",
         15727 => x"62",
         15728 => x"6d",
         15729 => x"9c",
         15730 => x"71",
         15731 => x"73",
         15732 => x"9f",
         15733 => x"77",
         15734 => x"79",
         15735 => x"7b",
         15736 => x"64",
         15737 => x"7f",
         15738 => x"81",
         15739 => x"a9",
         15740 => x"85",
         15741 => x"87",
         15742 => x"44",
         15743 => x"b2",
         15744 => x"8d",
         15745 => x"8f",
         15746 => x"91",
         15747 => x"7b",
         15748 => x"fd",
         15749 => x"ff",
         15750 => x"04",
         15751 => x"88",
         15752 => x"8a",
         15753 => x"11",
         15754 => x"02",
         15755 => x"a3",
         15756 => x"08",
         15757 => x"03",
         15758 => x"8e",
         15759 => x"d8",
         15760 => x"f2",
         15761 => x"f9",
         15762 => x"f4",
         15763 => x"f6",
         15764 => x"f7",
         15765 => x"fa",
         15766 => x"30",
         15767 => x"50",
         15768 => x"60",
         15769 => x"8a",
         15770 => x"c1",
         15771 => x"cf",
         15772 => x"c0",
         15773 => x"44",
         15774 => x"26",
         15775 => x"00",
         15776 => x"01",
         15777 => x"00",
         15778 => x"a0",
         15779 => x"00",
         15780 => x"10",
         15781 => x"20",
         15782 => x"30",
         15783 => x"40",
         15784 => x"51",
         15785 => x"59",
         15786 => x"5b",
         15787 => x"5d",
         15788 => x"5f",
         15789 => x"08",
         15790 => x"0e",
         15791 => x"bb",
         15792 => x"c9",
         15793 => x"cb",
         15794 => x"db",
         15795 => x"f9",
         15796 => x"eb",
         15797 => x"fb",
         15798 => x"08",
         15799 => x"08",
         15800 => x"08",
         15801 => x"04",
         15802 => x"b9",
         15803 => x"bc",
         15804 => x"01",
         15805 => x"d0",
         15806 => x"e0",
         15807 => x"e5",
         15808 => x"ec",
         15809 => x"01",
         15810 => x"4e",
         15811 => x"32",
         15812 => x"10",
         15813 => x"01",
         15814 => x"d0",
         15815 => x"30",
         15816 => x"60",
         15817 => x"67",
         15818 => x"75",
         15819 => x"80",
         15820 => x"00",
         15821 => x"41",
         15822 => x"00",
         15823 => x"00",
         15824 => x"68",
         15825 => x"00",
         15826 => x"00",
         15827 => x"00",
         15828 => x"70",
         15829 => x"00",
         15830 => x"00",
         15831 => x"00",
         15832 => x"78",
         15833 => x"00",
         15834 => x"00",
         15835 => x"00",
         15836 => x"80",
         15837 => x"00",
         15838 => x"00",
         15839 => x"00",
         15840 => x"88",
         15841 => x"00",
         15842 => x"00",
         15843 => x"00",
         15844 => x"90",
         15845 => x"00",
         15846 => x"00",
         15847 => x"00",
         15848 => x"98",
         15849 => x"00",
         15850 => x"00",
         15851 => x"00",
         15852 => x"a0",
         15853 => x"00",
         15854 => x"00",
         15855 => x"00",
         15856 => x"a8",
         15857 => x"00",
         15858 => x"00",
         15859 => x"00",
         15860 => x"b0",
         15861 => x"00",
         15862 => x"00",
         15863 => x"00",
         15864 => x"b4",
         15865 => x"00",
         15866 => x"00",
         15867 => x"00",
         15868 => x"b8",
         15869 => x"00",
         15870 => x"00",
         15871 => x"00",
         15872 => x"bc",
         15873 => x"00",
         15874 => x"00",
         15875 => x"00",
         15876 => x"c0",
         15877 => x"00",
         15878 => x"00",
         15879 => x"00",
         15880 => x"c4",
         15881 => x"00",
         15882 => x"00",
         15883 => x"00",
         15884 => x"c8",
         15885 => x"00",
         15886 => x"00",
         15887 => x"00",
         15888 => x"cc",
         15889 => x"00",
         15890 => x"00",
         15891 => x"00",
         15892 => x"d4",
         15893 => x"00",
         15894 => x"00",
         15895 => x"00",
         15896 => x"d8",
         15897 => x"00",
         15898 => x"00",
         15899 => x"00",
         15900 => x"e0",
         15901 => x"00",
         15902 => x"00",
         15903 => x"00",
         15904 => x"e8",
         15905 => x"00",
         15906 => x"00",
         15907 => x"00",
         15908 => x"f0",
         15909 => x"00",
         15910 => x"00",
         15911 => x"00",
         15912 => x"f8",
         15913 => x"00",
         15914 => x"00",
         15915 => x"00",
         15916 => x"fc",
         15917 => x"00",
         15918 => x"00",
         15919 => x"00",
         15920 => x"00",
         15921 => x"00",
         15922 => x"00",
         15923 => x"00",
         15924 => x"08",
         15925 => x"00",
         15926 => x"00",
         15927 => x"00",
         15928 => x"10",
         15929 => x"00",
         15930 => x"00",
         15931 => x"00",
         15932 => x"18",
         15933 => x"00",
         15934 => x"00",
         15935 => x"00",
         15936 => x"00",
         15937 => x"00",
         15938 => x"ff",
         15939 => x"00",
         15940 => x"ff",
         15941 => x"00",
         15942 => x"ff",
         15943 => x"00",
         15944 => x"00",
         15945 => x"00",
         15946 => x"ff",
         15947 => x"00",
         15948 => x"00",
         15949 => x"00",
         15950 => x"00",
         15951 => x"00",
         15952 => x"00",
         15953 => x"00",
         15954 => x"00",
         15955 => x"01",
         15956 => x"01",
         15957 => x"01",
         15958 => x"00",
         15959 => x"00",
         15960 => x"00",
         15961 => x"00",
         15962 => x"00",
         15963 => x"00",
         15964 => x"00",
         15965 => x"00",
         15966 => x"00",
         15967 => x"00",
         15968 => x"00",
         15969 => x"00",
         15970 => x"00",
         15971 => x"00",
         15972 => x"00",
         15973 => x"00",
         15974 => x"00",
         15975 => x"00",
         15976 => x"00",
         15977 => x"00",
         15978 => x"00",
         15979 => x"00",
         15980 => x"00",
         15981 => x"00",
         15982 => x"00",
         15983 => x"dc",
         15984 => x"00",
         15985 => x"e4",
         15986 => x"00",
         15987 => x"ec",
         15988 => x"00",
         15989 => x"80",
         15990 => x"fd",
         15991 => x"0d",
         15992 => x"5b",
         15993 => x"f0",
         15994 => x"74",
         15995 => x"78",
         15996 => x"6c",
         15997 => x"70",
         15998 => x"64",
         15999 => x"68",
         16000 => x"34",
         16001 => x"38",
         16002 => x"20",
         16003 => x"2e",
         16004 => x"f4",
         16005 => x"2f",
         16006 => x"f0",
         16007 => x"f0",
         16008 => x"83",
         16009 => x"f0",
         16010 => x"fd",
         16011 => x"0d",
         16012 => x"5b",
         16013 => x"f0",
         16014 => x"54",
         16015 => x"58",
         16016 => x"4c",
         16017 => x"50",
         16018 => x"44",
         16019 => x"48",
         16020 => x"34",
         16021 => x"38",
         16022 => x"20",
         16023 => x"2e",
         16024 => x"f4",
         16025 => x"2f",
         16026 => x"f0",
         16027 => x"f0",
         16028 => x"83",
         16029 => x"f0",
         16030 => x"fd",
         16031 => x"0d",
         16032 => x"7b",
         16033 => x"f0",
         16034 => x"54",
         16035 => x"58",
         16036 => x"4c",
         16037 => x"50",
         16038 => x"44",
         16039 => x"48",
         16040 => x"24",
         16041 => x"28",
         16042 => x"20",
         16043 => x"3e",
         16044 => x"e1",
         16045 => x"2f",
         16046 => x"f0",
         16047 => x"f0",
         16048 => x"88",
         16049 => x"f0",
         16050 => x"fa",
         16051 => x"f0",
         16052 => x"1b",
         16053 => x"f0",
         16054 => x"14",
         16055 => x"18",
         16056 => x"0c",
         16057 => x"10",
         16058 => x"04",
         16059 => x"08",
         16060 => x"f0",
         16061 => x"f0",
         16062 => x"f0",
         16063 => x"f0",
         16064 => x"f0",
         16065 => x"1c",
         16066 => x"f0",
         16067 => x"f0",
         16068 => x"83",
         16069 => x"f0",
         16070 => x"c9",
         16071 => x"cd",
         16072 => x"b3",
         16073 => x"f0",
         16074 => x"31",
         16075 => x"dd",
         16076 => x"56",
         16077 => x"b1",
         16078 => x"48",
         16079 => x"73",
         16080 => x"3b",
         16081 => x"a2",
         16082 => x"00",
         16083 => x"b9",
         16084 => x"c1",
         16085 => x"be",
         16086 => x"f0",
         16087 => x"f0",
         16088 => x"83",
         16089 => x"f0",
         16090 => x"00",
         16091 => x"00",
         16092 => x"00",
         16093 => x"00",
         16094 => x"00",
         16095 => x"00",
         16096 => x"00",
         16097 => x"00",
         16098 => x"00",
         16099 => x"00",
         16100 => x"00",
         16101 => x"00",
         16102 => x"00",
         16103 => x"00",
         16104 => x"00",
         16105 => x"00",
         16106 => x"00",
         16107 => x"00",
         16108 => x"00",
         16109 => x"00",
         16110 => x"00",
         16111 => x"00",
         16112 => x"00",
         16113 => x"00",
         16114 => x"00",
         16115 => x"00",
         16116 => x"00",
         16117 => x"00",
         16118 => x"30",
         16119 => x"00",
         16120 => x"38",
         16121 => x"00",
         16122 => x"3c",
         16123 => x"00",
         16124 => x"40",
         16125 => x"00",
         16126 => x"44",
         16127 => x"00",
         16128 => x"48",
         16129 => x"00",
         16130 => x"50",
         16131 => x"00",
         16132 => x"58",
         16133 => x"00",
         16134 => x"60",
         16135 => x"00",
         16136 => x"68",
         16137 => x"00",
         16138 => x"70",
         16139 => x"00",
         16140 => x"78",
         16141 => x"00",
         16142 => x"80",
         16143 => x"00",
         16144 => x"88",
         16145 => x"00",
         16146 => x"90",
         16147 => x"00",
         16148 => x"98",
         16149 => x"00",
         16150 => x"a0",
         16151 => x"00",
         16152 => x"a8",
         16153 => x"00",
         16154 => x"ac",
         16155 => x"00",
         16156 => x"b4",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"00",
         16166 => x"00",
         16167 => x"00",
         16168 => x"00",
         16169 => x"00",
         16170 => x"00",
         16171 => x"00",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"19",
         18159 => x"00",
         18160 => x"00",
         18161 => x"f3",
         18162 => x"f7",
         18163 => x"fb",
         18164 => x"ff",
         18165 => x"c3",
         18166 => x"e2",
         18167 => x"e6",
         18168 => x"f4",
         18169 => x"63",
         18170 => x"67",
         18171 => x"6a",
         18172 => x"2d",
         18173 => x"23",
         18174 => x"27",
         18175 => x"2c",
         18176 => x"49",
         18177 => x"03",
         18178 => x"07",
         18179 => x"0b",
         18180 => x"0f",
         18181 => x"13",
         18182 => x"17",
         18183 => x"52",
         18184 => x"3c",
         18185 => x"83",
         18186 => x"87",
         18187 => x"8b",
         18188 => x"8f",
         18189 => x"93",
         18190 => x"97",
         18191 => x"bc",
         18192 => x"c0",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"00",
         18199 => x"00",
         18200 => x"00",
         18201 => x"00",
         18202 => x"00",
         18203 => x"00",
         18204 => x"00",
         18205 => x"00",
         18206 => x"00",
         18207 => x"00",
         18208 => x"00",
         18209 => x"00",
         18210 => x"00",
         18211 => x"00",
         18212 => x"00",
         18213 => x"00",
         18214 => x"00",
         18215 => x"00",
         18216 => x"00",
         18217 => x"00",
         18218 => x"00",
         18219 => x"00",
         18220 => x"00",
         18221 => x"00",
         18222 => x"00",
         18223 => x"03",
         18224 => x"01",
         18225 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"0b",
             2 => x"e9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"83",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a6",
           270 => x"0b",
           271 => x"0b",
           272 => x"c6",
           273 => x"0b",
           274 => x"0b",
           275 => x"e6",
           276 => x"0b",
           277 => x"0b",
           278 => x"86",
           279 => x"0b",
           280 => x"0b",
           281 => x"a6",
           282 => x"0b",
           283 => x"0b",
           284 => x"c6",
           285 => x"0b",
           286 => x"0b",
           287 => x"e8",
           288 => x"0b",
           289 => x"0b",
           290 => x"8a",
           291 => x"0b",
           292 => x"0b",
           293 => x"ac",
           294 => x"0b",
           295 => x"0b",
           296 => x"ce",
           297 => x"0b",
           298 => x"0b",
           299 => x"f0",
           300 => x"0b",
           301 => x"0b",
           302 => x"92",
           303 => x"0b",
           304 => x"0b",
           305 => x"b4",
           306 => x"0b",
           307 => x"0b",
           308 => x"d6",
           309 => x"0b",
           310 => x"0b",
           311 => x"f8",
           312 => x"0b",
           313 => x"0b",
           314 => x"9a",
           315 => x"0b",
           316 => x"0b",
           317 => x"bc",
           318 => x"0b",
           319 => x"0b",
           320 => x"de",
           321 => x"0b",
           322 => x"0b",
           323 => x"80",
           324 => x"0b",
           325 => x"0b",
           326 => x"a2",
           327 => x"0b",
           328 => x"0b",
           329 => x"c4",
           330 => x"0b",
           331 => x"0b",
           332 => x"e6",
           333 => x"0b",
           334 => x"0b",
           335 => x"88",
           336 => x"0b",
           337 => x"0b",
           338 => x"aa",
           339 => x"0b",
           340 => x"0b",
           341 => x"cb",
           342 => x"0b",
           343 => x"0b",
           344 => x"ed",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"b9",
           386 => x"d6",
           387 => x"b9",
           388 => x"c0",
           389 => x"84",
           390 => x"a2",
           391 => x"b9",
           392 => x"c0",
           393 => x"84",
           394 => x"a0",
           395 => x"b9",
           396 => x"c0",
           397 => x"84",
           398 => x"a0",
           399 => x"b9",
           400 => x"c0",
           401 => x"84",
           402 => x"94",
           403 => x"b9",
           404 => x"c0",
           405 => x"84",
           406 => x"a1",
           407 => x"b9",
           408 => x"c0",
           409 => x"84",
           410 => x"af",
           411 => x"b9",
           412 => x"c0",
           413 => x"84",
           414 => x"ad",
           415 => x"b9",
           416 => x"c0",
           417 => x"84",
           418 => x"94",
           419 => x"b9",
           420 => x"c0",
           421 => x"84",
           422 => x"95",
           423 => x"b9",
           424 => x"c0",
           425 => x"84",
           426 => x"95",
           427 => x"b9",
           428 => x"c0",
           429 => x"84",
           430 => x"b1",
           431 => x"b9",
           432 => x"c0",
           433 => x"84",
           434 => x"80",
           435 => x"84",
           436 => x"80",
           437 => x"04",
           438 => x"0c",
           439 => x"2d",
           440 => x"08",
           441 => x"90",
           442 => x"d4",
           443 => x"a8",
           444 => x"d4",
           445 => x"80",
           446 => x"b9",
           447 => x"d3",
           448 => x"b9",
           449 => x"c0",
           450 => x"84",
           451 => x"82",
           452 => x"84",
           453 => x"80",
           454 => x"04",
           455 => x"0c",
           456 => x"2d",
           457 => x"08",
           458 => x"90",
           459 => x"d4",
           460 => x"9e",
           461 => x"d4",
           462 => x"80",
           463 => x"b9",
           464 => x"d7",
           465 => x"b9",
           466 => x"c0",
           467 => x"84",
           468 => x"82",
           469 => x"84",
           470 => x"80",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"90",
           476 => x"d4",
           477 => x"87",
           478 => x"d4",
           479 => x"80",
           480 => x"b9",
           481 => x"f1",
           482 => x"b9",
           483 => x"c0",
           484 => x"84",
           485 => x"82",
           486 => x"84",
           487 => x"80",
           488 => x"04",
           489 => x"0c",
           490 => x"2d",
           491 => x"08",
           492 => x"90",
           493 => x"d4",
           494 => x"a2",
           495 => x"d4",
           496 => x"80",
           497 => x"b9",
           498 => x"fe",
           499 => x"b9",
           500 => x"c0",
           501 => x"84",
           502 => x"83",
           503 => x"84",
           504 => x"80",
           505 => x"04",
           506 => x"0c",
           507 => x"2d",
           508 => x"08",
           509 => x"90",
           510 => x"d4",
           511 => x"fd",
           512 => x"d4",
           513 => x"80",
           514 => x"b9",
           515 => x"95",
           516 => x"b9",
           517 => x"c0",
           518 => x"84",
           519 => x"82",
           520 => x"84",
           521 => x"80",
           522 => x"04",
           523 => x"0c",
           524 => x"2d",
           525 => x"08",
           526 => x"90",
           527 => x"d4",
           528 => x"8e",
           529 => x"d4",
           530 => x"80",
           531 => x"b9",
           532 => x"f6",
           533 => x"b9",
           534 => x"c0",
           535 => x"84",
           536 => x"83",
           537 => x"84",
           538 => x"80",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"90",
           544 => x"d4",
           545 => x"e9",
           546 => x"d4",
           547 => x"80",
           548 => x"b9",
           549 => x"c6",
           550 => x"b9",
           551 => x"c0",
           552 => x"84",
           553 => x"83",
           554 => x"84",
           555 => x"80",
           556 => x"04",
           557 => x"0c",
           558 => x"2d",
           559 => x"08",
           560 => x"90",
           561 => x"d4",
           562 => x"c5",
           563 => x"d4",
           564 => x"80",
           565 => x"b9",
           566 => x"f3",
           567 => x"b9",
           568 => x"c0",
           569 => x"84",
           570 => x"81",
           571 => x"84",
           572 => x"80",
           573 => x"04",
           574 => x"0c",
           575 => x"2d",
           576 => x"08",
           577 => x"90",
           578 => x"d4",
           579 => x"aa",
           580 => x"d4",
           581 => x"80",
           582 => x"b9",
           583 => x"d1",
           584 => x"b9",
           585 => x"c0",
           586 => x"84",
           587 => x"80",
           588 => x"84",
           589 => x"80",
           590 => x"04",
           591 => x"0c",
           592 => x"84",
           593 => x"80",
           594 => x"04",
           595 => x"0c",
           596 => x"2d",
           597 => x"08",
           598 => x"90",
           599 => x"d4",
           600 => x"bc",
           601 => x"d4",
           602 => x"80",
           603 => x"b9",
           604 => x"f1",
           605 => x"b9",
           606 => x"c0",
           607 => x"84",
           608 => x"81",
           609 => x"84",
           610 => x"80",
           611 => x"04",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"04",
           621 => x"81",
           622 => x"83",
           623 => x"05",
           624 => x"10",
           625 => x"72",
           626 => x"51",
           627 => x"72",
           628 => x"06",
           629 => x"72",
           630 => x"10",
           631 => x"10",
           632 => x"ed",
           633 => x"53",
           634 => x"b9",
           635 => x"d5",
           636 => x"38",
           637 => x"84",
           638 => x"0b",
           639 => x"ec",
           640 => x"51",
           641 => x"04",
           642 => x"0d",
           643 => x"70",
           644 => x"08",
           645 => x"52",
           646 => x"08",
           647 => x"3f",
           648 => x"04",
           649 => x"78",
           650 => x"11",
           651 => x"81",
           652 => x"25",
           653 => x"55",
           654 => x"72",
           655 => x"81",
           656 => x"38",
           657 => x"74",
           658 => x"30",
           659 => x"9f",
           660 => x"55",
           661 => x"74",
           662 => x"71",
           663 => x"38",
           664 => x"fa",
           665 => x"c8",
           666 => x"b9",
           667 => x"2e",
           668 => x"b9",
           669 => x"70",
           670 => x"34",
           671 => x"8a",
           672 => x"70",
           673 => x"2a",
           674 => x"54",
           675 => x"cb",
           676 => x"34",
           677 => x"84",
           678 => x"88",
           679 => x"80",
           680 => x"c8",
           681 => x"0d",
           682 => x"0d",
           683 => x"02",
           684 => x"05",
           685 => x"fe",
           686 => x"3d",
           687 => x"7e",
           688 => x"e4",
           689 => x"3f",
           690 => x"80",
           691 => x"3d",
           692 => x"3d",
           693 => x"88",
           694 => x"52",
           695 => x"3f",
           696 => x"04",
           697 => x"61",
           698 => x"5d",
           699 => x"8c",
           700 => x"1e",
           701 => x"2a",
           702 => x"06",
           703 => x"ff",
           704 => x"2e",
           705 => x"80",
           706 => x"33",
           707 => x"2e",
           708 => x"81",
           709 => x"06",
           710 => x"80",
           711 => x"38",
           712 => x"7e",
           713 => x"a3",
           714 => x"32",
           715 => x"80",
           716 => x"55",
           717 => x"72",
           718 => x"38",
           719 => x"70",
           720 => x"06",
           721 => x"80",
           722 => x"7a",
           723 => x"5b",
           724 => x"76",
           725 => x"8c",
           726 => x"73",
           727 => x"0c",
           728 => x"04",
           729 => x"54",
           730 => x"10",
           731 => x"70",
           732 => x"98",
           733 => x"81",
           734 => x"8b",
           735 => x"98",
           736 => x"5b",
           737 => x"79",
           738 => x"38",
           739 => x"53",
           740 => x"38",
           741 => x"58",
           742 => x"f7",
           743 => x"39",
           744 => x"09",
           745 => x"38",
           746 => x"5a",
           747 => x"7c",
           748 => x"76",
           749 => x"ff",
           750 => x"52",
           751 => x"af",
           752 => x"57",
           753 => x"38",
           754 => x"7a",
           755 => x"81",
           756 => x"78",
           757 => x"70",
           758 => x"54",
           759 => x"e0",
           760 => x"80",
           761 => x"38",
           762 => x"83",
           763 => x"54",
           764 => x"73",
           765 => x"59",
           766 => x"27",
           767 => x"52",
           768 => x"eb",
           769 => x"33",
           770 => x"fe",
           771 => x"c7",
           772 => x"59",
           773 => x"88",
           774 => x"84",
           775 => x"7d",
           776 => x"06",
           777 => x"54",
           778 => x"5e",
           779 => x"51",
           780 => x"84",
           781 => x"81",
           782 => x"b9",
           783 => x"df",
           784 => x"72",
           785 => x"38",
           786 => x"08",
           787 => x"74",
           788 => x"05",
           789 => x"52",
           790 => x"ca",
           791 => x"c8",
           792 => x"b9",
           793 => x"38",
           794 => x"d8",
           795 => x"7b",
           796 => x"56",
           797 => x"8f",
           798 => x"80",
           799 => x"80",
           800 => x"90",
           801 => x"7a",
           802 => x"81",
           803 => x"73",
           804 => x"38",
           805 => x"80",
           806 => x"80",
           807 => x"90",
           808 => x"77",
           809 => x"29",
           810 => x"05",
           811 => x"2c",
           812 => x"2a",
           813 => x"54",
           814 => x"2e",
           815 => x"98",
           816 => x"ff",
           817 => x"78",
           818 => x"cc",
           819 => x"ff",
           820 => x"83",
           821 => x"2a",
           822 => x"74",
           823 => x"73",
           824 => x"f0",
           825 => x"31",
           826 => x"90",
           827 => x"80",
           828 => x"53",
           829 => x"85",
           830 => x"81",
           831 => x"54",
           832 => x"38",
           833 => x"81",
           834 => x"86",
           835 => x"85",
           836 => x"54",
           837 => x"38",
           838 => x"54",
           839 => x"38",
           840 => x"81",
           841 => x"80",
           842 => x"77",
           843 => x"80",
           844 => x"80",
           845 => x"2c",
           846 => x"80",
           847 => x"38",
           848 => x"51",
           849 => x"77",
           850 => x"80",
           851 => x"80",
           852 => x"2c",
           853 => x"73",
           854 => x"38",
           855 => x"53",
           856 => x"b2",
           857 => x"81",
           858 => x"81",
           859 => x"70",
           860 => x"55",
           861 => x"25",
           862 => x"52",
           863 => x"ef",
           864 => x"81",
           865 => x"81",
           866 => x"70",
           867 => x"55",
           868 => x"24",
           869 => x"87",
           870 => x"06",
           871 => x"80",
           872 => x"38",
           873 => x"2e",
           874 => x"76",
           875 => x"81",
           876 => x"80",
           877 => x"e2",
           878 => x"b9",
           879 => x"38",
           880 => x"1e",
           881 => x"5e",
           882 => x"7d",
           883 => x"2e",
           884 => x"ec",
           885 => x"06",
           886 => x"2e",
           887 => x"77",
           888 => x"80",
           889 => x"80",
           890 => x"2c",
           891 => x"80",
           892 => x"91",
           893 => x"a0",
           894 => x"3f",
           895 => x"90",
           896 => x"a0",
           897 => x"58",
           898 => x"87",
           899 => x"39",
           900 => x"07",
           901 => x"57",
           902 => x"84",
           903 => x"7e",
           904 => x"06",
           905 => x"55",
           906 => x"39",
           907 => x"05",
           908 => x"0a",
           909 => x"33",
           910 => x"72",
           911 => x"80",
           912 => x"80",
           913 => x"90",
           914 => x"5a",
           915 => x"5f",
           916 => x"70",
           917 => x"55",
           918 => x"38",
           919 => x"80",
           920 => x"80",
           921 => x"90",
           922 => x"5f",
           923 => x"fe",
           924 => x"52",
           925 => x"f7",
           926 => x"ff",
           927 => x"ff",
           928 => x"57",
           929 => x"ff",
           930 => x"38",
           931 => x"70",
           932 => x"33",
           933 => x"3f",
           934 => x"1a",
           935 => x"ff",
           936 => x"79",
           937 => x"2e",
           938 => x"7c",
           939 => x"81",
           940 => x"51",
           941 => x"e2",
           942 => x"0a",
           943 => x"0a",
           944 => x"80",
           945 => x"80",
           946 => x"90",
           947 => x"56",
           948 => x"87",
           949 => x"06",
           950 => x"7a",
           951 => x"fe",
           952 => x"60",
           953 => x"08",
           954 => x"41",
           955 => x"24",
           956 => x"7a",
           957 => x"06",
           958 => x"d8",
           959 => x"39",
           960 => x"7c",
           961 => x"76",
           962 => x"f8",
           963 => x"88",
           964 => x"7c",
           965 => x"76",
           966 => x"f8",
           967 => x"60",
           968 => x"08",
           969 => x"56",
           970 => x"72",
           971 => x"75",
           972 => x"3f",
           973 => x"08",
           974 => x"06",
           975 => x"90",
           976 => x"72",
           977 => x"fe",
           978 => x"80",
           979 => x"33",
           980 => x"f7",
           981 => x"ff",
           982 => x"84",
           983 => x"77",
           984 => x"58",
           985 => x"81",
           986 => x"51",
           987 => x"84",
           988 => x"83",
           989 => x"78",
           990 => x"2b",
           991 => x"39",
           992 => x"07",
           993 => x"5b",
           994 => x"38",
           995 => x"77",
           996 => x"80",
           997 => x"80",
           998 => x"2c",
           999 => x"80",
          1000 => x"d6",
          1001 => x"a0",
          1002 => x"3f",
          1003 => x"52",
          1004 => x"bb",
          1005 => x"2e",
          1006 => x"fa",
          1007 => x"52",
          1008 => x"ab",
          1009 => x"2a",
          1010 => x"7e",
          1011 => x"8c",
          1012 => x"39",
          1013 => x"78",
          1014 => x"2b",
          1015 => x"7d",
          1016 => x"57",
          1017 => x"73",
          1018 => x"ff",
          1019 => x"52",
          1020 => x"fb",
          1021 => x"06",
          1022 => x"2e",
          1023 => x"ff",
          1024 => x"52",
          1025 => x"51",
          1026 => x"74",
          1027 => x"7a",
          1028 => x"f1",
          1029 => x"39",
          1030 => x"98",
          1031 => x"2c",
          1032 => x"b7",
          1033 => x"ab",
          1034 => x"3f",
          1035 => x"52",
          1036 => x"bb",
          1037 => x"39",
          1038 => x"51",
          1039 => x"84",
          1040 => x"83",
          1041 => x"78",
          1042 => x"2b",
          1043 => x"f3",
          1044 => x"07",
          1045 => x"83",
          1046 => x"52",
          1047 => x"99",
          1048 => x"0d",
          1049 => x"08",
          1050 => x"74",
          1051 => x"3f",
          1052 => x"04",
          1053 => x"78",
          1054 => x"84",
          1055 => x"85",
          1056 => x"81",
          1057 => x"70",
          1058 => x"56",
          1059 => x"ff",
          1060 => x"2e",
          1061 => x"80",
          1062 => x"70",
          1063 => x"33",
          1064 => x"2e",
          1065 => x"d5",
          1066 => x"72",
          1067 => x"08",
          1068 => x"84",
          1069 => x"80",
          1070 => x"ff",
          1071 => x"81",
          1072 => x"53",
          1073 => x"88",
          1074 => x"ac",
          1075 => x"39",
          1076 => x"08",
          1077 => x"ac",
          1078 => x"51",
          1079 => x"55",
          1080 => x"b9",
          1081 => x"2e",
          1082 => x"57",
          1083 => x"84",
          1084 => x"88",
          1085 => x"fa",
          1086 => x"7a",
          1087 => x"0b",
          1088 => x"70",
          1089 => x"32",
          1090 => x"51",
          1091 => x"ff",
          1092 => x"2e",
          1093 => x"92",
          1094 => x"81",
          1095 => x"53",
          1096 => x"09",
          1097 => x"38",
          1098 => x"84",
          1099 => x"88",
          1100 => x"73",
          1101 => x"55",
          1102 => x"80",
          1103 => x"74",
          1104 => x"90",
          1105 => x"72",
          1106 => x"c8",
          1107 => x"e3",
          1108 => x"70",
          1109 => x"33",
          1110 => x"e3",
          1111 => x"ff",
          1112 => x"d5",
          1113 => x"73",
          1114 => x"83",
          1115 => x"fa",
          1116 => x"7a",
          1117 => x"70",
          1118 => x"32",
          1119 => x"56",
          1120 => x"56",
          1121 => x"73",
          1122 => x"06",
          1123 => x"2e",
          1124 => x"15",
          1125 => x"88",
          1126 => x"91",
          1127 => x"56",
          1128 => x"74",
          1129 => x"75",
          1130 => x"08",
          1131 => x"8c",
          1132 => x"56",
          1133 => x"c8",
          1134 => x"0d",
          1135 => x"76",
          1136 => x"51",
          1137 => x"54",
          1138 => x"56",
          1139 => x"08",
          1140 => x"15",
          1141 => x"8c",
          1142 => x"56",
          1143 => x"3d",
          1144 => x"11",
          1145 => x"ff",
          1146 => x"32",
          1147 => x"55",
          1148 => x"54",
          1149 => x"72",
          1150 => x"06",
          1151 => x"38",
          1152 => x"81",
          1153 => x"80",
          1154 => x"38",
          1155 => x"33",
          1156 => x"80",
          1157 => x"38",
          1158 => x"0c",
          1159 => x"81",
          1160 => x"0c",
          1161 => x"06",
          1162 => x"b9",
          1163 => x"3d",
          1164 => x"ff",
          1165 => x"72",
          1166 => x"8c",
          1167 => x"05",
          1168 => x"84",
          1169 => x"b9",
          1170 => x"3d",
          1171 => x"51",
          1172 => x"55",
          1173 => x"b9",
          1174 => x"84",
          1175 => x"80",
          1176 => x"38",
          1177 => x"70",
          1178 => x"52",
          1179 => x"08",
          1180 => x"38",
          1181 => x"53",
          1182 => x"34",
          1183 => x"84",
          1184 => x"87",
          1185 => x"74",
          1186 => x"72",
          1187 => x"ff",
          1188 => x"fd",
          1189 => x"77",
          1190 => x"54",
          1191 => x"05",
          1192 => x"70",
          1193 => x"12",
          1194 => x"81",
          1195 => x"51",
          1196 => x"81",
          1197 => x"70",
          1198 => x"84",
          1199 => x"85",
          1200 => x"fc",
          1201 => x"79",
          1202 => x"55",
          1203 => x"80",
          1204 => x"73",
          1205 => x"38",
          1206 => x"93",
          1207 => x"81",
          1208 => x"73",
          1209 => x"55",
          1210 => x"51",
          1211 => x"73",
          1212 => x"0c",
          1213 => x"04",
          1214 => x"73",
          1215 => x"38",
          1216 => x"53",
          1217 => x"ff",
          1218 => x"71",
          1219 => x"ff",
          1220 => x"80",
          1221 => x"ff",
          1222 => x"53",
          1223 => x"73",
          1224 => x"51",
          1225 => x"c7",
          1226 => x"0d",
          1227 => x"53",
          1228 => x"05",
          1229 => x"70",
          1230 => x"12",
          1231 => x"84",
          1232 => x"51",
          1233 => x"04",
          1234 => x"75",
          1235 => x"54",
          1236 => x"81",
          1237 => x"51",
          1238 => x"81",
          1239 => x"70",
          1240 => x"84",
          1241 => x"85",
          1242 => x"fd",
          1243 => x"78",
          1244 => x"55",
          1245 => x"80",
          1246 => x"71",
          1247 => x"53",
          1248 => x"81",
          1249 => x"ff",
          1250 => x"ef",
          1251 => x"b9",
          1252 => x"3d",
          1253 => x"3d",
          1254 => x"7a",
          1255 => x"72",
          1256 => x"38",
          1257 => x"70",
          1258 => x"33",
          1259 => x"71",
          1260 => x"06",
          1261 => x"14",
          1262 => x"2e",
          1263 => x"13",
          1264 => x"38",
          1265 => x"84",
          1266 => x"86",
          1267 => x"72",
          1268 => x"38",
          1269 => x"ff",
          1270 => x"2e",
          1271 => x"15",
          1272 => x"51",
          1273 => x"de",
          1274 => x"31",
          1275 => x"0c",
          1276 => x"04",
          1277 => x"c8",
          1278 => x"0d",
          1279 => x"0d",
          1280 => x"70",
          1281 => x"c1",
          1282 => x"c8",
          1283 => x"c8",
          1284 => x"52",
          1285 => x"ea",
          1286 => x"c8",
          1287 => x"b9",
          1288 => x"2e",
          1289 => x"b9",
          1290 => x"54",
          1291 => x"74",
          1292 => x"84",
          1293 => x"51",
          1294 => x"84",
          1295 => x"54",
          1296 => x"c8",
          1297 => x"0d",
          1298 => x"0d",
          1299 => x"71",
          1300 => x"54",
          1301 => x"9f",
          1302 => x"81",
          1303 => x"51",
          1304 => x"8c",
          1305 => x"52",
          1306 => x"09",
          1307 => x"38",
          1308 => x"75",
          1309 => x"70",
          1310 => x"0c",
          1311 => x"04",
          1312 => x"75",
          1313 => x"55",
          1314 => x"70",
          1315 => x"38",
          1316 => x"81",
          1317 => x"ff",
          1318 => x"f4",
          1319 => x"b9",
          1320 => x"3d",
          1321 => x"3d",
          1322 => x"58",
          1323 => x"76",
          1324 => x"38",
          1325 => x"f5",
          1326 => x"c8",
          1327 => x"12",
          1328 => x"2e",
          1329 => x"51",
          1330 => x"71",
          1331 => x"08",
          1332 => x"52",
          1333 => x"80",
          1334 => x"52",
          1335 => x"80",
          1336 => x"13",
          1337 => x"a0",
          1338 => x"71",
          1339 => x"54",
          1340 => x"74",
          1341 => x"38",
          1342 => x"9f",
          1343 => x"10",
          1344 => x"72",
          1345 => x"9f",
          1346 => x"06",
          1347 => x"75",
          1348 => x"1c",
          1349 => x"52",
          1350 => x"53",
          1351 => x"73",
          1352 => x"52",
          1353 => x"c8",
          1354 => x"0d",
          1355 => x"0d",
          1356 => x"80",
          1357 => x"30",
          1358 => x"80",
          1359 => x"2b",
          1360 => x"75",
          1361 => x"83",
          1362 => x"70",
          1363 => x"25",
          1364 => x"71",
          1365 => x"2a",
          1366 => x"06",
          1367 => x"80",
          1368 => x"84",
          1369 => x"71",
          1370 => x"75",
          1371 => x"8c",
          1372 => x"70",
          1373 => x"82",
          1374 => x"71",
          1375 => x"2a",
          1376 => x"81",
          1377 => x"82",
          1378 => x"75",
          1379 => x"b9",
          1380 => x"52",
          1381 => x"54",
          1382 => x"55",
          1383 => x"56",
          1384 => x"51",
          1385 => x"52",
          1386 => x"04",
          1387 => x"75",
          1388 => x"71",
          1389 => x"81",
          1390 => x"b9",
          1391 => x"29",
          1392 => x"84",
          1393 => x"53",
          1394 => x"04",
          1395 => x"78",
          1396 => x"a0",
          1397 => x"2e",
          1398 => x"51",
          1399 => x"84",
          1400 => x"53",
          1401 => x"73",
          1402 => x"38",
          1403 => x"bd",
          1404 => x"b9",
          1405 => x"52",
          1406 => x"9f",
          1407 => x"38",
          1408 => x"9f",
          1409 => x"81",
          1410 => x"2a",
          1411 => x"76",
          1412 => x"54",
          1413 => x"56",
          1414 => x"a8",
          1415 => x"74",
          1416 => x"74",
          1417 => x"78",
          1418 => x"11",
          1419 => x"81",
          1420 => x"06",
          1421 => x"ff",
          1422 => x"52",
          1423 => x"55",
          1424 => x"38",
          1425 => x"c8",
          1426 => x"0d",
          1427 => x"0d",
          1428 => x"7a",
          1429 => x"9f",
          1430 => x"7c",
          1431 => x"32",
          1432 => x"71",
          1433 => x"72",
          1434 => x"59",
          1435 => x"56",
          1436 => x"84",
          1437 => x"75",
          1438 => x"84",
          1439 => x"88",
          1440 => x"f7",
          1441 => x"7d",
          1442 => x"70",
          1443 => x"08",
          1444 => x"56",
          1445 => x"2e",
          1446 => x"8f",
          1447 => x"70",
          1448 => x"33",
          1449 => x"a0",
          1450 => x"73",
          1451 => x"f5",
          1452 => x"2e",
          1453 => x"d0",
          1454 => x"56",
          1455 => x"80",
          1456 => x"58",
          1457 => x"74",
          1458 => x"38",
          1459 => x"27",
          1460 => x"14",
          1461 => x"06",
          1462 => x"14",
          1463 => x"06",
          1464 => x"73",
          1465 => x"f9",
          1466 => x"ff",
          1467 => x"89",
          1468 => x"89",
          1469 => x"27",
          1470 => x"77",
          1471 => x"81",
          1472 => x"0c",
          1473 => x"56",
          1474 => x"26",
          1475 => x"78",
          1476 => x"38",
          1477 => x"75",
          1478 => x"56",
          1479 => x"c8",
          1480 => x"0d",
          1481 => x"16",
          1482 => x"70",
          1483 => x"59",
          1484 => x"09",
          1485 => x"ff",
          1486 => x"70",
          1487 => x"33",
          1488 => x"80",
          1489 => x"38",
          1490 => x"80",
          1491 => x"38",
          1492 => x"74",
          1493 => x"d0",
          1494 => x"56",
          1495 => x"73",
          1496 => x"38",
          1497 => x"c8",
          1498 => x"0d",
          1499 => x"81",
          1500 => x"0c",
          1501 => x"55",
          1502 => x"ca",
          1503 => x"84",
          1504 => x"8b",
          1505 => x"f7",
          1506 => x"7d",
          1507 => x"70",
          1508 => x"08",
          1509 => x"56",
          1510 => x"2e",
          1511 => x"8f",
          1512 => x"70",
          1513 => x"33",
          1514 => x"a0",
          1515 => x"73",
          1516 => x"f5",
          1517 => x"2e",
          1518 => x"d0",
          1519 => x"56",
          1520 => x"80",
          1521 => x"58",
          1522 => x"74",
          1523 => x"38",
          1524 => x"27",
          1525 => x"14",
          1526 => x"06",
          1527 => x"14",
          1528 => x"06",
          1529 => x"73",
          1530 => x"f9",
          1531 => x"ff",
          1532 => x"89",
          1533 => x"89",
          1534 => x"27",
          1535 => x"77",
          1536 => x"81",
          1537 => x"0c",
          1538 => x"56",
          1539 => x"26",
          1540 => x"78",
          1541 => x"38",
          1542 => x"75",
          1543 => x"56",
          1544 => x"c8",
          1545 => x"0d",
          1546 => x"16",
          1547 => x"70",
          1548 => x"59",
          1549 => x"09",
          1550 => x"ff",
          1551 => x"70",
          1552 => x"33",
          1553 => x"80",
          1554 => x"38",
          1555 => x"80",
          1556 => x"38",
          1557 => x"74",
          1558 => x"d0",
          1559 => x"56",
          1560 => x"73",
          1561 => x"38",
          1562 => x"c8",
          1563 => x"0d",
          1564 => x"81",
          1565 => x"0c",
          1566 => x"55",
          1567 => x"ca",
          1568 => x"84",
          1569 => x"8b",
          1570 => x"80",
          1571 => x"84",
          1572 => x"81",
          1573 => x"b9",
          1574 => x"ff",
          1575 => x"52",
          1576 => x"8c",
          1577 => x"10",
          1578 => x"05",
          1579 => x"04",
          1580 => x"51",
          1581 => x"83",
          1582 => x"83",
          1583 => x"ef",
          1584 => x"3d",
          1585 => x"ce",
          1586 => x"a8",
          1587 => x"0d",
          1588 => x"dc",
          1589 => x"3f",
          1590 => x"04",
          1591 => x"51",
          1592 => x"83",
          1593 => x"83",
          1594 => x"ef",
          1595 => x"3d",
          1596 => x"cf",
          1597 => x"fc",
          1598 => x"0d",
          1599 => x"b4",
          1600 => x"3f",
          1601 => x"04",
          1602 => x"51",
          1603 => x"83",
          1604 => x"83",
          1605 => x"ee",
          1606 => x"3d",
          1607 => x"d0",
          1608 => x"d0",
          1609 => x"0d",
          1610 => x"a4",
          1611 => x"3f",
          1612 => x"04",
          1613 => x"51",
          1614 => x"83",
          1615 => x"83",
          1616 => x"ee",
          1617 => x"3d",
          1618 => x"d0",
          1619 => x"a4",
          1620 => x"0d",
          1621 => x"f8",
          1622 => x"3f",
          1623 => x"04",
          1624 => x"51",
          1625 => x"83",
          1626 => x"83",
          1627 => x"ee",
          1628 => x"3d",
          1629 => x"d1",
          1630 => x"f8",
          1631 => x"0d",
          1632 => x"b8",
          1633 => x"3f",
          1634 => x"04",
          1635 => x"51",
          1636 => x"83",
          1637 => x"ec",
          1638 => x"02",
          1639 => x"e3",
          1640 => x"58",
          1641 => x"30",
          1642 => x"73",
          1643 => x"57",
          1644 => x"75",
          1645 => x"83",
          1646 => x"74",
          1647 => x"81",
          1648 => x"55",
          1649 => x"80",
          1650 => x"53",
          1651 => x"3d",
          1652 => x"82",
          1653 => x"84",
          1654 => x"57",
          1655 => x"08",
          1656 => x"d0",
          1657 => x"82",
          1658 => x"76",
          1659 => x"07",
          1660 => x"30",
          1661 => x"72",
          1662 => x"57",
          1663 => x"2e",
          1664 => x"c0",
          1665 => x"55",
          1666 => x"26",
          1667 => x"74",
          1668 => x"e8",
          1669 => x"8e",
          1670 => x"c8",
          1671 => x"d1",
          1672 => x"52",
          1673 => x"51",
          1674 => x"76",
          1675 => x"0c",
          1676 => x"04",
          1677 => x"08",
          1678 => x"88",
          1679 => x"c8",
          1680 => x"3d",
          1681 => x"84",
          1682 => x"52",
          1683 => x"9d",
          1684 => x"b9",
          1685 => x"84",
          1686 => x"ff",
          1687 => x"55",
          1688 => x"ff",
          1689 => x"19",
          1690 => x"59",
          1691 => x"e8",
          1692 => x"f4",
          1693 => x"b9",
          1694 => x"78",
          1695 => x"3f",
          1696 => x"08",
          1697 => x"f4",
          1698 => x"83",
          1699 => x"de",
          1700 => x"97",
          1701 => x"0d",
          1702 => x"05",
          1703 => x"58",
          1704 => x"80",
          1705 => x"7a",
          1706 => x"3f",
          1707 => x"08",
          1708 => x"80",
          1709 => x"76",
          1710 => x"38",
          1711 => x"c8",
          1712 => x"0d",
          1713 => x"84",
          1714 => x"61",
          1715 => x"84",
          1716 => x"7f",
          1717 => x"78",
          1718 => x"c8",
          1719 => x"c8",
          1720 => x"0d",
          1721 => x"0d",
          1722 => x"02",
          1723 => x"cf",
          1724 => x"73",
          1725 => x"5f",
          1726 => x"5d",
          1727 => x"2e",
          1728 => x"7a",
          1729 => x"fc",
          1730 => x"3f",
          1731 => x"51",
          1732 => x"80",
          1733 => x"27",
          1734 => x"90",
          1735 => x"38",
          1736 => x"82",
          1737 => x"18",
          1738 => x"27",
          1739 => x"72",
          1740 => x"d2",
          1741 => x"d1",
          1742 => x"84",
          1743 => x"53",
          1744 => x"ec",
          1745 => x"74",
          1746 => x"83",
          1747 => x"dd",
          1748 => x"56",
          1749 => x"80",
          1750 => x"18",
          1751 => x"53",
          1752 => x"7a",
          1753 => x"81",
          1754 => x"9f",
          1755 => x"38",
          1756 => x"73",
          1757 => x"ff",
          1758 => x"74",
          1759 => x"38",
          1760 => x"27",
          1761 => x"84",
          1762 => x"52",
          1763 => x"df",
          1764 => x"56",
          1765 => x"c2",
          1766 => x"94",
          1767 => x"3f",
          1768 => x"1c",
          1769 => x"51",
          1770 => x"84",
          1771 => x"98",
          1772 => x"2c",
          1773 => x"a0",
          1774 => x"38",
          1775 => x"82",
          1776 => x"1e",
          1777 => x"26",
          1778 => x"ff",
          1779 => x"c8",
          1780 => x"0d",
          1781 => x"98",
          1782 => x"3f",
          1783 => x"d5",
          1784 => x"54",
          1785 => x"87",
          1786 => x"26",
          1787 => x"fe",
          1788 => x"d2",
          1789 => x"91",
          1790 => x"84",
          1791 => x"53",
          1792 => x"ea",
          1793 => x"79",
          1794 => x"38",
          1795 => x"72",
          1796 => x"38",
          1797 => x"83",
          1798 => x"db",
          1799 => x"14",
          1800 => x"08",
          1801 => x"51",
          1802 => x"78",
          1803 => x"38",
          1804 => x"83",
          1805 => x"db",
          1806 => x"14",
          1807 => x"08",
          1808 => x"51",
          1809 => x"73",
          1810 => x"ff",
          1811 => x"53",
          1812 => x"df",
          1813 => x"52",
          1814 => x"51",
          1815 => x"84",
          1816 => x"ac",
          1817 => x"a0",
          1818 => x"3f",
          1819 => x"dd",
          1820 => x"39",
          1821 => x"08",
          1822 => x"e9",
          1823 => x"16",
          1824 => x"39",
          1825 => x"3f",
          1826 => x"08",
          1827 => x"53",
          1828 => x"a8",
          1829 => x"38",
          1830 => x"80",
          1831 => x"81",
          1832 => x"38",
          1833 => x"db",
          1834 => x"9b",
          1835 => x"b9",
          1836 => x"2b",
          1837 => x"70",
          1838 => x"30",
          1839 => x"70",
          1840 => x"07",
          1841 => x"06",
          1842 => x"59",
          1843 => x"72",
          1844 => x"e8",
          1845 => x"9b",
          1846 => x"b9",
          1847 => x"2b",
          1848 => x"70",
          1849 => x"30",
          1850 => x"70",
          1851 => x"07",
          1852 => x"06",
          1853 => x"59",
          1854 => x"80",
          1855 => x"a9",
          1856 => x"39",
          1857 => x"b9",
          1858 => x"3d",
          1859 => x"3d",
          1860 => x"96",
          1861 => x"aa",
          1862 => x"51",
          1863 => x"83",
          1864 => x"9d",
          1865 => x"51",
          1866 => x"72",
          1867 => x"81",
          1868 => x"71",
          1869 => x"72",
          1870 => x"81",
          1871 => x"71",
          1872 => x"72",
          1873 => x"81",
          1874 => x"71",
          1875 => x"72",
          1876 => x"81",
          1877 => x"71",
          1878 => x"72",
          1879 => x"81",
          1880 => x"71",
          1881 => x"72",
          1882 => x"81",
          1883 => x"71",
          1884 => x"72",
          1885 => x"81",
          1886 => x"71",
          1887 => x"88",
          1888 => x"53",
          1889 => x"a9",
          1890 => x"3d",
          1891 => x"51",
          1892 => x"83",
          1893 => x"9c",
          1894 => x"51",
          1895 => x"a9",
          1896 => x"3d",
          1897 => x"51",
          1898 => x"83",
          1899 => x"9c",
          1900 => x"51",
          1901 => x"72",
          1902 => x"06",
          1903 => x"2e",
          1904 => x"39",
          1905 => x"de",
          1906 => x"80",
          1907 => x"3f",
          1908 => x"d2",
          1909 => x"2a",
          1910 => x"51",
          1911 => x"2e",
          1912 => x"c2",
          1913 => x"9b",
          1914 => x"d4",
          1915 => x"ce",
          1916 => x"9b",
          1917 => x"86",
          1918 => x"06",
          1919 => x"80",
          1920 => x"38",
          1921 => x"81",
          1922 => x"3f",
          1923 => x"51",
          1924 => x"80",
          1925 => x"3f",
          1926 => x"70",
          1927 => x"52",
          1928 => x"fe",
          1929 => x"bd",
          1930 => x"9a",
          1931 => x"d4",
          1932 => x"8a",
          1933 => x"9a",
          1934 => x"84",
          1935 => x"06",
          1936 => x"80",
          1937 => x"38",
          1938 => x"81",
          1939 => x"3f",
          1940 => x"51",
          1941 => x"80",
          1942 => x"3f",
          1943 => x"70",
          1944 => x"52",
          1945 => x"fd",
          1946 => x"bd",
          1947 => x"9a",
          1948 => x"d4",
          1949 => x"c6",
          1950 => x"9a",
          1951 => x"82",
          1952 => x"06",
          1953 => x"80",
          1954 => x"38",
          1955 => x"ca",
          1956 => x"70",
          1957 => x"61",
          1958 => x"0c",
          1959 => x"60",
          1960 => x"8c",
          1961 => x"c8",
          1962 => x"06",
          1963 => x"59",
          1964 => x"84",
          1965 => x"d5",
          1966 => x"b8",
          1967 => x"43",
          1968 => x"51",
          1969 => x"7e",
          1970 => x"53",
          1971 => x"51",
          1972 => x"0b",
          1973 => x"bc",
          1974 => x"ff",
          1975 => x"79",
          1976 => x"f1",
          1977 => x"2e",
          1978 => x"78",
          1979 => x"5e",
          1980 => x"83",
          1981 => x"70",
          1982 => x"80",
          1983 => x"38",
          1984 => x"7b",
          1985 => x"81",
          1986 => x"81",
          1987 => x"5d",
          1988 => x"2e",
          1989 => x"5c",
          1990 => x"be",
          1991 => x"29",
          1992 => x"05",
          1993 => x"5b",
          1994 => x"84",
          1995 => x"84",
          1996 => x"54",
          1997 => x"08",
          1998 => x"da",
          1999 => x"c8",
          2000 => x"84",
          2001 => x"7d",
          2002 => x"80",
          2003 => x"70",
          2004 => x"5d",
          2005 => x"27",
          2006 => x"3d",
          2007 => x"80",
          2008 => x"38",
          2009 => x"7e",
          2010 => x"3f",
          2011 => x"08",
          2012 => x"c8",
          2013 => x"8d",
          2014 => x"b9",
          2015 => x"b8",
          2016 => x"05",
          2017 => x"3f",
          2018 => x"08",
          2019 => x"5c",
          2020 => x"2e",
          2021 => x"84",
          2022 => x"51",
          2023 => x"84",
          2024 => x"8f",
          2025 => x"38",
          2026 => x"3d",
          2027 => x"82",
          2028 => x"38",
          2029 => x"8c",
          2030 => x"81",
          2031 => x"38",
          2032 => x"53",
          2033 => x"52",
          2034 => x"dd",
          2035 => x"84",
          2036 => x"f8",
          2037 => x"67",
          2038 => x"90",
          2039 => x"90",
          2040 => x"7c",
          2041 => x"3f",
          2042 => x"08",
          2043 => x"08",
          2044 => x"70",
          2045 => x"25",
          2046 => x"42",
          2047 => x"83",
          2048 => x"81",
          2049 => x"06",
          2050 => x"2e",
          2051 => x"1b",
          2052 => x"06",
          2053 => x"ff",
          2054 => x"81",
          2055 => x"32",
          2056 => x"81",
          2057 => x"ff",
          2058 => x"38",
          2059 => x"94",
          2060 => x"d5",
          2061 => x"d1",
          2062 => x"80",
          2063 => x"52",
          2064 => x"bc",
          2065 => x"83",
          2066 => x"70",
          2067 => x"5b",
          2068 => x"91",
          2069 => x"83",
          2070 => x"84",
          2071 => x"82",
          2072 => x"84",
          2073 => x"80",
          2074 => x"0b",
          2075 => x"ee",
          2076 => x"d0",
          2077 => x"f8",
          2078 => x"82",
          2079 => x"84",
          2080 => x"80",
          2081 => x"84",
          2082 => x"51",
          2083 => x"0b",
          2084 => x"bc",
          2085 => x"ff",
          2086 => x"7d",
          2087 => x"81",
          2088 => x"38",
          2089 => x"d0",
          2090 => x"a1",
          2091 => x"0b",
          2092 => x"ee",
          2093 => x"d5",
          2094 => x"f8",
          2095 => x"a7",
          2096 => x"70",
          2097 => x"fc",
          2098 => x"39",
          2099 => x"0c",
          2100 => x"59",
          2101 => x"26",
          2102 => x"78",
          2103 => x"be",
          2104 => x"79",
          2105 => x"53",
          2106 => x"52",
          2107 => x"fb",
          2108 => x"7e",
          2109 => x"f4",
          2110 => x"84",
          2111 => x"c8",
          2112 => x"09",
          2113 => x"ae",
          2114 => x"9a",
          2115 => x"41",
          2116 => x"83",
          2117 => x"de",
          2118 => x"51",
          2119 => x"3f",
          2120 => x"83",
          2121 => x"7b",
          2122 => x"90",
          2123 => x"83",
          2124 => x"7c",
          2125 => x"3f",
          2126 => x"81",
          2127 => x"fa",
          2128 => x"f8",
          2129 => x"39",
          2130 => x"51",
          2131 => x"fa",
          2132 => x"8d",
          2133 => x"e8",
          2134 => x"a4",
          2135 => x"3f",
          2136 => x"04",
          2137 => x"51",
          2138 => x"d0",
          2139 => x"d0",
          2140 => x"ff",
          2141 => x"ff",
          2142 => x"ec",
          2143 => x"b9",
          2144 => x"2e",
          2145 => x"68",
          2146 => x"d4",
          2147 => x"3f",
          2148 => x"2d",
          2149 => x"08",
          2150 => x"a4",
          2151 => x"c8",
          2152 => x"d6",
          2153 => x"e1",
          2154 => x"39",
          2155 => x"84",
          2156 => x"80",
          2157 => x"cf",
          2158 => x"c8",
          2159 => x"f9",
          2160 => x"52",
          2161 => x"51",
          2162 => x"68",
          2163 => x"b8",
          2164 => x"11",
          2165 => x"05",
          2166 => x"3f",
          2167 => x"08",
          2168 => x"dc",
          2169 => x"fe",
          2170 => x"ff",
          2171 => x"e9",
          2172 => x"b9",
          2173 => x"d0",
          2174 => x"78",
          2175 => x"52",
          2176 => x"51",
          2177 => x"84",
          2178 => x"53",
          2179 => x"7e",
          2180 => x"3f",
          2181 => x"33",
          2182 => x"2e",
          2183 => x"78",
          2184 => x"d3",
          2185 => x"05",
          2186 => x"cf",
          2187 => x"fe",
          2188 => x"ff",
          2189 => x"e8",
          2190 => x"b9",
          2191 => x"2e",
          2192 => x"b8",
          2193 => x"11",
          2194 => x"05",
          2195 => x"3f",
          2196 => x"08",
          2197 => x"64",
          2198 => x"53",
          2199 => x"d7",
          2200 => x"a5",
          2201 => x"a8",
          2202 => x"f8",
          2203 => x"cf",
          2204 => x"48",
          2205 => x"78",
          2206 => x"c4",
          2207 => x"26",
          2208 => x"64",
          2209 => x"46",
          2210 => x"b8",
          2211 => x"11",
          2212 => x"05",
          2213 => x"3f",
          2214 => x"08",
          2215 => x"a0",
          2216 => x"fe",
          2217 => x"ff",
          2218 => x"e9",
          2219 => x"b9",
          2220 => x"2e",
          2221 => x"b8",
          2222 => x"11",
          2223 => x"05",
          2224 => x"3f",
          2225 => x"08",
          2226 => x"f4",
          2227 => x"c4",
          2228 => x"3f",
          2229 => x"59",
          2230 => x"83",
          2231 => x"70",
          2232 => x"5f",
          2233 => x"7d",
          2234 => x"7a",
          2235 => x"78",
          2236 => x"52",
          2237 => x"51",
          2238 => x"66",
          2239 => x"81",
          2240 => x"47",
          2241 => x"b8",
          2242 => x"11",
          2243 => x"05",
          2244 => x"3f",
          2245 => x"08",
          2246 => x"a4",
          2247 => x"fe",
          2248 => x"ff",
          2249 => x"e8",
          2250 => x"b9",
          2251 => x"2e",
          2252 => x"b8",
          2253 => x"11",
          2254 => x"05",
          2255 => x"3f",
          2256 => x"08",
          2257 => x"f8",
          2258 => x"f0",
          2259 => x"3f",
          2260 => x"67",
          2261 => x"38",
          2262 => x"70",
          2263 => x"33",
          2264 => x"81",
          2265 => x"39",
          2266 => x"84",
          2267 => x"80",
          2268 => x"93",
          2269 => x"c8",
          2270 => x"f6",
          2271 => x"3d",
          2272 => x"53",
          2273 => x"51",
          2274 => x"84",
          2275 => x"b1",
          2276 => x"33",
          2277 => x"d7",
          2278 => x"ed",
          2279 => x"a8",
          2280 => x"f8",
          2281 => x"cc",
          2282 => x"48",
          2283 => x"78",
          2284 => x"8c",
          2285 => x"26",
          2286 => x"68",
          2287 => x"d1",
          2288 => x"02",
          2289 => x"33",
          2290 => x"81",
          2291 => x"3d",
          2292 => x"53",
          2293 => x"51",
          2294 => x"84",
          2295 => x"80",
          2296 => x"38",
          2297 => x"80",
          2298 => x"79",
          2299 => x"05",
          2300 => x"fe",
          2301 => x"ff",
          2302 => x"e7",
          2303 => x"b9",
          2304 => x"bd",
          2305 => x"39",
          2306 => x"84",
          2307 => x"80",
          2308 => x"f3",
          2309 => x"c8",
          2310 => x"f5",
          2311 => x"3d",
          2312 => x"53",
          2313 => x"51",
          2314 => x"84",
          2315 => x"80",
          2316 => x"38",
          2317 => x"f8",
          2318 => x"80",
          2319 => x"c7",
          2320 => x"c8",
          2321 => x"84",
          2322 => x"46",
          2323 => x"51",
          2324 => x"68",
          2325 => x"78",
          2326 => x"38",
          2327 => x"79",
          2328 => x"5b",
          2329 => x"26",
          2330 => x"51",
          2331 => x"f4",
          2332 => x"3d",
          2333 => x"51",
          2334 => x"84",
          2335 => x"b9",
          2336 => x"05",
          2337 => x"f3",
          2338 => x"84",
          2339 => x"52",
          2340 => x"83",
          2341 => x"c8",
          2342 => x"f4",
          2343 => x"b9",
          2344 => x"e7",
          2345 => x"98",
          2346 => x"ff",
          2347 => x"ff",
          2348 => x"e5",
          2349 => x"b9",
          2350 => x"38",
          2351 => x"33",
          2352 => x"2e",
          2353 => x"83",
          2354 => x"49",
          2355 => x"fc",
          2356 => x"80",
          2357 => x"af",
          2358 => x"c8",
          2359 => x"83",
          2360 => x"5a",
          2361 => x"83",
          2362 => x"f2",
          2363 => x"b8",
          2364 => x"11",
          2365 => x"05",
          2366 => x"3f",
          2367 => x"08",
          2368 => x"38",
          2369 => x"5c",
          2370 => x"83",
          2371 => x"7a",
          2372 => x"30",
          2373 => x"9f",
          2374 => x"5c",
          2375 => x"80",
          2376 => x"7a",
          2377 => x"38",
          2378 => x"d8",
          2379 => x"c4",
          2380 => x"68",
          2381 => x"66",
          2382 => x"eb",
          2383 => x"d8",
          2384 => x"b0",
          2385 => x"39",
          2386 => x"0c",
          2387 => x"05",
          2388 => x"fe",
          2389 => x"ff",
          2390 => x"e2",
          2391 => x"b9",
          2392 => x"2e",
          2393 => x"64",
          2394 => x"59",
          2395 => x"45",
          2396 => x"f0",
          2397 => x"80",
          2398 => x"87",
          2399 => x"c8",
          2400 => x"f2",
          2401 => x"5e",
          2402 => x"05",
          2403 => x"82",
          2404 => x"7d",
          2405 => x"fe",
          2406 => x"ff",
          2407 => x"e1",
          2408 => x"b9",
          2409 => x"2e",
          2410 => x"64",
          2411 => x"ce",
          2412 => x"70",
          2413 => x"23",
          2414 => x"3d",
          2415 => x"53",
          2416 => x"51",
          2417 => x"84",
          2418 => x"ff",
          2419 => x"f0",
          2420 => x"fe",
          2421 => x"ff",
          2422 => x"e3",
          2423 => x"b9",
          2424 => x"2e",
          2425 => x"68",
          2426 => x"db",
          2427 => x"34",
          2428 => x"49",
          2429 => x"b8",
          2430 => x"11",
          2431 => x"05",
          2432 => x"3f",
          2433 => x"08",
          2434 => x"98",
          2435 => x"71",
          2436 => x"84",
          2437 => x"59",
          2438 => x"7a",
          2439 => x"81",
          2440 => x"38",
          2441 => x"d6",
          2442 => x"53",
          2443 => x"52",
          2444 => x"f5",
          2445 => x"39",
          2446 => x"51",
          2447 => x"f3",
          2448 => x"d8",
          2449 => x"ac",
          2450 => x"39",
          2451 => x"f0",
          2452 => x"80",
          2453 => x"ab",
          2454 => x"c8",
          2455 => x"b8",
          2456 => x"02",
          2457 => x"22",
          2458 => x"05",
          2459 => x"45",
          2460 => x"83",
          2461 => x"5c",
          2462 => x"80",
          2463 => x"f2",
          2464 => x"fc",
          2465 => x"f2",
          2466 => x"7b",
          2467 => x"38",
          2468 => x"08",
          2469 => x"39",
          2470 => x"51",
          2471 => x"64",
          2472 => x"39",
          2473 => x"51",
          2474 => x"64",
          2475 => x"39",
          2476 => x"33",
          2477 => x"2e",
          2478 => x"f2",
          2479 => x"fc",
          2480 => x"d8",
          2481 => x"ac",
          2482 => x"39",
          2483 => x"33",
          2484 => x"2e",
          2485 => x"f2",
          2486 => x"fc",
          2487 => x"f2",
          2488 => x"7d",
          2489 => x"38",
          2490 => x"08",
          2491 => x"39",
          2492 => x"33",
          2493 => x"2e",
          2494 => x"f2",
          2495 => x"fb",
          2496 => x"f2",
          2497 => x"7c",
          2498 => x"38",
          2499 => x"08",
          2500 => x"39",
          2501 => x"33",
          2502 => x"2e",
          2503 => x"f2",
          2504 => x"fb",
          2505 => x"f2",
          2506 => x"80",
          2507 => x"9c",
          2508 => x"b4",
          2509 => x"47",
          2510 => x"f3",
          2511 => x"0b",
          2512 => x"34",
          2513 => x"8c",
          2514 => x"57",
          2515 => x"52",
          2516 => x"d2",
          2517 => x"c8",
          2518 => x"77",
          2519 => x"87",
          2520 => x"75",
          2521 => x"3f",
          2522 => x"c8",
          2523 => x"0c",
          2524 => x"9c",
          2525 => x"57",
          2526 => x"52",
          2527 => x"a6",
          2528 => x"c8",
          2529 => x"77",
          2530 => x"87",
          2531 => x"75",
          2532 => x"3f",
          2533 => x"c8",
          2534 => x"0c",
          2535 => x"0b",
          2536 => x"84",
          2537 => x"83",
          2538 => x"94",
          2539 => x"bc",
          2540 => x"c7",
          2541 => x"02",
          2542 => x"05",
          2543 => x"84",
          2544 => x"89",
          2545 => x"13",
          2546 => x"0c",
          2547 => x"0c",
          2548 => x"3f",
          2549 => x"95",
          2550 => x"8d",
          2551 => x"3f",
          2552 => x"52",
          2553 => x"51",
          2554 => x"83",
          2555 => x"22",
          2556 => x"97",
          2557 => x"bc",
          2558 => x"c8",
          2559 => x"33",
          2560 => x"d0",
          2561 => x"3f",
          2562 => x"83",
          2563 => x"d0",
          2564 => x"52",
          2565 => x"51",
          2566 => x"90",
          2567 => x"83",
          2568 => x"c3",
          2569 => x"e7",
          2570 => x"fb",
          2571 => x"70",
          2572 => x"80",
          2573 => x"74",
          2574 => x"83",
          2575 => x"70",
          2576 => x"52",
          2577 => x"2e",
          2578 => x"91",
          2579 => x"70",
          2580 => x"ff",
          2581 => x"55",
          2582 => x"f1",
          2583 => x"ff",
          2584 => x"a2",
          2585 => x"38",
          2586 => x"81",
          2587 => x"38",
          2588 => x"70",
          2589 => x"53",
          2590 => x"a0",
          2591 => x"81",
          2592 => x"2e",
          2593 => x"80",
          2594 => x"81",
          2595 => x"39",
          2596 => x"ff",
          2597 => x"70",
          2598 => x"81",
          2599 => x"81",
          2600 => x"32",
          2601 => x"80",
          2602 => x"52",
          2603 => x"80",
          2604 => x"80",
          2605 => x"05",
          2606 => x"76",
          2607 => x"70",
          2608 => x"0c",
          2609 => x"04",
          2610 => x"c4",
          2611 => x"2e",
          2612 => x"81",
          2613 => x"72",
          2614 => x"ff",
          2615 => x"54",
          2616 => x"e4",
          2617 => x"e0",
          2618 => x"55",
          2619 => x"53",
          2620 => x"09",
          2621 => x"f8",
          2622 => x"fc",
          2623 => x"53",
          2624 => x"38",
          2625 => x"b9",
          2626 => x"3d",
          2627 => x"3d",
          2628 => x"72",
          2629 => x"3f",
          2630 => x"08",
          2631 => x"38",
          2632 => x"c8",
          2633 => x"0d",
          2634 => x"0d",
          2635 => x"33",
          2636 => x"53",
          2637 => x"8b",
          2638 => x"38",
          2639 => x"ff",
          2640 => x"52",
          2641 => x"81",
          2642 => x"13",
          2643 => x"52",
          2644 => x"80",
          2645 => x"13",
          2646 => x"52",
          2647 => x"80",
          2648 => x"13",
          2649 => x"52",
          2650 => x"80",
          2651 => x"13",
          2652 => x"52",
          2653 => x"26",
          2654 => x"8a",
          2655 => x"87",
          2656 => x"e7",
          2657 => x"38",
          2658 => x"c0",
          2659 => x"72",
          2660 => x"98",
          2661 => x"13",
          2662 => x"98",
          2663 => x"13",
          2664 => x"98",
          2665 => x"13",
          2666 => x"98",
          2667 => x"13",
          2668 => x"98",
          2669 => x"13",
          2670 => x"98",
          2671 => x"87",
          2672 => x"0c",
          2673 => x"98",
          2674 => x"0b",
          2675 => x"9c",
          2676 => x"71",
          2677 => x"0c",
          2678 => x"04",
          2679 => x"7f",
          2680 => x"98",
          2681 => x"7d",
          2682 => x"98",
          2683 => x"7d",
          2684 => x"c0",
          2685 => x"5c",
          2686 => x"34",
          2687 => x"b4",
          2688 => x"83",
          2689 => x"c0",
          2690 => x"5c",
          2691 => x"34",
          2692 => x"ac",
          2693 => x"85",
          2694 => x"c0",
          2695 => x"5c",
          2696 => x"34",
          2697 => x"a4",
          2698 => x"88",
          2699 => x"c0",
          2700 => x"5a",
          2701 => x"23",
          2702 => x"79",
          2703 => x"06",
          2704 => x"ff",
          2705 => x"86",
          2706 => x"85",
          2707 => x"84",
          2708 => x"83",
          2709 => x"82",
          2710 => x"7d",
          2711 => x"06",
          2712 => x"ec",
          2713 => x"a1",
          2714 => x"0d",
          2715 => x"0d",
          2716 => x"33",
          2717 => x"2e",
          2718 => x"51",
          2719 => x"3f",
          2720 => x"08",
          2721 => x"98",
          2722 => x"71",
          2723 => x"81",
          2724 => x"72",
          2725 => x"38",
          2726 => x"c8",
          2727 => x"0d",
          2728 => x"80",
          2729 => x"84",
          2730 => x"98",
          2731 => x"2c",
          2732 => x"ff",
          2733 => x"06",
          2734 => x"51",
          2735 => x"3f",
          2736 => x"08",
          2737 => x"98",
          2738 => x"71",
          2739 => x"38",
          2740 => x"3d",
          2741 => x"54",
          2742 => x"2b",
          2743 => x"80",
          2744 => x"84",
          2745 => x"98",
          2746 => x"2c",
          2747 => x"ff",
          2748 => x"73",
          2749 => x"14",
          2750 => x"73",
          2751 => x"71",
          2752 => x"0c",
          2753 => x"04",
          2754 => x"02",
          2755 => x"83",
          2756 => x"70",
          2757 => x"53",
          2758 => x"80",
          2759 => x"38",
          2760 => x"94",
          2761 => x"2a",
          2762 => x"53",
          2763 => x"80",
          2764 => x"71",
          2765 => x"81",
          2766 => x"70",
          2767 => x"81",
          2768 => x"53",
          2769 => x"8a",
          2770 => x"2a",
          2771 => x"71",
          2772 => x"81",
          2773 => x"87",
          2774 => x"52",
          2775 => x"86",
          2776 => x"94",
          2777 => x"72",
          2778 => x"b9",
          2779 => x"3d",
          2780 => x"91",
          2781 => x"06",
          2782 => x"97",
          2783 => x"32",
          2784 => x"72",
          2785 => x"38",
          2786 => x"81",
          2787 => x"80",
          2788 => x"87",
          2789 => x"08",
          2790 => x"70",
          2791 => x"54",
          2792 => x"38",
          2793 => x"3d",
          2794 => x"05",
          2795 => x"70",
          2796 => x"52",
          2797 => x"f2",
          2798 => x"3d",
          2799 => x"3d",
          2800 => x"80",
          2801 => x"56",
          2802 => x"77",
          2803 => x"38",
          2804 => x"f2",
          2805 => x"81",
          2806 => x"57",
          2807 => x"2e",
          2808 => x"87",
          2809 => x"08",
          2810 => x"70",
          2811 => x"54",
          2812 => x"2e",
          2813 => x"91",
          2814 => x"06",
          2815 => x"e3",
          2816 => x"32",
          2817 => x"72",
          2818 => x"38",
          2819 => x"81",
          2820 => x"cf",
          2821 => x"ff",
          2822 => x"c0",
          2823 => x"70",
          2824 => x"38",
          2825 => x"90",
          2826 => x"0c",
          2827 => x"33",
          2828 => x"ff",
          2829 => x"84",
          2830 => x"88",
          2831 => x"71",
          2832 => x"81",
          2833 => x"70",
          2834 => x"81",
          2835 => x"53",
          2836 => x"c1",
          2837 => x"2a",
          2838 => x"71",
          2839 => x"b5",
          2840 => x"94",
          2841 => x"96",
          2842 => x"06",
          2843 => x"70",
          2844 => x"39",
          2845 => x"87",
          2846 => x"08",
          2847 => x"8a",
          2848 => x"70",
          2849 => x"ab",
          2850 => x"9e",
          2851 => x"f2",
          2852 => x"c0",
          2853 => x"83",
          2854 => x"87",
          2855 => x"08",
          2856 => x"0c",
          2857 => x"98",
          2858 => x"90",
          2859 => x"9e",
          2860 => x"f2",
          2861 => x"c0",
          2862 => x"83",
          2863 => x"87",
          2864 => x"08",
          2865 => x"0c",
          2866 => x"b0",
          2867 => x"a0",
          2868 => x"9e",
          2869 => x"f2",
          2870 => x"c0",
          2871 => x"83",
          2872 => x"87",
          2873 => x"08",
          2874 => x"0c",
          2875 => x"c0",
          2876 => x"b0",
          2877 => x"9e",
          2878 => x"f2",
          2879 => x"c0",
          2880 => x"52",
          2881 => x"b8",
          2882 => x"9e",
          2883 => x"f2",
          2884 => x"c0",
          2885 => x"83",
          2886 => x"87",
          2887 => x"08",
          2888 => x"0c",
          2889 => x"f2",
          2890 => x"0b",
          2891 => x"90",
          2892 => x"80",
          2893 => x"52",
          2894 => x"fb",
          2895 => x"f2",
          2896 => x"0b",
          2897 => x"90",
          2898 => x"80",
          2899 => x"52",
          2900 => x"2e",
          2901 => x"52",
          2902 => x"ca",
          2903 => x"87",
          2904 => x"08",
          2905 => x"0a",
          2906 => x"52",
          2907 => x"83",
          2908 => x"71",
          2909 => x"34",
          2910 => x"c0",
          2911 => x"70",
          2912 => x"06",
          2913 => x"70",
          2914 => x"38",
          2915 => x"83",
          2916 => x"80",
          2917 => x"9e",
          2918 => x"a0",
          2919 => x"51",
          2920 => x"80",
          2921 => x"81",
          2922 => x"f2",
          2923 => x"0b",
          2924 => x"90",
          2925 => x"80",
          2926 => x"52",
          2927 => x"2e",
          2928 => x"52",
          2929 => x"ce",
          2930 => x"87",
          2931 => x"08",
          2932 => x"80",
          2933 => x"52",
          2934 => x"83",
          2935 => x"71",
          2936 => x"34",
          2937 => x"c0",
          2938 => x"70",
          2939 => x"06",
          2940 => x"70",
          2941 => x"38",
          2942 => x"83",
          2943 => x"80",
          2944 => x"9e",
          2945 => x"81",
          2946 => x"51",
          2947 => x"80",
          2948 => x"81",
          2949 => x"f2",
          2950 => x"0b",
          2951 => x"90",
          2952 => x"c0",
          2953 => x"52",
          2954 => x"2e",
          2955 => x"52",
          2956 => x"d2",
          2957 => x"87",
          2958 => x"08",
          2959 => x"06",
          2960 => x"70",
          2961 => x"38",
          2962 => x"83",
          2963 => x"87",
          2964 => x"08",
          2965 => x"70",
          2966 => x"51",
          2967 => x"d4",
          2968 => x"87",
          2969 => x"08",
          2970 => x"06",
          2971 => x"70",
          2972 => x"38",
          2973 => x"83",
          2974 => x"87",
          2975 => x"08",
          2976 => x"70",
          2977 => x"51",
          2978 => x"d6",
          2979 => x"87",
          2980 => x"08",
          2981 => x"51",
          2982 => x"80",
          2983 => x"81",
          2984 => x"f2",
          2985 => x"c0",
          2986 => x"87",
          2987 => x"83",
          2988 => x"83",
          2989 => x"81",
          2990 => x"39",
          2991 => x"83",
          2992 => x"ff",
          2993 => x"83",
          2994 => x"54",
          2995 => x"38",
          2996 => x"51",
          2997 => x"83",
          2998 => x"55",
          2999 => x"38",
          3000 => x"33",
          3001 => x"c6",
          3002 => x"cc",
          3003 => x"85",
          3004 => x"f2",
          3005 => x"74",
          3006 => x"83",
          3007 => x"54",
          3008 => x"38",
          3009 => x"33",
          3010 => x"a8",
          3011 => x"d7",
          3012 => x"84",
          3013 => x"f2",
          3014 => x"74",
          3015 => x"83",
          3016 => x"56",
          3017 => x"38",
          3018 => x"33",
          3019 => x"a6",
          3020 => x"d0",
          3021 => x"83",
          3022 => x"f2",
          3023 => x"75",
          3024 => x"83",
          3025 => x"54",
          3026 => x"38",
          3027 => x"51",
          3028 => x"83",
          3029 => x"52",
          3030 => x"51",
          3031 => x"3f",
          3032 => x"08",
          3033 => x"e4",
          3034 => x"9d",
          3035 => x"b4",
          3036 => x"da",
          3037 => x"b5",
          3038 => x"da",
          3039 => x"f4",
          3040 => x"b8",
          3041 => x"da",
          3042 => x"b4",
          3043 => x"f2",
          3044 => x"bd",
          3045 => x"75",
          3046 => x"3f",
          3047 => x"08",
          3048 => x"29",
          3049 => x"54",
          3050 => x"c8",
          3051 => x"da",
          3052 => x"b4",
          3053 => x"f2",
          3054 => x"74",
          3055 => x"f2",
          3056 => x"74",
          3057 => x"3d",
          3058 => x"f2",
          3059 => x"bd",
          3060 => x"75",
          3061 => x"3f",
          3062 => x"08",
          3063 => x"29",
          3064 => x"54",
          3065 => x"c8",
          3066 => x"db",
          3067 => x"b4",
          3068 => x"3d",
          3069 => x"f2",
          3070 => x"bd",
          3071 => x"75",
          3072 => x"3f",
          3073 => x"08",
          3074 => x"29",
          3075 => x"54",
          3076 => x"c8",
          3077 => x"db",
          3078 => x"b3",
          3079 => x"f2",
          3080 => x"74",
          3081 => x"9e",
          3082 => x"39",
          3083 => x"51",
          3084 => x"83",
          3085 => x"c0",
          3086 => x"f2",
          3087 => x"83",
          3088 => x"ff",
          3089 => x"83",
          3090 => x"52",
          3091 => x"51",
          3092 => x"3f",
          3093 => x"08",
          3094 => x"8c",
          3095 => x"a9",
          3096 => x"b4",
          3097 => x"3f",
          3098 => x"22",
          3099 => x"bc",
          3100 => x"95",
          3101 => x"bc",
          3102 => x"84",
          3103 => x"51",
          3104 => x"84",
          3105 => x"bd",
          3106 => x"76",
          3107 => x"54",
          3108 => x"08",
          3109 => x"e4",
          3110 => x"ed",
          3111 => x"cf",
          3112 => x"80",
          3113 => x"38",
          3114 => x"83",
          3115 => x"ff",
          3116 => x"83",
          3117 => x"54",
          3118 => x"fd",
          3119 => x"ec",
          3120 => x"f8",
          3121 => x"ac",
          3122 => x"d1",
          3123 => x"80",
          3124 => x"38",
          3125 => x"dc",
          3126 => x"bf",
          3127 => x"f2",
          3128 => x"74",
          3129 => x"d2",
          3130 => x"83",
          3131 => x"ff",
          3132 => x"83",
          3133 => x"54",
          3134 => x"fc",
          3135 => x"39",
          3136 => x"33",
          3137 => x"a4",
          3138 => x"fd",
          3139 => x"c9",
          3140 => x"80",
          3141 => x"38",
          3142 => x"f2",
          3143 => x"83",
          3144 => x"ff",
          3145 => x"83",
          3146 => x"55",
          3147 => x"fb",
          3148 => x"39",
          3149 => x"33",
          3150 => x"e4",
          3151 => x"c9",
          3152 => x"d7",
          3153 => x"80",
          3154 => x"38",
          3155 => x"f2",
          3156 => x"f2",
          3157 => x"54",
          3158 => x"84",
          3159 => x"a9",
          3160 => x"d3",
          3161 => x"80",
          3162 => x"38",
          3163 => x"f2",
          3164 => x"f2",
          3165 => x"54",
          3166 => x"a0",
          3167 => x"89",
          3168 => x"ce",
          3169 => x"80",
          3170 => x"38",
          3171 => x"f2",
          3172 => x"f2",
          3173 => x"54",
          3174 => x"bc",
          3175 => x"e9",
          3176 => x"cd",
          3177 => x"80",
          3178 => x"38",
          3179 => x"f2",
          3180 => x"f2",
          3181 => x"54",
          3182 => x"d8",
          3183 => x"c9",
          3184 => x"cc",
          3185 => x"80",
          3186 => x"38",
          3187 => x"f2",
          3188 => x"f2",
          3189 => x"54",
          3190 => x"f4",
          3191 => x"a9",
          3192 => x"cf",
          3193 => x"80",
          3194 => x"38",
          3195 => x"de",
          3196 => x"b0",
          3197 => x"d9",
          3198 => x"bc",
          3199 => x"f2",
          3200 => x"74",
          3201 => x"d8",
          3202 => x"ff",
          3203 => x"8e",
          3204 => x"71",
          3205 => x"38",
          3206 => x"83",
          3207 => x"52",
          3208 => x"83",
          3209 => x"ff",
          3210 => x"83",
          3211 => x"83",
          3212 => x"ff",
          3213 => x"83",
          3214 => x"83",
          3215 => x"ff",
          3216 => x"83",
          3217 => x"83",
          3218 => x"ff",
          3219 => x"83",
          3220 => x"83",
          3221 => x"ff",
          3222 => x"83",
          3223 => x"83",
          3224 => x"ff",
          3225 => x"83",
          3226 => x"71",
          3227 => x"04",
          3228 => x"c0",
          3229 => x"04",
          3230 => x"08",
          3231 => x"84",
          3232 => x"3d",
          3233 => x"08",
          3234 => x"5a",
          3235 => x"57",
          3236 => x"83",
          3237 => x"51",
          3238 => x"3f",
          3239 => x"08",
          3240 => x"8b",
          3241 => x"0b",
          3242 => x"08",
          3243 => x"f8",
          3244 => x"82",
          3245 => x"84",
          3246 => x"80",
          3247 => x"76",
          3248 => x"3f",
          3249 => x"08",
          3250 => x"55",
          3251 => x"b9",
          3252 => x"8e",
          3253 => x"c8",
          3254 => x"70",
          3255 => x"80",
          3256 => x"09",
          3257 => x"72",
          3258 => x"51",
          3259 => x"76",
          3260 => x"73",
          3261 => x"83",
          3262 => x"8c",
          3263 => x"51",
          3264 => x"3f",
          3265 => x"08",
          3266 => x"76",
          3267 => x"77",
          3268 => x"0c",
          3269 => x"04",
          3270 => x"51",
          3271 => x"3f",
          3272 => x"09",
          3273 => x"38",
          3274 => x"51",
          3275 => x"79",
          3276 => x"f5",
          3277 => x"08",
          3278 => x"c8",
          3279 => x"76",
          3280 => x"a8",
          3281 => x"c1",
          3282 => x"84",
          3283 => x"a9",
          3284 => x"d8",
          3285 => x"3d",
          3286 => x"08",
          3287 => x"72",
          3288 => x"5a",
          3289 => x"2e",
          3290 => x"80",
          3291 => x"59",
          3292 => x"10",
          3293 => x"bc",
          3294 => x"52",
          3295 => x"a9",
          3296 => x"c8",
          3297 => x"52",
          3298 => x"c0",
          3299 => x"b9",
          3300 => x"38",
          3301 => x"54",
          3302 => x"81",
          3303 => x"82",
          3304 => x"81",
          3305 => x"ff",
          3306 => x"82",
          3307 => x"38",
          3308 => x"84",
          3309 => x"aa",
          3310 => x"81",
          3311 => x"3d",
          3312 => x"53",
          3313 => x"51",
          3314 => x"84",
          3315 => x"80",
          3316 => x"ff",
          3317 => x"52",
          3318 => x"a6",
          3319 => x"c8",
          3320 => x"06",
          3321 => x"2e",
          3322 => x"16",
          3323 => x"06",
          3324 => x"76",
          3325 => x"38",
          3326 => x"78",
          3327 => x"56",
          3328 => x"fe",
          3329 => x"15",
          3330 => x"33",
          3331 => x"a0",
          3332 => x"06",
          3333 => x"75",
          3334 => x"38",
          3335 => x"3d",
          3336 => x"cd",
          3337 => x"b9",
          3338 => x"83",
          3339 => x"52",
          3340 => x"ea",
          3341 => x"c8",
          3342 => x"38",
          3343 => x"08",
          3344 => x"52",
          3345 => x"ce",
          3346 => x"b9",
          3347 => x"2e",
          3348 => x"51",
          3349 => x"3f",
          3350 => x"08",
          3351 => x"84",
          3352 => x"25",
          3353 => x"b9",
          3354 => x"05",
          3355 => x"55",
          3356 => x"77",
          3357 => x"81",
          3358 => x"f0",
          3359 => x"ab",
          3360 => x"ff",
          3361 => x"06",
          3362 => x"81",
          3363 => x"c8",
          3364 => x"0d",
          3365 => x"0d",
          3366 => x"b7",
          3367 => x"3d",
          3368 => x"5c",
          3369 => x"3d",
          3370 => x"b8",
          3371 => x"b4",
          3372 => x"74",
          3373 => x"83",
          3374 => x"56",
          3375 => x"2e",
          3376 => x"77",
          3377 => x"8d",
          3378 => x"77",
          3379 => x"78",
          3380 => x"77",
          3381 => x"fd",
          3382 => x"b4",
          3383 => x"80",
          3384 => x"3f",
          3385 => x"08",
          3386 => x"98",
          3387 => x"79",
          3388 => x"38",
          3389 => x"06",
          3390 => x"33",
          3391 => x"70",
          3392 => x"d1",
          3393 => x"98",
          3394 => x"2c",
          3395 => x"05",
          3396 => x"83",
          3397 => x"70",
          3398 => x"33",
          3399 => x"5d",
          3400 => x"58",
          3401 => x"57",
          3402 => x"80",
          3403 => x"75",
          3404 => x"38",
          3405 => x"0a",
          3406 => x"0a",
          3407 => x"2c",
          3408 => x"76",
          3409 => x"38",
          3410 => x"70",
          3411 => x"57",
          3412 => x"de",
          3413 => x"42",
          3414 => x"25",
          3415 => x"de",
          3416 => x"18",
          3417 => x"41",
          3418 => x"81",
          3419 => x"80",
          3420 => x"75",
          3421 => x"34",
          3422 => x"80",
          3423 => x"38",
          3424 => x"98",
          3425 => x"2c",
          3426 => x"33",
          3427 => x"70",
          3428 => x"98",
          3429 => x"82",
          3430 => x"d4",
          3431 => x"53",
          3432 => x"5d",
          3433 => x"78",
          3434 => x"38",
          3435 => x"84",
          3436 => x"39",
          3437 => x"ff",
          3438 => x"81",
          3439 => x"81",
          3440 => x"70",
          3441 => x"81",
          3442 => x"57",
          3443 => x"26",
          3444 => x"75",
          3445 => x"82",
          3446 => x"80",
          3447 => x"d4",
          3448 => x"57",
          3449 => x"ce",
          3450 => x"d0",
          3451 => x"70",
          3452 => x"78",
          3453 => x"bc",
          3454 => x"2e",
          3455 => x"fe",
          3456 => x"57",
          3457 => x"fe",
          3458 => x"e7",
          3459 => x"fd",
          3460 => x"57",
          3461 => x"38",
          3462 => x"84",
          3463 => x"d1",
          3464 => x"7e",
          3465 => x"0c",
          3466 => x"95",
          3467 => x"38",
          3468 => x"83",
          3469 => x"57",
          3470 => x"83",
          3471 => x"08",
          3472 => x"0b",
          3473 => x"34",
          3474 => x"d1",
          3475 => x"39",
          3476 => x"33",
          3477 => x"2e",
          3478 => x"84",
          3479 => x"52",
          3480 => x"b6",
          3481 => x"d1",
          3482 => x"05",
          3483 => x"d1",
          3484 => x"eb",
          3485 => x"8c",
          3486 => x"ff",
          3487 => x"88",
          3488 => x"55",
          3489 => x"fc",
          3490 => x"d5",
          3491 => x"81",
          3492 => x"84",
          3493 => x"7b",
          3494 => x"52",
          3495 => x"cf",
          3496 => x"39",
          3497 => x"8b",
          3498 => x"10",
          3499 => x"e4",
          3500 => x"57",
          3501 => x"83",
          3502 => x"d1",
          3503 => x"7c",
          3504 => x"88",
          3505 => x"8c",
          3506 => x"74",
          3507 => x"38",
          3508 => x"08",
          3509 => x"ff",
          3510 => x"84",
          3511 => x"52",
          3512 => x"b5",
          3513 => x"d5",
          3514 => x"88",
          3515 => x"ff",
          3516 => x"8c",
          3517 => x"5b",
          3518 => x"8c",
          3519 => x"ff",
          3520 => x"cc",
          3521 => x"ff",
          3522 => x"75",
          3523 => x"34",
          3524 => x"7c",
          3525 => x"f3",
          3526 => x"75",
          3527 => x"7c",
          3528 => x"f2",
          3529 => x"11",
          3530 => x"75",
          3531 => x"74",
          3532 => x"80",
          3533 => x"38",
          3534 => x"b7",
          3535 => x"b9",
          3536 => x"d1",
          3537 => x"b9",
          3538 => x"ff",
          3539 => x"53",
          3540 => x"51",
          3541 => x"3f",
          3542 => x"33",
          3543 => x"33",
          3544 => x"80",
          3545 => x"38",
          3546 => x"08",
          3547 => x"ff",
          3548 => x"84",
          3549 => x"52",
          3550 => x"b3",
          3551 => x"d5",
          3552 => x"88",
          3553 => x"e7",
          3554 => x"8c",
          3555 => x"55",
          3556 => x"8c",
          3557 => x"ff",
          3558 => x"39",
          3559 => x"33",
          3560 => x"06",
          3561 => x"33",
          3562 => x"75",
          3563 => x"af",
          3564 => x"ac",
          3565 => x"15",
          3566 => x"d1",
          3567 => x"16",
          3568 => x"55",
          3569 => x"3f",
          3570 => x"33",
          3571 => x"06",
          3572 => x"33",
          3573 => x"75",
          3574 => x"83",
          3575 => x"ac",
          3576 => x"15",
          3577 => x"d1",
          3578 => x"16",
          3579 => x"55",
          3580 => x"3f",
          3581 => x"33",
          3582 => x"06",
          3583 => x"33",
          3584 => x"77",
          3585 => x"a9",
          3586 => x"39",
          3587 => x"33",
          3588 => x"33",
          3589 => x"76",
          3590 => x"38",
          3591 => x"7a",
          3592 => x"34",
          3593 => x"70",
          3594 => x"81",
          3595 => x"57",
          3596 => x"24",
          3597 => x"84",
          3598 => x"52",
          3599 => x"b2",
          3600 => x"d1",
          3601 => x"98",
          3602 => x"2c",
          3603 => x"33",
          3604 => x"41",
          3605 => x"f9",
          3606 => x"d5",
          3607 => x"88",
          3608 => x"8b",
          3609 => x"80",
          3610 => x"80",
          3611 => x"98",
          3612 => x"88",
          3613 => x"5a",
          3614 => x"f8",
          3615 => x"d5",
          3616 => x"88",
          3617 => x"e7",
          3618 => x"80",
          3619 => x"80",
          3620 => x"98",
          3621 => x"88",
          3622 => x"5a",
          3623 => x"ff",
          3624 => x"bb",
          3625 => x"58",
          3626 => x"78",
          3627 => x"ac",
          3628 => x"33",
          3629 => x"b7",
          3630 => x"80",
          3631 => x"80",
          3632 => x"98",
          3633 => x"88",
          3634 => x"55",
          3635 => x"fe",
          3636 => x"16",
          3637 => x"33",
          3638 => x"d5",
          3639 => x"77",
          3640 => x"b1",
          3641 => x"81",
          3642 => x"81",
          3643 => x"70",
          3644 => x"d1",
          3645 => x"57",
          3646 => x"24",
          3647 => x"fe",
          3648 => x"d1",
          3649 => x"74",
          3650 => x"d3",
          3651 => x"ac",
          3652 => x"51",
          3653 => x"3f",
          3654 => x"33",
          3655 => x"76",
          3656 => x"34",
          3657 => x"06",
          3658 => x"84",
          3659 => x"7c",
          3660 => x"7f",
          3661 => x"ac",
          3662 => x"51",
          3663 => x"3f",
          3664 => x"52",
          3665 => x"8b",
          3666 => x"c8",
          3667 => x"06",
          3668 => x"cf",
          3669 => x"88",
          3670 => x"80",
          3671 => x"38",
          3672 => x"33",
          3673 => x"83",
          3674 => x"70",
          3675 => x"56",
          3676 => x"38",
          3677 => x"87",
          3678 => x"f2",
          3679 => x"18",
          3680 => x"5b",
          3681 => x"3f",
          3682 => x"08",
          3683 => x"f3",
          3684 => x"10",
          3685 => x"e0",
          3686 => x"57",
          3687 => x"8b",
          3688 => x"f3",
          3689 => x"75",
          3690 => x"38",
          3691 => x"33",
          3692 => x"2e",
          3693 => x"80",
          3694 => x"8c",
          3695 => x"84",
          3696 => x"7b",
          3697 => x"0c",
          3698 => x"04",
          3699 => x"33",
          3700 => x"2e",
          3701 => x"d5",
          3702 => x"88",
          3703 => x"8f",
          3704 => x"ac",
          3705 => x"51",
          3706 => x"3f",
          3707 => x"08",
          3708 => x"ff",
          3709 => x"84",
          3710 => x"ff",
          3711 => x"84",
          3712 => x"75",
          3713 => x"55",
          3714 => x"83",
          3715 => x"ff",
          3716 => x"80",
          3717 => x"8c",
          3718 => x"84",
          3719 => x"f5",
          3720 => x"7c",
          3721 => x"81",
          3722 => x"d1",
          3723 => x"74",
          3724 => x"38",
          3725 => x"08",
          3726 => x"ff",
          3727 => x"84",
          3728 => x"52",
          3729 => x"ae",
          3730 => x"d5",
          3731 => x"88",
          3732 => x"9b",
          3733 => x"8c",
          3734 => x"5d",
          3735 => x"8c",
          3736 => x"ff",
          3737 => x"cc",
          3738 => x"f0",
          3739 => x"99",
          3740 => x"84",
          3741 => x"80",
          3742 => x"88",
          3743 => x"b9",
          3744 => x"3d",
          3745 => x"d1",
          3746 => x"81",
          3747 => x"56",
          3748 => x"f4",
          3749 => x"d1",
          3750 => x"05",
          3751 => x"d1",
          3752 => x"16",
          3753 => x"d1",
          3754 => x"d5",
          3755 => x"88",
          3756 => x"bb",
          3757 => x"8c",
          3758 => x"2b",
          3759 => x"84",
          3760 => x"5a",
          3761 => x"76",
          3762 => x"ef",
          3763 => x"ac",
          3764 => x"51",
          3765 => x"3f",
          3766 => x"33",
          3767 => x"70",
          3768 => x"d1",
          3769 => x"57",
          3770 => x"7a",
          3771 => x"38",
          3772 => x"08",
          3773 => x"ff",
          3774 => x"74",
          3775 => x"29",
          3776 => x"05",
          3777 => x"84",
          3778 => x"5b",
          3779 => x"79",
          3780 => x"38",
          3781 => x"08",
          3782 => x"ff",
          3783 => x"74",
          3784 => x"29",
          3785 => x"05",
          3786 => x"84",
          3787 => x"5b",
          3788 => x"75",
          3789 => x"38",
          3790 => x"7b",
          3791 => x"17",
          3792 => x"84",
          3793 => x"52",
          3794 => x"ff",
          3795 => x"75",
          3796 => x"29",
          3797 => x"05",
          3798 => x"84",
          3799 => x"43",
          3800 => x"61",
          3801 => x"38",
          3802 => x"81",
          3803 => x"34",
          3804 => x"08",
          3805 => x"51",
          3806 => x"3f",
          3807 => x"0a",
          3808 => x"0a",
          3809 => x"2c",
          3810 => x"33",
          3811 => x"60",
          3812 => x"a7",
          3813 => x"39",
          3814 => x"33",
          3815 => x"06",
          3816 => x"60",
          3817 => x"38",
          3818 => x"33",
          3819 => x"27",
          3820 => x"98",
          3821 => x"2c",
          3822 => x"76",
          3823 => x"7b",
          3824 => x"33",
          3825 => x"75",
          3826 => x"29",
          3827 => x"05",
          3828 => x"84",
          3829 => x"52",
          3830 => x"78",
          3831 => x"81",
          3832 => x"84",
          3833 => x"77",
          3834 => x"7c",
          3835 => x"3d",
          3836 => x"84",
          3837 => x"57",
          3838 => x"8b",
          3839 => x"56",
          3840 => x"88",
          3841 => x"84",
          3842 => x"70",
          3843 => x"29",
          3844 => x"05",
          3845 => x"79",
          3846 => x"44",
          3847 => x"60",
          3848 => x"ef",
          3849 => x"2b",
          3850 => x"78",
          3851 => x"5c",
          3852 => x"7a",
          3853 => x"38",
          3854 => x"08",
          3855 => x"ff",
          3856 => x"75",
          3857 => x"29",
          3858 => x"05",
          3859 => x"84",
          3860 => x"57",
          3861 => x"75",
          3862 => x"38",
          3863 => x"08",
          3864 => x"ff",
          3865 => x"75",
          3866 => x"29",
          3867 => x"05",
          3868 => x"84",
          3869 => x"57",
          3870 => x"76",
          3871 => x"38",
          3872 => x"83",
          3873 => x"56",
          3874 => x"f4",
          3875 => x"51",
          3876 => x"3f",
          3877 => x"08",
          3878 => x"34",
          3879 => x"08",
          3880 => x"81",
          3881 => x"52",
          3882 => x"ad",
          3883 => x"d1",
          3884 => x"d1",
          3885 => x"56",
          3886 => x"f4",
          3887 => x"d5",
          3888 => x"88",
          3889 => x"a7",
          3890 => x"ac",
          3891 => x"51",
          3892 => x"3f",
          3893 => x"08",
          3894 => x"ff",
          3895 => x"84",
          3896 => x"ff",
          3897 => x"84",
          3898 => x"7a",
          3899 => x"55",
          3900 => x"51",
          3901 => x"3f",
          3902 => x"08",
          3903 => x"0c",
          3904 => x"08",
          3905 => x"76",
          3906 => x"34",
          3907 => x"38",
          3908 => x"84",
          3909 => x"52",
          3910 => x"33",
          3911 => x"a8",
          3912 => x"81",
          3913 => x"81",
          3914 => x"70",
          3915 => x"d1",
          3916 => x"57",
          3917 => x"24",
          3918 => x"d1",
          3919 => x"98",
          3920 => x"2c",
          3921 => x"06",
          3922 => x"58",
          3923 => x"ef",
          3924 => x"e4",
          3925 => x"b4",
          3926 => x"ee",
          3927 => x"f2",
          3928 => x"56",
          3929 => x"74",
          3930 => x"16",
          3931 => x"56",
          3932 => x"f0",
          3933 => x"83",
          3934 => x"83",
          3935 => x"55",
          3936 => x"ee",
          3937 => x"51",
          3938 => x"3f",
          3939 => x"08",
          3940 => x"fe",
          3941 => x"83",
          3942 => x"93",
          3943 => x"5f",
          3944 => x"39",
          3945 => x"d9",
          3946 => x"77",
          3947 => x"84",
          3948 => x"75",
          3949 => x"ac",
          3950 => x"39",
          3951 => x"aa",
          3952 => x"b9",
          3953 => x"d1",
          3954 => x"b9",
          3955 => x"ff",
          3956 => x"53",
          3957 => x"51",
          3958 => x"3f",
          3959 => x"d1",
          3960 => x"d1",
          3961 => x"57",
          3962 => x"2e",
          3963 => x"84",
          3964 => x"52",
          3965 => x"a6",
          3966 => x"d5",
          3967 => x"a0",
          3968 => x"eb",
          3969 => x"ac",
          3970 => x"51",
          3971 => x"3f",
          3972 => x"33",
          3973 => x"79",
          3974 => x"34",
          3975 => x"06",
          3976 => x"80",
          3977 => x"0b",
          3978 => x"34",
          3979 => x"d1",
          3980 => x"84",
          3981 => x"b4",
          3982 => x"75",
          3983 => x"e9",
          3984 => x"c8",
          3985 => x"88",
          3986 => x"c8",
          3987 => x"06",
          3988 => x"75",
          3989 => x"ff",
          3990 => x"81",
          3991 => x"ff",
          3992 => x"88",
          3993 => x"8c",
          3994 => x"5e",
          3995 => x"2e",
          3996 => x"84",
          3997 => x"52",
          3998 => x"a5",
          3999 => x"d5",
          4000 => x"a0",
          4001 => x"e7",
          4002 => x"ac",
          4003 => x"51",
          4004 => x"3f",
          4005 => x"33",
          4006 => x"76",
          4007 => x"34",
          4008 => x"06",
          4009 => x"75",
          4010 => x"fd",
          4011 => x"c8",
          4012 => x"88",
          4013 => x"c8",
          4014 => x"06",
          4015 => x"75",
          4016 => x"ff",
          4017 => x"ff",
          4018 => x"ff",
          4019 => x"88",
          4020 => x"8c",
          4021 => x"5e",
          4022 => x"2e",
          4023 => x"84",
          4024 => x"52",
          4025 => x"a5",
          4026 => x"d5",
          4027 => x"a0",
          4028 => x"fb",
          4029 => x"ac",
          4030 => x"51",
          4031 => x"3f",
          4032 => x"33",
          4033 => x"60",
          4034 => x"34",
          4035 => x"06",
          4036 => x"74",
          4037 => x"fa",
          4038 => x"b8",
          4039 => x"2b",
          4040 => x"83",
          4041 => x"81",
          4042 => x"52",
          4043 => x"dc",
          4044 => x"b9",
          4045 => x"0c",
          4046 => x"33",
          4047 => x"83",
          4048 => x"70",
          4049 => x"41",
          4050 => x"f4",
          4051 => x"53",
          4052 => x"51",
          4053 => x"3f",
          4054 => x"33",
          4055 => x"81",
          4056 => x"56",
          4057 => x"82",
          4058 => x"83",
          4059 => x"f4",
          4060 => x"3d",
          4061 => x"54",
          4062 => x"52",
          4063 => x"d8",
          4064 => x"f3",
          4065 => x"8a",
          4066 => x"88",
          4067 => x"b4",
          4068 => x"df",
          4069 => x"0b",
          4070 => x"34",
          4071 => x"d1",
          4072 => x"84",
          4073 => x"b4",
          4074 => x"93",
          4075 => x"84",
          4076 => x"51",
          4077 => x"3f",
          4078 => x"08",
          4079 => x"84",
          4080 => x"96",
          4081 => x"83",
          4082 => x"53",
          4083 => x"7a",
          4084 => x"f2",
          4085 => x"c8",
          4086 => x"b9",
          4087 => x"2e",
          4088 => x"e9",
          4089 => x"b9",
          4090 => x"ff",
          4091 => x"84",
          4092 => x"56",
          4093 => x"b9",
          4094 => x"80",
          4095 => x"b9",
          4096 => x"05",
          4097 => x"56",
          4098 => x"75",
          4099 => x"83",
          4100 => x"70",
          4101 => x"f2",
          4102 => x"08",
          4103 => x"59",
          4104 => x"38",
          4105 => x"87",
          4106 => x"f2",
          4107 => x"1a",
          4108 => x"55",
          4109 => x"3f",
          4110 => x"08",
          4111 => x"f3",
          4112 => x"10",
          4113 => x"e0",
          4114 => x"57",
          4115 => x"a0",
          4116 => x"70",
          4117 => x"5e",
          4118 => x"27",
          4119 => x"5d",
          4120 => x"09",
          4121 => x"df",
          4122 => x"ed",
          4123 => x"39",
          4124 => x"52",
          4125 => x"a5",
          4126 => x"f3",
          4127 => x"05",
          4128 => x"06",
          4129 => x"7a",
          4130 => x"38",
          4131 => x"f3",
          4132 => x"bd",
          4133 => x"80",
          4134 => x"83",
          4135 => x"70",
          4136 => x"fc",
          4137 => x"e0",
          4138 => x"70",
          4139 => x"57",
          4140 => x"3f",
          4141 => x"08",
          4142 => x"f3",
          4143 => x"10",
          4144 => x"e0",
          4145 => x"57",
          4146 => x"80",
          4147 => x"38",
          4148 => x"76",
          4149 => x"34",
          4150 => x"75",
          4151 => x"34",
          4152 => x"83",
          4153 => x"ff",
          4154 => x"77",
          4155 => x"f8",
          4156 => x"3d",
          4157 => x"c3",
          4158 => x"84",
          4159 => x"05",
          4160 => x"72",
          4161 => x"8d",
          4162 => x"2e",
          4163 => x"81",
          4164 => x"9e",
          4165 => x"2e",
          4166 => x"86",
          4167 => x"59",
          4168 => x"80",
          4169 => x"80",
          4170 => x"58",
          4171 => x"90",
          4172 => x"f8",
          4173 => x"83",
          4174 => x"75",
          4175 => x"23",
          4176 => x"33",
          4177 => x"71",
          4178 => x"71",
          4179 => x"71",
          4180 => x"56",
          4181 => x"78",
          4182 => x"38",
          4183 => x"84",
          4184 => x"74",
          4185 => x"05",
          4186 => x"74",
          4187 => x"75",
          4188 => x"38",
          4189 => x"33",
          4190 => x"17",
          4191 => x"55",
          4192 => x"0b",
          4193 => x"34",
          4194 => x"81",
          4195 => x"ff",
          4196 => x"ee",
          4197 => x"0d",
          4198 => x"a0",
          4199 => x"f8",
          4200 => x"10",
          4201 => x"f8",
          4202 => x"90",
          4203 => x"05",
          4204 => x"40",
          4205 => x"b0",
          4206 => x"b7",
          4207 => x"81",
          4208 => x"b7",
          4209 => x"81",
          4210 => x"f8",
          4211 => x"83",
          4212 => x"70",
          4213 => x"59",
          4214 => x"57",
          4215 => x"73",
          4216 => x"72",
          4217 => x"29",
          4218 => x"ff",
          4219 => x"ff",
          4220 => x"ff",
          4221 => x"ff",
          4222 => x"81",
          4223 => x"75",
          4224 => x"42",
          4225 => x"5c",
          4226 => x"8f",
          4227 => x"f8",
          4228 => x"31",
          4229 => x"29",
          4230 => x"76",
          4231 => x"7b",
          4232 => x"9c",
          4233 => x"55",
          4234 => x"26",
          4235 => x"80",
          4236 => x"05",
          4237 => x"f8",
          4238 => x"70",
          4239 => x"34",
          4240 => x"a7",
          4241 => x"86",
          4242 => x"70",
          4243 => x"33",
          4244 => x"06",
          4245 => x"33",
          4246 => x"06",
          4247 => x"22",
          4248 => x"5d",
          4249 => x"5e",
          4250 => x"74",
          4251 => x"df",
          4252 => x"ff",
          4253 => x"ff",
          4254 => x"29",
          4255 => x"54",
          4256 => x"fd",
          4257 => x"0b",
          4258 => x"34",
          4259 => x"f8",
          4260 => x"f8",
          4261 => x"98",
          4262 => x"2b",
          4263 => x"2b",
          4264 => x"7a",
          4265 => x"56",
          4266 => x"26",
          4267 => x"fd",
          4268 => x"fc",
          4269 => x"f8",
          4270 => x"81",
          4271 => x"10",
          4272 => x"f8",
          4273 => x"90",
          4274 => x"a7",
          4275 => x"5e",
          4276 => x"56",
          4277 => x"b0",
          4278 => x"84",
          4279 => x"70",
          4280 => x"84",
          4281 => x"70",
          4282 => x"83",
          4283 => x"70",
          4284 => x"06",
          4285 => x"60",
          4286 => x"41",
          4287 => x"40",
          4288 => x"73",
          4289 => x"72",
          4290 => x"70",
          4291 => x"57",
          4292 => x"ff",
          4293 => x"ff",
          4294 => x"29",
          4295 => x"ff",
          4296 => x"ff",
          4297 => x"29",
          4298 => x"5c",
          4299 => x"78",
          4300 => x"77",
          4301 => x"79",
          4302 => x"79",
          4303 => x"58",
          4304 => x"38",
          4305 => x"5c",
          4306 => x"38",
          4307 => x"74",
          4308 => x"29",
          4309 => x"39",
          4310 => x"87",
          4311 => x"53",
          4312 => x"34",
          4313 => x"85",
          4314 => x"73",
          4315 => x"80",
          4316 => x"f4",
          4317 => x"b0",
          4318 => x"8e",
          4319 => x"80",
          4320 => x"76",
          4321 => x"80",
          4322 => x"74",
          4323 => x"34",
          4324 => x"34",
          4325 => x"51",
          4326 => x"86",
          4327 => x"70",
          4328 => x"81",
          4329 => x"a0",
          4330 => x"77",
          4331 => x"54",
          4332 => x"34",
          4333 => x"80",
          4334 => x"c0",
          4335 => x"72",
          4336 => x"a0",
          4337 => x"70",
          4338 => x"07",
          4339 => x"86",
          4340 => x"34",
          4341 => x"f7",
          4342 => x"53",
          4343 => x"80",
          4344 => x"b7",
          4345 => x"0b",
          4346 => x"0c",
          4347 => x"04",
          4348 => x"33",
          4349 => x"0c",
          4350 => x"0d",
          4351 => x"33",
          4352 => x"b3",
          4353 => x"b7",
          4354 => x"59",
          4355 => x"75",
          4356 => x"da",
          4357 => x"bc",
          4358 => x"f9",
          4359 => x"f8",
          4360 => x"29",
          4361 => x"a0",
          4362 => x"f8",
          4363 => x"51",
          4364 => x"7c",
          4365 => x"83",
          4366 => x"83",
          4367 => x"53",
          4368 => x"72",
          4369 => x"c4",
          4370 => x"f6",
          4371 => x"55",
          4372 => x"f6",
          4373 => x"f8",
          4374 => x"70",
          4375 => x"7a",
          4376 => x"55",
          4377 => x"7a",
          4378 => x"38",
          4379 => x"72",
          4380 => x"34",
          4381 => x"22",
          4382 => x"ff",
          4383 => x"ba",
          4384 => x"57",
          4385 => x"82",
          4386 => x"b7",
          4387 => x"71",
          4388 => x"80",
          4389 => x"9f",
          4390 => x"84",
          4391 => x"14",
          4392 => x"e0",
          4393 => x"e0",
          4394 => x"70",
          4395 => x"33",
          4396 => x"05",
          4397 => x"14",
          4398 => x"b9",
          4399 => x"38",
          4400 => x"26",
          4401 => x"f8",
          4402 => x"98",
          4403 => x"55",
          4404 => x"e0",
          4405 => x"73",
          4406 => x"55",
          4407 => x"54",
          4408 => x"27",
          4409 => x"b7",
          4410 => x"05",
          4411 => x"f8",
          4412 => x"57",
          4413 => x"06",
          4414 => x"ff",
          4415 => x"73",
          4416 => x"fd",
          4417 => x"31",
          4418 => x"b7",
          4419 => x"71",
          4420 => x"57",
          4421 => x"a7",
          4422 => x"86",
          4423 => x"79",
          4424 => x"75",
          4425 => x"71",
          4426 => x"5c",
          4427 => x"75",
          4428 => x"38",
          4429 => x"16",
          4430 => x"14",
          4431 => x"b7",
          4432 => x"78",
          4433 => x"5a",
          4434 => x"81",
          4435 => x"77",
          4436 => x"59",
          4437 => x"84",
          4438 => x"84",
          4439 => x"71",
          4440 => x"56",
          4441 => x"72",
          4442 => x"38",
          4443 => x"84",
          4444 => x"8b",
          4445 => x"74",
          4446 => x"34",
          4447 => x"22",
          4448 => x"ff",
          4449 => x"ba",
          4450 => x"57",
          4451 => x"fd",
          4452 => x"80",
          4453 => x"38",
          4454 => x"06",
          4455 => x"f8",
          4456 => x"53",
          4457 => x"09",
          4458 => x"c8",
          4459 => x"31",
          4460 => x"b7",
          4461 => x"71",
          4462 => x"29",
          4463 => x"59",
          4464 => x"27",
          4465 => x"83",
          4466 => x"84",
          4467 => x"74",
          4468 => x"56",
          4469 => x"e0",
          4470 => x"75",
          4471 => x"05",
          4472 => x"13",
          4473 => x"2e",
          4474 => x"a0",
          4475 => x"16",
          4476 => x"70",
          4477 => x"34",
          4478 => x"72",
          4479 => x"f4",
          4480 => x"84",
          4481 => x"55",
          4482 => x"39",
          4483 => x"15",
          4484 => x"b7",
          4485 => x"74",
          4486 => x"bb",
          4487 => x"a9",
          4488 => x"0d",
          4489 => x"05",
          4490 => x"53",
          4491 => x"26",
          4492 => x"10",
          4493 => x"ec",
          4494 => x"08",
          4495 => x"bc",
          4496 => x"71",
          4497 => x"71",
          4498 => x"34",
          4499 => x"b9",
          4500 => x"3d",
          4501 => x"0b",
          4502 => x"34",
          4503 => x"33",
          4504 => x"06",
          4505 => x"80",
          4506 => x"ff",
          4507 => x"83",
          4508 => x"80",
          4509 => x"c8",
          4510 => x"0d",
          4511 => x"f8",
          4512 => x"31",
          4513 => x"9f",
          4514 => x"54",
          4515 => x"70",
          4516 => x"34",
          4517 => x"f8",
          4518 => x"05",
          4519 => x"33",
          4520 => x"56",
          4521 => x"25",
          4522 => x"53",
          4523 => x"f8",
          4524 => x"84",
          4525 => x"86",
          4526 => x"83",
          4527 => x"70",
          4528 => x"09",
          4529 => x"72",
          4530 => x"53",
          4531 => x"f8",
          4532 => x"0b",
          4533 => x"0c",
          4534 => x"04",
          4535 => x"33",
          4536 => x"b7",
          4537 => x"11",
          4538 => x"70",
          4539 => x"38",
          4540 => x"83",
          4541 => x"80",
          4542 => x"c8",
          4543 => x"0d",
          4544 => x"83",
          4545 => x"83",
          4546 => x"84",
          4547 => x"ff",
          4548 => x"71",
          4549 => x"b4",
          4550 => x"51",
          4551 => x"f8",
          4552 => x"39",
          4553 => x"02",
          4554 => x"51",
          4555 => x"b3",
          4556 => x"10",
          4557 => x"05",
          4558 => x"04",
          4559 => x"33",
          4560 => x"06",
          4561 => x"80",
          4562 => x"72",
          4563 => x"51",
          4564 => x"71",
          4565 => x"09",
          4566 => x"38",
          4567 => x"83",
          4568 => x"80",
          4569 => x"c8",
          4570 => x"0d",
          4571 => x"f4",
          4572 => x"06",
          4573 => x"70",
          4574 => x"34",
          4575 => x"b9",
          4576 => x"3d",
          4577 => x"f8",
          4578 => x"f0",
          4579 => x"83",
          4580 => x"e8",
          4581 => x"f4",
          4582 => x"06",
          4583 => x"70",
          4584 => x"34",
          4585 => x"f1",
          4586 => x"f4",
          4587 => x"84",
          4588 => x"83",
          4589 => x"83",
          4590 => x"81",
          4591 => x"07",
          4592 => x"f8",
          4593 => x"b4",
          4594 => x"f4",
          4595 => x"51",
          4596 => x"f4",
          4597 => x"39",
          4598 => x"33",
          4599 => x"85",
          4600 => x"83",
          4601 => x"ff",
          4602 => x"f8",
          4603 => x"fb",
          4604 => x"51",
          4605 => x"f4",
          4606 => x"39",
          4607 => x"33",
          4608 => x"81",
          4609 => x"83",
          4610 => x"fe",
          4611 => x"f8",
          4612 => x"f8",
          4613 => x"83",
          4614 => x"fe",
          4615 => x"f8",
          4616 => x"df",
          4617 => x"07",
          4618 => x"f8",
          4619 => x"cc",
          4620 => x"f4",
          4621 => x"06",
          4622 => x"70",
          4623 => x"34",
          4624 => x"83",
          4625 => x"81",
          4626 => x"e0",
          4627 => x"83",
          4628 => x"fe",
          4629 => x"f8",
          4630 => x"cf",
          4631 => x"07",
          4632 => x"f8",
          4633 => x"94",
          4634 => x"f4",
          4635 => x"06",
          4636 => x"70",
          4637 => x"34",
          4638 => x"83",
          4639 => x"81",
          4640 => x"70",
          4641 => x"34",
          4642 => x"83",
          4643 => x"81",
          4644 => x"07",
          4645 => x"f8",
          4646 => x"e0",
          4647 => x"0d",
          4648 => x"33",
          4649 => x"80",
          4650 => x"83",
          4651 => x"83",
          4652 => x"83",
          4653 => x"84",
          4654 => x"43",
          4655 => x"5b",
          4656 => x"2e",
          4657 => x"78",
          4658 => x"38",
          4659 => x"81",
          4660 => x"84",
          4661 => x"80",
          4662 => x"c0",
          4663 => x"f8",
          4664 => x"83",
          4665 => x"7c",
          4666 => x"34",
          4667 => x"04",
          4668 => x"09",
          4669 => x"38",
          4670 => x"b7",
          4671 => x"0b",
          4672 => x"34",
          4673 => x"f8",
          4674 => x"0b",
          4675 => x"34",
          4676 => x"f8",
          4677 => x"58",
          4678 => x"33",
          4679 => x"bb",
          4680 => x"b7",
          4681 => x"7b",
          4682 => x"7a",
          4683 => x"bc",
          4684 => x"d5",
          4685 => x"b7",
          4686 => x"0b",
          4687 => x"34",
          4688 => x"f8",
          4689 => x"f8",
          4690 => x"83",
          4691 => x"8f",
          4692 => x"80",
          4693 => x"be",
          4694 => x"84",
          4695 => x"80",
          4696 => x"f8",
          4697 => x"83",
          4698 => x"80",
          4699 => x"f6",
          4700 => x"cb",
          4701 => x"b8",
          4702 => x"84",
          4703 => x"56",
          4704 => x"54",
          4705 => x"52",
          4706 => x"51",
          4707 => x"3f",
          4708 => x"b8",
          4709 => x"5a",
          4710 => x"a5",
          4711 => x"84",
          4712 => x"70",
          4713 => x"83",
          4714 => x"ff",
          4715 => x"81",
          4716 => x"ff",
          4717 => x"c9",
          4718 => x"59",
          4719 => x"dd",
          4720 => x"a4",
          4721 => x"c1",
          4722 => x"b7",
          4723 => x"0b",
          4724 => x"34",
          4725 => x"f8",
          4726 => x"f8",
          4727 => x"83",
          4728 => x"8f",
          4729 => x"80",
          4730 => x"be",
          4731 => x"84",
          4732 => x"81",
          4733 => x"f8",
          4734 => x"83",
          4735 => x"81",
          4736 => x"f6",
          4737 => x"ac",
          4738 => x"9d",
          4739 => x"c8",
          4740 => x"e3",
          4741 => x"ff",
          4742 => x"59",
          4743 => x"51",
          4744 => x"3f",
          4745 => x"c8",
          4746 => x"a6",
          4747 => x"ac",
          4748 => x"83",
          4749 => x"fe",
          4750 => x"81",
          4751 => x"ff",
          4752 => x"d8",
          4753 => x"0d",
          4754 => x"05",
          4755 => x"84",
          4756 => x"83",
          4757 => x"83",
          4758 => x"72",
          4759 => x"86",
          4760 => x"11",
          4761 => x"22",
          4762 => x"5c",
          4763 => x"05",
          4764 => x"ff",
          4765 => x"ce",
          4766 => x"51",
          4767 => x"72",
          4768 => x"e9",
          4769 => x"2e",
          4770 => x"75",
          4771 => x"b9",
          4772 => x"2e",
          4773 => x"75",
          4774 => x"d5",
          4775 => x"bc",
          4776 => x"f8",
          4777 => x"f9",
          4778 => x"29",
          4779 => x"54",
          4780 => x"16",
          4781 => x"a0",
          4782 => x"84",
          4783 => x"83",
          4784 => x"83",
          4785 => x"72",
          4786 => x"5a",
          4787 => x"75",
          4788 => x"18",
          4789 => x"f8",
          4790 => x"29",
          4791 => x"83",
          4792 => x"86",
          4793 => x"18",
          4794 => x"bc",
          4795 => x"ff",
          4796 => x"f6",
          4797 => x"f9",
          4798 => x"29",
          4799 => x"57",
          4800 => x"f8",
          4801 => x"98",
          4802 => x"81",
          4803 => x"ff",
          4804 => x"73",
          4805 => x"99",
          4806 => x"bd",
          4807 => x"81",
          4808 => x"17",
          4809 => x"f8",
          4810 => x"b7",
          4811 => x"72",
          4812 => x"38",
          4813 => x"33",
          4814 => x"2e",
          4815 => x"80",
          4816 => x"c8",
          4817 => x"0d",
          4818 => x"2e",
          4819 => x"8d",
          4820 => x"38",
          4821 => x"09",
          4822 => x"c1",
          4823 => x"81",
          4824 => x"3f",
          4825 => x"f8",
          4826 => x"be",
          4827 => x"fa",
          4828 => x"84",
          4829 => x"33",
          4830 => x"89",
          4831 => x"06",
          4832 => x"80",
          4833 => x"a0",
          4834 => x"3f",
          4835 => x"81",
          4836 => x"54",
          4837 => x"ff",
          4838 => x"52",
          4839 => x"a5",
          4840 => x"70",
          4841 => x"54",
          4842 => x"27",
          4843 => x"fa",
          4844 => x"f8",
          4845 => x"f2",
          4846 => x"83",
          4847 => x"3f",
          4848 => x"b9",
          4849 => x"3d",
          4850 => x"80",
          4851 => x"81",
          4852 => x"38",
          4853 => x"33",
          4854 => x"06",
          4855 => x"53",
          4856 => x"73",
          4857 => x"f8",
          4858 => x"52",
          4859 => x"d5",
          4860 => x"f9",
          4861 => x"ff",
          4862 => x"05",
          4863 => x"a5",
          4864 => x"72",
          4865 => x"34",
          4866 => x"80",
          4867 => x"f9",
          4868 => x"81",
          4869 => x"3f",
          4870 => x"80",
          4871 => x"ef",
          4872 => x"86",
          4873 => x"0d",
          4874 => x"05",
          4875 => x"c4",
          4876 => x"75",
          4877 => x"b8",
          4878 => x"2e",
          4879 => x"78",
          4880 => x"b5",
          4881 => x"24",
          4882 => x"78",
          4883 => x"b9",
          4884 => x"2e",
          4885 => x"84",
          4886 => x"83",
          4887 => x"83",
          4888 => x"72",
          4889 => x"58",
          4890 => x"b7",
          4891 => x"86",
          4892 => x"17",
          4893 => x"bc",
          4894 => x"f9",
          4895 => x"f6",
          4896 => x"29",
          4897 => x"42",
          4898 => x"f8",
          4899 => x"83",
          4900 => x"60",
          4901 => x"05",
          4902 => x"f8",
          4903 => x"86",
          4904 => x"05",
          4905 => x"bc",
          4906 => x"ff",
          4907 => x"f6",
          4908 => x"f9",
          4909 => x"29",
          4910 => x"5d",
          4911 => x"f8",
          4912 => x"98",
          4913 => x"81",
          4914 => x"ff",
          4915 => x"76",
          4916 => x"b8",
          4917 => x"bd",
          4918 => x"86",
          4919 => x"19",
          4920 => x"f8",
          4921 => x"0b",
          4922 => x"0c",
          4923 => x"04",
          4924 => x"84",
          4925 => x"79",
          4926 => x"38",
          4927 => x"9b",
          4928 => x"80",
          4929 => x"cc",
          4930 => x"84",
          4931 => x"84",
          4932 => x"83",
          4933 => x"83",
          4934 => x"72",
          4935 => x"5e",
          4936 => x"b7",
          4937 => x"86",
          4938 => x"1d",
          4939 => x"bc",
          4940 => x"f9",
          4941 => x"f6",
          4942 => x"29",
          4943 => x"59",
          4944 => x"f8",
          4945 => x"83",
          4946 => x"76",
          4947 => x"5b",
          4948 => x"f4",
          4949 => x"b0",
          4950 => x"84",
          4951 => x"70",
          4952 => x"83",
          4953 => x"83",
          4954 => x"72",
          4955 => x"44",
          4956 => x"59",
          4957 => x"33",
          4958 => x"9a",
          4959 => x"1f",
          4960 => x"ff",
          4961 => x"77",
          4962 => x"38",
          4963 => x"f9",
          4964 => x"84",
          4965 => x"9c",
          4966 => x"78",
          4967 => x"b7",
          4968 => x"24",
          4969 => x"78",
          4970 => x"81",
          4971 => x"38",
          4972 => x"f8",
          4973 => x"0b",
          4974 => x"0c",
          4975 => x"04",
          4976 => x"82",
          4977 => x"19",
          4978 => x"26",
          4979 => x"84",
          4980 => x"81",
          4981 => x"77",
          4982 => x"34",
          4983 => x"cc",
          4984 => x"81",
          4985 => x"80",
          4986 => x"cc",
          4987 => x"0b",
          4988 => x"0c",
          4989 => x"04",
          4990 => x"fd",
          4991 => x"0b",
          4992 => x"0c",
          4993 => x"33",
          4994 => x"33",
          4995 => x"33",
          4996 => x"05",
          4997 => x"84",
          4998 => x"33",
          4999 => x"80",
          5000 => x"b7",
          5001 => x"f8",
          5002 => x"f8",
          5003 => x"71",
          5004 => x"5f",
          5005 => x"83",
          5006 => x"34",
          5007 => x"33",
          5008 => x"19",
          5009 => x"f8",
          5010 => x"a7",
          5011 => x"34",
          5012 => x"33",
          5013 => x"06",
          5014 => x"22",
          5015 => x"33",
          5016 => x"11",
          5017 => x"58",
          5018 => x"f4",
          5019 => x"98",
          5020 => x"81",
          5021 => x"89",
          5022 => x"81",
          5023 => x"3f",
          5024 => x"f8",
          5025 => x"ae",
          5026 => x"bc",
          5027 => x"f9",
          5028 => x"ff",
          5029 => x"f8",
          5030 => x"29",
          5031 => x"a0",
          5032 => x"f8",
          5033 => x"51",
          5034 => x"29",
          5035 => x"ff",
          5036 => x"f7",
          5037 => x"51",
          5038 => x"75",
          5039 => x"a4",
          5040 => x"ff",
          5041 => x"57",
          5042 => x"95",
          5043 => x"75",
          5044 => x"34",
          5045 => x"80",
          5046 => x"c8",
          5047 => x"84",
          5048 => x"80",
          5049 => x"ca",
          5050 => x"84",
          5051 => x"81",
          5052 => x"c4",
          5053 => x"84",
          5054 => x"9c",
          5055 => x"83",
          5056 => x"84",
          5057 => x"83",
          5058 => x"84",
          5059 => x"83",
          5060 => x"84",
          5061 => x"80",
          5062 => x"c4",
          5063 => x"84",
          5064 => x"9c",
          5065 => x"78",
          5066 => x"09",
          5067 => x"a7",
          5068 => x"f8",
          5069 => x"bc",
          5070 => x"ff",
          5071 => x"f9",
          5072 => x"ff",
          5073 => x"29",
          5074 => x"a0",
          5075 => x"f8",
          5076 => x"40",
          5077 => x"05",
          5078 => x"ff",
          5079 => x"ce",
          5080 => x"43",
          5081 => x"5c",
          5082 => x"85",
          5083 => x"81",
          5084 => x"1a",
          5085 => x"83",
          5086 => x"76",
          5087 => x"34",
          5088 => x"06",
          5089 => x"06",
          5090 => x"06",
          5091 => x"05",
          5092 => x"84",
          5093 => x"86",
          5094 => x"1e",
          5095 => x"bc",
          5096 => x"f9",
          5097 => x"f6",
          5098 => x"29",
          5099 => x"42",
          5100 => x"83",
          5101 => x"34",
          5102 => x"33",
          5103 => x"62",
          5104 => x"83",
          5105 => x"86",
          5106 => x"1a",
          5107 => x"bc",
          5108 => x"ff",
          5109 => x"f6",
          5110 => x"f9",
          5111 => x"29",
          5112 => x"5a",
          5113 => x"f8",
          5114 => x"84",
          5115 => x"34",
          5116 => x"81",
          5117 => x"58",
          5118 => x"95",
          5119 => x"b7",
          5120 => x"79",
          5121 => x"ff",
          5122 => x"83",
          5123 => x"83",
          5124 => x"70",
          5125 => x"58",
          5126 => x"fd",
          5127 => x"bb",
          5128 => x"38",
          5129 => x"83",
          5130 => x"bf",
          5131 => x"38",
          5132 => x"33",
          5133 => x"f9",
          5134 => x"19",
          5135 => x"26",
          5136 => x"75",
          5137 => x"c5",
          5138 => x"77",
          5139 => x"0b",
          5140 => x"34",
          5141 => x"51",
          5142 => x"80",
          5143 => x"c8",
          5144 => x"0d",
          5145 => x"f8",
          5146 => x"bc",
          5147 => x"ff",
          5148 => x"f9",
          5149 => x"ff",
          5150 => x"29",
          5151 => x"a0",
          5152 => x"f8",
          5153 => x"41",
          5154 => x"05",
          5155 => x"ff",
          5156 => x"ce",
          5157 => x"45",
          5158 => x"5b",
          5159 => x"82",
          5160 => x"5c",
          5161 => x"06",
          5162 => x"06",
          5163 => x"06",
          5164 => x"05",
          5165 => x"84",
          5166 => x"86",
          5167 => x"1b",
          5168 => x"bc",
          5169 => x"f9",
          5170 => x"f6",
          5171 => x"29",
          5172 => x"5e",
          5173 => x"83",
          5174 => x"34",
          5175 => x"33",
          5176 => x"1e",
          5177 => x"f8",
          5178 => x"a7",
          5179 => x"34",
          5180 => x"33",
          5181 => x"06",
          5182 => x"22",
          5183 => x"33",
          5184 => x"11",
          5185 => x"40",
          5186 => x"f4",
          5187 => x"9a",
          5188 => x"81",
          5189 => x"ff",
          5190 => x"7e",
          5191 => x"ac",
          5192 => x"bd",
          5193 => x"92",
          5194 => x"19",
          5195 => x"f8",
          5196 => x"1c",
          5197 => x"06",
          5198 => x"83",
          5199 => x"38",
          5200 => x"33",
          5201 => x"33",
          5202 => x"33",
          5203 => x"06",
          5204 => x"06",
          5205 => x"06",
          5206 => x"05",
          5207 => x"5b",
          5208 => x"b7",
          5209 => x"a7",
          5210 => x"34",
          5211 => x"33",
          5212 => x"33",
          5213 => x"22",
          5214 => x"12",
          5215 => x"56",
          5216 => x"f8",
          5217 => x"83",
          5218 => x"76",
          5219 => x"5a",
          5220 => x"f4",
          5221 => x"b0",
          5222 => x"84",
          5223 => x"70",
          5224 => x"83",
          5225 => x"83",
          5226 => x"72",
          5227 => x"5b",
          5228 => x"59",
          5229 => x"33",
          5230 => x"18",
          5231 => x"05",
          5232 => x"06",
          5233 => x"7f",
          5234 => x"38",
          5235 => x"f9",
          5236 => x"39",
          5237 => x"b8",
          5238 => x"0b",
          5239 => x"0c",
          5240 => x"04",
          5241 => x"17",
          5242 => x"b7",
          5243 => x"7a",
          5244 => x"f9",
          5245 => x"ff",
          5246 => x"05",
          5247 => x"39",
          5248 => x"b8",
          5249 => x"0b",
          5250 => x"0c",
          5251 => x"04",
          5252 => x"17",
          5253 => x"b7",
          5254 => x"7c",
          5255 => x"f8",
          5256 => x"bc",
          5257 => x"f9",
          5258 => x"5b",
          5259 => x"f4",
          5260 => x"cc",
          5261 => x"dc",
          5262 => x"05",
          5263 => x"c7",
          5264 => x"c8",
          5265 => x"fb",
          5266 => x"b8",
          5267 => x"11",
          5268 => x"84",
          5269 => x"79",
          5270 => x"06",
          5271 => x"ca",
          5272 => x"84",
          5273 => x"23",
          5274 => x"83",
          5275 => x"33",
          5276 => x"c4",
          5277 => x"34",
          5278 => x"33",
          5279 => x"33",
          5280 => x"33",
          5281 => x"f9",
          5282 => x"b7",
          5283 => x"f8",
          5284 => x"f8",
          5285 => x"72",
          5286 => x"5d",
          5287 => x"c4",
          5288 => x"86",
          5289 => x"05",
          5290 => x"bc",
          5291 => x"f9",
          5292 => x"f6",
          5293 => x"29",
          5294 => x"5b",
          5295 => x"f8",
          5296 => x"83",
          5297 => x"76",
          5298 => x"41",
          5299 => x"f4",
          5300 => x"a7",
          5301 => x"34",
          5302 => x"33",
          5303 => x"06",
          5304 => x"22",
          5305 => x"33",
          5306 => x"11",
          5307 => x"42",
          5308 => x"f4",
          5309 => x"9a",
          5310 => x"1c",
          5311 => x"06",
          5312 => x"7b",
          5313 => x"38",
          5314 => x"33",
          5315 => x"e2",
          5316 => x"56",
          5317 => x"f9",
          5318 => x"84",
          5319 => x"84",
          5320 => x"40",
          5321 => x"f3",
          5322 => x"b7",
          5323 => x"75",
          5324 => x"78",
          5325 => x"ea",
          5326 => x"0b",
          5327 => x"0c",
          5328 => x"04",
          5329 => x"33",
          5330 => x"34",
          5331 => x"33",
          5332 => x"34",
          5333 => x"33",
          5334 => x"f8",
          5335 => x"b9",
          5336 => x"f8",
          5337 => x"b0",
          5338 => x"f9",
          5339 => x"b1",
          5340 => x"f7",
          5341 => x"b2",
          5342 => x"39",
          5343 => x"33",
          5344 => x"2e",
          5345 => x"84",
          5346 => x"5d",
          5347 => x"09",
          5348 => x"85",
          5349 => x"f9",
          5350 => x"55",
          5351 => x"33",
          5352 => x"9b",
          5353 => x"84",
          5354 => x"70",
          5355 => x"ed",
          5356 => x"51",
          5357 => x"3f",
          5358 => x"08",
          5359 => x"83",
          5360 => x"57",
          5361 => x"60",
          5362 => x"cd",
          5363 => x"83",
          5364 => x"fe",
          5365 => x"fe",
          5366 => x"0b",
          5367 => x"33",
          5368 => x"81",
          5369 => x"77",
          5370 => x"ad",
          5371 => x"84",
          5372 => x"81",
          5373 => x"41",
          5374 => x"8a",
          5375 => x"10",
          5376 => x"a4",
          5377 => x"08",
          5378 => x"c9",
          5379 => x"80",
          5380 => x"38",
          5381 => x"33",
          5382 => x"33",
          5383 => x"70",
          5384 => x"2c",
          5385 => x"42",
          5386 => x"75",
          5387 => x"34",
          5388 => x"84",
          5389 => x"56",
          5390 => x"8e",
          5391 => x"b9",
          5392 => x"05",
          5393 => x"06",
          5394 => x"33",
          5395 => x"75",
          5396 => x"c5",
          5397 => x"f8",
          5398 => x"bd",
          5399 => x"83",
          5400 => x"83",
          5401 => x"70",
          5402 => x"5d",
          5403 => x"2e",
          5404 => x"ff",
          5405 => x"83",
          5406 => x"fd",
          5407 => x"0b",
          5408 => x"34",
          5409 => x"33",
          5410 => x"33",
          5411 => x"57",
          5412 => x"fd",
          5413 => x"17",
          5414 => x"f8",
          5415 => x"f9",
          5416 => x"c9",
          5417 => x"80",
          5418 => x"38",
          5419 => x"33",
          5420 => x"33",
          5421 => x"70",
          5422 => x"2c",
          5423 => x"41",
          5424 => x"75",
          5425 => x"34",
          5426 => x"84",
          5427 => x"5b",
          5428 => x"fc",
          5429 => x"b9",
          5430 => x"60",
          5431 => x"81",
          5432 => x"38",
          5433 => x"33",
          5434 => x"33",
          5435 => x"33",
          5436 => x"12",
          5437 => x"80",
          5438 => x"f6",
          5439 => x"5a",
          5440 => x"29",
          5441 => x"ff",
          5442 => x"f7",
          5443 => x"ff",
          5444 => x"42",
          5445 => x"7e",
          5446 => x"2e",
          5447 => x"80",
          5448 => x"cd",
          5449 => x"39",
          5450 => x"33",
          5451 => x"2e",
          5452 => x"84",
          5453 => x"58",
          5454 => x"09",
          5455 => x"d9",
          5456 => x"83",
          5457 => x"fb",
          5458 => x"b8",
          5459 => x"75",
          5460 => x"be",
          5461 => x"9d",
          5462 => x"f9",
          5463 => x"05",
          5464 => x"33",
          5465 => x"5e",
          5466 => x"25",
          5467 => x"57",
          5468 => x"f9",
          5469 => x"39",
          5470 => x"33",
          5471 => x"2e",
          5472 => x"84",
          5473 => x"83",
          5474 => x"42",
          5475 => x"b7",
          5476 => x"11",
          5477 => x"75",
          5478 => x"38",
          5479 => x"83",
          5480 => x"fa",
          5481 => x"e4",
          5482 => x"e8",
          5483 => x"0b",
          5484 => x"33",
          5485 => x"76",
          5486 => x"38",
          5487 => x"b9",
          5488 => x"22",
          5489 => x"e3",
          5490 => x"e8",
          5491 => x"17",
          5492 => x"06",
          5493 => x"33",
          5494 => x"da",
          5495 => x"84",
          5496 => x"5f",
          5497 => x"2e",
          5498 => x"b9",
          5499 => x"75",
          5500 => x"38",
          5501 => x"52",
          5502 => x"06",
          5503 => x"3f",
          5504 => x"84",
          5505 => x"57",
          5506 => x"8e",
          5507 => x"b9",
          5508 => x"05",
          5509 => x"06",
          5510 => x"33",
          5511 => x"81",
          5512 => x"b7",
          5513 => x"81",
          5514 => x"11",
          5515 => x"5b",
          5516 => x"77",
          5517 => x"38",
          5518 => x"83",
          5519 => x"76",
          5520 => x"ff",
          5521 => x"77",
          5522 => x"38",
          5523 => x"83",
          5524 => x"84",
          5525 => x"ff",
          5526 => x"7a",
          5527 => x"b4",
          5528 => x"75",
          5529 => x"34",
          5530 => x"84",
          5531 => x"5f",
          5532 => x"8a",
          5533 => x"b9",
          5534 => x"b7",
          5535 => x"5b",
          5536 => x"f9",
          5537 => x"f8",
          5538 => x"b7",
          5539 => x"81",
          5540 => x"f8",
          5541 => x"74",
          5542 => x"a7",
          5543 => x"83",
          5544 => x"5f",
          5545 => x"29",
          5546 => x"ff",
          5547 => x"f7",
          5548 => x"52",
          5549 => x"5d",
          5550 => x"84",
          5551 => x"83",
          5552 => x"70",
          5553 => x"57",
          5554 => x"8e",
          5555 => x"b7",
          5556 => x"76",
          5557 => x"d6",
          5558 => x"56",
          5559 => x"f6",
          5560 => x"ff",
          5561 => x"31",
          5562 => x"60",
          5563 => x"38",
          5564 => x"33",
          5565 => x"27",
          5566 => x"ff",
          5567 => x"83",
          5568 => x"7e",
          5569 => x"83",
          5570 => x"57",
          5571 => x"76",
          5572 => x"38",
          5573 => x"81",
          5574 => x"ff",
          5575 => x"29",
          5576 => x"79",
          5577 => x"a0",
          5578 => x"a7",
          5579 => x"81",
          5580 => x"81",
          5581 => x"71",
          5582 => x"58",
          5583 => x"7f",
          5584 => x"38",
          5585 => x"1a",
          5586 => x"17",
          5587 => x"b7",
          5588 => x"7b",
          5589 => x"5d",
          5590 => x"81",
          5591 => x"7c",
          5592 => x"5e",
          5593 => x"84",
          5594 => x"84",
          5595 => x"71",
          5596 => x"43",
          5597 => x"77",
          5598 => x"9d",
          5599 => x"17",
          5600 => x"b7",
          5601 => x"7b",
          5602 => x"5d",
          5603 => x"81",
          5604 => x"7c",
          5605 => x"5e",
          5606 => x"84",
          5607 => x"84",
          5608 => x"71",
          5609 => x"43",
          5610 => x"7f",
          5611 => x"99",
          5612 => x"39",
          5613 => x"33",
          5614 => x"2e",
          5615 => x"80",
          5616 => x"9d",
          5617 => x"b1",
          5618 => x"39",
          5619 => x"b7",
          5620 => x"11",
          5621 => x"33",
          5622 => x"58",
          5623 => x"94",
          5624 => x"9c",
          5625 => x"78",
          5626 => x"06",
          5627 => x"83",
          5628 => x"58",
          5629 => x"06",
          5630 => x"33",
          5631 => x"5c",
          5632 => x"81",
          5633 => x"b7",
          5634 => x"7a",
          5635 => x"89",
          5636 => x"ff",
          5637 => x"76",
          5638 => x"38",
          5639 => x"61",
          5640 => x"57",
          5641 => x"38",
          5642 => x"1b",
          5643 => x"62",
          5644 => x"a0",
          5645 => x"1f",
          5646 => x"a7",
          5647 => x"79",
          5648 => x"51",
          5649 => x"ac",
          5650 => x"06",
          5651 => x"a4",
          5652 => x"f4",
          5653 => x"2b",
          5654 => x"07",
          5655 => x"07",
          5656 => x"7f",
          5657 => x"57",
          5658 => x"9e",
          5659 => x"70",
          5660 => x"0c",
          5661 => x"84",
          5662 => x"79",
          5663 => x"38",
          5664 => x"33",
          5665 => x"33",
          5666 => x"81",
          5667 => x"81",
          5668 => x"f8",
          5669 => x"73",
          5670 => x"59",
          5671 => x"77",
          5672 => x"38",
          5673 => x"1b",
          5674 => x"62",
          5675 => x"75",
          5676 => x"57",
          5677 => x"f4",
          5678 => x"f8",
          5679 => x"98",
          5680 => x"5a",
          5681 => x"e0",
          5682 => x"78",
          5683 => x"5a",
          5684 => x"57",
          5685 => x"f4",
          5686 => x"0b",
          5687 => x"34",
          5688 => x"81",
          5689 => x"81",
          5690 => x"77",
          5691 => x"f4",
          5692 => x"1f",
          5693 => x"06",
          5694 => x"8a",
          5695 => x"f4",
          5696 => x"f0",
          5697 => x"2b",
          5698 => x"71",
          5699 => x"58",
          5700 => x"80",
          5701 => x"81",
          5702 => x"80",
          5703 => x"f8",
          5704 => x"18",
          5705 => x"06",
          5706 => x"b6",
          5707 => x"fa",
          5708 => x"84",
          5709 => x"33",
          5710 => x"f8",
          5711 => x"b7",
          5712 => x"f8",
          5713 => x"b7",
          5714 => x"5c",
          5715 => x"ee",
          5716 => x"f4",
          5717 => x"56",
          5718 => x"f4",
          5719 => x"70",
          5720 => x"59",
          5721 => x"39",
          5722 => x"33",
          5723 => x"85",
          5724 => x"83",
          5725 => x"e5",
          5726 => x"f4",
          5727 => x"06",
          5728 => x"75",
          5729 => x"34",
          5730 => x"f8",
          5731 => x"f9",
          5732 => x"56",
          5733 => x"f4",
          5734 => x"83",
          5735 => x"81",
          5736 => x"07",
          5737 => x"f8",
          5738 => x"b1",
          5739 => x"0b",
          5740 => x"34",
          5741 => x"81",
          5742 => x"56",
          5743 => x"83",
          5744 => x"81",
          5745 => x"75",
          5746 => x"34",
          5747 => x"83",
          5748 => x"81",
          5749 => x"07",
          5750 => x"f8",
          5751 => x"fd",
          5752 => x"f4",
          5753 => x"06",
          5754 => x"56",
          5755 => x"f4",
          5756 => x"39",
          5757 => x"33",
          5758 => x"80",
          5759 => x"75",
          5760 => x"34",
          5761 => x"83",
          5762 => x"81",
          5763 => x"07",
          5764 => x"f8",
          5765 => x"c5",
          5766 => x"f4",
          5767 => x"06",
          5768 => x"75",
          5769 => x"34",
          5770 => x"83",
          5771 => x"81",
          5772 => x"07",
          5773 => x"f8",
          5774 => x"a1",
          5775 => x"f4",
          5776 => x"06",
          5777 => x"75",
          5778 => x"34",
          5779 => x"83",
          5780 => x"81",
          5781 => x"75",
          5782 => x"34",
          5783 => x"83",
          5784 => x"80",
          5785 => x"75",
          5786 => x"34",
          5787 => x"83",
          5788 => x"80",
          5789 => x"75",
          5790 => x"34",
          5791 => x"83",
          5792 => x"81",
          5793 => x"d0",
          5794 => x"83",
          5795 => x"fd",
          5796 => x"f8",
          5797 => x"bf",
          5798 => x"56",
          5799 => x"f4",
          5800 => x"39",
          5801 => x"f8",
          5802 => x"52",
          5803 => x"c9",
          5804 => x"39",
          5805 => x"33",
          5806 => x"34",
          5807 => x"33",
          5808 => x"34",
          5809 => x"33",
          5810 => x"f8",
          5811 => x"0b",
          5812 => x"0c",
          5813 => x"81",
          5814 => x"cb",
          5815 => x"84",
          5816 => x"9c",
          5817 => x"77",
          5818 => x"34",
          5819 => x"33",
          5820 => x"06",
          5821 => x"56",
          5822 => x"84",
          5823 => x"9c",
          5824 => x"53",
          5825 => x"fe",
          5826 => x"84",
          5827 => x"a1",
          5828 => x"c8",
          5829 => x"c4",
          5830 => x"84",
          5831 => x"80",
          5832 => x"c8",
          5833 => x"0d",
          5834 => x"f8",
          5835 => x"e9",
          5836 => x"c9",
          5837 => x"5c",
          5838 => x"b8",
          5839 => x"10",
          5840 => x"5d",
          5841 => x"05",
          5842 => x"9c",
          5843 => x"0b",
          5844 => x"34",
          5845 => x"0b",
          5846 => x"34",
          5847 => x"51",
          5848 => x"83",
          5849 => x"70",
          5850 => x"58",
          5851 => x"e6",
          5852 => x"0b",
          5853 => x"34",
          5854 => x"51",
          5855 => x"ef",
          5856 => x"51",
          5857 => x"3f",
          5858 => x"83",
          5859 => x"ff",
          5860 => x"70",
          5861 => x"06",
          5862 => x"f2",
          5863 => x"52",
          5864 => x"39",
          5865 => x"33",
          5866 => x"27",
          5867 => x"75",
          5868 => x"34",
          5869 => x"83",
          5870 => x"ff",
          5871 => x"70",
          5872 => x"06",
          5873 => x"f0",
          5874 => x"f8",
          5875 => x"05",
          5876 => x"33",
          5877 => x"59",
          5878 => x"25",
          5879 => x"75",
          5880 => x"39",
          5881 => x"33",
          5882 => x"06",
          5883 => x"77",
          5884 => x"38",
          5885 => x"33",
          5886 => x"33",
          5887 => x"06",
          5888 => x"33",
          5889 => x"11",
          5890 => x"80",
          5891 => x"f6",
          5892 => x"71",
          5893 => x"70",
          5894 => x"06",
          5895 => x"33",
          5896 => x"42",
          5897 => x"81",
          5898 => x"38",
          5899 => x"ff",
          5900 => x"5c",
          5901 => x"24",
          5902 => x"84",
          5903 => x"56",
          5904 => x"83",
          5905 => x"16",
          5906 => x"f8",
          5907 => x"81",
          5908 => x"11",
          5909 => x"76",
          5910 => x"38",
          5911 => x"33",
          5912 => x"27",
          5913 => x"ff",
          5914 => x"83",
          5915 => x"7b",
          5916 => x"83",
          5917 => x"57",
          5918 => x"76",
          5919 => x"38",
          5920 => x"81",
          5921 => x"ff",
          5922 => x"29",
          5923 => x"79",
          5924 => x"a0",
          5925 => x"a7",
          5926 => x"81",
          5927 => x"81",
          5928 => x"71",
          5929 => x"42",
          5930 => x"7e",
          5931 => x"38",
          5932 => x"1a",
          5933 => x"17",
          5934 => x"b7",
          5935 => x"7b",
          5936 => x"5d",
          5937 => x"81",
          5938 => x"7d",
          5939 => x"5f",
          5940 => x"84",
          5941 => x"84",
          5942 => x"71",
          5943 => x"59",
          5944 => x"77",
          5945 => x"b1",
          5946 => x"17",
          5947 => x"b7",
          5948 => x"7b",
          5949 => x"5d",
          5950 => x"81",
          5951 => x"7d",
          5952 => x"5f",
          5953 => x"84",
          5954 => x"84",
          5955 => x"71",
          5956 => x"59",
          5957 => x"75",
          5958 => x"99",
          5959 => x"39",
          5960 => x"17",
          5961 => x"b7",
          5962 => x"7b",
          5963 => x"f8",
          5964 => x"bc",
          5965 => x"f6",
          5966 => x"bb",
          5967 => x"5f",
          5968 => x"39",
          5969 => x"38",
          5970 => x"33",
          5971 => x"06",
          5972 => x"42",
          5973 => x"27",
          5974 => x"5a",
          5975 => x"f6",
          5976 => x"ff",
          5977 => x"58",
          5978 => x"27",
          5979 => x"57",
          5980 => x"f8",
          5981 => x"bc",
          5982 => x"ff",
          5983 => x"52",
          5984 => x"78",
          5985 => x"38",
          5986 => x"83",
          5987 => x"eb",
          5988 => x"f8",
          5989 => x"05",
          5990 => x"33",
          5991 => x"40",
          5992 => x"25",
          5993 => x"75",
          5994 => x"39",
          5995 => x"09",
          5996 => x"c0",
          5997 => x"f9",
          5998 => x"ff",
          5999 => x"f8",
          6000 => x"5d",
          6001 => x"ff",
          6002 => x"06",
          6003 => x"f6",
          6004 => x"1d",
          6005 => x"f8",
          6006 => x"93",
          6007 => x"56",
          6008 => x"f6",
          6009 => x"39",
          6010 => x"56",
          6011 => x"f8",
          6012 => x"39",
          6013 => x"56",
          6014 => x"f5",
          6015 => x"76",
          6016 => x"58",
          6017 => x"f4",
          6018 => x"81",
          6019 => x"75",
          6020 => x"ec",
          6021 => x"70",
          6022 => x"34",
          6023 => x"33",
          6024 => x"05",
          6025 => x"76",
          6026 => x"f4",
          6027 => x"7b",
          6028 => x"83",
          6029 => x"f1",
          6030 => x"0b",
          6031 => x"34",
          6032 => x"7e",
          6033 => x"23",
          6034 => x"80",
          6035 => x"f6",
          6036 => x"39",
          6037 => x"f8",
          6038 => x"a7",
          6039 => x"fa",
          6040 => x"84",
          6041 => x"33",
          6042 => x"0b",
          6043 => x"34",
          6044 => x"fd",
          6045 => x"97",
          6046 => x"b7",
          6047 => x"54",
          6048 => x"90",
          6049 => x"db",
          6050 => x"0b",
          6051 => x"0c",
          6052 => x"04",
          6053 => x"51",
          6054 => x"80",
          6055 => x"c8",
          6056 => x"0d",
          6057 => x"0d",
          6058 => x"33",
          6059 => x"83",
          6060 => x"70",
          6061 => x"83",
          6062 => x"33",
          6063 => x"59",
          6064 => x"80",
          6065 => x"14",
          6066 => x"f7",
          6067 => x"59",
          6068 => x"c8",
          6069 => x"0d",
          6070 => x"a8",
          6071 => x"53",
          6072 => x"91",
          6073 => x"32",
          6074 => x"07",
          6075 => x"9f",
          6076 => x"5e",
          6077 => x"f7",
          6078 => x"59",
          6079 => x"81",
          6080 => x"06",
          6081 => x"54",
          6082 => x"70",
          6083 => x"25",
          6084 => x"5c",
          6085 => x"2e",
          6086 => x"84",
          6087 => x"83",
          6088 => x"83",
          6089 => x"72",
          6090 => x"86",
          6091 => x"05",
          6092 => x"22",
          6093 => x"71",
          6094 => x"70",
          6095 => x"06",
          6096 => x"33",
          6097 => x"58",
          6098 => x"83",
          6099 => x"f0",
          6100 => x"8e",
          6101 => x"80",
          6102 => x"98",
          6103 => x"c0",
          6104 => x"56",
          6105 => x"f6",
          6106 => x"80",
          6107 => x"76",
          6108 => x"15",
          6109 => x"70",
          6110 => x"55",
          6111 => x"74",
          6112 => x"80",
          6113 => x"e8",
          6114 => x"81",
          6115 => x"f6",
          6116 => x"58",
          6117 => x"76",
          6118 => x"38",
          6119 => x"2e",
          6120 => x"74",
          6121 => x"15",
          6122 => x"ff",
          6123 => x"81",
          6124 => x"cd",
          6125 => x"f7",
          6126 => x"83",
          6127 => x"33",
          6128 => x"15",
          6129 => x"70",
          6130 => x"55",
          6131 => x"27",
          6132 => x"83",
          6133 => x"70",
          6134 => x"80",
          6135 => x"54",
          6136 => x"a0",
          6137 => x"ff",
          6138 => x"2a",
          6139 => x"81",
          6140 => x"58",
          6141 => x"85",
          6142 => x"0b",
          6143 => x"34",
          6144 => x"06",
          6145 => x"2e",
          6146 => x"81",
          6147 => x"a2",
          6148 => x"83",
          6149 => x"83",
          6150 => x"83",
          6151 => x"70",
          6152 => x"33",
          6153 => x"33",
          6154 => x"5e",
          6155 => x"83",
          6156 => x"33",
          6157 => x"ff",
          6158 => x"83",
          6159 => x"33",
          6160 => x"2e",
          6161 => x"83",
          6162 => x"33",
          6163 => x"ff",
          6164 => x"83",
          6165 => x"33",
          6166 => x"ec",
          6167 => x"ff",
          6168 => x"81",
          6169 => x"38",
          6170 => x"16",
          6171 => x"81",
          6172 => x"38",
          6173 => x"06",
          6174 => x"ff",
          6175 => x"38",
          6176 => x"16",
          6177 => x"74",
          6178 => x"38",
          6179 => x"08",
          6180 => x"87",
          6181 => x"08",
          6182 => x"73",
          6183 => x"38",
          6184 => x"c0",
          6185 => x"83",
          6186 => x"58",
          6187 => x"81",
          6188 => x"54",
          6189 => x"fe",
          6190 => x"83",
          6191 => x"77",
          6192 => x"34",
          6193 => x"53",
          6194 => x"82",
          6195 => x"10",
          6196 => x"ec",
          6197 => x"08",
          6198 => x"d0",
          6199 => x"80",
          6200 => x"83",
          6201 => x"c0",
          6202 => x"5e",
          6203 => x"27",
          6204 => x"80",
          6205 => x"ce",
          6206 => x"72",
          6207 => x"38",
          6208 => x"83",
          6209 => x"87",
          6210 => x"08",
          6211 => x"0c",
          6212 => x"06",
          6213 => x"2e",
          6214 => x"f8",
          6215 => x"54",
          6216 => x"14",
          6217 => x"81",
          6218 => x"a5",
          6219 => x"a8",
          6220 => x"80",
          6221 => x"38",
          6222 => x"83",
          6223 => x"c3",
          6224 => x"f0",
          6225 => x"39",
          6226 => x"e0",
          6227 => x"56",
          6228 => x"7c",
          6229 => x"38",
          6230 => x"09",
          6231 => x"b4",
          6232 => x"2e",
          6233 => x"79",
          6234 => x"d7",
          6235 => x"ff",
          6236 => x"77",
          6237 => x"2b",
          6238 => x"80",
          6239 => x"73",
          6240 => x"38",
          6241 => x"81",
          6242 => x"10",
          6243 => x"87",
          6244 => x"98",
          6245 => x"57",
          6246 => x"73",
          6247 => x"78",
          6248 => x"79",
          6249 => x"11",
          6250 => x"05",
          6251 => x"05",
          6252 => x"56",
          6253 => x"c0",
          6254 => x"83",
          6255 => x"57",
          6256 => x"80",
          6257 => x"2e",
          6258 => x"79",
          6259 => x"59",
          6260 => x"82",
          6261 => x"39",
          6262 => x"fa",
          6263 => x"0b",
          6264 => x"33",
          6265 => x"81",
          6266 => x"38",
          6267 => x"70",
          6268 => x"25",
          6269 => x"59",
          6270 => x"38",
          6271 => x"09",
          6272 => x"cc",
          6273 => x"2e",
          6274 => x"80",
          6275 => x"10",
          6276 => x"d4",
          6277 => x"5d",
          6278 => x"2e",
          6279 => x"81",
          6280 => x"ff",
          6281 => x"93",
          6282 => x"38",
          6283 => x"33",
          6284 => x"2e",
          6285 => x"84",
          6286 => x"55",
          6287 => x"38",
          6288 => x"06",
          6289 => x"cc",
          6290 => x"84",
          6291 => x"8f",
          6292 => x"be",
          6293 => x"f0",
          6294 => x"39",
          6295 => x"2e",
          6296 => x"f7",
          6297 => x"81",
          6298 => x"83",
          6299 => x"34",
          6300 => x"80",
          6301 => x"90",
          6302 => x"0b",
          6303 => x"15",
          6304 => x"83",
          6305 => x"34",
          6306 => x"74",
          6307 => x"53",
          6308 => x"2e",
          6309 => x"83",
          6310 => x"33",
          6311 => x"27",
          6312 => x"77",
          6313 => x"54",
          6314 => x"09",
          6315 => x"fc",
          6316 => x"9c",
          6317 => x"05",
          6318 => x"9c",
          6319 => x"74",
          6320 => x"e8",
          6321 => x"98",
          6322 => x"f7",
          6323 => x"81",
          6324 => x"fb",
          6325 => x"0b",
          6326 => x"15",
          6327 => x"39",
          6328 => x"a1",
          6329 => x"81",
          6330 => x"fa",
          6331 => x"83",
          6332 => x"80",
          6333 => x"a1",
          6334 => x"a8",
          6335 => x"a2",
          6336 => x"f7",
          6337 => x"f7",
          6338 => x"5d",
          6339 => x"5e",
          6340 => x"39",
          6341 => x"09",
          6342 => x"cb",
          6343 => x"7a",
          6344 => x"ce",
          6345 => x"2e",
          6346 => x"fc",
          6347 => x"93",
          6348 => x"34",
          6349 => x"f8",
          6350 => x"0b",
          6351 => x"33",
          6352 => x"83",
          6353 => x"73",
          6354 => x"34",
          6355 => x"ac",
          6356 => x"84",
          6357 => x"58",
          6358 => x"38",
          6359 => x"84",
          6360 => x"ff",
          6361 => x"39",
          6362 => x"f7",
          6363 => x"2e",
          6364 => x"84",
          6365 => x"a8",
          6366 => x"39",
          6367 => x"33",
          6368 => x"06",
          6369 => x"5a",
          6370 => x"27",
          6371 => x"55",
          6372 => x"f6",
          6373 => x"ff",
          6374 => x"55",
          6375 => x"27",
          6376 => x"54",
          6377 => x"f8",
          6378 => x"bc",
          6379 => x"ff",
          6380 => x"05",
          6381 => x"27",
          6382 => x"53",
          6383 => x"f9",
          6384 => x"f6",
          6385 => x"52",
          6386 => x"ba",
          6387 => x"59",
          6388 => x"72",
          6389 => x"39",
          6390 => x"52",
          6391 => x"51",
          6392 => x"3f",
          6393 => x"f7",
          6394 => x"f7",
          6395 => x"fc",
          6396 => x"3d",
          6397 => x"f5",
          6398 => x"3d",
          6399 => x"3d",
          6400 => x"83",
          6401 => x"53",
          6402 => x"05",
          6403 => x"34",
          6404 => x"08",
          6405 => x"71",
          6406 => x"83",
          6407 => x"55",
          6408 => x"81",
          6409 => x"0b",
          6410 => x"e8",
          6411 => x"98",
          6412 => x"f3",
          6413 => x"80",
          6414 => x"53",
          6415 => x"9c",
          6416 => x"c0",
          6417 => x"51",
          6418 => x"f6",
          6419 => x"33",
          6420 => x"9c",
          6421 => x"74",
          6422 => x"38",
          6423 => x"2e",
          6424 => x"c0",
          6425 => x"51",
          6426 => x"73",
          6427 => x"38",
          6428 => x"ff",
          6429 => x"38",
          6430 => x"9c",
          6431 => x"90",
          6432 => x"c0",
          6433 => x"52",
          6434 => x"9c",
          6435 => x"72",
          6436 => x"81",
          6437 => x"c0",
          6438 => x"52",
          6439 => x"27",
          6440 => x"81",
          6441 => x"38",
          6442 => x"a4",
          6443 => x"75",
          6444 => x"ff",
          6445 => x"ff",
          6446 => x"ff",
          6447 => x"75",
          6448 => x"38",
          6449 => x"06",
          6450 => x"d5",
          6451 => x"2e",
          6452 => x"84",
          6453 => x"88",
          6454 => x"81",
          6455 => x"c8",
          6456 => x"0d",
          6457 => x"0d",
          6458 => x"05",
          6459 => x"56",
          6460 => x"83",
          6461 => x"73",
          6462 => x"fc",
          6463 => x"70",
          6464 => x"07",
          6465 => x"57",
          6466 => x"34",
          6467 => x"51",
          6468 => x"34",
          6469 => x"56",
          6470 => x"34",
          6471 => x"34",
          6472 => x"08",
          6473 => x"13",
          6474 => x"d4",
          6475 => x"e1",
          6476 => x"0b",
          6477 => x"08",
          6478 => x"0b",
          6479 => x"80",
          6480 => x"80",
          6481 => x"c0",
          6482 => x"83",
          6483 => x"55",
          6484 => x"05",
          6485 => x"98",
          6486 => x"87",
          6487 => x"08",
          6488 => x"2e",
          6489 => x"14",
          6490 => x"98",
          6491 => x"52",
          6492 => x"87",
          6493 => x"fe",
          6494 => x"87",
          6495 => x"08",
          6496 => x"70",
          6497 => x"c8",
          6498 => x"71",
          6499 => x"c0",
          6500 => x"98",
          6501 => x"ce",
          6502 => x"87",
          6503 => x"08",
          6504 => x"98",
          6505 => x"74",
          6506 => x"38",
          6507 => x"87",
          6508 => x"08",
          6509 => x"73",
          6510 => x"71",
          6511 => x"db",
          6512 => x"98",
          6513 => x"72",
          6514 => x"38",
          6515 => x"55",
          6516 => x"81",
          6517 => x"53",
          6518 => x"80",
          6519 => x"81",
          6520 => x"71",
          6521 => x"74",
          6522 => x"ff",
          6523 => x"aa",
          6524 => x"14",
          6525 => x"11",
          6526 => x"70",
          6527 => x"38",
          6528 => x"05",
          6529 => x"70",
          6530 => x"34",
          6531 => x"f0",
          6532 => x"b9",
          6533 => x"3d",
          6534 => x"0b",
          6535 => x"0c",
          6536 => x"04",
          6537 => x"39",
          6538 => x"79",
          6539 => x"a3",
          6540 => x"56",
          6541 => x"f3",
          6542 => x"88",
          6543 => x"80",
          6544 => x"79",
          6545 => x"51",
          6546 => x"75",
          6547 => x"72",
          6548 => x"70",
          6549 => x"75",
          6550 => x"71",
          6551 => x"72",
          6552 => x"7a",
          6553 => x"08",
          6554 => x"84",
          6555 => x"54",
          6556 => x"73",
          6557 => x"70",
          6558 => x"52",
          6559 => x"81",
          6560 => x"72",
          6561 => x"38",
          6562 => x"08",
          6563 => x"15",
          6564 => x"d4",
          6565 => x"e2",
          6566 => x"0b",
          6567 => x"08",
          6568 => x"0b",
          6569 => x"80",
          6570 => x"80",
          6571 => x"c0",
          6572 => x"83",
          6573 => x"55",
          6574 => x"05",
          6575 => x"98",
          6576 => x"87",
          6577 => x"08",
          6578 => x"2e",
          6579 => x"14",
          6580 => x"98",
          6581 => x"52",
          6582 => x"87",
          6583 => x"fe",
          6584 => x"87",
          6585 => x"08",
          6586 => x"70",
          6587 => x"c8",
          6588 => x"71",
          6589 => x"c0",
          6590 => x"98",
          6591 => x"ce",
          6592 => x"87",
          6593 => x"08",
          6594 => x"98",
          6595 => x"74",
          6596 => x"38",
          6597 => x"87",
          6598 => x"08",
          6599 => x"73",
          6600 => x"71",
          6601 => x"db",
          6602 => x"98",
          6603 => x"72",
          6604 => x"38",
          6605 => x"55",
          6606 => x"81",
          6607 => x"53",
          6608 => x"a1",
          6609 => x"ff",
          6610 => x"fe",
          6611 => x"51",
          6612 => x"06",
          6613 => x"2e",
          6614 => x"57",
          6615 => x"c8",
          6616 => x"0d",
          6617 => x"e8",
          6618 => x"0d",
          6619 => x"08",
          6620 => x"71",
          6621 => x"83",
          6622 => x"56",
          6623 => x"81",
          6624 => x"0b",
          6625 => x"e8",
          6626 => x"98",
          6627 => x"f3",
          6628 => x"80",
          6629 => x"54",
          6630 => x"9c",
          6631 => x"c0",
          6632 => x"53",
          6633 => x"f6",
          6634 => x"33",
          6635 => x"9c",
          6636 => x"70",
          6637 => x"38",
          6638 => x"2e",
          6639 => x"c0",
          6640 => x"51",
          6641 => x"74",
          6642 => x"38",
          6643 => x"ff",
          6644 => x"38",
          6645 => x"9c",
          6646 => x"90",
          6647 => x"c0",
          6648 => x"52",
          6649 => x"9c",
          6650 => x"72",
          6651 => x"81",
          6652 => x"c0",
          6653 => x"55",
          6654 => x"27",
          6655 => x"81",
          6656 => x"38",
          6657 => x"a4",
          6658 => x"71",
          6659 => x"ff",
          6660 => x"ff",
          6661 => x"ff",
          6662 => x"75",
          6663 => x"38",
          6664 => x"06",
          6665 => x"d5",
          6666 => x"80",
          6667 => x"e4",
          6668 => x"d0",
          6669 => x"3d",
          6670 => x"3d",
          6671 => x"b8",
          6672 => x"31",
          6673 => x"83",
          6674 => x"70",
          6675 => x"11",
          6676 => x"12",
          6677 => x"2b",
          6678 => x"07",
          6679 => x"33",
          6680 => x"71",
          6681 => x"90",
          6682 => x"54",
          6683 => x"5d",
          6684 => x"56",
          6685 => x"71",
          6686 => x"38",
          6687 => x"11",
          6688 => x"33",
          6689 => x"71",
          6690 => x"76",
          6691 => x"81",
          6692 => x"98",
          6693 => x"2b",
          6694 => x"5c",
          6695 => x"52",
          6696 => x"83",
          6697 => x"13",
          6698 => x"33",
          6699 => x"71",
          6700 => x"75",
          6701 => x"2a",
          6702 => x"57",
          6703 => x"34",
          6704 => x"06",
          6705 => x"13",
          6706 => x"b8",
          6707 => x"84",
          6708 => x"13",
          6709 => x"2b",
          6710 => x"2a",
          6711 => x"54",
          6712 => x"14",
          6713 => x"14",
          6714 => x"b8",
          6715 => x"80",
          6716 => x"34",
          6717 => x"13",
          6718 => x"b8",
          6719 => x"84",
          6720 => x"85",
          6721 => x"b9",
          6722 => x"70",
          6723 => x"33",
          6724 => x"07",
          6725 => x"07",
          6726 => x"58",
          6727 => x"74",
          6728 => x"81",
          6729 => x"3d",
          6730 => x"12",
          6731 => x"33",
          6732 => x"71",
          6733 => x"75",
          6734 => x"33",
          6735 => x"71",
          6736 => x"70",
          6737 => x"58",
          6738 => x"58",
          6739 => x"12",
          6740 => x"12",
          6741 => x"b8",
          6742 => x"84",
          6743 => x"12",
          6744 => x"2b",
          6745 => x"07",
          6746 => x"52",
          6747 => x"12",
          6748 => x"33",
          6749 => x"07",
          6750 => x"52",
          6751 => x"77",
          6752 => x"72",
          6753 => x"84",
          6754 => x"15",
          6755 => x"12",
          6756 => x"2b",
          6757 => x"ff",
          6758 => x"2a",
          6759 => x"52",
          6760 => x"77",
          6761 => x"84",
          6762 => x"70",
          6763 => x"81",
          6764 => x"8b",
          6765 => x"2b",
          6766 => x"70",
          6767 => x"33",
          6768 => x"07",
          6769 => x"8f",
          6770 => x"77",
          6771 => x"2a",
          6772 => x"54",
          6773 => x"54",
          6774 => x"14",
          6775 => x"14",
          6776 => x"b8",
          6777 => x"70",
          6778 => x"33",
          6779 => x"71",
          6780 => x"74",
          6781 => x"81",
          6782 => x"88",
          6783 => x"ff",
          6784 => x"88",
          6785 => x"53",
          6786 => x"54",
          6787 => x"34",
          6788 => x"34",
          6789 => x"08",
          6790 => x"11",
          6791 => x"33",
          6792 => x"71",
          6793 => x"74",
          6794 => x"81",
          6795 => x"98",
          6796 => x"2b",
          6797 => x"5d",
          6798 => x"53",
          6799 => x"25",
          6800 => x"71",
          6801 => x"33",
          6802 => x"07",
          6803 => x"07",
          6804 => x"59",
          6805 => x"75",
          6806 => x"16",
          6807 => x"b8",
          6808 => x"70",
          6809 => x"33",
          6810 => x"71",
          6811 => x"74",
          6812 => x"33",
          6813 => x"71",
          6814 => x"70",
          6815 => x"5c",
          6816 => x"56",
          6817 => x"82",
          6818 => x"83",
          6819 => x"3d",
          6820 => x"3d",
          6821 => x"b9",
          6822 => x"58",
          6823 => x"8f",
          6824 => x"2e",
          6825 => x"51",
          6826 => x"89",
          6827 => x"84",
          6828 => x"84",
          6829 => x"a0",
          6830 => x"b9",
          6831 => x"80",
          6832 => x"52",
          6833 => x"51",
          6834 => x"3f",
          6835 => x"08",
          6836 => x"34",
          6837 => x"16",
          6838 => x"b8",
          6839 => x"84",
          6840 => x"0b",
          6841 => x"84",
          6842 => x"56",
          6843 => x"34",
          6844 => x"17",
          6845 => x"b8",
          6846 => x"b4",
          6847 => x"fe",
          6848 => x"70",
          6849 => x"06",
          6850 => x"58",
          6851 => x"74",
          6852 => x"73",
          6853 => x"84",
          6854 => x"70",
          6855 => x"84",
          6856 => x"05",
          6857 => x"55",
          6858 => x"34",
          6859 => x"15",
          6860 => x"39",
          6861 => x"7b",
          6862 => x"81",
          6863 => x"27",
          6864 => x"12",
          6865 => x"05",
          6866 => x"ff",
          6867 => x"70",
          6868 => x"06",
          6869 => x"08",
          6870 => x"85",
          6871 => x"88",
          6872 => x"52",
          6873 => x"55",
          6874 => x"54",
          6875 => x"80",
          6876 => x"10",
          6877 => x"70",
          6878 => x"33",
          6879 => x"07",
          6880 => x"ff",
          6881 => x"70",
          6882 => x"06",
          6883 => x"56",
          6884 => x"54",
          6885 => x"27",
          6886 => x"80",
          6887 => x"75",
          6888 => x"84",
          6889 => x"13",
          6890 => x"2b",
          6891 => x"75",
          6892 => x"81",
          6893 => x"85",
          6894 => x"54",
          6895 => x"83",
          6896 => x"70",
          6897 => x"33",
          6898 => x"07",
          6899 => x"ff",
          6900 => x"5d",
          6901 => x"70",
          6902 => x"38",
          6903 => x"51",
          6904 => x"82",
          6905 => x"51",
          6906 => x"82",
          6907 => x"75",
          6908 => x"38",
          6909 => x"83",
          6910 => x"74",
          6911 => x"07",
          6912 => x"5b",
          6913 => x"5a",
          6914 => x"78",
          6915 => x"84",
          6916 => x"15",
          6917 => x"53",
          6918 => x"14",
          6919 => x"14",
          6920 => x"b8",
          6921 => x"70",
          6922 => x"33",
          6923 => x"07",
          6924 => x"8f",
          6925 => x"74",
          6926 => x"ff",
          6927 => x"88",
          6928 => x"53",
          6929 => x"52",
          6930 => x"34",
          6931 => x"06",
          6932 => x"12",
          6933 => x"b8",
          6934 => x"75",
          6935 => x"81",
          6936 => x"b9",
          6937 => x"19",
          6938 => x"87",
          6939 => x"8b",
          6940 => x"2b",
          6941 => x"58",
          6942 => x"57",
          6943 => x"34",
          6944 => x"34",
          6945 => x"08",
          6946 => x"78",
          6947 => x"33",
          6948 => x"71",
          6949 => x"70",
          6950 => x"54",
          6951 => x"86",
          6952 => x"87",
          6953 => x"b9",
          6954 => x"19",
          6955 => x"85",
          6956 => x"8b",
          6957 => x"2b",
          6958 => x"58",
          6959 => x"52",
          6960 => x"34",
          6961 => x"34",
          6962 => x"08",
          6963 => x"78",
          6964 => x"33",
          6965 => x"71",
          6966 => x"70",
          6967 => x"5c",
          6968 => x"84",
          6969 => x"85",
          6970 => x"b9",
          6971 => x"84",
          6972 => x"84",
          6973 => x"8b",
          6974 => x"86",
          6975 => x"15",
          6976 => x"2b",
          6977 => x"07",
          6978 => x"17",
          6979 => x"33",
          6980 => x"07",
          6981 => x"5a",
          6982 => x"54",
          6983 => x"12",
          6984 => x"12",
          6985 => x"b8",
          6986 => x"84",
          6987 => x"12",
          6988 => x"2b",
          6989 => x"07",
          6990 => x"14",
          6991 => x"33",
          6992 => x"07",
          6993 => x"58",
          6994 => x"56",
          6995 => x"70",
          6996 => x"76",
          6997 => x"84",
          6998 => x"18",
          6999 => x"12",
          7000 => x"2b",
          7001 => x"ff",
          7002 => x"2a",
          7003 => x"57",
          7004 => x"74",
          7005 => x"84",
          7006 => x"18",
          7007 => x"fe",
          7008 => x"3d",
          7009 => x"b9",
          7010 => x"58",
          7011 => x"a0",
          7012 => x"77",
          7013 => x"84",
          7014 => x"89",
          7015 => x"77",
          7016 => x"3f",
          7017 => x"08",
          7018 => x"0c",
          7019 => x"04",
          7020 => x"0b",
          7021 => x"0c",
          7022 => x"84",
          7023 => x"82",
          7024 => x"76",
          7025 => x"f4",
          7026 => x"b4",
          7027 => x"b8",
          7028 => x"75",
          7029 => x"81",
          7030 => x"b9",
          7031 => x"76",
          7032 => x"81",
          7033 => x"34",
          7034 => x"08",
          7035 => x"17",
          7036 => x"87",
          7037 => x"b9",
          7038 => x"b9",
          7039 => x"05",
          7040 => x"07",
          7041 => x"ff",
          7042 => x"2a",
          7043 => x"56",
          7044 => x"34",
          7045 => x"34",
          7046 => x"22",
          7047 => x"10",
          7048 => x"08",
          7049 => x"55",
          7050 => x"15",
          7051 => x"83",
          7052 => x"54",
          7053 => x"fe",
          7054 => x"e3",
          7055 => x"0d",
          7056 => x"5f",
          7057 => x"b9",
          7058 => x"45",
          7059 => x"2e",
          7060 => x"7e",
          7061 => x"af",
          7062 => x"2e",
          7063 => x"81",
          7064 => x"27",
          7065 => x"fb",
          7066 => x"82",
          7067 => x"ff",
          7068 => x"58",
          7069 => x"ff",
          7070 => x"31",
          7071 => x"83",
          7072 => x"70",
          7073 => x"11",
          7074 => x"12",
          7075 => x"2b",
          7076 => x"31",
          7077 => x"ff",
          7078 => x"10",
          7079 => x"73",
          7080 => x"11",
          7081 => x"12",
          7082 => x"2b",
          7083 => x"2b",
          7084 => x"53",
          7085 => x"44",
          7086 => x"44",
          7087 => x"52",
          7088 => x"80",
          7089 => x"fd",
          7090 => x"33",
          7091 => x"71",
          7092 => x"70",
          7093 => x"19",
          7094 => x"12",
          7095 => x"2b",
          7096 => x"07",
          7097 => x"56",
          7098 => x"74",
          7099 => x"38",
          7100 => x"82",
          7101 => x"1b",
          7102 => x"2e",
          7103 => x"60",
          7104 => x"f9",
          7105 => x"58",
          7106 => x"87",
          7107 => x"18",
          7108 => x"24",
          7109 => x"76",
          7110 => x"81",
          7111 => x"8b",
          7112 => x"2b",
          7113 => x"70",
          7114 => x"33",
          7115 => x"71",
          7116 => x"47",
          7117 => x"53",
          7118 => x"80",
          7119 => x"ba",
          7120 => x"82",
          7121 => x"12",
          7122 => x"2b",
          7123 => x"07",
          7124 => x"11",
          7125 => x"33",
          7126 => x"71",
          7127 => x"7e",
          7128 => x"33",
          7129 => x"71",
          7130 => x"70",
          7131 => x"57",
          7132 => x"41",
          7133 => x"59",
          7134 => x"1d",
          7135 => x"1d",
          7136 => x"b8",
          7137 => x"84",
          7138 => x"12",
          7139 => x"2b",
          7140 => x"07",
          7141 => x"14",
          7142 => x"33",
          7143 => x"07",
          7144 => x"5f",
          7145 => x"40",
          7146 => x"77",
          7147 => x"7b",
          7148 => x"84",
          7149 => x"16",
          7150 => x"12",
          7151 => x"2b",
          7152 => x"ff",
          7153 => x"2a",
          7154 => x"59",
          7155 => x"79",
          7156 => x"84",
          7157 => x"70",
          7158 => x"33",
          7159 => x"71",
          7160 => x"83",
          7161 => x"05",
          7162 => x"15",
          7163 => x"2b",
          7164 => x"2a",
          7165 => x"5d",
          7166 => x"55",
          7167 => x"75",
          7168 => x"84",
          7169 => x"70",
          7170 => x"81",
          7171 => x"8b",
          7172 => x"2b",
          7173 => x"82",
          7174 => x"15",
          7175 => x"2b",
          7176 => x"2a",
          7177 => x"5d",
          7178 => x"55",
          7179 => x"34",
          7180 => x"34",
          7181 => x"08",
          7182 => x"11",
          7183 => x"33",
          7184 => x"07",
          7185 => x"56",
          7186 => x"42",
          7187 => x"7e",
          7188 => x"51",
          7189 => x"3f",
          7190 => x"08",
          7191 => x"61",
          7192 => x"70",
          7193 => x"06",
          7194 => x"7a",
          7195 => x"b6",
          7196 => x"73",
          7197 => x"0c",
          7198 => x"04",
          7199 => x"0b",
          7200 => x"0c",
          7201 => x"84",
          7202 => x"82",
          7203 => x"60",
          7204 => x"f4",
          7205 => x"e8",
          7206 => x"b8",
          7207 => x"7e",
          7208 => x"81",
          7209 => x"b9",
          7210 => x"60",
          7211 => x"81",
          7212 => x"34",
          7213 => x"08",
          7214 => x"1d",
          7215 => x"87",
          7216 => x"b9",
          7217 => x"b9",
          7218 => x"05",
          7219 => x"07",
          7220 => x"ff",
          7221 => x"2a",
          7222 => x"57",
          7223 => x"34",
          7224 => x"34",
          7225 => x"22",
          7226 => x"10",
          7227 => x"08",
          7228 => x"55",
          7229 => x"15",
          7230 => x"83",
          7231 => x"b9",
          7232 => x"7e",
          7233 => x"76",
          7234 => x"8c",
          7235 => x"7f",
          7236 => x"df",
          7237 => x"f4",
          7238 => x"b9",
          7239 => x"b9",
          7240 => x"3d",
          7241 => x"1c",
          7242 => x"08",
          7243 => x"71",
          7244 => x"7f",
          7245 => x"81",
          7246 => x"88",
          7247 => x"ff",
          7248 => x"88",
          7249 => x"5b",
          7250 => x"7b",
          7251 => x"1c",
          7252 => x"b9",
          7253 => x"7c",
          7254 => x"58",
          7255 => x"34",
          7256 => x"34",
          7257 => x"08",
          7258 => x"33",
          7259 => x"71",
          7260 => x"70",
          7261 => x"ff",
          7262 => x"05",
          7263 => x"ff",
          7264 => x"2a",
          7265 => x"57",
          7266 => x"63",
          7267 => x"34",
          7268 => x"06",
          7269 => x"83",
          7270 => x"b9",
          7271 => x"5b",
          7272 => x"60",
          7273 => x"61",
          7274 => x"08",
          7275 => x"51",
          7276 => x"7e",
          7277 => x"39",
          7278 => x"70",
          7279 => x"06",
          7280 => x"ac",
          7281 => x"ff",
          7282 => x"31",
          7283 => x"ff",
          7284 => x"33",
          7285 => x"71",
          7286 => x"70",
          7287 => x"1b",
          7288 => x"12",
          7289 => x"2b",
          7290 => x"07",
          7291 => x"54",
          7292 => x"54",
          7293 => x"f9",
          7294 => x"bc",
          7295 => x"24",
          7296 => x"80",
          7297 => x"8f",
          7298 => x"ff",
          7299 => x"61",
          7300 => x"dd",
          7301 => x"39",
          7302 => x"0b",
          7303 => x"0c",
          7304 => x"84",
          7305 => x"82",
          7306 => x"7e",
          7307 => x"f4",
          7308 => x"cc",
          7309 => x"b8",
          7310 => x"7a",
          7311 => x"81",
          7312 => x"b9",
          7313 => x"7e",
          7314 => x"81",
          7315 => x"34",
          7316 => x"08",
          7317 => x"19",
          7318 => x"87",
          7319 => x"b9",
          7320 => x"b9",
          7321 => x"05",
          7322 => x"07",
          7323 => x"ff",
          7324 => x"2a",
          7325 => x"44",
          7326 => x"05",
          7327 => x"89",
          7328 => x"b9",
          7329 => x"10",
          7330 => x"b9",
          7331 => x"f8",
          7332 => x"7e",
          7333 => x"34",
          7334 => x"05",
          7335 => x"39",
          7336 => x"83",
          7337 => x"83",
          7338 => x"5b",
          7339 => x"fb",
          7340 => x"f2",
          7341 => x"2e",
          7342 => x"7e",
          7343 => x"3f",
          7344 => x"84",
          7345 => x"95",
          7346 => x"76",
          7347 => x"33",
          7348 => x"71",
          7349 => x"83",
          7350 => x"11",
          7351 => x"87",
          7352 => x"8b",
          7353 => x"2b",
          7354 => x"84",
          7355 => x"15",
          7356 => x"2b",
          7357 => x"2a",
          7358 => x"56",
          7359 => x"53",
          7360 => x"78",
          7361 => x"34",
          7362 => x"05",
          7363 => x"b8",
          7364 => x"84",
          7365 => x"12",
          7366 => x"2b",
          7367 => x"07",
          7368 => x"14",
          7369 => x"33",
          7370 => x"07",
          7371 => x"5b",
          7372 => x"5d",
          7373 => x"73",
          7374 => x"34",
          7375 => x"05",
          7376 => x"b8",
          7377 => x"33",
          7378 => x"71",
          7379 => x"81",
          7380 => x"70",
          7381 => x"5c",
          7382 => x"7d",
          7383 => x"1e",
          7384 => x"b8",
          7385 => x"82",
          7386 => x"12",
          7387 => x"2b",
          7388 => x"07",
          7389 => x"33",
          7390 => x"71",
          7391 => x"70",
          7392 => x"5c",
          7393 => x"57",
          7394 => x"7c",
          7395 => x"1d",
          7396 => x"b8",
          7397 => x"70",
          7398 => x"33",
          7399 => x"71",
          7400 => x"74",
          7401 => x"33",
          7402 => x"71",
          7403 => x"70",
          7404 => x"47",
          7405 => x"5c",
          7406 => x"82",
          7407 => x"83",
          7408 => x"b9",
          7409 => x"1f",
          7410 => x"83",
          7411 => x"88",
          7412 => x"57",
          7413 => x"83",
          7414 => x"58",
          7415 => x"84",
          7416 => x"bd",
          7417 => x"b9",
          7418 => x"84",
          7419 => x"ff",
          7420 => x"5f",
          7421 => x"84",
          7422 => x"84",
          7423 => x"a0",
          7424 => x"b9",
          7425 => x"80",
          7426 => x"52",
          7427 => x"51",
          7428 => x"3f",
          7429 => x"08",
          7430 => x"34",
          7431 => x"17",
          7432 => x"b8",
          7433 => x"84",
          7434 => x"0b",
          7435 => x"84",
          7436 => x"54",
          7437 => x"34",
          7438 => x"15",
          7439 => x"b8",
          7440 => x"b4",
          7441 => x"fe",
          7442 => x"70",
          7443 => x"06",
          7444 => x"45",
          7445 => x"61",
          7446 => x"60",
          7447 => x"84",
          7448 => x"70",
          7449 => x"84",
          7450 => x"05",
          7451 => x"5d",
          7452 => x"34",
          7453 => x"1c",
          7454 => x"e7",
          7455 => x"54",
          7456 => x"86",
          7457 => x"1a",
          7458 => x"2b",
          7459 => x"07",
          7460 => x"1c",
          7461 => x"33",
          7462 => x"07",
          7463 => x"5c",
          7464 => x"59",
          7465 => x"84",
          7466 => x"61",
          7467 => x"84",
          7468 => x"70",
          7469 => x"33",
          7470 => x"71",
          7471 => x"83",
          7472 => x"05",
          7473 => x"87",
          7474 => x"88",
          7475 => x"88",
          7476 => x"48",
          7477 => x"59",
          7478 => x"86",
          7479 => x"64",
          7480 => x"84",
          7481 => x"1d",
          7482 => x"12",
          7483 => x"2b",
          7484 => x"ff",
          7485 => x"2a",
          7486 => x"58",
          7487 => x"7f",
          7488 => x"84",
          7489 => x"70",
          7490 => x"81",
          7491 => x"8b",
          7492 => x"2b",
          7493 => x"70",
          7494 => x"33",
          7495 => x"07",
          7496 => x"8f",
          7497 => x"77",
          7498 => x"2a",
          7499 => x"5a",
          7500 => x"44",
          7501 => x"17",
          7502 => x"17",
          7503 => x"b8",
          7504 => x"70",
          7505 => x"33",
          7506 => x"71",
          7507 => x"74",
          7508 => x"81",
          7509 => x"88",
          7510 => x"ff",
          7511 => x"88",
          7512 => x"5e",
          7513 => x"41",
          7514 => x"34",
          7515 => x"05",
          7516 => x"ff",
          7517 => x"fa",
          7518 => x"15",
          7519 => x"33",
          7520 => x"71",
          7521 => x"79",
          7522 => x"33",
          7523 => x"71",
          7524 => x"70",
          7525 => x"5e",
          7526 => x"5d",
          7527 => x"34",
          7528 => x"34",
          7529 => x"08",
          7530 => x"11",
          7531 => x"33",
          7532 => x"71",
          7533 => x"74",
          7534 => x"33",
          7535 => x"71",
          7536 => x"70",
          7537 => x"56",
          7538 => x"42",
          7539 => x"60",
          7540 => x"75",
          7541 => x"34",
          7542 => x"08",
          7543 => x"81",
          7544 => x"88",
          7545 => x"ff",
          7546 => x"88",
          7547 => x"58",
          7548 => x"34",
          7549 => x"34",
          7550 => x"08",
          7551 => x"33",
          7552 => x"71",
          7553 => x"83",
          7554 => x"05",
          7555 => x"12",
          7556 => x"2b",
          7557 => x"2b",
          7558 => x"06",
          7559 => x"88",
          7560 => x"5f",
          7561 => x"42",
          7562 => x"82",
          7563 => x"83",
          7564 => x"b9",
          7565 => x"1f",
          7566 => x"12",
          7567 => x"2b",
          7568 => x"07",
          7569 => x"33",
          7570 => x"71",
          7571 => x"81",
          7572 => x"70",
          7573 => x"54",
          7574 => x"59",
          7575 => x"7c",
          7576 => x"1d",
          7577 => x"b8",
          7578 => x"82",
          7579 => x"12",
          7580 => x"2b",
          7581 => x"07",
          7582 => x"11",
          7583 => x"33",
          7584 => x"71",
          7585 => x"78",
          7586 => x"33",
          7587 => x"71",
          7588 => x"70",
          7589 => x"57",
          7590 => x"42",
          7591 => x"5a",
          7592 => x"84",
          7593 => x"85",
          7594 => x"b9",
          7595 => x"17",
          7596 => x"85",
          7597 => x"8b",
          7598 => x"2b",
          7599 => x"86",
          7600 => x"15",
          7601 => x"2b",
          7602 => x"2a",
          7603 => x"52",
          7604 => x"57",
          7605 => x"34",
          7606 => x"34",
          7607 => x"08",
          7608 => x"81",
          7609 => x"88",
          7610 => x"ff",
          7611 => x"88",
          7612 => x"5e",
          7613 => x"34",
          7614 => x"34",
          7615 => x"08",
          7616 => x"11",
          7617 => x"33",
          7618 => x"71",
          7619 => x"74",
          7620 => x"81",
          7621 => x"88",
          7622 => x"88",
          7623 => x"45",
          7624 => x"55",
          7625 => x"34",
          7626 => x"34",
          7627 => x"08",
          7628 => x"33",
          7629 => x"71",
          7630 => x"83",
          7631 => x"05",
          7632 => x"83",
          7633 => x"88",
          7634 => x"88",
          7635 => x"45",
          7636 => x"55",
          7637 => x"1a",
          7638 => x"1a",
          7639 => x"b8",
          7640 => x"82",
          7641 => x"12",
          7642 => x"2b",
          7643 => x"62",
          7644 => x"2b",
          7645 => x"5d",
          7646 => x"05",
          7647 => x"c3",
          7648 => x"b8",
          7649 => x"05",
          7650 => x"1c",
          7651 => x"ff",
          7652 => x"5f",
          7653 => x"86",
          7654 => x"1a",
          7655 => x"2b",
          7656 => x"07",
          7657 => x"1c",
          7658 => x"33",
          7659 => x"07",
          7660 => x"40",
          7661 => x"41",
          7662 => x"84",
          7663 => x"61",
          7664 => x"84",
          7665 => x"70",
          7666 => x"33",
          7667 => x"71",
          7668 => x"83",
          7669 => x"05",
          7670 => x"87",
          7671 => x"88",
          7672 => x"88",
          7673 => x"5f",
          7674 => x"41",
          7675 => x"86",
          7676 => x"64",
          7677 => x"84",
          7678 => x"1d",
          7679 => x"12",
          7680 => x"2b",
          7681 => x"ff",
          7682 => x"2a",
          7683 => x"55",
          7684 => x"7c",
          7685 => x"84",
          7686 => x"70",
          7687 => x"81",
          7688 => x"8b",
          7689 => x"2b",
          7690 => x"70",
          7691 => x"33",
          7692 => x"07",
          7693 => x"8f",
          7694 => x"77",
          7695 => x"2a",
          7696 => x"49",
          7697 => x"58",
          7698 => x"1e",
          7699 => x"1e",
          7700 => x"b8",
          7701 => x"70",
          7702 => x"33",
          7703 => x"71",
          7704 => x"74",
          7705 => x"81",
          7706 => x"88",
          7707 => x"ff",
          7708 => x"88",
          7709 => x"49",
          7710 => x"5e",
          7711 => x"34",
          7712 => x"34",
          7713 => x"ff",
          7714 => x"83",
          7715 => x"52",
          7716 => x"3f",
          7717 => x"08",
          7718 => x"c8",
          7719 => x"93",
          7720 => x"73",
          7721 => x"c8",
          7722 => x"b5",
          7723 => x"51",
          7724 => x"61",
          7725 => x"27",
          7726 => x"f0",
          7727 => x"3d",
          7728 => x"29",
          7729 => x"08",
          7730 => x"80",
          7731 => x"77",
          7732 => x"38",
          7733 => x"c8",
          7734 => x"0d",
          7735 => x"e4",
          7736 => x"b9",
          7737 => x"84",
          7738 => x"80",
          7739 => x"77",
          7740 => x"84",
          7741 => x"51",
          7742 => x"3f",
          7743 => x"c8",
          7744 => x"0d",
          7745 => x"f4",
          7746 => x"b8",
          7747 => x"0b",
          7748 => x"23",
          7749 => x"53",
          7750 => x"ff",
          7751 => x"b6",
          7752 => x"b9",
          7753 => x"76",
          7754 => x"0b",
          7755 => x"84",
          7756 => x"54",
          7757 => x"34",
          7758 => x"15",
          7759 => x"b8",
          7760 => x"86",
          7761 => x"0b",
          7762 => x"84",
          7763 => x"84",
          7764 => x"ff",
          7765 => x"80",
          7766 => x"ff",
          7767 => x"88",
          7768 => x"55",
          7769 => x"17",
          7770 => x"17",
          7771 => x"b4",
          7772 => x"10",
          7773 => x"b8",
          7774 => x"05",
          7775 => x"82",
          7776 => x"0b",
          7777 => x"77",
          7778 => x"2e",
          7779 => x"fe",
          7780 => x"3d",
          7781 => x"05",
          7782 => x"52",
          7783 => x"87",
          7784 => x"c4",
          7785 => x"71",
          7786 => x"0c",
          7787 => x"04",
          7788 => x"02",
          7789 => x"52",
          7790 => x"81",
          7791 => x"71",
          7792 => x"3f",
          7793 => x"08",
          7794 => x"53",
          7795 => x"72",
          7796 => x"13",
          7797 => x"c4",
          7798 => x"72",
          7799 => x"0c",
          7800 => x"04",
          7801 => x"7c",
          7802 => x"8c",
          7803 => x"33",
          7804 => x"59",
          7805 => x"74",
          7806 => x"84",
          7807 => x"33",
          7808 => x"06",
          7809 => x"73",
          7810 => x"58",
          7811 => x"c0",
          7812 => x"78",
          7813 => x"76",
          7814 => x"3f",
          7815 => x"08",
          7816 => x"55",
          7817 => x"a7",
          7818 => x"98",
          7819 => x"73",
          7820 => x"78",
          7821 => x"74",
          7822 => x"06",
          7823 => x"2e",
          7824 => x"54",
          7825 => x"84",
          7826 => x"8b",
          7827 => x"84",
          7828 => x"19",
          7829 => x"06",
          7830 => x"79",
          7831 => x"ac",
          7832 => x"f7",
          7833 => x"7e",
          7834 => x"05",
          7835 => x"5a",
          7836 => x"81",
          7837 => x"26",
          7838 => x"b9",
          7839 => x"54",
          7840 => x"54",
          7841 => x"bd",
          7842 => x"85",
          7843 => x"98",
          7844 => x"53",
          7845 => x"51",
          7846 => x"84",
          7847 => x"81",
          7848 => x"74",
          7849 => x"38",
          7850 => x"8c",
          7851 => x"e2",
          7852 => x"26",
          7853 => x"fc",
          7854 => x"54",
          7855 => x"83",
          7856 => x"73",
          7857 => x"b9",
          7858 => x"3d",
          7859 => x"80",
          7860 => x"70",
          7861 => x"5a",
          7862 => x"78",
          7863 => x"38",
          7864 => x"3d",
          7865 => x"84",
          7866 => x"33",
          7867 => x"9f",
          7868 => x"53",
          7869 => x"71",
          7870 => x"38",
          7871 => x"12",
          7872 => x"81",
          7873 => x"53",
          7874 => x"85",
          7875 => x"98",
          7876 => x"53",
          7877 => x"96",
          7878 => x"25",
          7879 => x"83",
          7880 => x"84",
          7881 => x"b9",
          7882 => x"3d",
          7883 => x"80",
          7884 => x"73",
          7885 => x"0c",
          7886 => x"04",
          7887 => x"0c",
          7888 => x"b9",
          7889 => x"3d",
          7890 => x"84",
          7891 => x"92",
          7892 => x"54",
          7893 => x"71",
          7894 => x"2a",
          7895 => x"51",
          7896 => x"8a",
          7897 => x"98",
          7898 => x"74",
          7899 => x"c0",
          7900 => x"51",
          7901 => x"81",
          7902 => x"c0",
          7903 => x"52",
          7904 => x"06",
          7905 => x"2e",
          7906 => x"71",
          7907 => x"54",
          7908 => x"ff",
          7909 => x"3d",
          7910 => x"80",
          7911 => x"33",
          7912 => x"57",
          7913 => x"09",
          7914 => x"38",
          7915 => x"75",
          7916 => x"87",
          7917 => x"80",
          7918 => x"33",
          7919 => x"3f",
          7920 => x"08",
          7921 => x"38",
          7922 => x"84",
          7923 => x"8c",
          7924 => x"81",
          7925 => x"08",
          7926 => x"70",
          7927 => x"33",
          7928 => x"ff",
          7929 => x"84",
          7930 => x"77",
          7931 => x"06",
          7932 => x"b9",
          7933 => x"19",
          7934 => x"08",
          7935 => x"08",
          7936 => x"08",
          7937 => x"08",
          7938 => x"5b",
          7939 => x"ff",
          7940 => x"18",
          7941 => x"82",
          7942 => x"06",
          7943 => x"81",
          7944 => x"53",
          7945 => x"18",
          7946 => x"b7",
          7947 => x"33",
          7948 => x"83",
          7949 => x"06",
          7950 => x"84",
          7951 => x"76",
          7952 => x"81",
          7953 => x"38",
          7954 => x"84",
          7955 => x"57",
          7956 => x"81",
          7957 => x"ff",
          7958 => x"f4",
          7959 => x"0b",
          7960 => x"34",
          7961 => x"84",
          7962 => x"80",
          7963 => x"80",
          7964 => x"19",
          7965 => x"0b",
          7966 => x"80",
          7967 => x"19",
          7968 => x"0b",
          7969 => x"34",
          7970 => x"84",
          7971 => x"80",
          7972 => x"9e",
          7973 => x"e1",
          7974 => x"19",
          7975 => x"08",
          7976 => x"a0",
          7977 => x"88",
          7978 => x"84",
          7979 => x"74",
          7980 => x"75",
          7981 => x"34",
          7982 => x"5b",
          7983 => x"19",
          7984 => x"08",
          7985 => x"a4",
          7986 => x"88",
          7987 => x"84",
          7988 => x"7a",
          7989 => x"75",
          7990 => x"34",
          7991 => x"55",
          7992 => x"19",
          7993 => x"08",
          7994 => x"b4",
          7995 => x"81",
          7996 => x"79",
          7997 => x"33",
          7998 => x"3f",
          7999 => x"34",
          8000 => x"52",
          8001 => x"51",
          8002 => x"84",
          8003 => x"80",
          8004 => x"38",
          8005 => x"f3",
          8006 => x"60",
          8007 => x"56",
          8008 => x"27",
          8009 => x"17",
          8010 => x"8c",
          8011 => x"77",
          8012 => x"0c",
          8013 => x"04",
          8014 => x"56",
          8015 => x"2e",
          8016 => x"74",
          8017 => x"a5",
          8018 => x"2e",
          8019 => x"dd",
          8020 => x"2a",
          8021 => x"2a",
          8022 => x"05",
          8023 => x"5b",
          8024 => x"79",
          8025 => x"83",
          8026 => x"7b",
          8027 => x"81",
          8028 => x"38",
          8029 => x"53",
          8030 => x"81",
          8031 => x"f8",
          8032 => x"b9",
          8033 => x"2e",
          8034 => x"59",
          8035 => x"b4",
          8036 => x"ff",
          8037 => x"83",
          8038 => x"b8",
          8039 => x"1c",
          8040 => x"a8",
          8041 => x"53",
          8042 => x"b4",
          8043 => x"2e",
          8044 => x"0b",
          8045 => x"71",
          8046 => x"74",
          8047 => x"81",
          8048 => x"38",
          8049 => x"53",
          8050 => x"81",
          8051 => x"f8",
          8052 => x"b9",
          8053 => x"2e",
          8054 => x"59",
          8055 => x"b4",
          8056 => x"fe",
          8057 => x"83",
          8058 => x"b8",
          8059 => x"88",
          8060 => x"78",
          8061 => x"84",
          8062 => x"59",
          8063 => x"fe",
          8064 => x"9f",
          8065 => x"b9",
          8066 => x"3d",
          8067 => x"88",
          8068 => x"08",
          8069 => x"17",
          8070 => x"b5",
          8071 => x"83",
          8072 => x"5c",
          8073 => x"7b",
          8074 => x"06",
          8075 => x"81",
          8076 => x"b8",
          8077 => x"17",
          8078 => x"a8",
          8079 => x"c8",
          8080 => x"85",
          8081 => x"81",
          8082 => x"18",
          8083 => x"df",
          8084 => x"83",
          8085 => x"05",
          8086 => x"11",
          8087 => x"71",
          8088 => x"84",
          8089 => x"57",
          8090 => x"0d",
          8091 => x"2e",
          8092 => x"fd",
          8093 => x"87",
          8094 => x"08",
          8095 => x"17",
          8096 => x"b5",
          8097 => x"83",
          8098 => x"5c",
          8099 => x"7b",
          8100 => x"06",
          8101 => x"81",
          8102 => x"b8",
          8103 => x"17",
          8104 => x"c0",
          8105 => x"c8",
          8106 => x"85",
          8107 => x"81",
          8108 => x"18",
          8109 => x"f7",
          8110 => x"2b",
          8111 => x"77",
          8112 => x"83",
          8113 => x"12",
          8114 => x"2b",
          8115 => x"07",
          8116 => x"70",
          8117 => x"2b",
          8118 => x"80",
          8119 => x"80",
          8120 => x"b9",
          8121 => x"5c",
          8122 => x"56",
          8123 => x"04",
          8124 => x"17",
          8125 => x"17",
          8126 => x"18",
          8127 => x"f6",
          8128 => x"5a",
          8129 => x"08",
          8130 => x"81",
          8131 => x"38",
          8132 => x"08",
          8133 => x"b4",
          8134 => x"18",
          8135 => x"b9",
          8136 => x"5e",
          8137 => x"08",
          8138 => x"38",
          8139 => x"55",
          8140 => x"09",
          8141 => x"f7",
          8142 => x"b4",
          8143 => x"18",
          8144 => x"7b",
          8145 => x"33",
          8146 => x"3f",
          8147 => x"df",
          8148 => x"b4",
          8149 => x"b8",
          8150 => x"81",
          8151 => x"5c",
          8152 => x"84",
          8153 => x"7b",
          8154 => x"06",
          8155 => x"84",
          8156 => x"83",
          8157 => x"17",
          8158 => x"08",
          8159 => x"a0",
          8160 => x"8b",
          8161 => x"33",
          8162 => x"2e",
          8163 => x"84",
          8164 => x"5b",
          8165 => x"81",
          8166 => x"08",
          8167 => x"70",
          8168 => x"33",
          8169 => x"bb",
          8170 => x"84",
          8171 => x"7b",
          8172 => x"06",
          8173 => x"84",
          8174 => x"83",
          8175 => x"17",
          8176 => x"08",
          8177 => x"c8",
          8178 => x"7d",
          8179 => x"27",
          8180 => x"82",
          8181 => x"74",
          8182 => x"81",
          8183 => x"38",
          8184 => x"17",
          8185 => x"08",
          8186 => x"52",
          8187 => x"51",
          8188 => x"7a",
          8189 => x"39",
          8190 => x"17",
          8191 => x"17",
          8192 => x"18",
          8193 => x"f4",
          8194 => x"5a",
          8195 => x"08",
          8196 => x"81",
          8197 => x"38",
          8198 => x"08",
          8199 => x"b4",
          8200 => x"18",
          8201 => x"b9",
          8202 => x"55",
          8203 => x"08",
          8204 => x"38",
          8205 => x"55",
          8206 => x"09",
          8207 => x"84",
          8208 => x"b4",
          8209 => x"18",
          8210 => x"7d",
          8211 => x"33",
          8212 => x"3f",
          8213 => x"ec",
          8214 => x"b4",
          8215 => x"18",
          8216 => x"7b",
          8217 => x"33",
          8218 => x"3f",
          8219 => x"81",
          8220 => x"bb",
          8221 => x"39",
          8222 => x"60",
          8223 => x"57",
          8224 => x"81",
          8225 => x"38",
          8226 => x"08",
          8227 => x"78",
          8228 => x"78",
          8229 => x"74",
          8230 => x"80",
          8231 => x"2e",
          8232 => x"77",
          8233 => x"0c",
          8234 => x"04",
          8235 => x"a8",
          8236 => x"58",
          8237 => x"1a",
          8238 => x"76",
          8239 => x"b6",
          8240 => x"33",
          8241 => x"7c",
          8242 => x"81",
          8243 => x"38",
          8244 => x"53",
          8245 => x"81",
          8246 => x"f2",
          8247 => x"b9",
          8248 => x"2e",
          8249 => x"58",
          8250 => x"b4",
          8251 => x"58",
          8252 => x"38",
          8253 => x"fe",
          8254 => x"7b",
          8255 => x"06",
          8256 => x"b8",
          8257 => x"88",
          8258 => x"b9",
          8259 => x"0b",
          8260 => x"77",
          8261 => x"0c",
          8262 => x"04",
          8263 => x"09",
          8264 => x"ff",
          8265 => x"2a",
          8266 => x"05",
          8267 => x"b4",
          8268 => x"5c",
          8269 => x"85",
          8270 => x"19",
          8271 => x"5d",
          8272 => x"09",
          8273 => x"bd",
          8274 => x"77",
          8275 => x"52",
          8276 => x"51",
          8277 => x"84",
          8278 => x"80",
          8279 => x"ff",
          8280 => x"77",
          8281 => x"79",
          8282 => x"b7",
          8283 => x"2b",
          8284 => x"79",
          8285 => x"83",
          8286 => x"98",
          8287 => x"06",
          8288 => x"06",
          8289 => x"5e",
          8290 => x"34",
          8291 => x"56",
          8292 => x"34",
          8293 => x"5a",
          8294 => x"34",
          8295 => x"5b",
          8296 => x"34",
          8297 => x"1a",
          8298 => x"39",
          8299 => x"16",
          8300 => x"a8",
          8301 => x"b4",
          8302 => x"59",
          8303 => x"2e",
          8304 => x"0b",
          8305 => x"71",
          8306 => x"74",
          8307 => x"81",
          8308 => x"38",
          8309 => x"53",
          8310 => x"81",
          8311 => x"f0",
          8312 => x"b9",
          8313 => x"2e",
          8314 => x"58",
          8315 => x"b4",
          8316 => x"58",
          8317 => x"38",
          8318 => x"06",
          8319 => x"81",
          8320 => x"06",
          8321 => x"7a",
          8322 => x"2e",
          8323 => x"84",
          8324 => x"06",
          8325 => x"06",
          8326 => x"5a",
          8327 => x"81",
          8328 => x"34",
          8329 => x"a8",
          8330 => x"56",
          8331 => x"1a",
          8332 => x"74",
          8333 => x"dd",
          8334 => x"74",
          8335 => x"70",
          8336 => x"33",
          8337 => x"9b",
          8338 => x"84",
          8339 => x"7f",
          8340 => x"06",
          8341 => x"84",
          8342 => x"83",
          8343 => x"19",
          8344 => x"1b",
          8345 => x"1b",
          8346 => x"c8",
          8347 => x"56",
          8348 => x"27",
          8349 => x"19",
          8350 => x"82",
          8351 => x"38",
          8352 => x"53",
          8353 => x"19",
          8354 => x"d8",
          8355 => x"c8",
          8356 => x"85",
          8357 => x"81",
          8358 => x"1a",
          8359 => x"83",
          8360 => x"ff",
          8361 => x"05",
          8362 => x"56",
          8363 => x"38",
          8364 => x"76",
          8365 => x"06",
          8366 => x"07",
          8367 => x"76",
          8368 => x"83",
          8369 => x"cb",
          8370 => x"76",
          8371 => x"70",
          8372 => x"33",
          8373 => x"8b",
          8374 => x"84",
          8375 => x"7c",
          8376 => x"06",
          8377 => x"84",
          8378 => x"83",
          8379 => x"19",
          8380 => x"1b",
          8381 => x"1b",
          8382 => x"c8",
          8383 => x"40",
          8384 => x"27",
          8385 => x"82",
          8386 => x"74",
          8387 => x"81",
          8388 => x"38",
          8389 => x"1e",
          8390 => x"81",
          8391 => x"ee",
          8392 => x"5a",
          8393 => x"81",
          8394 => x"b8",
          8395 => x"81",
          8396 => x"57",
          8397 => x"81",
          8398 => x"c8",
          8399 => x"09",
          8400 => x"ae",
          8401 => x"c8",
          8402 => x"34",
          8403 => x"70",
          8404 => x"31",
          8405 => x"84",
          8406 => x"5f",
          8407 => x"74",
          8408 => x"f0",
          8409 => x"33",
          8410 => x"2e",
          8411 => x"fc",
          8412 => x"54",
          8413 => x"76",
          8414 => x"33",
          8415 => x"3f",
          8416 => x"d0",
          8417 => x"76",
          8418 => x"70",
          8419 => x"33",
          8420 => x"cf",
          8421 => x"84",
          8422 => x"7c",
          8423 => x"06",
          8424 => x"84",
          8425 => x"83",
          8426 => x"19",
          8427 => x"1b",
          8428 => x"1b",
          8429 => x"c8",
          8430 => x"40",
          8431 => x"27",
          8432 => x"82",
          8433 => x"74",
          8434 => x"81",
          8435 => x"38",
          8436 => x"1e",
          8437 => x"81",
          8438 => x"ed",
          8439 => x"5a",
          8440 => x"81",
          8441 => x"53",
          8442 => x"19",
          8443 => x"f3",
          8444 => x"fd",
          8445 => x"76",
          8446 => x"06",
          8447 => x"83",
          8448 => x"59",
          8449 => x"b8",
          8450 => x"88",
          8451 => x"b9",
          8452 => x"fa",
          8453 => x"fd",
          8454 => x"76",
          8455 => x"fc",
          8456 => x"b8",
          8457 => x"33",
          8458 => x"8f",
          8459 => x"f0",
          8460 => x"42",
          8461 => x"58",
          8462 => x"7d",
          8463 => x"75",
          8464 => x"7d",
          8465 => x"79",
          8466 => x"7d",
          8467 => x"7a",
          8468 => x"fa",
          8469 => x"3d",
          8470 => x"71",
          8471 => x"5a",
          8472 => x"38",
          8473 => x"57",
          8474 => x"80",
          8475 => x"9c",
          8476 => x"80",
          8477 => x"19",
          8478 => x"54",
          8479 => x"80",
          8480 => x"7b",
          8481 => x"38",
          8482 => x"16",
          8483 => x"08",
          8484 => x"38",
          8485 => x"77",
          8486 => x"38",
          8487 => x"51",
          8488 => x"84",
          8489 => x"80",
          8490 => x"38",
          8491 => x"b9",
          8492 => x"2e",
          8493 => x"b9",
          8494 => x"70",
          8495 => x"07",
          8496 => x"7b",
          8497 => x"55",
          8498 => x"aa",
          8499 => x"2e",
          8500 => x"ff",
          8501 => x"55",
          8502 => x"c8",
          8503 => x"0d",
          8504 => x"ff",
          8505 => x"b9",
          8506 => x"ca",
          8507 => x"79",
          8508 => x"3f",
          8509 => x"84",
          8510 => x"27",
          8511 => x"b9",
          8512 => x"84",
          8513 => x"ff",
          8514 => x"9c",
          8515 => x"b9",
          8516 => x"c4",
          8517 => x"fe",
          8518 => x"1b",
          8519 => x"08",
          8520 => x"38",
          8521 => x"52",
          8522 => x"eb",
          8523 => x"84",
          8524 => x"81",
          8525 => x"38",
          8526 => x"08",
          8527 => x"70",
          8528 => x"25",
          8529 => x"84",
          8530 => x"54",
          8531 => x"55",
          8532 => x"38",
          8533 => x"08",
          8534 => x"38",
          8535 => x"54",
          8536 => x"fe",
          8537 => x"9c",
          8538 => x"fe",
          8539 => x"70",
          8540 => x"96",
          8541 => x"2e",
          8542 => x"ff",
          8543 => x"78",
          8544 => x"3f",
          8545 => x"08",
          8546 => x"08",
          8547 => x"b9",
          8548 => x"80",
          8549 => x"55",
          8550 => x"38",
          8551 => x"38",
          8552 => x"0c",
          8553 => x"fe",
          8554 => x"08",
          8555 => x"78",
          8556 => x"ff",
          8557 => x"0c",
          8558 => x"81",
          8559 => x"84",
          8560 => x"55",
          8561 => x"c8",
          8562 => x"0d",
          8563 => x"84",
          8564 => x"8c",
          8565 => x"84",
          8566 => x"58",
          8567 => x"73",
          8568 => x"b8",
          8569 => x"7a",
          8570 => x"f5",
          8571 => x"b9",
          8572 => x"ff",
          8573 => x"b9",
          8574 => x"b9",
          8575 => x"3d",
          8576 => x"56",
          8577 => x"ff",
          8578 => x"55",
          8579 => x"f8",
          8580 => x"7c",
          8581 => x"55",
          8582 => x"80",
          8583 => x"df",
          8584 => x"06",
          8585 => x"d7",
          8586 => x"19",
          8587 => x"08",
          8588 => x"df",
          8589 => x"56",
          8590 => x"80",
          8591 => x"85",
          8592 => x"0b",
          8593 => x"5a",
          8594 => x"27",
          8595 => x"17",
          8596 => x"0c",
          8597 => x"0c",
          8598 => x"53",
          8599 => x"80",
          8600 => x"73",
          8601 => x"98",
          8602 => x"83",
          8603 => x"b8",
          8604 => x"0c",
          8605 => x"84",
          8606 => x"8a",
          8607 => x"82",
          8608 => x"c8",
          8609 => x"0d",
          8610 => x"08",
          8611 => x"2e",
          8612 => x"8a",
          8613 => x"89",
          8614 => x"73",
          8615 => x"38",
          8616 => x"53",
          8617 => x"14",
          8618 => x"59",
          8619 => x"8d",
          8620 => x"22",
          8621 => x"b0",
          8622 => x"5a",
          8623 => x"19",
          8624 => x"39",
          8625 => x"51",
          8626 => x"84",
          8627 => x"55",
          8628 => x"08",
          8629 => x"38",
          8630 => x"b9",
          8631 => x"ff",
          8632 => x"17",
          8633 => x"b9",
          8634 => x"27",
          8635 => x"73",
          8636 => x"73",
          8637 => x"38",
          8638 => x"81",
          8639 => x"c8",
          8640 => x"0d",
          8641 => x"0d",
          8642 => x"90",
          8643 => x"05",
          8644 => x"f0",
          8645 => x"27",
          8646 => x"0b",
          8647 => x"98",
          8648 => x"84",
          8649 => x"2e",
          8650 => x"83",
          8651 => x"7a",
          8652 => x"15",
          8653 => x"57",
          8654 => x"38",
          8655 => x"88",
          8656 => x"55",
          8657 => x"81",
          8658 => x"98",
          8659 => x"90",
          8660 => x"1b",
          8661 => x"18",
          8662 => x"75",
          8663 => x"0c",
          8664 => x"04",
          8665 => x"0c",
          8666 => x"ff",
          8667 => x"2a",
          8668 => x"da",
          8669 => x"76",
          8670 => x"3f",
          8671 => x"08",
          8672 => x"81",
          8673 => x"c8",
          8674 => x"38",
          8675 => x"b9",
          8676 => x"2e",
          8677 => x"19",
          8678 => x"c8",
          8679 => x"91",
          8680 => x"2e",
          8681 => x"94",
          8682 => x"76",
          8683 => x"3f",
          8684 => x"08",
          8685 => x"84",
          8686 => x"80",
          8687 => x"38",
          8688 => x"b9",
          8689 => x"2e",
          8690 => x"81",
          8691 => x"c8",
          8692 => x"ff",
          8693 => x"b9",
          8694 => x"1a",
          8695 => x"7d",
          8696 => x"fe",
          8697 => x"08",
          8698 => x"56",
          8699 => x"78",
          8700 => x"8a",
          8701 => x"71",
          8702 => x"08",
          8703 => x"7b",
          8704 => x"b8",
          8705 => x"80",
          8706 => x"80",
          8707 => x"05",
          8708 => x"15",
          8709 => x"38",
          8710 => x"19",
          8711 => x"75",
          8712 => x"38",
          8713 => x"1c",
          8714 => x"81",
          8715 => x"e4",
          8716 => x"b9",
          8717 => x"e7",
          8718 => x"56",
          8719 => x"98",
          8720 => x"0b",
          8721 => x"0c",
          8722 => x"04",
          8723 => x"19",
          8724 => x"19",
          8725 => x"1a",
          8726 => x"e4",
          8727 => x"b9",
          8728 => x"f3",
          8729 => x"c8",
          8730 => x"34",
          8731 => x"a8",
          8732 => x"55",
          8733 => x"08",
          8734 => x"38",
          8735 => x"5c",
          8736 => x"09",
          8737 => x"db",
          8738 => x"b4",
          8739 => x"1a",
          8740 => x"75",
          8741 => x"33",
          8742 => x"3f",
          8743 => x"8a",
          8744 => x"74",
          8745 => x"06",
          8746 => x"2e",
          8747 => x"a7",
          8748 => x"18",
          8749 => x"9c",
          8750 => x"05",
          8751 => x"58",
          8752 => x"fd",
          8753 => x"19",
          8754 => x"29",
          8755 => x"05",
          8756 => x"5c",
          8757 => x"81",
          8758 => x"c8",
          8759 => x"0d",
          8760 => x"0d",
          8761 => x"5c",
          8762 => x"5a",
          8763 => x"70",
          8764 => x"58",
          8765 => x"80",
          8766 => x"38",
          8767 => x"75",
          8768 => x"b4",
          8769 => x"2e",
          8770 => x"83",
          8771 => x"58",
          8772 => x"2e",
          8773 => x"81",
          8774 => x"54",
          8775 => x"19",
          8776 => x"33",
          8777 => x"3f",
          8778 => x"08",
          8779 => x"38",
          8780 => x"57",
          8781 => x"0c",
          8782 => x"82",
          8783 => x"1c",
          8784 => x"58",
          8785 => x"2e",
          8786 => x"8b",
          8787 => x"06",
          8788 => x"06",
          8789 => x"86",
          8790 => x"81",
          8791 => x"30",
          8792 => x"70",
          8793 => x"25",
          8794 => x"07",
          8795 => x"57",
          8796 => x"38",
          8797 => x"06",
          8798 => x"88",
          8799 => x"38",
          8800 => x"81",
          8801 => x"ff",
          8802 => x"7b",
          8803 => x"3f",
          8804 => x"08",
          8805 => x"c8",
          8806 => x"38",
          8807 => x"56",
          8808 => x"38",
          8809 => x"c8",
          8810 => x"0d",
          8811 => x"b4",
          8812 => x"7e",
          8813 => x"33",
          8814 => x"3f",
          8815 => x"b9",
          8816 => x"2e",
          8817 => x"fe",
          8818 => x"b9",
          8819 => x"1a",
          8820 => x"08",
          8821 => x"31",
          8822 => x"08",
          8823 => x"a0",
          8824 => x"fe",
          8825 => x"19",
          8826 => x"82",
          8827 => x"06",
          8828 => x"81",
          8829 => x"08",
          8830 => x"05",
          8831 => x"81",
          8832 => x"e0",
          8833 => x"57",
          8834 => x"79",
          8835 => x"81",
          8836 => x"38",
          8837 => x"81",
          8838 => x"80",
          8839 => x"8d",
          8840 => x"81",
          8841 => x"90",
          8842 => x"ac",
          8843 => x"5e",
          8844 => x"2e",
          8845 => x"ff",
          8846 => x"fe",
          8847 => x"56",
          8848 => x"09",
          8849 => x"be",
          8850 => x"84",
          8851 => x"98",
          8852 => x"84",
          8853 => x"94",
          8854 => x"77",
          8855 => x"39",
          8856 => x"57",
          8857 => x"09",
          8858 => x"38",
          8859 => x"9b",
          8860 => x"1a",
          8861 => x"2b",
          8862 => x"41",
          8863 => x"38",
          8864 => x"81",
          8865 => x"29",
          8866 => x"5a",
          8867 => x"5b",
          8868 => x"17",
          8869 => x"81",
          8870 => x"33",
          8871 => x"07",
          8872 => x"7a",
          8873 => x"c5",
          8874 => x"fe",
          8875 => x"38",
          8876 => x"05",
          8877 => x"75",
          8878 => x"1a",
          8879 => x"57",
          8880 => x"cc",
          8881 => x"70",
          8882 => x"06",
          8883 => x"80",
          8884 => x"79",
          8885 => x"fe",
          8886 => x"10",
          8887 => x"80",
          8888 => x"1d",
          8889 => x"06",
          8890 => x"9d",
          8891 => x"ff",
          8892 => x"38",
          8893 => x"fe",
          8894 => x"a8",
          8895 => x"8b",
          8896 => x"2a",
          8897 => x"29",
          8898 => x"81",
          8899 => x"40",
          8900 => x"81",
          8901 => x"19",
          8902 => x"76",
          8903 => x"7e",
          8904 => x"38",
          8905 => x"1d",
          8906 => x"b9",
          8907 => x"3d",
          8908 => x"3d",
          8909 => x"08",
          8910 => x"52",
          8911 => x"cf",
          8912 => x"c8",
          8913 => x"b9",
          8914 => x"80",
          8915 => x"70",
          8916 => x"0b",
          8917 => x"b8",
          8918 => x"1c",
          8919 => x"58",
          8920 => x"76",
          8921 => x"38",
          8922 => x"78",
          8923 => x"78",
          8924 => x"06",
          8925 => x"81",
          8926 => x"b8",
          8927 => x"1b",
          8928 => x"e0",
          8929 => x"c8",
          8930 => x"85",
          8931 => x"81",
          8932 => x"1c",
          8933 => x"76",
          8934 => x"9c",
          8935 => x"33",
          8936 => x"80",
          8937 => x"38",
          8938 => x"bf",
          8939 => x"ff",
          8940 => x"77",
          8941 => x"76",
          8942 => x"80",
          8943 => x"83",
          8944 => x"55",
          8945 => x"81",
          8946 => x"80",
          8947 => x"8f",
          8948 => x"38",
          8949 => x"78",
          8950 => x"8b",
          8951 => x"2a",
          8952 => x"29",
          8953 => x"81",
          8954 => x"57",
          8955 => x"81",
          8956 => x"19",
          8957 => x"76",
          8958 => x"7f",
          8959 => x"38",
          8960 => x"81",
          8961 => x"a7",
          8962 => x"a0",
          8963 => x"78",
          8964 => x"5a",
          8965 => x"81",
          8966 => x"71",
          8967 => x"1a",
          8968 => x"40",
          8969 => x"81",
          8970 => x"80",
          8971 => x"81",
          8972 => x"0b",
          8973 => x"80",
          8974 => x"f5",
          8975 => x"b9",
          8976 => x"84",
          8977 => x"80",
          8978 => x"38",
          8979 => x"c8",
          8980 => x"0d",
          8981 => x"b4",
          8982 => x"7d",
          8983 => x"33",
          8984 => x"3f",
          8985 => x"b9",
          8986 => x"2e",
          8987 => x"fe",
          8988 => x"b9",
          8989 => x"1c",
          8990 => x"08",
          8991 => x"31",
          8992 => x"08",
          8993 => x"a0",
          8994 => x"fd",
          8995 => x"1b",
          8996 => x"82",
          8997 => x"06",
          8998 => x"81",
          8999 => x"08",
          9000 => x"05",
          9001 => x"81",
          9002 => x"db",
          9003 => x"57",
          9004 => x"77",
          9005 => x"39",
          9006 => x"70",
          9007 => x"06",
          9008 => x"fe",
          9009 => x"86",
          9010 => x"5a",
          9011 => x"93",
          9012 => x"33",
          9013 => x"06",
          9014 => x"08",
          9015 => x"0c",
          9016 => x"76",
          9017 => x"38",
          9018 => x"74",
          9019 => x"7b",
          9020 => x"3f",
          9021 => x"08",
          9022 => x"c8",
          9023 => x"fc",
          9024 => x"c8",
          9025 => x"2e",
          9026 => x"81",
          9027 => x"0b",
          9028 => x"fe",
          9029 => x"19",
          9030 => x"77",
          9031 => x"06",
          9032 => x"1b",
          9033 => x"33",
          9034 => x"71",
          9035 => x"59",
          9036 => x"ff",
          9037 => x"33",
          9038 => x"8d",
          9039 => x"5b",
          9040 => x"59",
          9041 => x"c8",
          9042 => x"05",
          9043 => x"71",
          9044 => x"2b",
          9045 => x"57",
          9046 => x"80",
          9047 => x"81",
          9048 => x"84",
          9049 => x"81",
          9050 => x"84",
          9051 => x"7a",
          9052 => x"70",
          9053 => x"81",
          9054 => x"81",
          9055 => x"75",
          9056 => x"08",
          9057 => x"06",
          9058 => x"76",
          9059 => x"58",
          9060 => x"ff",
          9061 => x"33",
          9062 => x"81",
          9063 => x"75",
          9064 => x"38",
          9065 => x"8d",
          9066 => x"60",
          9067 => x"41",
          9068 => x"b4",
          9069 => x"70",
          9070 => x"5e",
          9071 => x"39",
          9072 => x"b9",
          9073 => x"3d",
          9074 => x"83",
          9075 => x"ff",
          9076 => x"ff",
          9077 => x"39",
          9078 => x"68",
          9079 => x"ab",
          9080 => x"a0",
          9081 => x"5d",
          9082 => x"74",
          9083 => x"74",
          9084 => x"70",
          9085 => x"5d",
          9086 => x"8e",
          9087 => x"70",
          9088 => x"22",
          9089 => x"74",
          9090 => x"3d",
          9091 => x"40",
          9092 => x"58",
          9093 => x"70",
          9094 => x"33",
          9095 => x"05",
          9096 => x"15",
          9097 => x"38",
          9098 => x"05",
          9099 => x"06",
          9100 => x"80",
          9101 => x"38",
          9102 => x"ab",
          9103 => x"0b",
          9104 => x"5b",
          9105 => x"7b",
          9106 => x"7a",
          9107 => x"55",
          9108 => x"05",
          9109 => x"70",
          9110 => x"34",
          9111 => x"74",
          9112 => x"7b",
          9113 => x"38",
          9114 => x"56",
          9115 => x"2e",
          9116 => x"82",
          9117 => x"8f",
          9118 => x"06",
          9119 => x"76",
          9120 => x"83",
          9121 => x"72",
          9122 => x"06",
          9123 => x"57",
          9124 => x"87",
          9125 => x"a0",
          9126 => x"ff",
          9127 => x"80",
          9128 => x"78",
          9129 => x"ca",
          9130 => x"84",
          9131 => x"05",
          9132 => x"b0",
          9133 => x"55",
          9134 => x"84",
          9135 => x"55",
          9136 => x"ff",
          9137 => x"78",
          9138 => x"59",
          9139 => x"38",
          9140 => x"80",
          9141 => x"76",
          9142 => x"80",
          9143 => x"38",
          9144 => x"74",
          9145 => x"38",
          9146 => x"75",
          9147 => x"a2",
          9148 => x"70",
          9149 => x"74",
          9150 => x"81",
          9151 => x"81",
          9152 => x"55",
          9153 => x"8e",
          9154 => x"78",
          9155 => x"81",
          9156 => x"57",
          9157 => x"77",
          9158 => x"27",
          9159 => x"7d",
          9160 => x"3f",
          9161 => x"08",
          9162 => x"1b",
          9163 => x"7b",
          9164 => x"38",
          9165 => x"80",
          9166 => x"e7",
          9167 => x"c8",
          9168 => x"b9",
          9169 => x"2e",
          9170 => x"82",
          9171 => x"80",
          9172 => x"ab",
          9173 => x"08",
          9174 => x"80",
          9175 => x"57",
          9176 => x"2a",
          9177 => x"81",
          9178 => x"2e",
          9179 => x"52",
          9180 => x"fe",
          9181 => x"84",
          9182 => x"1b",
          9183 => x"7d",
          9184 => x"3f",
          9185 => x"08",
          9186 => x"c8",
          9187 => x"38",
          9188 => x"08",
          9189 => x"59",
          9190 => x"56",
          9191 => x"18",
          9192 => x"85",
          9193 => x"18",
          9194 => x"77",
          9195 => x"06",
          9196 => x"81",
          9197 => x"b8",
          9198 => x"18",
          9199 => x"a4",
          9200 => x"c8",
          9201 => x"85",
          9202 => x"81",
          9203 => x"19",
          9204 => x"76",
          9205 => x"1e",
          9206 => x"56",
          9207 => x"e5",
          9208 => x"38",
          9209 => x"80",
          9210 => x"56",
          9211 => x"2e",
          9212 => x"81",
          9213 => x"7b",
          9214 => x"38",
          9215 => x"51",
          9216 => x"84",
          9217 => x"56",
          9218 => x"08",
          9219 => x"88",
          9220 => x"75",
          9221 => x"89",
          9222 => x"75",
          9223 => x"ff",
          9224 => x"81",
          9225 => x"1e",
          9226 => x"1c",
          9227 => x"af",
          9228 => x"33",
          9229 => x"7f",
          9230 => x"81",
          9231 => x"b8",
          9232 => x"1c",
          9233 => x"9c",
          9234 => x"c8",
          9235 => x"85",
          9236 => x"81",
          9237 => x"1d",
          9238 => x"75",
          9239 => x"a0",
          9240 => x"08",
          9241 => x"76",
          9242 => x"58",
          9243 => x"55",
          9244 => x"8b",
          9245 => x"08",
          9246 => x"55",
          9247 => x"05",
          9248 => x"70",
          9249 => x"34",
          9250 => x"74",
          9251 => x"1e",
          9252 => x"33",
          9253 => x"5a",
          9254 => x"34",
          9255 => x"1d",
          9256 => x"75",
          9257 => x"0c",
          9258 => x"04",
          9259 => x"70",
          9260 => x"07",
          9261 => x"74",
          9262 => x"74",
          9263 => x"7d",
          9264 => x"3f",
          9265 => x"08",
          9266 => x"c8",
          9267 => x"fd",
          9268 => x"bd",
          9269 => x"b4",
          9270 => x"7c",
          9271 => x"33",
          9272 => x"3f",
          9273 => x"08",
          9274 => x"81",
          9275 => x"38",
          9276 => x"08",
          9277 => x"b4",
          9278 => x"19",
          9279 => x"74",
          9280 => x"27",
          9281 => x"18",
          9282 => x"82",
          9283 => x"38",
          9284 => x"08",
          9285 => x"39",
          9286 => x"90",
          9287 => x"31",
          9288 => x"51",
          9289 => x"84",
          9290 => x"58",
          9291 => x"08",
          9292 => x"79",
          9293 => x"08",
          9294 => x"57",
          9295 => x"75",
          9296 => x"05",
          9297 => x"05",
          9298 => x"76",
          9299 => x"ff",
          9300 => x"59",
          9301 => x"e4",
          9302 => x"ff",
          9303 => x"43",
          9304 => x"08",
          9305 => x"b4",
          9306 => x"2e",
          9307 => x"1c",
          9308 => x"76",
          9309 => x"06",
          9310 => x"81",
          9311 => x"b8",
          9312 => x"1c",
          9313 => x"dc",
          9314 => x"c8",
          9315 => x"85",
          9316 => x"81",
          9317 => x"1d",
          9318 => x"75",
          9319 => x"8c",
          9320 => x"1f",
          9321 => x"ff",
          9322 => x"5f",
          9323 => x"34",
          9324 => x"1c",
          9325 => x"1c",
          9326 => x"1c",
          9327 => x"1c",
          9328 => x"29",
          9329 => x"77",
          9330 => x"76",
          9331 => x"2e",
          9332 => x"10",
          9333 => x"81",
          9334 => x"56",
          9335 => x"18",
          9336 => x"55",
          9337 => x"81",
          9338 => x"76",
          9339 => x"75",
          9340 => x"85",
          9341 => x"ff",
          9342 => x"58",
          9343 => x"cb",
          9344 => x"ff",
          9345 => x"b3",
          9346 => x"1f",
          9347 => x"58",
          9348 => x"81",
          9349 => x"7b",
          9350 => x"83",
          9351 => x"52",
          9352 => x"e1",
          9353 => x"c8",
          9354 => x"b9",
          9355 => x"f1",
          9356 => x"05",
          9357 => x"a9",
          9358 => x"39",
          9359 => x"1c",
          9360 => x"1c",
          9361 => x"1d",
          9362 => x"d0",
          9363 => x"56",
          9364 => x"08",
          9365 => x"84",
          9366 => x"83",
          9367 => x"1c",
          9368 => x"08",
          9369 => x"c8",
          9370 => x"60",
          9371 => x"27",
          9372 => x"82",
          9373 => x"61",
          9374 => x"81",
          9375 => x"38",
          9376 => x"1c",
          9377 => x"08",
          9378 => x"52",
          9379 => x"51",
          9380 => x"77",
          9381 => x"39",
          9382 => x"08",
          9383 => x"43",
          9384 => x"e5",
          9385 => x"06",
          9386 => x"fb",
          9387 => x"70",
          9388 => x"80",
          9389 => x"38",
          9390 => x"7c",
          9391 => x"5d",
          9392 => x"81",
          9393 => x"08",
          9394 => x"81",
          9395 => x"cf",
          9396 => x"b9",
          9397 => x"2e",
          9398 => x"bc",
          9399 => x"c8",
          9400 => x"34",
          9401 => x"a8",
          9402 => x"55",
          9403 => x"08",
          9404 => x"82",
          9405 => x"7e",
          9406 => x"38",
          9407 => x"08",
          9408 => x"39",
          9409 => x"41",
          9410 => x"2e",
          9411 => x"fc",
          9412 => x"1a",
          9413 => x"39",
          9414 => x"56",
          9415 => x"fc",
          9416 => x"fd",
          9417 => x"b4",
          9418 => x"1d",
          9419 => x"61",
          9420 => x"33",
          9421 => x"3f",
          9422 => x"81",
          9423 => x"08",
          9424 => x"05",
          9425 => x"81",
          9426 => x"ce",
          9427 => x"e3",
          9428 => x"0d",
          9429 => x"08",
          9430 => x"80",
          9431 => x"34",
          9432 => x"80",
          9433 => x"38",
          9434 => x"ff",
          9435 => x"38",
          9436 => x"60",
          9437 => x"70",
          9438 => x"5b",
          9439 => x"78",
          9440 => x"77",
          9441 => x"70",
          9442 => x"5b",
          9443 => x"82",
          9444 => x"d0",
          9445 => x"83",
          9446 => x"58",
          9447 => x"ff",
          9448 => x"38",
          9449 => x"76",
          9450 => x"5d",
          9451 => x"79",
          9452 => x"30",
          9453 => x"70",
          9454 => x"5a",
          9455 => x"18",
          9456 => x"80",
          9457 => x"34",
          9458 => x"1f",
          9459 => x"9c",
          9460 => x"70",
          9461 => x"58",
          9462 => x"a0",
          9463 => x"74",
          9464 => x"bc",
          9465 => x"32",
          9466 => x"72",
          9467 => x"55",
          9468 => x"8b",
          9469 => x"72",
          9470 => x"38",
          9471 => x"81",
          9472 => x"81",
          9473 => x"77",
          9474 => x"59",
          9475 => x"58",
          9476 => x"ff",
          9477 => x"18",
          9478 => x"80",
          9479 => x"34",
          9480 => x"53",
          9481 => x"77",
          9482 => x"bf",
          9483 => x"34",
          9484 => x"17",
          9485 => x"80",
          9486 => x"34",
          9487 => x"8c",
          9488 => x"53",
          9489 => x"73",
          9490 => x"9c",
          9491 => x"8b",
          9492 => x"1e",
          9493 => x"08",
          9494 => x"11",
          9495 => x"33",
          9496 => x"71",
          9497 => x"81",
          9498 => x"72",
          9499 => x"75",
          9500 => x"64",
          9501 => x"16",
          9502 => x"33",
          9503 => x"07",
          9504 => x"40",
          9505 => x"55",
          9506 => x"23",
          9507 => x"98",
          9508 => x"88",
          9509 => x"54",
          9510 => x"23",
          9511 => x"04",
          9512 => x"fe",
          9513 => x"1d",
          9514 => x"ff",
          9515 => x"5b",
          9516 => x"52",
          9517 => x"74",
          9518 => x"91",
          9519 => x"b9",
          9520 => x"ff",
          9521 => x"81",
          9522 => x"ad",
          9523 => x"27",
          9524 => x"74",
          9525 => x"73",
          9526 => x"97",
          9527 => x"78",
          9528 => x"0b",
          9529 => x"56",
          9530 => x"75",
          9531 => x"5c",
          9532 => x"fd",
          9533 => x"ba",
          9534 => x"76",
          9535 => x"07",
          9536 => x"80",
          9537 => x"55",
          9538 => x"f9",
          9539 => x"34",
          9540 => x"58",
          9541 => x"1f",
          9542 => x"cd",
          9543 => x"89",
          9544 => x"57",
          9545 => x"2e",
          9546 => x"7c",
          9547 => x"57",
          9548 => x"14",
          9549 => x"11",
          9550 => x"99",
          9551 => x"9c",
          9552 => x"11",
          9553 => x"88",
          9554 => x"38",
          9555 => x"53",
          9556 => x"5e",
          9557 => x"8a",
          9558 => x"70",
          9559 => x"06",
          9560 => x"78",
          9561 => x"5a",
          9562 => x"81",
          9563 => x"71",
          9564 => x"5e",
          9565 => x"56",
          9566 => x"38",
          9567 => x"72",
          9568 => x"cc",
          9569 => x"30",
          9570 => x"70",
          9571 => x"53",
          9572 => x"fc",
          9573 => x"3d",
          9574 => x"08",
          9575 => x"5c",
          9576 => x"33",
          9577 => x"74",
          9578 => x"38",
          9579 => x"80",
          9580 => x"df",
          9581 => x"2e",
          9582 => x"98",
          9583 => x"1d",
          9584 => x"96",
          9585 => x"41",
          9586 => x"75",
          9587 => x"38",
          9588 => x"16",
          9589 => x"57",
          9590 => x"81",
          9591 => x"55",
          9592 => x"df",
          9593 => x"0c",
          9594 => x"81",
          9595 => x"ff",
          9596 => x"8b",
          9597 => x"18",
          9598 => x"23",
          9599 => x"73",
          9600 => x"06",
          9601 => x"70",
          9602 => x"27",
          9603 => x"07",
          9604 => x"55",
          9605 => x"38",
          9606 => x"2e",
          9607 => x"74",
          9608 => x"b2",
          9609 => x"e4",
          9610 => x"e4",
          9611 => x"ff",
          9612 => x"56",
          9613 => x"81",
          9614 => x"75",
          9615 => x"81",
          9616 => x"70",
          9617 => x"56",
          9618 => x"ee",
          9619 => x"ff",
          9620 => x"81",
          9621 => x"81",
          9622 => x"fd",
          9623 => x"18",
          9624 => x"23",
          9625 => x"70",
          9626 => x"52",
          9627 => x"57",
          9628 => x"fe",
          9629 => x"cb",
          9630 => x"80",
          9631 => x"30",
          9632 => x"73",
          9633 => x"58",
          9634 => x"2e",
          9635 => x"14",
          9636 => x"80",
          9637 => x"55",
          9638 => x"dd",
          9639 => x"dc",
          9640 => x"70",
          9641 => x"07",
          9642 => x"72",
          9643 => x"88",
          9644 => x"33",
          9645 => x"3d",
          9646 => x"74",
          9647 => x"90",
          9648 => x"83",
          9649 => x"51",
          9650 => x"3f",
          9651 => x"08",
          9652 => x"06",
          9653 => x"8d",
          9654 => x"73",
          9655 => x"0c",
          9656 => x"04",
          9657 => x"33",
          9658 => x"06",
          9659 => x"80",
          9660 => x"38",
          9661 => x"80",
          9662 => x"34",
          9663 => x"51",
          9664 => x"84",
          9665 => x"84",
          9666 => x"93",
          9667 => x"81",
          9668 => x"32",
          9669 => x"80",
          9670 => x"41",
          9671 => x"7d",
          9672 => x"38",
          9673 => x"80",
          9674 => x"55",
          9675 => x"af",
          9676 => x"72",
          9677 => x"70",
          9678 => x"25",
          9679 => x"54",
          9680 => x"38",
          9681 => x"9f",
          9682 => x"2b",
          9683 => x"2e",
          9684 => x"76",
          9685 => x"d1",
          9686 => x"59",
          9687 => x"a7",
          9688 => x"78",
          9689 => x"70",
          9690 => x"32",
          9691 => x"9f",
          9692 => x"56",
          9693 => x"7c",
          9694 => x"38",
          9695 => x"ff",
          9696 => x"dd",
          9697 => x"77",
          9698 => x"76",
          9699 => x"2e",
          9700 => x"80",
          9701 => x"83",
          9702 => x"72",
          9703 => x"56",
          9704 => x"82",
          9705 => x"83",
          9706 => x"53",
          9707 => x"82",
          9708 => x"80",
          9709 => x"77",
          9710 => x"70",
          9711 => x"78",
          9712 => x"38",
          9713 => x"fe",
          9714 => x"17",
          9715 => x"2e",
          9716 => x"14",
          9717 => x"54",
          9718 => x"09",
          9719 => x"38",
          9720 => x"1d",
          9721 => x"74",
          9722 => x"56",
          9723 => x"53",
          9724 => x"72",
          9725 => x"88",
          9726 => x"22",
          9727 => x"57",
          9728 => x"80",
          9729 => x"38",
          9730 => x"83",
          9731 => x"ae",
          9732 => x"70",
          9733 => x"5a",
          9734 => x"2e",
          9735 => x"72",
          9736 => x"72",
          9737 => x"26",
          9738 => x"59",
          9739 => x"70",
          9740 => x"07",
          9741 => x"7c",
          9742 => x"54",
          9743 => x"2e",
          9744 => x"7c",
          9745 => x"83",
          9746 => x"2e",
          9747 => x"83",
          9748 => x"77",
          9749 => x"76",
          9750 => x"8b",
          9751 => x"81",
          9752 => x"18",
          9753 => x"77",
          9754 => x"81",
          9755 => x"53",
          9756 => x"38",
          9757 => x"57",
          9758 => x"2e",
          9759 => x"7c",
          9760 => x"e3",
          9761 => x"06",
          9762 => x"2e",
          9763 => x"7d",
          9764 => x"74",
          9765 => x"e3",
          9766 => x"2a",
          9767 => x"75",
          9768 => x"81",
          9769 => x"80",
          9770 => x"79",
          9771 => x"7d",
          9772 => x"06",
          9773 => x"2e",
          9774 => x"88",
          9775 => x"ab",
          9776 => x"51",
          9777 => x"84",
          9778 => x"ab",
          9779 => x"54",
          9780 => x"08",
          9781 => x"ac",
          9782 => x"c8",
          9783 => x"09",
          9784 => x"f7",
          9785 => x"2a",
          9786 => x"79",
          9787 => x"f0",
          9788 => x"2a",
          9789 => x"78",
          9790 => x"7b",
          9791 => x"56",
          9792 => x"16",
          9793 => x"57",
          9794 => x"81",
          9795 => x"79",
          9796 => x"40",
          9797 => x"7c",
          9798 => x"38",
          9799 => x"fd",
          9800 => x"83",
          9801 => x"8a",
          9802 => x"22",
          9803 => x"2e",
          9804 => x"fc",
          9805 => x"22",
          9806 => x"2e",
          9807 => x"fc",
          9808 => x"10",
          9809 => x"7b",
          9810 => x"a0",
          9811 => x"ae",
          9812 => x"26",
          9813 => x"54",
          9814 => x"81",
          9815 => x"81",
          9816 => x"73",
          9817 => x"79",
          9818 => x"77",
          9819 => x"7b",
          9820 => x"3f",
          9821 => x"08",
          9822 => x"56",
          9823 => x"c8",
          9824 => x"38",
          9825 => x"81",
          9826 => x"fa",
          9827 => x"1c",
          9828 => x"2a",
          9829 => x"5d",
          9830 => x"83",
          9831 => x"1c",
          9832 => x"06",
          9833 => x"d3",
          9834 => x"d2",
          9835 => x"88",
          9836 => x"33",
          9837 => x"54",
          9838 => x"82",
          9839 => x"88",
          9840 => x"08",
          9841 => x"fe",
          9842 => x"22",
          9843 => x"2e",
          9844 => x"76",
          9845 => x"fb",
          9846 => x"ab",
          9847 => x"07",
          9848 => x"5a",
          9849 => x"7d",
          9850 => x"fc",
          9851 => x"06",
          9852 => x"8c",
          9853 => x"06",
          9854 => x"79",
          9855 => x"fd",
          9856 => x"0b",
          9857 => x"7c",
          9858 => x"81",
          9859 => x"38",
          9860 => x"80",
          9861 => x"34",
          9862 => x"b9",
          9863 => x"3d",
          9864 => x"80",
          9865 => x"38",
          9866 => x"27",
          9867 => x"ff",
          9868 => x"7b",
          9869 => x"38",
          9870 => x"7d",
          9871 => x"5c",
          9872 => x"39",
          9873 => x"5a",
          9874 => x"74",
          9875 => x"f6",
          9876 => x"c8",
          9877 => x"ff",
          9878 => x"2a",
          9879 => x"55",
          9880 => x"c4",
          9881 => x"ff",
          9882 => x"d8",
          9883 => x"54",
          9884 => x"26",
          9885 => x"74",
          9886 => x"85",
          9887 => x"f0",
          9888 => x"f0",
          9889 => x"ff",
          9890 => x"59",
          9891 => x"80",
          9892 => x"75",
          9893 => x"81",
          9894 => x"70",
          9895 => x"56",
          9896 => x"ee",
          9897 => x"ff",
          9898 => x"80",
          9899 => x"bf",
          9900 => x"99",
          9901 => x"7d",
          9902 => x"81",
          9903 => x"53",
          9904 => x"59",
          9905 => x"93",
          9906 => x"07",
          9907 => x"06",
          9908 => x"83",
          9909 => x"58",
          9910 => x"7b",
          9911 => x"59",
          9912 => x"81",
          9913 => x"16",
          9914 => x"39",
          9915 => x"b3",
          9916 => x"f0",
          9917 => x"ff",
          9918 => x"78",
          9919 => x"ae",
          9920 => x"7a",
          9921 => x"1d",
          9922 => x"5b",
          9923 => x"34",
          9924 => x"d2",
          9925 => x"14",
          9926 => x"15",
          9927 => x"2b",
          9928 => x"07",
          9929 => x"1f",
          9930 => x"fd",
          9931 => x"1b",
          9932 => x"88",
          9933 => x"72",
          9934 => x"1b",
          9935 => x"05",
          9936 => x"79",
          9937 => x"5b",
          9938 => x"79",
          9939 => x"1d",
          9940 => x"76",
          9941 => x"09",
          9942 => x"a3",
          9943 => x"39",
          9944 => x"81",
          9945 => x"f6",
          9946 => x"0b",
          9947 => x"0c",
          9948 => x"04",
          9949 => x"67",
          9950 => x"05",
          9951 => x"33",
          9952 => x"80",
          9953 => x"7e",
          9954 => x"5b",
          9955 => x"2e",
          9956 => x"79",
          9957 => x"5b",
          9958 => x"26",
          9959 => x"ba",
          9960 => x"38",
          9961 => x"75",
          9962 => x"c7",
          9963 => x"a4",
          9964 => x"76",
          9965 => x"38",
          9966 => x"84",
          9967 => x"70",
          9968 => x"8c",
          9969 => x"2e",
          9970 => x"76",
          9971 => x"81",
          9972 => x"33",
          9973 => x"80",
          9974 => x"81",
          9975 => x"ff",
          9976 => x"84",
          9977 => x"81",
          9978 => x"81",
          9979 => x"7c",
          9980 => x"96",
          9981 => x"34",
          9982 => x"84",
          9983 => x"33",
          9984 => x"81",
          9985 => x"33",
          9986 => x"a4",
          9987 => x"c8",
          9988 => x"06",
          9989 => x"41",
          9990 => x"7f",
          9991 => x"78",
          9992 => x"38",
          9993 => x"81",
          9994 => x"58",
          9995 => x"38",
          9996 => x"83",
          9997 => x"0b",
          9998 => x"7a",
          9999 => x"81",
         10000 => x"b8",
         10001 => x"81",
         10002 => x"58",
         10003 => x"3f",
         10004 => x"08",
         10005 => x"38",
         10006 => x"59",
         10007 => x"0c",
         10008 => x"99",
         10009 => x"17",
         10010 => x"18",
         10011 => x"2b",
         10012 => x"83",
         10013 => x"d4",
         10014 => x"a5",
         10015 => x"26",
         10016 => x"b9",
         10017 => x"42",
         10018 => x"38",
         10019 => x"84",
         10020 => x"38",
         10021 => x"81",
         10022 => x"38",
         10023 => x"33",
         10024 => x"33",
         10025 => x"07",
         10026 => x"84",
         10027 => x"81",
         10028 => x"38",
         10029 => x"33",
         10030 => x"33",
         10031 => x"07",
         10032 => x"a4",
         10033 => x"17",
         10034 => x"82",
         10035 => x"90",
         10036 => x"2b",
         10037 => x"33",
         10038 => x"88",
         10039 => x"71",
         10040 => x"45",
         10041 => x"56",
         10042 => x"0c",
         10043 => x"33",
         10044 => x"80",
         10045 => x"ff",
         10046 => x"ff",
         10047 => x"59",
         10048 => x"81",
         10049 => x"38",
         10050 => x"06",
         10051 => x"80",
         10052 => x"5a",
         10053 => x"8a",
         10054 => x"59",
         10055 => x"87",
         10056 => x"18",
         10057 => x"61",
         10058 => x"80",
         10059 => x"80",
         10060 => x"71",
         10061 => x"56",
         10062 => x"18",
         10063 => x"8f",
         10064 => x"8d",
         10065 => x"98",
         10066 => x"17",
         10067 => x"18",
         10068 => x"2b",
         10069 => x"74",
         10070 => x"d8",
         10071 => x"33",
         10072 => x"71",
         10073 => x"88",
         10074 => x"14",
         10075 => x"07",
         10076 => x"33",
         10077 => x"44",
         10078 => x"42",
         10079 => x"17",
         10080 => x"18",
         10081 => x"2b",
         10082 => x"8d",
         10083 => x"2e",
         10084 => x"7d",
         10085 => x"2a",
         10086 => x"75",
         10087 => x"38",
         10088 => x"7a",
         10089 => x"ed",
         10090 => x"b9",
         10091 => x"84",
         10092 => x"80",
         10093 => x"38",
         10094 => x"08",
         10095 => x"ff",
         10096 => x"38",
         10097 => x"83",
         10098 => x"83",
         10099 => x"75",
         10100 => x"85",
         10101 => x"5d",
         10102 => x"9c",
         10103 => x"a4",
         10104 => x"1d",
         10105 => x"0c",
         10106 => x"1a",
         10107 => x"7c",
         10108 => x"87",
         10109 => x"22",
         10110 => x"7b",
         10111 => x"e0",
         10112 => x"ac",
         10113 => x"19",
         10114 => x"2e",
         10115 => x"10",
         10116 => x"2a",
         10117 => x"05",
         10118 => x"ff",
         10119 => x"59",
         10120 => x"a0",
         10121 => x"b8",
         10122 => x"94",
         10123 => x"0b",
         10124 => x"ff",
         10125 => x"18",
         10126 => x"2e",
         10127 => x"7c",
         10128 => x"d1",
         10129 => x"05",
         10130 => x"d1",
         10131 => x"86",
         10132 => x"d1",
         10133 => x"18",
         10134 => x"98",
         10135 => x"58",
         10136 => x"c8",
         10137 => x"0d",
         10138 => x"84",
         10139 => x"97",
         10140 => x"76",
         10141 => x"70",
         10142 => x"57",
         10143 => x"89",
         10144 => x"82",
         10145 => x"ff",
         10146 => x"5d",
         10147 => x"2e",
         10148 => x"80",
         10149 => x"e5",
         10150 => x"5c",
         10151 => x"5a",
         10152 => x"81",
         10153 => x"79",
         10154 => x"5b",
         10155 => x"12",
         10156 => x"77",
         10157 => x"38",
         10158 => x"81",
         10159 => x"55",
         10160 => x"58",
         10161 => x"89",
         10162 => x"70",
         10163 => x"58",
         10164 => x"70",
         10165 => x"55",
         10166 => x"09",
         10167 => x"38",
         10168 => x"38",
         10169 => x"70",
         10170 => x"07",
         10171 => x"07",
         10172 => x"7a",
         10173 => x"98",
         10174 => x"84",
         10175 => x"83",
         10176 => x"98",
         10177 => x"f9",
         10178 => x"80",
         10179 => x"38",
         10180 => x"81",
         10181 => x"58",
         10182 => x"38",
         10183 => x"c0",
         10184 => x"33",
         10185 => x"81",
         10186 => x"81",
         10187 => x"81",
         10188 => x"eb",
         10189 => x"70",
         10190 => x"07",
         10191 => x"77",
         10192 => x"75",
         10193 => x"83",
         10194 => x"3d",
         10195 => x"83",
         10196 => x"16",
         10197 => x"5b",
         10198 => x"a5",
         10199 => x"16",
         10200 => x"17",
         10201 => x"2b",
         10202 => x"07",
         10203 => x"33",
         10204 => x"88",
         10205 => x"1b",
         10206 => x"52",
         10207 => x"40",
         10208 => x"70",
         10209 => x"0c",
         10210 => x"17",
         10211 => x"80",
         10212 => x"38",
         10213 => x"1d",
         10214 => x"70",
         10215 => x"71",
         10216 => x"71",
         10217 => x"f0",
         10218 => x"1c",
         10219 => x"43",
         10220 => x"08",
         10221 => x"7a",
         10222 => x"fb",
         10223 => x"83",
         10224 => x"0b",
         10225 => x"7a",
         10226 => x"7a",
         10227 => x"38",
         10228 => x"53",
         10229 => x"81",
         10230 => x"ff",
         10231 => x"84",
         10232 => x"76",
         10233 => x"ff",
         10234 => x"74",
         10235 => x"84",
         10236 => x"38",
         10237 => x"7f",
         10238 => x"2b",
         10239 => x"83",
         10240 => x"d4",
         10241 => x"81",
         10242 => x"80",
         10243 => x"33",
         10244 => x"81",
         10245 => x"b7",
         10246 => x"eb",
         10247 => x"70",
         10248 => x"07",
         10249 => x"7f",
         10250 => x"81",
         10251 => x"38",
         10252 => x"81",
         10253 => x"80",
         10254 => x"bd",
         10255 => x"58",
         10256 => x"09",
         10257 => x"38",
         10258 => x"76",
         10259 => x"38",
         10260 => x"f8",
         10261 => x"1a",
         10262 => x"5a",
         10263 => x"fe",
         10264 => x"a8",
         10265 => x"80",
         10266 => x"e4",
         10267 => x"58",
         10268 => x"05",
         10269 => x"70",
         10270 => x"33",
         10271 => x"ff",
         10272 => x"56",
         10273 => x"2e",
         10274 => x"75",
         10275 => x"38",
         10276 => x"8a",
         10277 => x"fc",
         10278 => x"7b",
         10279 => x"5d",
         10280 => x"81",
         10281 => x"71",
         10282 => x"1b",
         10283 => x"40",
         10284 => x"85",
         10285 => x"80",
         10286 => x"82",
         10287 => x"39",
         10288 => x"fa",
         10289 => x"84",
         10290 => x"97",
         10291 => x"75",
         10292 => x"2e",
         10293 => x"85",
         10294 => x"18",
         10295 => x"40",
         10296 => x"b7",
         10297 => x"84",
         10298 => x"97",
         10299 => x"83",
         10300 => x"18",
         10301 => x"5c",
         10302 => x"70",
         10303 => x"33",
         10304 => x"05",
         10305 => x"71",
         10306 => x"5b",
         10307 => x"77",
         10308 => x"d1",
         10309 => x"2e",
         10310 => x"0b",
         10311 => x"83",
         10312 => x"5a",
         10313 => x"81",
         10314 => x"7a",
         10315 => x"5c",
         10316 => x"31",
         10317 => x"58",
         10318 => x"80",
         10319 => x"38",
         10320 => x"e1",
         10321 => x"77",
         10322 => x"59",
         10323 => x"81",
         10324 => x"39",
         10325 => x"33",
         10326 => x"33",
         10327 => x"07",
         10328 => x"81",
         10329 => x"06",
         10330 => x"81",
         10331 => x"5a",
         10332 => x"78",
         10333 => x"83",
         10334 => x"7a",
         10335 => x"81",
         10336 => x"38",
         10337 => x"53",
         10338 => x"81",
         10339 => x"ff",
         10340 => x"84",
         10341 => x"80",
         10342 => x"ff",
         10343 => x"77",
         10344 => x"79",
         10345 => x"79",
         10346 => x"84",
         10347 => x"84",
         10348 => x"71",
         10349 => x"57",
         10350 => x"d4",
         10351 => x"81",
         10352 => x"38",
         10353 => x"11",
         10354 => x"33",
         10355 => x"71",
         10356 => x"81",
         10357 => x"72",
         10358 => x"75",
         10359 => x"5e",
         10360 => x"42",
         10361 => x"84",
         10362 => x"d2",
         10363 => x"06",
         10364 => x"84",
         10365 => x"11",
         10366 => x"33",
         10367 => x"71",
         10368 => x"81",
         10369 => x"72",
         10370 => x"75",
         10371 => x"47",
         10372 => x"5c",
         10373 => x"86",
         10374 => x"f2",
         10375 => x"06",
         10376 => x"84",
         10377 => x"11",
         10378 => x"33",
         10379 => x"71",
         10380 => x"81",
         10381 => x"72",
         10382 => x"75",
         10383 => x"94",
         10384 => x"84",
         10385 => x"11",
         10386 => x"33",
         10387 => x"71",
         10388 => x"81",
         10389 => x"72",
         10390 => x"75",
         10391 => x"62",
         10392 => x"59",
         10393 => x"5c",
         10394 => x"5b",
         10395 => x"77",
         10396 => x"a0",
         10397 => x"5d",
         10398 => x"a0",
         10399 => x"18",
         10400 => x"a8",
         10401 => x"0c",
         10402 => x"18",
         10403 => x"39",
         10404 => x"f8",
         10405 => x"7a",
         10406 => x"f2",
         10407 => x"54",
         10408 => x"53",
         10409 => x"53",
         10410 => x"52",
         10411 => x"b3",
         10412 => x"c8",
         10413 => x"09",
         10414 => x"a4",
         10415 => x"c8",
         10416 => x"34",
         10417 => x"a8",
         10418 => x"40",
         10419 => x"08",
         10420 => x"82",
         10421 => x"60",
         10422 => x"8d",
         10423 => x"c8",
         10424 => x"a0",
         10425 => x"74",
         10426 => x"91",
         10427 => x"81",
         10428 => x"e4",
         10429 => x"58",
         10430 => x"80",
         10431 => x"80",
         10432 => x"71",
         10433 => x"5f",
         10434 => x"7d",
         10435 => x"88",
         10436 => x"61",
         10437 => x"80",
         10438 => x"11",
         10439 => x"33",
         10440 => x"71",
         10441 => x"81",
         10442 => x"72",
         10443 => x"75",
         10444 => x"ac",
         10445 => x"7d",
         10446 => x"43",
         10447 => x"40",
         10448 => x"75",
         10449 => x"2e",
         10450 => x"82",
         10451 => x"39",
         10452 => x"f2",
         10453 => x"3d",
         10454 => x"83",
         10455 => x"39",
         10456 => x"f5",
         10457 => x"bf",
         10458 => x"b4",
         10459 => x"18",
         10460 => x"78",
         10461 => x"33",
         10462 => x"e7",
         10463 => x"39",
         10464 => x"02",
         10465 => x"33",
         10466 => x"93",
         10467 => x"5d",
         10468 => x"40",
         10469 => x"80",
         10470 => x"70",
         10471 => x"33",
         10472 => x"55",
         10473 => x"2e",
         10474 => x"73",
         10475 => x"ba",
         10476 => x"38",
         10477 => x"33",
         10478 => x"24",
         10479 => x"73",
         10480 => x"d1",
         10481 => x"08",
         10482 => x"80",
         10483 => x"80",
         10484 => x"54",
         10485 => x"86",
         10486 => x"34",
         10487 => x"75",
         10488 => x"7c",
         10489 => x"38",
         10490 => x"3d",
         10491 => x"05",
         10492 => x"3f",
         10493 => x"08",
         10494 => x"b9",
         10495 => x"3d",
         10496 => x"0b",
         10497 => x"0c",
         10498 => x"04",
         10499 => x"11",
         10500 => x"06",
         10501 => x"73",
         10502 => x"38",
         10503 => x"81",
         10504 => x"05",
         10505 => x"79",
         10506 => x"38",
         10507 => x"83",
         10508 => x"5f",
         10509 => x"7e",
         10510 => x"70",
         10511 => x"33",
         10512 => x"05",
         10513 => x"9f",
         10514 => x"55",
         10515 => x"89",
         10516 => x"70",
         10517 => x"56",
         10518 => x"16",
         10519 => x"26",
         10520 => x"16",
         10521 => x"06",
         10522 => x"30",
         10523 => x"58",
         10524 => x"2e",
         10525 => x"85",
         10526 => x"be",
         10527 => x"32",
         10528 => x"72",
         10529 => x"79",
         10530 => x"54",
         10531 => x"92",
         10532 => x"84",
         10533 => x"83",
         10534 => x"99",
         10535 => x"fe",
         10536 => x"83",
         10537 => x"7a",
         10538 => x"54",
         10539 => x"e6",
         10540 => x"02",
         10541 => x"fb",
         10542 => x"59",
         10543 => x"80",
         10544 => x"74",
         10545 => x"54",
         10546 => x"05",
         10547 => x"84",
         10548 => x"ed",
         10549 => x"b9",
         10550 => x"84",
         10551 => x"80",
         10552 => x"80",
         10553 => x"56",
         10554 => x"c8",
         10555 => x"0d",
         10556 => x"6d",
         10557 => x"70",
         10558 => x"9a",
         10559 => x"c8",
         10560 => x"b9",
         10561 => x"2e",
         10562 => x"77",
         10563 => x"7c",
         10564 => x"ca",
         10565 => x"2e",
         10566 => x"76",
         10567 => x"ea",
         10568 => x"07",
         10569 => x"bb",
         10570 => x"2a",
         10571 => x"7a",
         10572 => x"d1",
         10573 => x"11",
         10574 => x"33",
         10575 => x"07",
         10576 => x"42",
         10577 => x"56",
         10578 => x"84",
         10579 => x"0b",
         10580 => x"80",
         10581 => x"34",
         10582 => x"17",
         10583 => x"0b",
         10584 => x"66",
         10585 => x"8b",
         10586 => x"67",
         10587 => x"0b",
         10588 => x"80",
         10589 => x"34",
         10590 => x"7c",
         10591 => x"a9",
         10592 => x"80",
         10593 => x"34",
         10594 => x"1c",
         10595 => x"9e",
         10596 => x"0b",
         10597 => x"7e",
         10598 => x"83",
         10599 => x"80",
         10600 => x"38",
         10601 => x"08",
         10602 => x"53",
         10603 => x"81",
         10604 => x"38",
         10605 => x"7c",
         10606 => x"38",
         10607 => x"79",
         10608 => x"39",
         10609 => x"05",
         10610 => x"2b",
         10611 => x"80",
         10612 => x"38",
         10613 => x"06",
         10614 => x"fe",
         10615 => x"fe",
         10616 => x"80",
         10617 => x"70",
         10618 => x"06",
         10619 => x"82",
         10620 => x"81",
         10621 => x"5e",
         10622 => x"89",
         10623 => x"06",
         10624 => x"f6",
         10625 => x"2a",
         10626 => x"75",
         10627 => x"38",
         10628 => x"07",
         10629 => x"11",
         10630 => x"0c",
         10631 => x"0c",
         10632 => x"33",
         10633 => x"71",
         10634 => x"73",
         10635 => x"40",
         10636 => x"83",
         10637 => x"38",
         10638 => x"0c",
         10639 => x"11",
         10640 => x"33",
         10641 => x"71",
         10642 => x"81",
         10643 => x"72",
         10644 => x"75",
         10645 => x"70",
         10646 => x"0c",
         10647 => x"51",
         10648 => x"57",
         10649 => x"1a",
         10650 => x"23",
         10651 => x"34",
         10652 => x"1a",
         10653 => x"9c",
         10654 => x"85",
         10655 => x"55",
         10656 => x"84",
         10657 => x"80",
         10658 => x"38",
         10659 => x"0c",
         10660 => x"70",
         10661 => x"52",
         10662 => x"30",
         10663 => x"80",
         10664 => x"79",
         10665 => x"92",
         10666 => x"76",
         10667 => x"7d",
         10668 => x"86",
         10669 => x"78",
         10670 => x"db",
         10671 => x"c8",
         10672 => x"b9",
         10673 => x"26",
         10674 => x"57",
         10675 => x"08",
         10676 => x"cb",
         10677 => x"31",
         10678 => x"02",
         10679 => x"33",
         10680 => x"7d",
         10681 => x"82",
         10682 => x"55",
         10683 => x"fc",
         10684 => x"57",
         10685 => x"fb",
         10686 => x"57",
         10687 => x"fb",
         10688 => x"57",
         10689 => x"fb",
         10690 => x"51",
         10691 => x"84",
         10692 => x"78",
         10693 => x"57",
         10694 => x"38",
         10695 => x"7a",
         10696 => x"57",
         10697 => x"39",
         10698 => x"94",
         10699 => x"98",
         10700 => x"2b",
         10701 => x"5d",
         10702 => x"fc",
         10703 => x"7c",
         10704 => x"bd",
         10705 => x"79",
         10706 => x"cb",
         10707 => x"c8",
         10708 => x"b9",
         10709 => x"2e",
         10710 => x"84",
         10711 => x"81",
         10712 => x"38",
         10713 => x"08",
         10714 => x"99",
         10715 => x"74",
         10716 => x"ff",
         10717 => x"84",
         10718 => x"83",
         10719 => x"17",
         10720 => x"94",
         10721 => x"56",
         10722 => x"27",
         10723 => x"81",
         10724 => x"0c",
         10725 => x"81",
         10726 => x"84",
         10727 => x"55",
         10728 => x"ff",
         10729 => x"d9",
         10730 => x"94",
         10731 => x"0b",
         10732 => x"fb",
         10733 => x"16",
         10734 => x"33",
         10735 => x"71",
         10736 => x"7e",
         10737 => x"5b",
         10738 => x"17",
         10739 => x"8f",
         10740 => x"0b",
         10741 => x"80",
         10742 => x"17",
         10743 => x"a0",
         10744 => x"34",
         10745 => x"5e",
         10746 => x"17",
         10747 => x"9b",
         10748 => x"33",
         10749 => x"2e",
         10750 => x"fb",
         10751 => x"a9",
         10752 => x"7f",
         10753 => x"57",
         10754 => x"08",
         10755 => x"38",
         10756 => x"5a",
         10757 => x"09",
         10758 => x"38",
         10759 => x"53",
         10760 => x"81",
         10761 => x"ff",
         10762 => x"84",
         10763 => x"80",
         10764 => x"ff",
         10765 => x"76",
         10766 => x"7e",
         10767 => x"1d",
         10768 => x"57",
         10769 => x"fb",
         10770 => x"79",
         10771 => x"39",
         10772 => x"16",
         10773 => x"16",
         10774 => x"17",
         10775 => x"ff",
         10776 => x"84",
         10777 => x"7d",
         10778 => x"06",
         10779 => x"84",
         10780 => x"83",
         10781 => x"16",
         10782 => x"08",
         10783 => x"c8",
         10784 => x"74",
         10785 => x"27",
         10786 => x"82",
         10787 => x"74",
         10788 => x"81",
         10789 => x"38",
         10790 => x"16",
         10791 => x"08",
         10792 => x"52",
         10793 => x"51",
         10794 => x"3f",
         10795 => x"ec",
         10796 => x"1a",
         10797 => x"f8",
         10798 => x"98",
         10799 => x"f8",
         10800 => x"83",
         10801 => x"79",
         10802 => x"9a",
         10803 => x"19",
         10804 => x"fe",
         10805 => x"5a",
         10806 => x"f9",
         10807 => x"1a",
         10808 => x"29",
         10809 => x"05",
         10810 => x"80",
         10811 => x"38",
         10812 => x"15",
         10813 => x"76",
         10814 => x"39",
         10815 => x"0c",
         10816 => x"e4",
         10817 => x"80",
         10818 => x"da",
         10819 => x"c8",
         10820 => x"79",
         10821 => x"39",
         10822 => x"5b",
         10823 => x"f0",
         10824 => x"65",
         10825 => x"40",
         10826 => x"7e",
         10827 => x"79",
         10828 => x"38",
         10829 => x"75",
         10830 => x"38",
         10831 => x"74",
         10832 => x"38",
         10833 => x"84",
         10834 => x"59",
         10835 => x"84",
         10836 => x"55",
         10837 => x"55",
         10838 => x"38",
         10839 => x"55",
         10840 => x"38",
         10841 => x"81",
         10842 => x"56",
         10843 => x"81",
         10844 => x"1a",
         10845 => x"08",
         10846 => x"56",
         10847 => x"81",
         10848 => x"80",
         10849 => x"38",
         10850 => x"83",
         10851 => x"7a",
         10852 => x"8a",
         10853 => x"05",
         10854 => x"06",
         10855 => x"38",
         10856 => x"38",
         10857 => x"55",
         10858 => x"84",
         10859 => x"ff",
         10860 => x"38",
         10861 => x"0c",
         10862 => x"1a",
         10863 => x"9c",
         10864 => x"05",
         10865 => x"60",
         10866 => x"38",
         10867 => x"70",
         10868 => x"1b",
         10869 => x"56",
         10870 => x"83",
         10871 => x"15",
         10872 => x"59",
         10873 => x"2e",
         10874 => x"77",
         10875 => x"75",
         10876 => x"75",
         10877 => x"77",
         10878 => x"7c",
         10879 => x"33",
         10880 => x"e0",
         10881 => x"c8",
         10882 => x"38",
         10883 => x"33",
         10884 => x"80",
         10885 => x"b4",
         10886 => x"31",
         10887 => x"27",
         10888 => x"80",
         10889 => x"1e",
         10890 => x"58",
         10891 => x"81",
         10892 => x"77",
         10893 => x"59",
         10894 => x"55",
         10895 => x"77",
         10896 => x"7b",
         10897 => x"08",
         10898 => x"78",
         10899 => x"08",
         10900 => x"94",
         10901 => x"5c",
         10902 => x"38",
         10903 => x"84",
         10904 => x"92",
         10905 => x"74",
         10906 => x"0c",
         10907 => x"04",
         10908 => x"8e",
         10909 => x"08",
         10910 => x"ff",
         10911 => x"71",
         10912 => x"7b",
         10913 => x"38",
         10914 => x"56",
         10915 => x"77",
         10916 => x"80",
         10917 => x"33",
         10918 => x"5f",
         10919 => x"09",
         10920 => x"e4",
         10921 => x"76",
         10922 => x"52",
         10923 => x"51",
         10924 => x"3f",
         10925 => x"08",
         10926 => x"38",
         10927 => x"5b",
         10928 => x"0c",
         10929 => x"38",
         10930 => x"08",
         10931 => x"11",
         10932 => x"58",
         10933 => x"59",
         10934 => x"fe",
         10935 => x"70",
         10936 => x"33",
         10937 => x"05",
         10938 => x"16",
         10939 => x"2e",
         10940 => x"74",
         10941 => x"56",
         10942 => x"81",
         10943 => x"ff",
         10944 => x"da",
         10945 => x"39",
         10946 => x"19",
         10947 => x"19",
         10948 => x"1a",
         10949 => x"ff",
         10950 => x"81",
         10951 => x"c8",
         10952 => x"09",
         10953 => x"9c",
         10954 => x"c8",
         10955 => x"34",
         10956 => x"a8",
         10957 => x"84",
         10958 => x"5c",
         10959 => x"1a",
         10960 => x"e1",
         10961 => x"33",
         10962 => x"2e",
         10963 => x"fe",
         10964 => x"54",
         10965 => x"a0",
         10966 => x"53",
         10967 => x"19",
         10968 => x"9d",
         10969 => x"5b",
         10970 => x"76",
         10971 => x"94",
         10972 => x"fe",
         10973 => x"1a",
         10974 => x"51",
         10975 => x"3f",
         10976 => x"08",
         10977 => x"39",
         10978 => x"51",
         10979 => x"3f",
         10980 => x"08",
         10981 => x"74",
         10982 => x"74",
         10983 => x"57",
         10984 => x"81",
         10985 => x"34",
         10986 => x"b9",
         10987 => x"3d",
         10988 => x"0b",
         10989 => x"82",
         10990 => x"c8",
         10991 => x"0d",
         10992 => x"0d",
         10993 => x"66",
         10994 => x"5a",
         10995 => x"89",
         10996 => x"2e",
         10997 => x"08",
         10998 => x"2e",
         10999 => x"33",
         11000 => x"2e",
         11001 => x"16",
         11002 => x"22",
         11003 => x"78",
         11004 => x"38",
         11005 => x"41",
         11006 => x"82",
         11007 => x"1a",
         11008 => x"82",
         11009 => x"1a",
         11010 => x"2a",
         11011 => x"58",
         11012 => x"80",
         11013 => x"38",
         11014 => x"7b",
         11015 => x"7b",
         11016 => x"38",
         11017 => x"7a",
         11018 => x"81",
         11019 => x"ff",
         11020 => x"82",
         11021 => x"8a",
         11022 => x"05",
         11023 => x"06",
         11024 => x"aa",
         11025 => x"9e",
         11026 => x"08",
         11027 => x"2e",
         11028 => x"74",
         11029 => x"a1",
         11030 => x"2e",
         11031 => x"74",
         11032 => x"88",
         11033 => x"38",
         11034 => x"0c",
         11035 => x"16",
         11036 => x"08",
         11037 => x"38",
         11038 => x"fe",
         11039 => x"08",
         11040 => x"58",
         11041 => x"85",
         11042 => x"16",
         11043 => x"29",
         11044 => x"05",
         11045 => x"80",
         11046 => x"38",
         11047 => x"89",
         11048 => x"77",
         11049 => x"98",
         11050 => x"5f",
         11051 => x"85",
         11052 => x"31",
         11053 => x"7b",
         11054 => x"81",
         11055 => x"ff",
         11056 => x"84",
         11057 => x"85",
         11058 => x"b4",
         11059 => x"31",
         11060 => x"78",
         11061 => x"84",
         11062 => x"18",
         11063 => x"1f",
         11064 => x"74",
         11065 => x"56",
         11066 => x"81",
         11067 => x"ff",
         11068 => x"ef",
         11069 => x"75",
         11070 => x"77",
         11071 => x"7a",
         11072 => x"08",
         11073 => x"79",
         11074 => x"08",
         11075 => x"94",
         11076 => x"1e",
         11077 => x"57",
         11078 => x"75",
         11079 => x"74",
         11080 => x"1b",
         11081 => x"85",
         11082 => x"33",
         11083 => x"c0",
         11084 => x"90",
         11085 => x"56",
         11086 => x"c8",
         11087 => x"0d",
         11088 => x"b9",
         11089 => x"3d",
         11090 => x"16",
         11091 => x"82",
         11092 => x"56",
         11093 => x"60",
         11094 => x"59",
         11095 => x"ff",
         11096 => x"71",
         11097 => x"7a",
         11098 => x"38",
         11099 => x"57",
         11100 => x"78",
         11101 => x"80",
         11102 => x"33",
         11103 => x"5f",
         11104 => x"09",
         11105 => x"d5",
         11106 => x"77",
         11107 => x"52",
         11108 => x"51",
         11109 => x"3f",
         11110 => x"08",
         11111 => x"38",
         11112 => x"5c",
         11113 => x"0c",
         11114 => x"38",
         11115 => x"08",
         11116 => x"11",
         11117 => x"05",
         11118 => x"58",
         11119 => x"95",
         11120 => x"81",
         11121 => x"75",
         11122 => x"57",
         11123 => x"56",
         11124 => x"60",
         11125 => x"83",
         11126 => x"a3",
         11127 => x"b4",
         11128 => x"b8",
         11129 => x"81",
         11130 => x"40",
         11131 => x"3f",
         11132 => x"b9",
         11133 => x"2e",
         11134 => x"ff",
         11135 => x"b9",
         11136 => x"17",
         11137 => x"08",
         11138 => x"31",
         11139 => x"08",
         11140 => x"a0",
         11141 => x"fe",
         11142 => x"16",
         11143 => x"82",
         11144 => x"06",
         11145 => x"81",
         11146 => x"08",
         11147 => x"05",
         11148 => x"81",
         11149 => x"ff",
         11150 => x"7e",
         11151 => x"39",
         11152 => x"57",
         11153 => x"77",
         11154 => x"83",
         11155 => x"7f",
         11156 => x"60",
         11157 => x"0c",
         11158 => x"58",
         11159 => x"9c",
         11160 => x"fd",
         11161 => x"1a",
         11162 => x"51",
         11163 => x"3f",
         11164 => x"08",
         11165 => x"c8",
         11166 => x"38",
         11167 => x"58",
         11168 => x"76",
         11169 => x"ff",
         11170 => x"84",
         11171 => x"55",
         11172 => x"08",
         11173 => x"e4",
         11174 => x"b4",
         11175 => x"b8",
         11176 => x"81",
         11177 => x"57",
         11178 => x"3f",
         11179 => x"08",
         11180 => x"84",
         11181 => x"83",
         11182 => x"16",
         11183 => x"08",
         11184 => x"a0",
         11185 => x"fd",
         11186 => x"16",
         11187 => x"82",
         11188 => x"06",
         11189 => x"81",
         11190 => x"08",
         11191 => x"05",
         11192 => x"81",
         11193 => x"ff",
         11194 => x"60",
         11195 => x"39",
         11196 => x"51",
         11197 => x"3f",
         11198 => x"08",
         11199 => x"74",
         11200 => x"74",
         11201 => x"57",
         11202 => x"81",
         11203 => x"08",
         11204 => x"70",
         11205 => x"33",
         11206 => x"96",
         11207 => x"b9",
         11208 => x"c6",
         11209 => x"c8",
         11210 => x"34",
         11211 => x"a8",
         11212 => x"55",
         11213 => x"08",
         11214 => x"38",
         11215 => x"58",
         11216 => x"09",
         11217 => x"8b",
         11218 => x"b4",
         11219 => x"17",
         11220 => x"76",
         11221 => x"33",
         11222 => x"87",
         11223 => x"b4",
         11224 => x"1b",
         11225 => x"fd",
         11226 => x"0b",
         11227 => x"81",
         11228 => x"c8",
         11229 => x"0d",
         11230 => x"91",
         11231 => x"0b",
         11232 => x"0c",
         11233 => x"04",
         11234 => x"7d",
         11235 => x"77",
         11236 => x"38",
         11237 => x"75",
         11238 => x"38",
         11239 => x"74",
         11240 => x"38",
         11241 => x"84",
         11242 => x"59",
         11243 => x"83",
         11244 => x"55",
         11245 => x"56",
         11246 => x"38",
         11247 => x"70",
         11248 => x"06",
         11249 => x"80",
         11250 => x"38",
         11251 => x"08",
         11252 => x"17",
         11253 => x"ac",
         11254 => x"33",
         11255 => x"bc",
         11256 => x"78",
         11257 => x"52",
         11258 => x"51",
         11259 => x"3f",
         11260 => x"08",
         11261 => x"38",
         11262 => x"56",
         11263 => x"0c",
         11264 => x"38",
         11265 => x"8b",
         11266 => x"07",
         11267 => x"8b",
         11268 => x"08",
         11269 => x"70",
         11270 => x"06",
         11271 => x"7a",
         11272 => x"7a",
         11273 => x"79",
         11274 => x"9c",
         11275 => x"96",
         11276 => x"5b",
         11277 => x"81",
         11278 => x"18",
         11279 => x"7b",
         11280 => x"2a",
         11281 => x"18",
         11282 => x"2a",
         11283 => x"18",
         11284 => x"2a",
         11285 => x"18",
         11286 => x"34",
         11287 => x"18",
         11288 => x"98",
         11289 => x"cc",
         11290 => x"34",
         11291 => x"18",
         11292 => x"93",
         11293 => x"5b",
         11294 => x"1c",
         11295 => x"ff",
         11296 => x"84",
         11297 => x"90",
         11298 => x"bf",
         11299 => x"79",
         11300 => x"75",
         11301 => x"0c",
         11302 => x"04",
         11303 => x"17",
         11304 => x"17",
         11305 => x"18",
         11306 => x"ff",
         11307 => x"81",
         11308 => x"c8",
         11309 => x"38",
         11310 => x"08",
         11311 => x"b4",
         11312 => x"18",
         11313 => x"b9",
         11314 => x"55",
         11315 => x"08",
         11316 => x"38",
         11317 => x"55",
         11318 => x"09",
         11319 => x"81",
         11320 => x"b4",
         11321 => x"18",
         11322 => x"7a",
         11323 => x"33",
         11324 => x"ef",
         11325 => x"fd",
         11326 => x"90",
         11327 => x"94",
         11328 => x"88",
         11329 => x"95",
         11330 => x"18",
         11331 => x"7b",
         11332 => x"2a",
         11333 => x"18",
         11334 => x"2a",
         11335 => x"18",
         11336 => x"2a",
         11337 => x"18",
         11338 => x"34",
         11339 => x"18",
         11340 => x"98",
         11341 => x"cc",
         11342 => x"34",
         11343 => x"18",
         11344 => x"93",
         11345 => x"5b",
         11346 => x"1c",
         11347 => x"ff",
         11348 => x"84",
         11349 => x"90",
         11350 => x"bf",
         11351 => x"79",
         11352 => x"fe",
         11353 => x"16",
         11354 => x"90",
         11355 => x"b9",
         11356 => x"06",
         11357 => x"ba",
         11358 => x"08",
         11359 => x"b4",
         11360 => x"0d",
         11361 => x"55",
         11362 => x"84",
         11363 => x"54",
         11364 => x"08",
         11365 => x"56",
         11366 => x"9e",
         11367 => x"53",
         11368 => x"96",
         11369 => x"52",
         11370 => x"8e",
         11371 => x"22",
         11372 => x"58",
         11373 => x"2e",
         11374 => x"52",
         11375 => x"54",
         11376 => x"75",
         11377 => x"84",
         11378 => x"89",
         11379 => x"81",
         11380 => x"ff",
         11381 => x"84",
         11382 => x"81",
         11383 => x"da",
         11384 => x"08",
         11385 => x"39",
         11386 => x"ff",
         11387 => x"57",
         11388 => x"2e",
         11389 => x"70",
         11390 => x"33",
         11391 => x"52",
         11392 => x"2e",
         11393 => x"ee",
         11394 => x"2e",
         11395 => x"d1",
         11396 => x"80",
         11397 => x"38",
         11398 => x"a4",
         11399 => x"84",
         11400 => x"8c",
         11401 => x"8b",
         11402 => x"c8",
         11403 => x"0d",
         11404 => x"d0",
         11405 => x"ff",
         11406 => x"53",
         11407 => x"91",
         11408 => x"73",
         11409 => x"d0",
         11410 => x"73",
         11411 => x"f5",
         11412 => x"83",
         11413 => x"58",
         11414 => x"56",
         11415 => x"81",
         11416 => x"75",
         11417 => x"57",
         11418 => x"12",
         11419 => x"70",
         11420 => x"38",
         11421 => x"81",
         11422 => x"54",
         11423 => x"51",
         11424 => x"89",
         11425 => x"70",
         11426 => x"54",
         11427 => x"70",
         11428 => x"51",
         11429 => x"09",
         11430 => x"38",
         11431 => x"38",
         11432 => x"70",
         11433 => x"07",
         11434 => x"07",
         11435 => x"76",
         11436 => x"38",
         11437 => x"1b",
         11438 => x"78",
         11439 => x"38",
         11440 => x"cf",
         11441 => x"24",
         11442 => x"76",
         11443 => x"c3",
         11444 => x"0d",
         11445 => x"3d",
         11446 => x"99",
         11447 => x"94",
         11448 => x"c8",
         11449 => x"b9",
         11450 => x"2e",
         11451 => x"84",
         11452 => x"98",
         11453 => x"7a",
         11454 => x"98",
         11455 => x"51",
         11456 => x"84",
         11457 => x"55",
         11458 => x"08",
         11459 => x"02",
         11460 => x"33",
         11461 => x"58",
         11462 => x"24",
         11463 => x"02",
         11464 => x"70",
         11465 => x"06",
         11466 => x"80",
         11467 => x"7a",
         11468 => x"33",
         11469 => x"71",
         11470 => x"73",
         11471 => x"5b",
         11472 => x"83",
         11473 => x"76",
         11474 => x"74",
         11475 => x"0c",
         11476 => x"04",
         11477 => x"08",
         11478 => x"81",
         11479 => x"38",
         11480 => x"b9",
         11481 => x"3d",
         11482 => x"16",
         11483 => x"33",
         11484 => x"71",
         11485 => x"79",
         11486 => x"0c",
         11487 => x"39",
         11488 => x"12",
         11489 => x"84",
         11490 => x"98",
         11491 => x"ff",
         11492 => x"80",
         11493 => x"80",
         11494 => x"5d",
         11495 => x"34",
         11496 => x"e4",
         11497 => x"05",
         11498 => x"3d",
         11499 => x"3f",
         11500 => x"08",
         11501 => x"c8",
         11502 => x"38",
         11503 => x"3d",
         11504 => x"98",
         11505 => x"dd",
         11506 => x"80",
         11507 => x"5b",
         11508 => x"2e",
         11509 => x"80",
         11510 => x"3d",
         11511 => x"52",
         11512 => x"a4",
         11513 => x"b9",
         11514 => x"84",
         11515 => x"83",
         11516 => x"80",
         11517 => x"58",
         11518 => x"08",
         11519 => x"38",
         11520 => x"08",
         11521 => x"5f",
         11522 => x"c7",
         11523 => x"76",
         11524 => x"52",
         11525 => x"51",
         11526 => x"3f",
         11527 => x"08",
         11528 => x"38",
         11529 => x"59",
         11530 => x"0c",
         11531 => x"38",
         11532 => x"08",
         11533 => x"9a",
         11534 => x"88",
         11535 => x"70",
         11536 => x"59",
         11537 => x"83",
         11538 => x"38",
         11539 => x"3d",
         11540 => x"7a",
         11541 => x"b7",
         11542 => x"c8",
         11543 => x"b9",
         11544 => x"9f",
         11545 => x"7a",
         11546 => x"f5",
         11547 => x"c8",
         11548 => x"b9",
         11549 => x"38",
         11550 => x"08",
         11551 => x"9a",
         11552 => x"88",
         11553 => x"70",
         11554 => x"59",
         11555 => x"83",
         11556 => x"38",
         11557 => x"a4",
         11558 => x"c8",
         11559 => x"51",
         11560 => x"3f",
         11561 => x"08",
         11562 => x"c8",
         11563 => x"ff",
         11564 => x"84",
         11565 => x"38",
         11566 => x"38",
         11567 => x"fd",
         11568 => x"7a",
         11569 => x"89",
         11570 => x"82",
         11571 => x"57",
         11572 => x"90",
         11573 => x"56",
         11574 => x"17",
         11575 => x"57",
         11576 => x"38",
         11577 => x"75",
         11578 => x"95",
         11579 => x"2e",
         11580 => x"17",
         11581 => x"ff",
         11582 => x"3d",
         11583 => x"19",
         11584 => x"59",
         11585 => x"33",
         11586 => x"eb",
         11587 => x"80",
         11588 => x"11",
         11589 => x"7e",
         11590 => x"3d",
         11591 => x"fd",
         11592 => x"60",
         11593 => x"38",
         11594 => x"d1",
         11595 => x"10",
         11596 => x"b8",
         11597 => x"70",
         11598 => x"59",
         11599 => x"7a",
         11600 => x"81",
         11601 => x"70",
         11602 => x"5a",
         11603 => x"82",
         11604 => x"78",
         11605 => x"80",
         11606 => x"27",
         11607 => x"16",
         11608 => x"7c",
         11609 => x"5e",
         11610 => x"57",
         11611 => x"ee",
         11612 => x"70",
         11613 => x"34",
         11614 => x"09",
         11615 => x"df",
         11616 => x"80",
         11617 => x"84",
         11618 => x"80",
         11619 => x"04",
         11620 => x"94",
         11621 => x"98",
         11622 => x"2b",
         11623 => x"59",
         11624 => x"f0",
         11625 => x"33",
         11626 => x"71",
         11627 => x"90",
         11628 => x"07",
         11629 => x"0c",
         11630 => x"52",
         11631 => x"a0",
         11632 => x"b9",
         11633 => x"84",
         11634 => x"80",
         11635 => x"38",
         11636 => x"81",
         11637 => x"08",
         11638 => x"70",
         11639 => x"33",
         11640 => x"88",
         11641 => x"59",
         11642 => x"08",
         11643 => x"84",
         11644 => x"83",
         11645 => x"16",
         11646 => x"08",
         11647 => x"c8",
         11648 => x"74",
         11649 => x"27",
         11650 => x"82",
         11651 => x"74",
         11652 => x"81",
         11653 => x"38",
         11654 => x"16",
         11655 => x"08",
         11656 => x"52",
         11657 => x"51",
         11658 => x"3f",
         11659 => x"dd",
         11660 => x"80",
         11661 => x"11",
         11662 => x"7b",
         11663 => x"84",
         11664 => x"70",
         11665 => x"e5",
         11666 => x"08",
         11667 => x"59",
         11668 => x"7e",
         11669 => x"81",
         11670 => x"38",
         11671 => x"80",
         11672 => x"18",
         11673 => x"5a",
         11674 => x"70",
         11675 => x"34",
         11676 => x"fe",
         11677 => x"e5",
         11678 => x"81",
         11679 => x"79",
         11680 => x"81",
         11681 => x"7f",
         11682 => x"38",
         11683 => x"82",
         11684 => x"34",
         11685 => x"c8",
         11686 => x"3d",
         11687 => x"3d",
         11688 => x"58",
         11689 => x"74",
         11690 => x"38",
         11691 => x"73",
         11692 => x"38",
         11693 => x"72",
         11694 => x"38",
         11695 => x"84",
         11696 => x"59",
         11697 => x"83",
         11698 => x"53",
         11699 => x"53",
         11700 => x"38",
         11701 => x"53",
         11702 => x"38",
         11703 => x"56",
         11704 => x"81",
         11705 => x"15",
         11706 => x"58",
         11707 => x"81",
         11708 => x"8a",
         11709 => x"89",
         11710 => x"56",
         11711 => x"81",
         11712 => x"52",
         11713 => x"fd",
         11714 => x"84",
         11715 => x"ff",
         11716 => x"70",
         11717 => x"fd",
         11718 => x"84",
         11719 => x"73",
         11720 => x"38",
         11721 => x"06",
         11722 => x"0c",
         11723 => x"98",
         11724 => x"58",
         11725 => x"2e",
         11726 => x"75",
         11727 => x"d9",
         11728 => x"31",
         11729 => x"17",
         11730 => x"90",
         11731 => x"81",
         11732 => x"51",
         11733 => x"80",
         11734 => x"38",
         11735 => x"51",
         11736 => x"3f",
         11737 => x"08",
         11738 => x"c8",
         11739 => x"81",
         11740 => x"ff",
         11741 => x"81",
         11742 => x"b4",
         11743 => x"73",
         11744 => x"27",
         11745 => x"73",
         11746 => x"ff",
         11747 => x"0b",
         11748 => x"81",
         11749 => x"b9",
         11750 => x"3d",
         11751 => x"15",
         11752 => x"2a",
         11753 => x"58",
         11754 => x"38",
         11755 => x"08",
         11756 => x"58",
         11757 => x"09",
         11758 => x"b6",
         11759 => x"16",
         11760 => x"08",
         11761 => x"27",
         11762 => x"8c",
         11763 => x"15",
         11764 => x"07",
         11765 => x"16",
         11766 => x"ff",
         11767 => x"80",
         11768 => x"9c",
         11769 => x"2e",
         11770 => x"9c",
         11771 => x"0b",
         11772 => x"0c",
         11773 => x"04",
         11774 => x"16",
         11775 => x"08",
         11776 => x"2e",
         11777 => x"73",
         11778 => x"73",
         11779 => x"c2",
         11780 => x"39",
         11781 => x"08",
         11782 => x"08",
         11783 => x"0c",
         11784 => x"06",
         11785 => x"2e",
         11786 => x"fe",
         11787 => x"08",
         11788 => x"55",
         11789 => x"27",
         11790 => x"8a",
         11791 => x"71",
         11792 => x"08",
         11793 => x"2a",
         11794 => x"53",
         11795 => x"80",
         11796 => x"15",
         11797 => x"e9",
         11798 => x"74",
         11799 => x"b7",
         11800 => x"c8",
         11801 => x"8a",
         11802 => x"33",
         11803 => x"a2",
         11804 => x"c8",
         11805 => x"53",
         11806 => x"38",
         11807 => x"54",
         11808 => x"39",
         11809 => x"51",
         11810 => x"3f",
         11811 => x"08",
         11812 => x"c8",
         11813 => x"98",
         11814 => x"c8",
         11815 => x"fd",
         11816 => x"b9",
         11817 => x"16",
         11818 => x"16",
         11819 => x"39",
         11820 => x"16",
         11821 => x"84",
         11822 => x"8b",
         11823 => x"f6",
         11824 => x"56",
         11825 => x"80",
         11826 => x"80",
         11827 => x"fc",
         11828 => x"3d",
         11829 => x"c5",
         11830 => x"b9",
         11831 => x"84",
         11832 => x"80",
         11833 => x"80",
         11834 => x"54",
         11835 => x"c8",
         11836 => x"0d",
         11837 => x"0c",
         11838 => x"51",
         11839 => x"3f",
         11840 => x"08",
         11841 => x"c8",
         11842 => x"38",
         11843 => x"70",
         11844 => x"59",
         11845 => x"af",
         11846 => x"33",
         11847 => x"81",
         11848 => x"79",
         11849 => x"c5",
         11850 => x"08",
         11851 => x"9a",
         11852 => x"88",
         11853 => x"70",
         11854 => x"5a",
         11855 => x"83",
         11856 => x"77",
         11857 => x"7a",
         11858 => x"22",
         11859 => x"74",
         11860 => x"ff",
         11861 => x"84",
         11862 => x"55",
         11863 => x"8d",
         11864 => x"2e",
         11865 => x"80",
         11866 => x"fe",
         11867 => x"80",
         11868 => x"f6",
         11869 => x"33",
         11870 => x"71",
         11871 => x"90",
         11872 => x"07",
         11873 => x"5a",
         11874 => x"39",
         11875 => x"78",
         11876 => x"74",
         11877 => x"38",
         11878 => x"72",
         11879 => x"38",
         11880 => x"71",
         11881 => x"38",
         11882 => x"84",
         11883 => x"52",
         11884 => x"94",
         11885 => x"71",
         11886 => x"38",
         11887 => x"73",
         11888 => x"0c",
         11889 => x"04",
         11890 => x"51",
         11891 => x"3f",
         11892 => x"08",
         11893 => x"71",
         11894 => x"75",
         11895 => x"d7",
         11896 => x"0d",
         11897 => x"55",
         11898 => x"80",
         11899 => x"74",
         11900 => x"80",
         11901 => x"73",
         11902 => x"80",
         11903 => x"86",
         11904 => x"16",
         11905 => x"72",
         11906 => x"97",
         11907 => x"72",
         11908 => x"75",
         11909 => x"76",
         11910 => x"f3",
         11911 => x"74",
         11912 => x"bd",
         11913 => x"c8",
         11914 => x"b9",
         11915 => x"2e",
         11916 => x"b9",
         11917 => x"38",
         11918 => x"51",
         11919 => x"3f",
         11920 => x"51",
         11921 => x"3f",
         11922 => x"08",
         11923 => x"30",
         11924 => x"9f",
         11925 => x"c8",
         11926 => x"57",
         11927 => x"b9",
         11928 => x"3d",
         11929 => x"77",
         11930 => x"53",
         11931 => x"3f",
         11932 => x"51",
         11933 => x"3f",
         11934 => x"08",
         11935 => x"30",
         11936 => x"9f",
         11937 => x"c8",
         11938 => x"57",
         11939 => x"75",
         11940 => x"ff",
         11941 => x"84",
         11942 => x"84",
         11943 => x"8a",
         11944 => x"81",
         11945 => x"fe",
         11946 => x"84",
         11947 => x"81",
         11948 => x"fe",
         11949 => x"75",
         11950 => x"fe",
         11951 => x"3d",
         11952 => x"80",
         11953 => x"70",
         11954 => x"52",
         11955 => x"3f",
         11956 => x"08",
         11957 => x"c8",
         11958 => x"8a",
         11959 => x"b9",
         11960 => x"3d",
         11961 => x"52",
         11962 => x"b5",
         11963 => x"b9",
         11964 => x"84",
         11965 => x"e5",
         11966 => x"cb",
         11967 => x"98",
         11968 => x"80",
         11969 => x"38",
         11970 => x"d1",
         11971 => x"75",
         11972 => x"bd",
         11973 => x"b9",
         11974 => x"3d",
         11975 => x"0b",
         11976 => x"0c",
         11977 => x"04",
         11978 => x"66",
         11979 => x"80",
         11980 => x"ec",
         11981 => x"3d",
         11982 => x"3f",
         11983 => x"08",
         11984 => x"c8",
         11985 => x"7f",
         11986 => x"08",
         11987 => x"fe",
         11988 => x"08",
         11989 => x"57",
         11990 => x"8d",
         11991 => x"0c",
         11992 => x"c8",
         11993 => x"0d",
         11994 => x"c8",
         11995 => x"5a",
         11996 => x"2e",
         11997 => x"77",
         11998 => x"84",
         11999 => x"5a",
         12000 => x"80",
         12001 => x"81",
         12002 => x"5d",
         12003 => x"08",
         12004 => x"ef",
         12005 => x"33",
         12006 => x"7c",
         12007 => x"81",
         12008 => x"b8",
         12009 => x"17",
         12010 => x"fc",
         12011 => x"b9",
         12012 => x"2e",
         12013 => x"5a",
         12014 => x"b4",
         12015 => x"7e",
         12016 => x"80",
         12017 => x"33",
         12018 => x"2e",
         12019 => x"77",
         12020 => x"83",
         12021 => x"12",
         12022 => x"2b",
         12023 => x"07",
         12024 => x"70",
         12025 => x"2b",
         12026 => x"80",
         12027 => x"80",
         12028 => x"30",
         12029 => x"63",
         12030 => x"05",
         12031 => x"62",
         12032 => x"41",
         12033 => x"52",
         12034 => x"5e",
         12035 => x"f2",
         12036 => x"0c",
         12037 => x"0c",
         12038 => x"81",
         12039 => x"84",
         12040 => x"84",
         12041 => x"95",
         12042 => x"81",
         12043 => x"08",
         12044 => x"70",
         12045 => x"33",
         12046 => x"fc",
         12047 => x"5e",
         12048 => x"08",
         12049 => x"84",
         12050 => x"83",
         12051 => x"17",
         12052 => x"08",
         12053 => x"c8",
         12054 => x"74",
         12055 => x"27",
         12056 => x"82",
         12057 => x"74",
         12058 => x"81",
         12059 => x"38",
         12060 => x"17",
         12061 => x"08",
         12062 => x"52",
         12063 => x"51",
         12064 => x"3f",
         12065 => x"97",
         12066 => x"42",
         12067 => x"56",
         12068 => x"51",
         12069 => x"3f",
         12070 => x"08",
         12071 => x"e8",
         12072 => x"c8",
         12073 => x"80",
         12074 => x"b9",
         12075 => x"70",
         12076 => x"08",
         12077 => x"7c",
         12078 => x"62",
         12079 => x"5c",
         12080 => x"76",
         12081 => x"7a",
         12082 => x"94",
         12083 => x"17",
         12084 => x"58",
         12085 => x"34",
         12086 => x"77",
         12087 => x"81",
         12088 => x"33",
         12089 => x"07",
         12090 => x"80",
         12091 => x"1d",
         12092 => x"ff",
         12093 => x"5f",
         12094 => x"55",
         12095 => x"38",
         12096 => x"77",
         12097 => x"39",
         12098 => x"5a",
         12099 => x"7a",
         12100 => x"84",
         12101 => x"07",
         12102 => x"18",
         12103 => x"39",
         12104 => x"5a",
         12105 => x"3d",
         12106 => x"89",
         12107 => x"2e",
         12108 => x"08",
         12109 => x"2e",
         12110 => x"33",
         12111 => x"2e",
         12112 => x"15",
         12113 => x"22",
         12114 => x"78",
         12115 => x"38",
         12116 => x"5a",
         12117 => x"38",
         12118 => x"56",
         12119 => x"38",
         12120 => x"70",
         12121 => x"06",
         12122 => x"55",
         12123 => x"80",
         12124 => x"17",
         12125 => x"8c",
         12126 => x"b7",
         12127 => x"d5",
         12128 => x"08",
         12129 => x"54",
         12130 => x"88",
         12131 => x"08",
         12132 => x"38",
         12133 => x"0b",
         12134 => x"94",
         12135 => x"18",
         12136 => x"c0",
         12137 => x"90",
         12138 => x"80",
         12139 => x"75",
         12140 => x"75",
         12141 => x"b9",
         12142 => x"3d",
         12143 => x"54",
         12144 => x"80",
         12145 => x"52",
         12146 => x"fe",
         12147 => x"b9",
         12148 => x"84",
         12149 => x"80",
         12150 => x"38",
         12151 => x"08",
         12152 => x"d8",
         12153 => x"c8",
         12154 => x"82",
         12155 => x"53",
         12156 => x"51",
         12157 => x"3f",
         12158 => x"08",
         12159 => x"9c",
         12160 => x"11",
         12161 => x"57",
         12162 => x"74",
         12163 => x"38",
         12164 => x"17",
         12165 => x"33",
         12166 => x"73",
         12167 => x"78",
         12168 => x"26",
         12169 => x"9c",
         12170 => x"33",
         12171 => x"e2",
         12172 => x"c8",
         12173 => x"54",
         12174 => x"38",
         12175 => x"55",
         12176 => x"39",
         12177 => x"18",
         12178 => x"73",
         12179 => x"88",
         12180 => x"c7",
         12181 => x"08",
         12182 => x"fe",
         12183 => x"84",
         12184 => x"ff",
         12185 => x"38",
         12186 => x"08",
         12187 => x"be",
         12188 => x"ae",
         12189 => x"84",
         12190 => x"9c",
         12191 => x"81",
         12192 => x"b9",
         12193 => x"18",
         12194 => x"58",
         12195 => x"0b",
         12196 => x"08",
         12197 => x"38",
         12198 => x"08",
         12199 => x"27",
         12200 => x"74",
         12201 => x"38",
         12202 => x"52",
         12203 => x"83",
         12204 => x"b9",
         12205 => x"84",
         12206 => x"80",
         12207 => x"52",
         12208 => x"fc",
         12209 => x"b9",
         12210 => x"84",
         12211 => x"80",
         12212 => x"38",
         12213 => x"08",
         12214 => x"dc",
         12215 => x"c8",
         12216 => x"80",
         12217 => x"53",
         12218 => x"51",
         12219 => x"3f",
         12220 => x"08",
         12221 => x"9c",
         12222 => x"11",
         12223 => x"57",
         12224 => x"74",
         12225 => x"81",
         12226 => x"0c",
         12227 => x"81",
         12228 => x"84",
         12229 => x"54",
         12230 => x"ff",
         12231 => x"55",
         12232 => x"17",
         12233 => x"f3",
         12234 => x"fe",
         12235 => x"0b",
         12236 => x"59",
         12237 => x"39",
         12238 => x"39",
         12239 => x"18",
         12240 => x"fe",
         12241 => x"b9",
         12242 => x"18",
         12243 => x"fd",
         12244 => x"0b",
         12245 => x"59",
         12246 => x"39",
         12247 => x"08",
         12248 => x"81",
         12249 => x"39",
         12250 => x"82",
         12251 => x"ff",
         12252 => x"a8",
         12253 => x"b7",
         12254 => x"b9",
         12255 => x"84",
         12256 => x"80",
         12257 => x"75",
         12258 => x"0c",
         12259 => x"04",
         12260 => x"3d",
         12261 => x"3d",
         12262 => x"ff",
         12263 => x"84",
         12264 => x"56",
         12265 => x"08",
         12266 => x"81",
         12267 => x"70",
         12268 => x"06",
         12269 => x"56",
         12270 => x"76",
         12271 => x"80",
         12272 => x"38",
         12273 => x"05",
         12274 => x"06",
         12275 => x"56",
         12276 => x"38",
         12277 => x"08",
         12278 => x"9a",
         12279 => x"88",
         12280 => x"33",
         12281 => x"57",
         12282 => x"2e",
         12283 => x"76",
         12284 => x"06",
         12285 => x"2e",
         12286 => x"87",
         12287 => x"08",
         12288 => x"83",
         12289 => x"7a",
         12290 => x"c8",
         12291 => x"3d",
         12292 => x"ff",
         12293 => x"84",
         12294 => x"56",
         12295 => x"08",
         12296 => x"84",
         12297 => x"52",
         12298 => x"91",
         12299 => x"b9",
         12300 => x"84",
         12301 => x"a0",
         12302 => x"84",
         12303 => x"a7",
         12304 => x"95",
         12305 => x"17",
         12306 => x"2b",
         12307 => x"07",
         12308 => x"5d",
         12309 => x"39",
         12310 => x"08",
         12311 => x"38",
         12312 => x"08",
         12313 => x"78",
         12314 => x"3d",
         12315 => x"57",
         12316 => x"80",
         12317 => x"52",
         12318 => x"8b",
         12319 => x"b9",
         12320 => x"84",
         12321 => x"80",
         12322 => x"75",
         12323 => x"07",
         12324 => x"5a",
         12325 => x"9a",
         12326 => x"2e",
         12327 => x"79",
         12328 => x"81",
         12329 => x"38",
         12330 => x"7b",
         12331 => x"38",
         12332 => x"fd",
         12333 => x"51",
         12334 => x"3f",
         12335 => x"08",
         12336 => x"0c",
         12337 => x"04",
         12338 => x"98",
         12339 => x"80",
         12340 => x"08",
         12341 => x"b9",
         12342 => x"33",
         12343 => x"74",
         12344 => x"81",
         12345 => x"38",
         12346 => x"53",
         12347 => x"81",
         12348 => x"fe",
         12349 => x"84",
         12350 => x"80",
         12351 => x"ff",
         12352 => x"75",
         12353 => x"77",
         12354 => x"38",
         12355 => x"58",
         12356 => x"81",
         12357 => x"34",
         12358 => x"7c",
         12359 => x"38",
         12360 => x"51",
         12361 => x"3f",
         12362 => x"08",
         12363 => x"c8",
         12364 => x"ff",
         12365 => x"84",
         12366 => x"06",
         12367 => x"82",
         12368 => x"39",
         12369 => x"17",
         12370 => x"52",
         12371 => x"51",
         12372 => x"3f",
         12373 => x"b9",
         12374 => x"2e",
         12375 => x"ff",
         12376 => x"b9",
         12377 => x"18",
         12378 => x"08",
         12379 => x"31",
         12380 => x"08",
         12381 => x"a0",
         12382 => x"fe",
         12383 => x"17",
         12384 => x"82",
         12385 => x"06",
         12386 => x"81",
         12387 => x"08",
         12388 => x"05",
         12389 => x"81",
         12390 => x"fe",
         12391 => x"79",
         12392 => x"39",
         12393 => x"78",
         12394 => x"38",
         12395 => x"51",
         12396 => x"3f",
         12397 => x"08",
         12398 => x"c8",
         12399 => x"80",
         12400 => x"b9",
         12401 => x"2e",
         12402 => x"84",
         12403 => x"ff",
         12404 => x"38",
         12405 => x"52",
         12406 => x"fd",
         12407 => x"b9",
         12408 => x"38",
         12409 => x"fe",
         12410 => x"08",
         12411 => x"75",
         12412 => x"b0",
         12413 => x"94",
         12414 => x"17",
         12415 => x"5c",
         12416 => x"34",
         12417 => x"7a",
         12418 => x"38",
         12419 => x"a2",
         12420 => x"fd",
         12421 => x"b9",
         12422 => x"fd",
         12423 => x"56",
         12424 => x"e3",
         12425 => x"53",
         12426 => x"bc",
         12427 => x"3d",
         12428 => x"c0",
         12429 => x"c8",
         12430 => x"b9",
         12431 => x"2e",
         12432 => x"84",
         12433 => x"9f",
         12434 => x"7d",
         12435 => x"93",
         12436 => x"5a",
         12437 => x"3f",
         12438 => x"08",
         12439 => x"c8",
         12440 => x"88",
         12441 => x"c8",
         12442 => x"0d",
         12443 => x"c8",
         12444 => x"09",
         12445 => x"38",
         12446 => x"05",
         12447 => x"2a",
         12448 => x"58",
         12449 => x"ff",
         12450 => x"5f",
         12451 => x"3d",
         12452 => x"ff",
         12453 => x"84",
         12454 => x"75",
         12455 => x"b9",
         12456 => x"38",
         12457 => x"b9",
         12458 => x"2e",
         12459 => x"84",
         12460 => x"ff",
         12461 => x"38",
         12462 => x"38",
         12463 => x"c8",
         12464 => x"33",
         12465 => x"7a",
         12466 => x"fe",
         12467 => x"08",
         12468 => x"56",
         12469 => x"79",
         12470 => x"8a",
         12471 => x"71",
         12472 => x"08",
         12473 => x"7a",
         12474 => x"b8",
         12475 => x"80",
         12476 => x"80",
         12477 => x"05",
         12478 => x"15",
         12479 => x"38",
         12480 => x"17",
         12481 => x"75",
         12482 => x"38",
         12483 => x"1b",
         12484 => x"81",
         12485 => x"fe",
         12486 => x"84",
         12487 => x"81",
         12488 => x"18",
         12489 => x"82",
         12490 => x"39",
         12491 => x"17",
         12492 => x"17",
         12493 => x"18",
         12494 => x"fe",
         12495 => x"81",
         12496 => x"c8",
         12497 => x"84",
         12498 => x"83",
         12499 => x"17",
         12500 => x"08",
         12501 => x"a0",
         12502 => x"fe",
         12503 => x"17",
         12504 => x"82",
         12505 => x"06",
         12506 => x"75",
         12507 => x"08",
         12508 => x"05",
         12509 => x"81",
         12510 => x"fe",
         12511 => x"fe",
         12512 => x"56",
         12513 => x"58",
         12514 => x"27",
         12515 => x"7b",
         12516 => x"27",
         12517 => x"74",
         12518 => x"fe",
         12519 => x"84",
         12520 => x"5a",
         12521 => x"08",
         12522 => x"96",
         12523 => x"c8",
         12524 => x"fd",
         12525 => x"b9",
         12526 => x"2e",
         12527 => x"80",
         12528 => x"76",
         12529 => x"b0",
         12530 => x"c8",
         12531 => x"38",
         12532 => x"fe",
         12533 => x"08",
         12534 => x"77",
         12535 => x"38",
         12536 => x"18",
         12537 => x"33",
         12538 => x"7b",
         12539 => x"79",
         12540 => x"26",
         12541 => x"75",
         12542 => x"0c",
         12543 => x"04",
         12544 => x"55",
         12545 => x"ff",
         12546 => x"56",
         12547 => x"09",
         12548 => x"f0",
         12549 => x"b8",
         12550 => x"a0",
         12551 => x"05",
         12552 => x"16",
         12553 => x"38",
         12554 => x"0b",
         12555 => x"7d",
         12556 => x"80",
         12557 => x"7d",
         12558 => x"ce",
         12559 => x"80",
         12560 => x"a1",
         12561 => x"1a",
         12562 => x"0b",
         12563 => x"34",
         12564 => x"ff",
         12565 => x"56",
         12566 => x"17",
         12567 => x"2a",
         12568 => x"d3",
         12569 => x"33",
         12570 => x"2e",
         12571 => x"7d",
         12572 => x"80",
         12573 => x"1b",
         12574 => x"74",
         12575 => x"56",
         12576 => x"81",
         12577 => x"ff",
         12578 => x"ef",
         12579 => x"ae",
         12580 => x"17",
         12581 => x"71",
         12582 => x"06",
         12583 => x"78",
         12584 => x"34",
         12585 => x"5b",
         12586 => x"17",
         12587 => x"55",
         12588 => x"80",
         12589 => x"5b",
         12590 => x"1c",
         12591 => x"ff",
         12592 => x"84",
         12593 => x"56",
         12594 => x"08",
         12595 => x"69",
         12596 => x"c8",
         12597 => x"34",
         12598 => x"08",
         12599 => x"a1",
         12600 => x"34",
         12601 => x"99",
         12602 => x"6a",
         12603 => x"9a",
         12604 => x"88",
         12605 => x"9b",
         12606 => x"33",
         12607 => x"2e",
         12608 => x"69",
         12609 => x"8b",
         12610 => x"57",
         12611 => x"18",
         12612 => x"fe",
         12613 => x"84",
         12614 => x"56",
         12615 => x"c8",
         12616 => x"0d",
         12617 => x"2a",
         12618 => x"ec",
         12619 => x"88",
         12620 => x"80",
         12621 => x"fe",
         12622 => x"90",
         12623 => x"80",
         12624 => x"7a",
         12625 => x"74",
         12626 => x"34",
         12627 => x"0b",
         12628 => x"b8",
         12629 => x"56",
         12630 => x"7b",
         12631 => x"77",
         12632 => x"77",
         12633 => x"7b",
         12634 => x"69",
         12635 => x"8b",
         12636 => x"57",
         12637 => x"18",
         12638 => x"fe",
         12639 => x"84",
         12640 => x"56",
         12641 => x"d1",
         12642 => x"3d",
         12643 => x"70",
         12644 => x"79",
         12645 => x"38",
         12646 => x"05",
         12647 => x"9f",
         12648 => x"75",
         12649 => x"b8",
         12650 => x"38",
         12651 => x"81",
         12652 => x"53",
         12653 => x"fc",
         12654 => x"3d",
         12655 => x"b4",
         12656 => x"c8",
         12657 => x"b9",
         12658 => x"2e",
         12659 => x"84",
         12660 => x"b1",
         12661 => x"7f",
         12662 => x"b2",
         12663 => x"a5",
         12664 => x"59",
         12665 => x"3f",
         12666 => x"08",
         12667 => x"c8",
         12668 => x"02",
         12669 => x"33",
         12670 => x"5d",
         12671 => x"ce",
         12672 => x"92",
         12673 => x"08",
         12674 => x"75",
         12675 => x"57",
         12676 => x"81",
         12677 => x"ff",
         12678 => x"ef",
         12679 => x"58",
         12680 => x"58",
         12681 => x"70",
         12682 => x"33",
         12683 => x"05",
         12684 => x"15",
         12685 => x"38",
         12686 => x"52",
         12687 => x"9e",
         12688 => x"b9",
         12689 => x"84",
         12690 => x"85",
         12691 => x"a8",
         12692 => x"81",
         12693 => x"0b",
         12694 => x"0c",
         12695 => x"04",
         12696 => x"11",
         12697 => x"06",
         12698 => x"74",
         12699 => x"38",
         12700 => x"81",
         12701 => x"05",
         12702 => x"7a",
         12703 => x"38",
         12704 => x"83",
         12705 => x"08",
         12706 => x"5f",
         12707 => x"70",
         12708 => x"33",
         12709 => x"05",
         12710 => x"9f",
         12711 => x"56",
         12712 => x"89",
         12713 => x"70",
         12714 => x"57",
         12715 => x"17",
         12716 => x"26",
         12717 => x"17",
         12718 => x"06",
         12719 => x"30",
         12720 => x"59",
         12721 => x"2e",
         12722 => x"85",
         12723 => x"be",
         12724 => x"32",
         12725 => x"72",
         12726 => x"7a",
         12727 => x"55",
         12728 => x"95",
         12729 => x"84",
         12730 => x"7b",
         12731 => x"c2",
         12732 => x"7e",
         12733 => x"96",
         12734 => x"24",
         12735 => x"79",
         12736 => x"53",
         12737 => x"fc",
         12738 => x"3d",
         12739 => x"e4",
         12740 => x"c8",
         12741 => x"b9",
         12742 => x"b2",
         12743 => x"39",
         12744 => x"08",
         12745 => x"06",
         12746 => x"77",
         12747 => x"a8",
         12748 => x"c8",
         12749 => x"b9",
         12750 => x"92",
         12751 => x"93",
         12752 => x"02",
         12753 => x"cd",
         12754 => x"5a",
         12755 => x"05",
         12756 => x"70",
         12757 => x"34",
         12758 => x"79",
         12759 => x"80",
         12760 => x"8b",
         12761 => x"18",
         12762 => x"2a",
         12763 => x"56",
         12764 => x"75",
         12765 => x"76",
         12766 => x"7f",
         12767 => x"83",
         12768 => x"18",
         12769 => x"2a",
         12770 => x"5c",
         12771 => x"81",
         12772 => x"3d",
         12773 => x"81",
         12774 => x"9b",
         12775 => x"1a",
         12776 => x"2b",
         12777 => x"41",
         12778 => x"7d",
         12779 => x"e0",
         12780 => x"9c",
         12781 => x"05",
         12782 => x"7d",
         12783 => x"38",
         12784 => x"76",
         12785 => x"19",
         12786 => x"5e",
         12787 => x"82",
         12788 => x"7a",
         12789 => x"17",
         12790 => x"aa",
         12791 => x"33",
         12792 => x"bc",
         12793 => x"75",
         12794 => x"52",
         12795 => x"51",
         12796 => x"3f",
         12797 => x"08",
         12798 => x"38",
         12799 => x"5c",
         12800 => x"0c",
         12801 => x"80",
         12802 => x"56",
         12803 => x"38",
         12804 => x"5a",
         12805 => x"09",
         12806 => x"38",
         12807 => x"ff",
         12808 => x"56",
         12809 => x"18",
         12810 => x"2a",
         12811 => x"f3",
         12812 => x"33",
         12813 => x"2e",
         12814 => x"93",
         12815 => x"2a",
         12816 => x"ec",
         12817 => x"88",
         12818 => x"80",
         12819 => x"7f",
         12820 => x"83",
         12821 => x"08",
         12822 => x"b2",
         12823 => x"5c",
         12824 => x"2e",
         12825 => x"52",
         12826 => x"fb",
         12827 => x"b9",
         12828 => x"84",
         12829 => x"80",
         12830 => x"16",
         12831 => x"08",
         12832 => x"b4",
         12833 => x"2e",
         12834 => x"16",
         12835 => x"5f",
         12836 => x"09",
         12837 => x"a8",
         12838 => x"76",
         12839 => x"52",
         12840 => x"51",
         12841 => x"3f",
         12842 => x"08",
         12843 => x"38",
         12844 => x"58",
         12845 => x"0c",
         12846 => x"aa",
         12847 => x"08",
         12848 => x"34",
         12849 => x"17",
         12850 => x"08",
         12851 => x"38",
         12852 => x"51",
         12853 => x"3f",
         12854 => x"08",
         12855 => x"c8",
         12856 => x"ff",
         12857 => x"56",
         12858 => x"f9",
         12859 => x"56",
         12860 => x"38",
         12861 => x"e5",
         12862 => x"b9",
         12863 => x"b9",
         12864 => x"3d",
         12865 => x"0b",
         12866 => x"0c",
         12867 => x"04",
         12868 => x"94",
         12869 => x"98",
         12870 => x"2b",
         12871 => x"58",
         12872 => x"8d",
         12873 => x"c8",
         12874 => x"fb",
         12875 => x"b9",
         12876 => x"2e",
         12877 => x"75",
         12878 => x"0c",
         12879 => x"04",
         12880 => x"16",
         12881 => x"52",
         12882 => x"51",
         12883 => x"3f",
         12884 => x"b9",
         12885 => x"2e",
         12886 => x"fe",
         12887 => x"b9",
         12888 => x"17",
         12889 => x"08",
         12890 => x"31",
         12891 => x"08",
         12892 => x"a0",
         12893 => x"fe",
         12894 => x"16",
         12895 => x"82",
         12896 => x"06",
         12897 => x"81",
         12898 => x"08",
         12899 => x"05",
         12900 => x"81",
         12901 => x"fe",
         12902 => x"79",
         12903 => x"39",
         12904 => x"17",
         12905 => x"17",
         12906 => x"18",
         12907 => x"fe",
         12908 => x"81",
         12909 => x"c8",
         12910 => x"38",
         12911 => x"08",
         12912 => x"b4",
         12913 => x"18",
         12914 => x"b9",
         12915 => x"55",
         12916 => x"08",
         12917 => x"38",
         12918 => x"5d",
         12919 => x"09",
         12920 => x"81",
         12921 => x"b4",
         12922 => x"18",
         12923 => x"7a",
         12924 => x"33",
         12925 => x"eb",
         12926 => x"fb",
         12927 => x"3d",
         12928 => x"df",
         12929 => x"84",
         12930 => x"05",
         12931 => x"82",
         12932 => x"cc",
         12933 => x"3d",
         12934 => x"d8",
         12935 => x"c8",
         12936 => x"b9",
         12937 => x"2e",
         12938 => x"84",
         12939 => x"96",
         12940 => x"78",
         12941 => x"96",
         12942 => x"51",
         12943 => x"3f",
         12944 => x"08",
         12945 => x"c8",
         12946 => x"02",
         12947 => x"33",
         12948 => x"54",
         12949 => x"d2",
         12950 => x"06",
         12951 => x"8b",
         12952 => x"06",
         12953 => x"07",
         12954 => x"55",
         12955 => x"34",
         12956 => x"0b",
         12957 => x"78",
         12958 => x"9a",
         12959 => x"c8",
         12960 => x"c8",
         12961 => x"0d",
         12962 => x"0d",
         12963 => x"53",
         12964 => x"05",
         12965 => x"51",
         12966 => x"3f",
         12967 => x"08",
         12968 => x"c8",
         12969 => x"8a",
         12970 => x"b9",
         12971 => x"3d",
         12972 => x"5a",
         12973 => x"3d",
         12974 => x"ff",
         12975 => x"84",
         12976 => x"55",
         12977 => x"08",
         12978 => x"80",
         12979 => x"81",
         12980 => x"86",
         12981 => x"38",
         12982 => x"22",
         12983 => x"71",
         12984 => x"59",
         12985 => x"96",
         12986 => x"88",
         12987 => x"97",
         12988 => x"90",
         12989 => x"98",
         12990 => x"98",
         12991 => x"99",
         12992 => x"57",
         12993 => x"18",
         12994 => x"fe",
         12995 => x"84",
         12996 => x"84",
         12997 => x"96",
         12998 => x"e8",
         12999 => x"6d",
         13000 => x"53",
         13001 => x"05",
         13002 => x"51",
         13003 => x"3f",
         13004 => x"08",
         13005 => x"08",
         13006 => x"b9",
         13007 => x"80",
         13008 => x"57",
         13009 => x"8b",
         13010 => x"76",
         13011 => x"78",
         13012 => x"76",
         13013 => x"07",
         13014 => x"5b",
         13015 => x"81",
         13016 => x"70",
         13017 => x"58",
         13018 => x"81",
         13019 => x"a4",
         13020 => x"56",
         13021 => x"16",
         13022 => x"82",
         13023 => x"16",
         13024 => x"55",
         13025 => x"09",
         13026 => x"98",
         13027 => x"76",
         13028 => x"52",
         13029 => x"51",
         13030 => x"3f",
         13031 => x"08",
         13032 => x"38",
         13033 => x"59",
         13034 => x"0c",
         13035 => x"bd",
         13036 => x"33",
         13037 => x"c3",
         13038 => x"2e",
         13039 => x"e4",
         13040 => x"2e",
         13041 => x"56",
         13042 => x"05",
         13043 => x"82",
         13044 => x"90",
         13045 => x"2b",
         13046 => x"33",
         13047 => x"88",
         13048 => x"71",
         13049 => x"5f",
         13050 => x"59",
         13051 => x"b9",
         13052 => x"3d",
         13053 => x"5e",
         13054 => x"52",
         13055 => x"52",
         13056 => x"8b",
         13057 => x"c8",
         13058 => x"b9",
         13059 => x"2e",
         13060 => x"76",
         13061 => x"81",
         13062 => x"38",
         13063 => x"80",
         13064 => x"39",
         13065 => x"16",
         13066 => x"16",
         13067 => x"17",
         13068 => x"fe",
         13069 => x"77",
         13070 => x"c8",
         13071 => x"09",
         13072 => x"e8",
         13073 => x"c8",
         13074 => x"34",
         13075 => x"a8",
         13076 => x"84",
         13077 => x"5a",
         13078 => x"17",
         13079 => x"ad",
         13080 => x"33",
         13081 => x"2e",
         13082 => x"fe",
         13083 => x"54",
         13084 => x"a0",
         13085 => x"53",
         13086 => x"16",
         13087 => x"db",
         13088 => x"59",
         13089 => x"53",
         13090 => x"81",
         13091 => x"fe",
         13092 => x"84",
         13093 => x"80",
         13094 => x"38",
         13095 => x"75",
         13096 => x"fe",
         13097 => x"84",
         13098 => x"57",
         13099 => x"08",
         13100 => x"84",
         13101 => x"84",
         13102 => x"66",
         13103 => x"79",
         13104 => x"7c",
         13105 => x"56",
         13106 => x"34",
         13107 => x"8a",
         13108 => x"38",
         13109 => x"57",
         13110 => x"34",
         13111 => x"fc",
         13112 => x"18",
         13113 => x"33",
         13114 => x"79",
         13115 => x"38",
         13116 => x"79",
         13117 => x"39",
         13118 => x"82",
         13119 => x"ff",
         13120 => x"a2",
         13121 => x"9c",
         13122 => x"b9",
         13123 => x"84",
         13124 => x"82",
         13125 => x"3d",
         13126 => x"57",
         13127 => x"70",
         13128 => x"34",
         13129 => x"74",
         13130 => x"a3",
         13131 => x"33",
         13132 => x"06",
         13133 => x"5a",
         13134 => x"81",
         13135 => x"3d",
         13136 => x"5c",
         13137 => x"06",
         13138 => x"55",
         13139 => x"38",
         13140 => x"74",
         13141 => x"26",
         13142 => x"74",
         13143 => x"3f",
         13144 => x"84",
         13145 => x"51",
         13146 => x"84",
         13147 => x"83",
         13148 => x"57",
         13149 => x"81",
         13150 => x"e6",
         13151 => x"e6",
         13152 => x"81",
         13153 => x"56",
         13154 => x"2e",
         13155 => x"74",
         13156 => x"2e",
         13157 => x"18",
         13158 => x"81",
         13159 => x"57",
         13160 => x"2e",
         13161 => x"77",
         13162 => x"06",
         13163 => x"81",
         13164 => x"78",
         13165 => x"81",
         13166 => x"81",
         13167 => x"89",
         13168 => x"38",
         13169 => x"27",
         13170 => x"88",
         13171 => x"7b",
         13172 => x"5d",
         13173 => x"5a",
         13174 => x"81",
         13175 => x"81",
         13176 => x"08",
         13177 => x"81",
         13178 => x"58",
         13179 => x"9f",
         13180 => x"38",
         13181 => x"57",
         13182 => x"81",
         13183 => x"38",
         13184 => x"99",
         13185 => x"05",
         13186 => x"70",
         13187 => x"7a",
         13188 => x"81",
         13189 => x"ff",
         13190 => x"ed",
         13191 => x"80",
         13192 => x"95",
         13193 => x"56",
         13194 => x"3f",
         13195 => x"08",
         13196 => x"c8",
         13197 => x"b4",
         13198 => x"75",
         13199 => x"0c",
         13200 => x"04",
         13201 => x"74",
         13202 => x"3f",
         13203 => x"08",
         13204 => x"06",
         13205 => x"f8",
         13206 => x"75",
         13207 => x"0c",
         13208 => x"04",
         13209 => x"33",
         13210 => x"39",
         13211 => x"51",
         13212 => x"3f",
         13213 => x"08",
         13214 => x"c8",
         13215 => x"38",
         13216 => x"82",
         13217 => x"6c",
         13218 => x"55",
         13219 => x"05",
         13220 => x"70",
         13221 => x"34",
         13222 => x"74",
         13223 => x"5d",
         13224 => x"1e",
         13225 => x"fe",
         13226 => x"84",
         13227 => x"55",
         13228 => x"87",
         13229 => x"27",
         13230 => x"86",
         13231 => x"39",
         13232 => x"08",
         13233 => x"81",
         13234 => x"38",
         13235 => x"75",
         13236 => x"38",
         13237 => x"53",
         13238 => x"fe",
         13239 => x"84",
         13240 => x"57",
         13241 => x"08",
         13242 => x"81",
         13243 => x"38",
         13244 => x"08",
         13245 => x"5a",
         13246 => x"57",
         13247 => x"18",
         13248 => x"b2",
         13249 => x"33",
         13250 => x"2e",
         13251 => x"81",
         13252 => x"54",
         13253 => x"18",
         13254 => x"33",
         13255 => x"c4",
         13256 => x"c8",
         13257 => x"85",
         13258 => x"81",
         13259 => x"19",
         13260 => x"78",
         13261 => x"9c",
         13262 => x"33",
         13263 => x"74",
         13264 => x"81",
         13265 => x"30",
         13266 => x"78",
         13267 => x"74",
         13268 => x"d7",
         13269 => x"5a",
         13270 => x"a5",
         13271 => x"75",
         13272 => x"a1",
         13273 => x"c8",
         13274 => x"b9",
         13275 => x"2e",
         13276 => x"87",
         13277 => x"2e",
         13278 => x"76",
         13279 => x"b9",
         13280 => x"57",
         13281 => x"70",
         13282 => x"34",
         13283 => x"74",
         13284 => x"56",
         13285 => x"17",
         13286 => x"7e",
         13287 => x"76",
         13288 => x"58",
         13289 => x"81",
         13290 => x"ff",
         13291 => x"80",
         13292 => x"38",
         13293 => x"05",
         13294 => x"70",
         13295 => x"34",
         13296 => x"74",
         13297 => x"d6",
         13298 => x"e5",
         13299 => x"5d",
         13300 => x"1e",
         13301 => x"fe",
         13302 => x"84",
         13303 => x"55",
         13304 => x"81",
         13305 => x"39",
         13306 => x"18",
         13307 => x"52",
         13308 => x"51",
         13309 => x"3f",
         13310 => x"08",
         13311 => x"81",
         13312 => x"38",
         13313 => x"08",
         13314 => x"b4",
         13315 => x"19",
         13316 => x"7b",
         13317 => x"27",
         13318 => x"18",
         13319 => x"82",
         13320 => x"84",
         13321 => x"59",
         13322 => x"74",
         13323 => x"75",
         13324 => x"d1",
         13325 => x"c8",
         13326 => x"b9",
         13327 => x"2e",
         13328 => x"fe",
         13329 => x"70",
         13330 => x"80",
         13331 => x"38",
         13332 => x"81",
         13333 => x"08",
         13334 => x"05",
         13335 => x"81",
         13336 => x"fe",
         13337 => x"fd",
         13338 => x"3d",
         13339 => x"02",
         13340 => x"cb",
         13341 => x"5b",
         13342 => x"76",
         13343 => x"38",
         13344 => x"74",
         13345 => x"38",
         13346 => x"73",
         13347 => x"38",
         13348 => x"84",
         13349 => x"59",
         13350 => x"81",
         13351 => x"54",
         13352 => x"81",
         13353 => x"17",
         13354 => x"81",
         13355 => x"80",
         13356 => x"38",
         13357 => x"81",
         13358 => x"17",
         13359 => x"2a",
         13360 => x"5d",
         13361 => x"81",
         13362 => x"8a",
         13363 => x"89",
         13364 => x"7c",
         13365 => x"59",
         13366 => x"3f",
         13367 => x"06",
         13368 => x"72",
         13369 => x"84",
         13370 => x"05",
         13371 => x"79",
         13372 => x"55",
         13373 => x"27",
         13374 => x"19",
         13375 => x"83",
         13376 => x"77",
         13377 => x"80",
         13378 => x"76",
         13379 => x"87",
         13380 => x"7f",
         13381 => x"14",
         13382 => x"83",
         13383 => x"84",
         13384 => x"81",
         13385 => x"38",
         13386 => x"08",
         13387 => x"d8",
         13388 => x"c8",
         13389 => x"38",
         13390 => x"78",
         13391 => x"38",
         13392 => x"09",
         13393 => x"38",
         13394 => x"54",
         13395 => x"c8",
         13396 => x"0d",
         13397 => x"84",
         13398 => x"90",
         13399 => x"81",
         13400 => x"fe",
         13401 => x"84",
         13402 => x"81",
         13403 => x"fe",
         13404 => x"77",
         13405 => x"fe",
         13406 => x"80",
         13407 => x"38",
         13408 => x"58",
         13409 => x"ab",
         13410 => x"54",
         13411 => x"80",
         13412 => x"53",
         13413 => x"51",
         13414 => x"3f",
         13415 => x"08",
         13416 => x"c8",
         13417 => x"38",
         13418 => x"ff",
         13419 => x"5e",
         13420 => x"7e",
         13421 => x"0c",
         13422 => x"2e",
         13423 => x"7a",
         13424 => x"79",
         13425 => x"90",
         13426 => x"c0",
         13427 => x"90",
         13428 => x"15",
         13429 => x"94",
         13430 => x"5a",
         13431 => x"fe",
         13432 => x"7d",
         13433 => x"0c",
         13434 => x"81",
         13435 => x"84",
         13436 => x"54",
         13437 => x"ff",
         13438 => x"39",
         13439 => x"59",
         13440 => x"82",
         13441 => x"39",
         13442 => x"c0",
         13443 => x"5e",
         13444 => x"84",
         13445 => x"e3",
         13446 => x"3d",
         13447 => x"08",
         13448 => x"81",
         13449 => x"44",
         13450 => x"0b",
         13451 => x"70",
         13452 => x"79",
         13453 => x"8a",
         13454 => x"81",
         13455 => x"70",
         13456 => x"56",
         13457 => x"85",
         13458 => x"ed",
         13459 => x"2e",
         13460 => x"84",
         13461 => x"56",
         13462 => x"84",
         13463 => x"10",
         13464 => x"90",
         13465 => x"56",
         13466 => x"2e",
         13467 => x"75",
         13468 => x"84",
         13469 => x"33",
         13470 => x"12",
         13471 => x"5d",
         13472 => x"51",
         13473 => x"3f",
         13474 => x"08",
         13475 => x"70",
         13476 => x"56",
         13477 => x"84",
         13478 => x"82",
         13479 => x"40",
         13480 => x"84",
         13481 => x"3d",
         13482 => x"83",
         13483 => x"fe",
         13484 => x"84",
         13485 => x"84",
         13486 => x"55",
         13487 => x"84",
         13488 => x"82",
         13489 => x"84",
         13490 => x"15",
         13491 => x"74",
         13492 => x"7e",
         13493 => x"38",
         13494 => x"26",
         13495 => x"7e",
         13496 => x"26",
         13497 => x"ff",
         13498 => x"55",
         13499 => x"38",
         13500 => x"a6",
         13501 => x"2a",
         13502 => x"77",
         13503 => x"5b",
         13504 => x"85",
         13505 => x"30",
         13506 => x"77",
         13507 => x"91",
         13508 => x"b0",
         13509 => x"2e",
         13510 => x"81",
         13511 => x"60",
         13512 => x"fe",
         13513 => x"81",
         13514 => x"c8",
         13515 => x"38",
         13516 => x"05",
         13517 => x"fe",
         13518 => x"88",
         13519 => x"56",
         13520 => x"82",
         13521 => x"09",
         13522 => x"f8",
         13523 => x"29",
         13524 => x"b2",
         13525 => x"58",
         13526 => x"82",
         13527 => x"b6",
         13528 => x"33",
         13529 => x"71",
         13530 => x"88",
         13531 => x"14",
         13532 => x"07",
         13533 => x"33",
         13534 => x"ba",
         13535 => x"33",
         13536 => x"71",
         13537 => x"88",
         13538 => x"14",
         13539 => x"07",
         13540 => x"33",
         13541 => x"a2",
         13542 => x"a3",
         13543 => x"3d",
         13544 => x"54",
         13545 => x"41",
         13546 => x"4d",
         13547 => x"ff",
         13548 => x"90",
         13549 => x"7a",
         13550 => x"82",
         13551 => x"81",
         13552 => x"06",
         13553 => x"80",
         13554 => x"38",
         13555 => x"45",
         13556 => x"89",
         13557 => x"06",
         13558 => x"f4",
         13559 => x"70",
         13560 => x"43",
         13561 => x"83",
         13562 => x"38",
         13563 => x"78",
         13564 => x"81",
         13565 => x"ec",
         13566 => x"74",
         13567 => x"38",
         13568 => x"98",
         13569 => x"ec",
         13570 => x"82",
         13571 => x"57",
         13572 => x"80",
         13573 => x"76",
         13574 => x"38",
         13575 => x"51",
         13576 => x"3f",
         13577 => x"08",
         13578 => x"55",
         13579 => x"08",
         13580 => x"96",
         13581 => x"84",
         13582 => x"10",
         13583 => x"08",
         13584 => x"72",
         13585 => x"57",
         13586 => x"ff",
         13587 => x"5d",
         13588 => x"47",
         13589 => x"11",
         13590 => x"11",
         13591 => x"6b",
         13592 => x"58",
         13593 => x"62",
         13594 => x"b8",
         13595 => x"5d",
         13596 => x"16",
         13597 => x"56",
         13598 => x"26",
         13599 => x"78",
         13600 => x"31",
         13601 => x"68",
         13602 => x"fd",
         13603 => x"84",
         13604 => x"40",
         13605 => x"89",
         13606 => x"82",
         13607 => x"06",
         13608 => x"83",
         13609 => x"84",
         13610 => x"27",
         13611 => x"7a",
         13612 => x"77",
         13613 => x"80",
         13614 => x"ef",
         13615 => x"fe",
         13616 => x"57",
         13617 => x"c8",
         13618 => x"0d",
         13619 => x"0c",
         13620 => x"fb",
         13621 => x"0b",
         13622 => x"0c",
         13623 => x"84",
         13624 => x"04",
         13625 => x"11",
         13626 => x"06",
         13627 => x"74",
         13628 => x"38",
         13629 => x"81",
         13630 => x"05",
         13631 => x"7a",
         13632 => x"38",
         13633 => x"e5",
         13634 => x"7d",
         13635 => x"5b",
         13636 => x"05",
         13637 => x"70",
         13638 => x"33",
         13639 => x"45",
         13640 => x"99",
         13641 => x"e0",
         13642 => x"ff",
         13643 => x"ff",
         13644 => x"64",
         13645 => x"38",
         13646 => x"81",
         13647 => x"46",
         13648 => x"9f",
         13649 => x"76",
         13650 => x"81",
         13651 => x"78",
         13652 => x"75",
         13653 => x"30",
         13654 => x"9f",
         13655 => x"5d",
         13656 => x"80",
         13657 => x"38",
         13658 => x"1f",
         13659 => x"7c",
         13660 => x"38",
         13661 => x"e0",
         13662 => x"f8",
         13663 => x"52",
         13664 => x"ca",
         13665 => x"57",
         13666 => x"08",
         13667 => x"61",
         13668 => x"06",
         13669 => x"08",
         13670 => x"83",
         13671 => x"6c",
         13672 => x"7e",
         13673 => x"9c",
         13674 => x"31",
         13675 => x"39",
         13676 => x"d2",
         13677 => x"24",
         13678 => x"7b",
         13679 => x"0c",
         13680 => x"39",
         13681 => x"48",
         13682 => x"80",
         13683 => x"38",
         13684 => x"30",
         13685 => x"fc",
         13686 => x"b9",
         13687 => x"f5",
         13688 => x"7a",
         13689 => x"18",
         13690 => x"7b",
         13691 => x"38",
         13692 => x"84",
         13693 => x"9f",
         13694 => x"b9",
         13695 => x"80",
         13696 => x"2e",
         13697 => x"9f",
         13698 => x"8b",
         13699 => x"06",
         13700 => x"7a",
         13701 => x"84",
         13702 => x"55",
         13703 => x"81",
         13704 => x"ff",
         13705 => x"f4",
         13706 => x"83",
         13707 => x"57",
         13708 => x"81",
         13709 => x"76",
         13710 => x"58",
         13711 => x"55",
         13712 => x"60",
         13713 => x"74",
         13714 => x"61",
         13715 => x"77",
         13716 => x"34",
         13717 => x"ff",
         13718 => x"61",
         13719 => x"6a",
         13720 => x"7b",
         13721 => x"34",
         13722 => x"05",
         13723 => x"32",
         13724 => x"48",
         13725 => x"05",
         13726 => x"2a",
         13727 => x"68",
         13728 => x"34",
         13729 => x"83",
         13730 => x"86",
         13731 => x"83",
         13732 => x"55",
         13733 => x"05",
         13734 => x"2a",
         13735 => x"94",
         13736 => x"61",
         13737 => x"bf",
         13738 => x"34",
         13739 => x"05",
         13740 => x"9a",
         13741 => x"61",
         13742 => x"7e",
         13743 => x"34",
         13744 => x"48",
         13745 => x"05",
         13746 => x"2a",
         13747 => x"9e",
         13748 => x"98",
         13749 => x"d4",
         13750 => x"d4",
         13751 => x"05",
         13752 => x"2e",
         13753 => x"80",
         13754 => x"34",
         13755 => x"05",
         13756 => x"a9",
         13757 => x"cc",
         13758 => x"34",
         13759 => x"ff",
         13760 => x"61",
         13761 => x"74",
         13762 => x"6a",
         13763 => x"34",
         13764 => x"a4",
         13765 => x"61",
         13766 => x"93",
         13767 => x"83",
         13768 => x"57",
         13769 => x"81",
         13770 => x"76",
         13771 => x"58",
         13772 => x"55",
         13773 => x"60",
         13774 => x"49",
         13775 => x"34",
         13776 => x"05",
         13777 => x"6b",
         13778 => x"7e",
         13779 => x"79",
         13780 => x"8f",
         13781 => x"84",
         13782 => x"fa",
         13783 => x"17",
         13784 => x"2e",
         13785 => x"69",
         13786 => x"80",
         13787 => x"05",
         13788 => x"15",
         13789 => x"38",
         13790 => x"5b",
         13791 => x"86",
         13792 => x"ff",
         13793 => x"62",
         13794 => x"38",
         13795 => x"61",
         13796 => x"2a",
         13797 => x"74",
         13798 => x"05",
         13799 => x"90",
         13800 => x"64",
         13801 => x"46",
         13802 => x"2a",
         13803 => x"34",
         13804 => x"59",
         13805 => x"83",
         13806 => x"78",
         13807 => x"60",
         13808 => x"fe",
         13809 => x"84",
         13810 => x"85",
         13811 => x"80",
         13812 => x"80",
         13813 => x"05",
         13814 => x"15",
         13815 => x"38",
         13816 => x"7a",
         13817 => x"76",
         13818 => x"81",
         13819 => x"80",
         13820 => x"38",
         13821 => x"83",
         13822 => x"66",
         13823 => x"75",
         13824 => x"38",
         13825 => x"54",
         13826 => x"52",
         13827 => x"c4",
         13828 => x"b9",
         13829 => x"9b",
         13830 => x"76",
         13831 => x"5b",
         13832 => x"8c",
         13833 => x"2e",
         13834 => x"58",
         13835 => x"ff",
         13836 => x"84",
         13837 => x"2e",
         13838 => x"58",
         13839 => x"38",
         13840 => x"81",
         13841 => x"81",
         13842 => x"80",
         13843 => x"80",
         13844 => x"05",
         13845 => x"19",
         13846 => x"38",
         13847 => x"34",
         13848 => x"34",
         13849 => x"05",
         13850 => x"34",
         13851 => x"05",
         13852 => x"82",
         13853 => x"67",
         13854 => x"77",
         13855 => x"34",
         13856 => x"fd",
         13857 => x"1f",
         13858 => x"9a",
         13859 => x"85",
         13860 => x"b9",
         13861 => x"2a",
         13862 => x"76",
         13863 => x"34",
         13864 => x"08",
         13865 => x"34",
         13866 => x"c6",
         13867 => x"61",
         13868 => x"34",
         13869 => x"c8",
         13870 => x"b9",
         13871 => x"83",
         13872 => x"62",
         13873 => x"05",
         13874 => x"2a",
         13875 => x"83",
         13876 => x"62",
         13877 => x"77",
         13878 => x"05",
         13879 => x"2a",
         13880 => x"83",
         13881 => x"81",
         13882 => x"60",
         13883 => x"fe",
         13884 => x"81",
         13885 => x"c8",
         13886 => x"38",
         13887 => x"52",
         13888 => x"c3",
         13889 => x"57",
         13890 => x"08",
         13891 => x"84",
         13892 => x"84",
         13893 => x"9f",
         13894 => x"b9",
         13895 => x"62",
         13896 => x"39",
         13897 => x"16",
         13898 => x"c4",
         13899 => x"38",
         13900 => x"57",
         13901 => x"e6",
         13902 => x"58",
         13903 => x"9d",
         13904 => x"26",
         13905 => x"e6",
         13906 => x"10",
         13907 => x"22",
         13908 => x"74",
         13909 => x"38",
         13910 => x"ee",
         13911 => x"78",
         13912 => x"c2",
         13913 => x"c8",
         13914 => x"84",
         13915 => x"89",
         13916 => x"a0",
         13917 => x"84",
         13918 => x"fc",
         13919 => x"58",
         13920 => x"f0",
         13921 => x"f5",
         13922 => x"57",
         13923 => x"84",
         13924 => x"83",
         13925 => x"f8",
         13926 => x"f8",
         13927 => x"81",
         13928 => x"f4",
         13929 => x"57",
         13930 => x"68",
         13931 => x"63",
         13932 => x"af",
         13933 => x"f4",
         13934 => x"61",
         13935 => x"75",
         13936 => x"68",
         13937 => x"34",
         13938 => x"5b",
         13939 => x"05",
         13940 => x"2a",
         13941 => x"a3",
         13942 => x"c6",
         13943 => x"80",
         13944 => x"80",
         13945 => x"05",
         13946 => x"80",
         13947 => x"80",
         13948 => x"c6",
         13949 => x"61",
         13950 => x"7c",
         13951 => x"7b",
         13952 => x"34",
         13953 => x"59",
         13954 => x"05",
         13955 => x"2a",
         13956 => x"a7",
         13957 => x"61",
         13958 => x"80",
         13959 => x"34",
         13960 => x"05",
         13961 => x"af",
         13962 => x"61",
         13963 => x"80",
         13964 => x"34",
         13965 => x"05",
         13966 => x"b3",
         13967 => x"80",
         13968 => x"05",
         13969 => x"80",
         13970 => x"93",
         13971 => x"05",
         13972 => x"59",
         13973 => x"70",
         13974 => x"33",
         13975 => x"05",
         13976 => x"15",
         13977 => x"2e",
         13978 => x"76",
         13979 => x"58",
         13980 => x"81",
         13981 => x"ff",
         13982 => x"da",
         13983 => x"39",
         13984 => x"53",
         13985 => x"51",
         13986 => x"3f",
         13987 => x"b9",
         13988 => x"b0",
         13989 => x"29",
         13990 => x"77",
         13991 => x"05",
         13992 => x"84",
         13993 => x"53",
         13994 => x"51",
         13995 => x"3f",
         13996 => x"81",
         13997 => x"c8",
         13998 => x"0d",
         13999 => x"0c",
         14000 => x"34",
         14001 => x"6a",
         14002 => x"4c",
         14003 => x"70",
         14004 => x"34",
         14005 => x"ff",
         14006 => x"34",
         14007 => x"05",
         14008 => x"86",
         14009 => x"61",
         14010 => x"ff",
         14011 => x"34",
         14012 => x"05",
         14013 => x"8a",
         14014 => x"65",
         14015 => x"f9",
         14016 => x"54",
         14017 => x"60",
         14018 => x"fe",
         14019 => x"84",
         14020 => x"57",
         14021 => x"81",
         14022 => x"ff",
         14023 => x"f4",
         14024 => x"80",
         14025 => x"81",
         14026 => x"7b",
         14027 => x"75",
         14028 => x"57",
         14029 => x"75",
         14030 => x"57",
         14031 => x"75",
         14032 => x"61",
         14033 => x"34",
         14034 => x"83",
         14035 => x"80",
         14036 => x"e6",
         14037 => x"e1",
         14038 => x"05",
         14039 => x"05",
         14040 => x"83",
         14041 => x"7a",
         14042 => x"78",
         14043 => x"05",
         14044 => x"2a",
         14045 => x"83",
         14046 => x"7a",
         14047 => x"7f",
         14048 => x"05",
         14049 => x"83",
         14050 => x"76",
         14051 => x"05",
         14052 => x"83",
         14053 => x"76",
         14054 => x"05",
         14055 => x"69",
         14056 => x"6b",
         14057 => x"87",
         14058 => x"52",
         14059 => x"bd",
         14060 => x"54",
         14061 => x"60",
         14062 => x"fe",
         14063 => x"69",
         14064 => x"f7",
         14065 => x"3d",
         14066 => x"5b",
         14067 => x"61",
         14068 => x"57",
         14069 => x"25",
         14070 => x"3d",
         14071 => x"f8",
         14072 => x"53",
         14073 => x"51",
         14074 => x"3f",
         14075 => x"09",
         14076 => x"38",
         14077 => x"55",
         14078 => x"90",
         14079 => x"70",
         14080 => x"34",
         14081 => x"74",
         14082 => x"38",
         14083 => x"cd",
         14084 => x"34",
         14085 => x"83",
         14086 => x"74",
         14087 => x"0c",
         14088 => x"04",
         14089 => x"7b",
         14090 => x"b3",
         14091 => x"57",
         14092 => x"80",
         14093 => x"17",
         14094 => x"76",
         14095 => x"88",
         14096 => x"17",
         14097 => x"59",
         14098 => x"81",
         14099 => x"bb",
         14100 => x"74",
         14101 => x"81",
         14102 => x"0c",
         14103 => x"04",
         14104 => x"05",
         14105 => x"8c",
         14106 => x"08",
         14107 => x"d1",
         14108 => x"32",
         14109 => x"72",
         14110 => x"70",
         14111 => x"0c",
         14112 => x"1b",
         14113 => x"56",
         14114 => x"52",
         14115 => x"94",
         14116 => x"39",
         14117 => x"02",
         14118 => x"33",
         14119 => x"58",
         14120 => x"57",
         14121 => x"70",
         14122 => x"34",
         14123 => x"74",
         14124 => x"3d",
         14125 => x"77",
         14126 => x"f7",
         14127 => x"80",
         14128 => x"c0",
         14129 => x"17",
         14130 => x"59",
         14131 => x"81",
         14132 => x"bb",
         14133 => x"74",
         14134 => x"81",
         14135 => x"0c",
         14136 => x"75",
         14137 => x"9f",
         14138 => x"11",
         14139 => x"c0",
         14140 => x"08",
         14141 => x"c9",
         14142 => x"c8",
         14143 => x"7c",
         14144 => x"38",
         14145 => x"b9",
         14146 => x"3d",
         14147 => x"3d",
         14148 => x"55",
         14149 => x"05",
         14150 => x"51",
         14151 => x"3f",
         14152 => x"70",
         14153 => x"07",
         14154 => x"30",
         14155 => x"56",
         14156 => x"8d",
         14157 => x"fd",
         14158 => x"81",
         14159 => x"b9",
         14160 => x"3d",
         14161 => x"3d",
         14162 => x"84",
         14163 => x"22",
         14164 => x"52",
         14165 => x"26",
         14166 => x"83",
         14167 => x"52",
         14168 => x"c8",
         14169 => x"0d",
         14170 => x"ff",
         14171 => x"70",
         14172 => x"09",
         14173 => x"38",
         14174 => x"e4",
         14175 => x"8c",
         14176 => x"71",
         14177 => x"81",
         14178 => x"ff",
         14179 => x"54",
         14180 => x"26",
         14181 => x"10",
         14182 => x"05",
         14183 => x"51",
         14184 => x"80",
         14185 => x"ff",
         14186 => x"c8",
         14187 => x"3d",
         14188 => x"3d",
         14189 => x"05",
         14190 => x"05",
         14191 => x"53",
         14192 => x"70",
         14193 => x"8c",
         14194 => x"72",
         14195 => x"0c",
         14196 => x"04",
         14197 => x"2e",
         14198 => x"ef",
         14199 => x"ff",
         14200 => x"70",
         14201 => x"8c",
         14202 => x"84",
         14203 => x"51",
         14204 => x"04",
         14205 => x"77",
         14206 => x"ff",
         14207 => x"e1",
         14208 => x"ff",
         14209 => x"e9",
         14210 => x"75",
         14211 => x"80",
         14212 => x"70",
         14213 => x"22",
         14214 => x"70",
         14215 => x"7a",
         14216 => x"56",
         14217 => x"b7",
         14218 => x"82",
         14219 => x"72",
         14220 => x"54",
         14221 => x"06",
         14222 => x"54",
         14223 => x"b1",
         14224 => x"38",
         14225 => x"70",
         14226 => x"52",
         14227 => x"30",
         14228 => x"75",
         14229 => x"53",
         14230 => x"80",
         14231 => x"75",
         14232 => x"b9",
         14233 => x"3d",
         14234 => x"ed",
         14235 => x"a2",
         14236 => x"26",
         14237 => x"10",
         14238 => x"e0",
         14239 => x"08",
         14240 => x"16",
         14241 => x"ff",
         14242 => x"75",
         14243 => x"ff",
         14244 => x"83",
         14245 => x"57",
         14246 => x"88",
         14247 => x"ff",
         14248 => x"51",
         14249 => x"16",
         14250 => x"ff",
         14251 => x"db",
         14252 => x"70",
         14253 => x"06",
         14254 => x"39",
         14255 => x"83",
         14256 => x"57",
         14257 => x"f0",
         14258 => x"ff",
         14259 => x"51",
         14260 => x"75",
         14261 => x"06",
         14262 => x"70",
         14263 => x"06",
         14264 => x"ff",
         14265 => x"73",
         14266 => x"05",
         14267 => x"52",
         14268 => x"00",
         14269 => x"ff",
         14270 => x"ff",
         14271 => x"00",
         14272 => x"ff",
         14273 => x"19",
         14274 => x"19",
         14275 => x"19",
         14276 => x"19",
         14277 => x"19",
         14278 => x"19",
         14279 => x"19",
         14280 => x"19",
         14281 => x"19",
         14282 => x"19",
         14283 => x"19",
         14284 => x"19",
         14285 => x"19",
         14286 => x"18",
         14287 => x"18",
         14288 => x"18",
         14289 => x"18",
         14290 => x"18",
         14291 => x"18",
         14292 => x"18",
         14293 => x"1e",
         14294 => x"1f",
         14295 => x"1f",
         14296 => x"1f",
         14297 => x"1f",
         14298 => x"1f",
         14299 => x"1f",
         14300 => x"1f",
         14301 => x"1f",
         14302 => x"1f",
         14303 => x"1f",
         14304 => x"1f",
         14305 => x"1f",
         14306 => x"1f",
         14307 => x"1f",
         14308 => x"1f",
         14309 => x"1f",
         14310 => x"1f",
         14311 => x"1f",
         14312 => x"1f",
         14313 => x"1f",
         14314 => x"1f",
         14315 => x"1f",
         14316 => x"1f",
         14317 => x"1f",
         14318 => x"1f",
         14319 => x"1f",
         14320 => x"1f",
         14321 => x"1f",
         14322 => x"1f",
         14323 => x"1f",
         14324 => x"1f",
         14325 => x"1f",
         14326 => x"1f",
         14327 => x"1f",
         14328 => x"1f",
         14329 => x"1f",
         14330 => x"1f",
         14331 => x"1f",
         14332 => x"1f",
         14333 => x"1f",
         14334 => x"1f",
         14335 => x"1f",
         14336 => x"24",
         14337 => x"1f",
         14338 => x"1f",
         14339 => x"1f",
         14340 => x"1f",
         14341 => x"1f",
         14342 => x"1f",
         14343 => x"1f",
         14344 => x"1f",
         14345 => x"1f",
         14346 => x"1f",
         14347 => x"1f",
         14348 => x"1f",
         14349 => x"1f",
         14350 => x"1f",
         14351 => x"1f",
         14352 => x"1f",
         14353 => x"24",
         14354 => x"23",
         14355 => x"1f",
         14356 => x"22",
         14357 => x"24",
         14358 => x"23",
         14359 => x"22",
         14360 => x"21",
         14361 => x"1f",
         14362 => x"1f",
         14363 => x"1f",
         14364 => x"1f",
         14365 => x"1f",
         14366 => x"1f",
         14367 => x"1f",
         14368 => x"1f",
         14369 => x"1f",
         14370 => x"1f",
         14371 => x"1f",
         14372 => x"1f",
         14373 => x"1f",
         14374 => x"1f",
         14375 => x"1f",
         14376 => x"1f",
         14377 => x"1f",
         14378 => x"1f",
         14379 => x"1f",
         14380 => x"1f",
         14381 => x"1f",
         14382 => x"1f",
         14383 => x"1f",
         14384 => x"1f",
         14385 => x"1f",
         14386 => x"1f",
         14387 => x"1f",
         14388 => x"1f",
         14389 => x"1f",
         14390 => x"1f",
         14391 => x"1f",
         14392 => x"1f",
         14393 => x"1f",
         14394 => x"1f",
         14395 => x"1f",
         14396 => x"1f",
         14397 => x"1f",
         14398 => x"1f",
         14399 => x"1f",
         14400 => x"1f",
         14401 => x"1f",
         14402 => x"1f",
         14403 => x"1f",
         14404 => x"1f",
         14405 => x"1f",
         14406 => x"1f",
         14407 => x"1f",
         14408 => x"1f",
         14409 => x"1f",
         14410 => x"1f",
         14411 => x"1f",
         14412 => x"1f",
         14413 => x"21",
         14414 => x"21",
         14415 => x"1f",
         14416 => x"1f",
         14417 => x"1f",
         14418 => x"1f",
         14419 => x"1f",
         14420 => x"1f",
         14421 => x"1f",
         14422 => x"1f",
         14423 => x"21",
         14424 => x"21",
         14425 => x"1f",
         14426 => x"21",
         14427 => x"1f",
         14428 => x"21",
         14429 => x"21",
         14430 => x"21",
         14431 => x"32",
         14432 => x"32",
         14433 => x"32",
         14434 => x"32",
         14435 => x"32",
         14436 => x"32",
         14437 => x"3b",
         14438 => x"3a",
         14439 => x"39",
         14440 => x"36",
         14441 => x"3a",
         14442 => x"34",
         14443 => x"37",
         14444 => x"36",
         14445 => x"39",
         14446 => x"36",
         14447 => x"37",
         14448 => x"39",
         14449 => x"34",
         14450 => x"39",
         14451 => x"38",
         14452 => x"37",
         14453 => x"34",
         14454 => x"34",
         14455 => x"37",
         14456 => x"36",
         14457 => x"36",
         14458 => x"36",
         14459 => x"46",
         14460 => x"46",
         14461 => x"46",
         14462 => x"46",
         14463 => x"46",
         14464 => x"47",
         14465 => x"46",
         14466 => x"47",
         14467 => x"47",
         14468 => x"47",
         14469 => x"47",
         14470 => x"47",
         14471 => x"47",
         14472 => x"47",
         14473 => x"47",
         14474 => x"47",
         14475 => x"47",
         14476 => x"47",
         14477 => x"47",
         14478 => x"47",
         14479 => x"47",
         14480 => x"47",
         14481 => x"47",
         14482 => x"47",
         14483 => x"47",
         14484 => x"47",
         14485 => x"47",
         14486 => x"47",
         14487 => x"47",
         14488 => x"47",
         14489 => x"47",
         14490 => x"47",
         14491 => x"47",
         14492 => x"47",
         14493 => x"47",
         14494 => x"47",
         14495 => x"47",
         14496 => x"48",
         14497 => x"48",
         14498 => x"48",
         14499 => x"48",
         14500 => x"47",
         14501 => x"48",
         14502 => x"48",
         14503 => x"47",
         14504 => x"47",
         14505 => x"47",
         14506 => x"48",
         14507 => x"48",
         14508 => x"47",
         14509 => x"47",
         14510 => x"47",
         14511 => x"47",
         14512 => x"47",
         14513 => x"47",
         14514 => x"47",
         14515 => x"47",
         14516 => x"54",
         14517 => x"55",
         14518 => x"55",
         14519 => x"54",
         14520 => x"54",
         14521 => x"54",
         14522 => x"54",
         14523 => x"56",
         14524 => x"52",
         14525 => x"55",
         14526 => x"57",
         14527 => x"52",
         14528 => x"52",
         14529 => x"52",
         14530 => x"52",
         14531 => x"52",
         14532 => x"52",
         14533 => x"55",
         14534 => x"57",
         14535 => x"56",
         14536 => x"52",
         14537 => x"52",
         14538 => x"52",
         14539 => x"52",
         14540 => x"52",
         14541 => x"52",
         14542 => x"52",
         14543 => x"52",
         14544 => x"52",
         14545 => x"52",
         14546 => x"52",
         14547 => x"52",
         14548 => x"52",
         14549 => x"52",
         14550 => x"52",
         14551 => x"52",
         14552 => x"52",
         14553 => x"52",
         14554 => x"52",
         14555 => x"55",
         14556 => x"52",
         14557 => x"52",
         14558 => x"52",
         14559 => x"54",
         14560 => x"53",
         14561 => x"53",
         14562 => x"52",
         14563 => x"52",
         14564 => x"52",
         14565 => x"52",
         14566 => x"53",
         14567 => x"52",
         14568 => x"53",
         14569 => x"59",
         14570 => x"59",
         14571 => x"59",
         14572 => x"59",
         14573 => x"59",
         14574 => x"59",
         14575 => x"59",
         14576 => x"58",
         14577 => x"59",
         14578 => x"59",
         14579 => x"59",
         14580 => x"59",
         14581 => x"59",
         14582 => x"59",
         14583 => x"59",
         14584 => x"59",
         14585 => x"59",
         14586 => x"59",
         14587 => x"59",
         14588 => x"59",
         14589 => x"59",
         14590 => x"59",
         14591 => x"59",
         14592 => x"59",
         14593 => x"59",
         14594 => x"59",
         14595 => x"59",
         14596 => x"59",
         14597 => x"59",
         14598 => x"59",
         14599 => x"59",
         14600 => x"5a",
         14601 => x"59",
         14602 => x"59",
         14603 => x"59",
         14604 => x"5a",
         14605 => x"5a",
         14606 => x"5a",
         14607 => x"59",
         14608 => x"5a",
         14609 => x"5a",
         14610 => x"5a",
         14611 => x"5a",
         14612 => x"5a",
         14613 => x"59",
         14614 => x"59",
         14615 => x"59",
         14616 => x"59",
         14617 => x"59",
         14618 => x"59",
         14619 => x"63",
         14620 => x"61",
         14621 => x"61",
         14622 => x"61",
         14623 => x"61",
         14624 => x"61",
         14625 => x"61",
         14626 => x"61",
         14627 => x"61",
         14628 => x"61",
         14629 => x"61",
         14630 => x"61",
         14631 => x"61",
         14632 => x"61",
         14633 => x"5e",
         14634 => x"61",
         14635 => x"61",
         14636 => x"61",
         14637 => x"61",
         14638 => x"61",
         14639 => x"61",
         14640 => x"63",
         14641 => x"61",
         14642 => x"61",
         14643 => x"63",
         14644 => x"61",
         14645 => x"63",
         14646 => x"5e",
         14647 => x"63",
         14648 => x"de",
         14649 => x"de",
         14650 => x"de",
         14651 => x"de",
         14652 => x"de",
         14653 => x"de",
         14654 => x"de",
         14655 => x"de",
         14656 => x"de",
         14657 => x"0e",
         14658 => x"0b",
         14659 => x"0b",
         14660 => x"0f",
         14661 => x"0b",
         14662 => x"0b",
         14663 => x"0b",
         14664 => x"0b",
         14665 => x"0b",
         14666 => x"0b",
         14667 => x"0b",
         14668 => x"0d",
         14669 => x"0b",
         14670 => x"0f",
         14671 => x"0f",
         14672 => x"0b",
         14673 => x"0b",
         14674 => x"0b",
         14675 => x"0b",
         14676 => x"0b",
         14677 => x"0b",
         14678 => x"0b",
         14679 => x"0b",
         14680 => x"0b",
         14681 => x"0b",
         14682 => x"0b",
         14683 => x"0b",
         14684 => x"0b",
         14685 => x"0b",
         14686 => x"0b",
         14687 => x"0b",
         14688 => x"0b",
         14689 => x"0b",
         14690 => x"0b",
         14691 => x"0b",
         14692 => x"0b",
         14693 => x"0b",
         14694 => x"0b",
         14695 => x"0b",
         14696 => x"0b",
         14697 => x"0b",
         14698 => x"0b",
         14699 => x"0b",
         14700 => x"0b",
         14701 => x"0b",
         14702 => x"0b",
         14703 => x"0b",
         14704 => x"0b",
         14705 => x"0b",
         14706 => x"0b",
         14707 => x"0b",
         14708 => x"0f",
         14709 => x"0b",
         14710 => x"0b",
         14711 => x"0b",
         14712 => x"0b",
         14713 => x"0e",
         14714 => x"0b",
         14715 => x"0b",
         14716 => x"0b",
         14717 => x"0b",
         14718 => x"0b",
         14719 => x"0b",
         14720 => x"0b",
         14721 => x"0b",
         14722 => x"0b",
         14723 => x"0b",
         14724 => x"0e",
         14725 => x"0e",
         14726 => x"0e",
         14727 => x"0e",
         14728 => x"0e",
         14729 => x"0b",
         14730 => x"0e",
         14731 => x"0b",
         14732 => x"0b",
         14733 => x"0e",
         14734 => x"0b",
         14735 => x"0b",
         14736 => x"0c",
         14737 => x"0e",
         14738 => x"0b",
         14739 => x"0b",
         14740 => x"0f",
         14741 => x"0b",
         14742 => x"0c",
         14743 => x"0b",
         14744 => x"0b",
         14745 => x"0e",
         14746 => x"6e",
         14747 => x"00",
         14748 => x"6f",
         14749 => x"00",
         14750 => x"6e",
         14751 => x"00",
         14752 => x"6f",
         14753 => x"00",
         14754 => x"78",
         14755 => x"00",
         14756 => x"6c",
         14757 => x"00",
         14758 => x"6f",
         14759 => x"00",
         14760 => x"69",
         14761 => x"00",
         14762 => x"75",
         14763 => x"00",
         14764 => x"62",
         14765 => x"68",
         14766 => x"77",
         14767 => x"64",
         14768 => x"65",
         14769 => x"64",
         14770 => x"65",
         14771 => x"6c",
         14772 => x"00",
         14773 => x"70",
         14774 => x"73",
         14775 => x"74",
         14776 => x"73",
         14777 => x"00",
         14778 => x"66",
         14779 => x"00",
         14780 => x"73",
         14781 => x"00",
         14782 => x"73",
         14783 => x"30",
         14784 => x"61",
         14785 => x"00",
         14786 => x"61",
         14787 => x"00",
         14788 => x"6c",
         14789 => x"00",
         14790 => x"00",
         14791 => x"6b",
         14792 => x"6e",
         14793 => x"72",
         14794 => x"00",
         14795 => x"72",
         14796 => x"74",
         14797 => x"20",
         14798 => x"6f",
         14799 => x"63",
         14800 => x"00",
         14801 => x"6f",
         14802 => x"6e",
         14803 => x"70",
         14804 => x"66",
         14805 => x"73",
         14806 => x"00",
         14807 => x"73",
         14808 => x"69",
         14809 => x"6e",
         14810 => x"65",
         14811 => x"79",
         14812 => x"00",
         14813 => x"6c",
         14814 => x"73",
         14815 => x"63",
         14816 => x"2e",
         14817 => x"6d",
         14818 => x"74",
         14819 => x"70",
         14820 => x"74",
         14821 => x"20",
         14822 => x"63",
         14823 => x"65",
         14824 => x"00",
         14825 => x"72",
         14826 => x"20",
         14827 => x"72",
         14828 => x"2e",
         14829 => x"20",
         14830 => x"70",
         14831 => x"62",
         14832 => x"66",
         14833 => x"73",
         14834 => x"65",
         14835 => x"6f",
         14836 => x"20",
         14837 => x"64",
         14838 => x"2e",
         14839 => x"73",
         14840 => x"6f",
         14841 => x"6e",
         14842 => x"65",
         14843 => x"00",
         14844 => x"69",
         14845 => x"6e",
         14846 => x"65",
         14847 => x"73",
         14848 => x"76",
         14849 => x"64",
         14850 => x"00",
         14851 => x"20",
         14852 => x"77",
         14853 => x"65",
         14854 => x"6f",
         14855 => x"74",
         14856 => x"00",
         14857 => x"6c",
         14858 => x"61",
         14859 => x"65",
         14860 => x"76",
         14861 => x"64",
         14862 => x"00",
         14863 => x"6c",
         14864 => x"6c",
         14865 => x"64",
         14866 => x"78",
         14867 => x"73",
         14868 => x"00",
         14869 => x"63",
         14870 => x"20",
         14871 => x"69",
         14872 => x"00",
         14873 => x"76",
         14874 => x"64",
         14875 => x"6c",
         14876 => x"6d",
         14877 => x"00",
         14878 => x"20",
         14879 => x"68",
         14880 => x"75",
         14881 => x"00",
         14882 => x"20",
         14883 => x"65",
         14884 => x"75",
         14885 => x"00",
         14886 => x"73",
         14887 => x"6f",
         14888 => x"65",
         14889 => x"2e",
         14890 => x"74",
         14891 => x"61",
         14892 => x"72",
         14893 => x"2e",
         14894 => x"73",
         14895 => x"72",
         14896 => x"00",
         14897 => x"63",
         14898 => x"73",
         14899 => x"00",
         14900 => x"6c",
         14901 => x"79",
         14902 => x"20",
         14903 => x"61",
         14904 => x"6c",
         14905 => x"79",
         14906 => x"2f",
         14907 => x"2e",
         14908 => x"00",
         14909 => x"61",
         14910 => x"00",
         14911 => x"38",
         14912 => x"00",
         14913 => x"20",
         14914 => x"32",
         14915 => x"00",
         14916 => x"00",
         14917 => x"00",
         14918 => x"00",
         14919 => x"34",
         14920 => x"00",
         14921 => x"20",
         14922 => x"20",
         14923 => x"00",
         14924 => x"53",
         14925 => x"20",
         14926 => x"28",
         14927 => x"2f",
         14928 => x"32",
         14929 => x"00",
         14930 => x"2e",
         14931 => x"00",
         14932 => x"50",
         14933 => x"72",
         14934 => x"25",
         14935 => x"29",
         14936 => x"20",
         14937 => x"2a",
         14938 => x"00",
         14939 => x"3a",
         14940 => x"20",
         14941 => x"73",
         14942 => x"64",
         14943 => x"73",
         14944 => x"20",
         14945 => x"20",
         14946 => x"20",
         14947 => x"20",
         14948 => x"6c",
         14949 => x"00",
         14950 => x"20",
         14951 => x"70",
         14952 => x"64",
         14953 => x"73",
         14954 => x"20",
         14955 => x"20",
         14956 => x"20",
         14957 => x"20",
         14958 => x"6c",
         14959 => x"00",
         14960 => x"55",
         14961 => x"74",
         14962 => x"75",
         14963 => x"48",
         14964 => x"6c",
         14965 => x"00",
         14966 => x"52",
         14967 => x"54",
         14968 => x"6e",
         14969 => x"72",
         14970 => x"00",
         14971 => x"52",
         14972 => x"52",
         14973 => x"6e",
         14974 => x"72",
         14975 => x"00",
         14976 => x"52",
         14977 => x"54",
         14978 => x"6e",
         14979 => x"72",
         14980 => x"00",
         14981 => x"52",
         14982 => x"52",
         14983 => x"6e",
         14984 => x"72",
         14985 => x"00",
         14986 => x"43",
         14987 => x"57",
         14988 => x"6e",
         14989 => x"72",
         14990 => x"00",
         14991 => x"43",
         14992 => x"52",
         14993 => x"6e",
         14994 => x"72",
         14995 => x"00",
         14996 => x"32",
         14997 => x"74",
         14998 => x"75",
         14999 => x"00",
         15000 => x"6d",
         15001 => x"69",
         15002 => x"72",
         15003 => x"74",
         15004 => x"74",
         15005 => x"67",
         15006 => x"20",
         15007 => x"65",
         15008 => x"2e",
         15009 => x"61",
         15010 => x"6e",
         15011 => x"69",
         15012 => x"2e",
         15013 => x"00",
         15014 => x"74",
         15015 => x"65",
         15016 => x"61",
         15017 => x"00",
         15018 => x"53",
         15019 => x"75",
         15020 => x"74",
         15021 => x"69",
         15022 => x"20",
         15023 => x"69",
         15024 => x"69",
         15025 => x"73",
         15026 => x"64",
         15027 => x"72",
         15028 => x"2c",
         15029 => x"65",
         15030 => x"20",
         15031 => x"74",
         15032 => x"6e",
         15033 => x"6c",
         15034 => x"00",
         15035 => x"00",
         15036 => x"3a",
         15037 => x"00",
         15038 => x"00",
         15039 => x"64",
         15040 => x"6d",
         15041 => x"64",
         15042 => x"00",
         15043 => x"55",
         15044 => x"6e",
         15045 => x"3a",
         15046 => x"5c",
         15047 => x"25",
         15048 => x"00",
         15049 => x"6c",
         15050 => x"65",
         15051 => x"74",
         15052 => x"2e",
         15053 => x"00",
         15054 => x"73",
         15055 => x"74",
         15056 => x"20",
         15057 => x"6c",
         15058 => x"74",
         15059 => x"2e",
         15060 => x"00",
         15061 => x"6c",
         15062 => x"67",
         15063 => x"64",
         15064 => x"20",
         15065 => x"6c",
         15066 => x"2e",
         15067 => x"00",
         15068 => x"6c",
         15069 => x"65",
         15070 => x"6e",
         15071 => x"63",
         15072 => x"20",
         15073 => x"29",
         15074 => x"00",
         15075 => x"65",
         15076 => x"69",
         15077 => x"63",
         15078 => x"20",
         15079 => x"30",
         15080 => x"20",
         15081 => x"0a",
         15082 => x"38",
         15083 => x"25",
         15084 => x"58",
         15085 => x"00",
         15086 => x"38",
         15087 => x"25",
         15088 => x"2d",
         15089 => x"6d",
         15090 => x"69",
         15091 => x"2e",
         15092 => x"00",
         15093 => x"38",
         15094 => x"25",
         15095 => x"29",
         15096 => x"30",
         15097 => x"28",
         15098 => x"78",
         15099 => x"00",
         15100 => x"70",
         15101 => x"67",
         15102 => x"00",
         15103 => x"38",
         15104 => x"25",
         15105 => x"2d",
         15106 => x"65",
         15107 => x"6e",
         15108 => x"2e",
         15109 => x"00",
         15110 => x"6d",
         15111 => x"65",
         15112 => x"79",
         15113 => x"6f",
         15114 => x"65",
         15115 => x"00",
         15116 => x"3a",
         15117 => x"5c",
         15118 => x"00",
         15119 => x"6d",
         15120 => x"20",
         15121 => x"61",
         15122 => x"65",
         15123 => x"63",
         15124 => x"6f",
         15125 => x"72",
         15126 => x"73",
         15127 => x"6f",
         15128 => x"6e",
         15129 => x"00",
         15130 => x"3f",
         15131 => x"2f",
         15132 => x"25",
         15133 => x"64",
         15134 => x"3a",
         15135 => x"25",
         15136 => x"0a",
         15137 => x"43",
         15138 => x"6e",
         15139 => x"75",
         15140 => x"69",
         15141 => x"00",
         15142 => x"44",
         15143 => x"63",
         15144 => x"69",
         15145 => x"65",
         15146 => x"74",
         15147 => x"00",
         15148 => x"64",
         15149 => x"73",
         15150 => x"00",
         15151 => x"20",
         15152 => x"55",
         15153 => x"73",
         15154 => x"56",
         15155 => x"6f",
         15156 => x"64",
         15157 => x"73",
         15158 => x"20",
         15159 => x"58",
         15160 => x"00",
         15161 => x"20",
         15162 => x"55",
         15163 => x"6d",
         15164 => x"20",
         15165 => x"72",
         15166 => x"64",
         15167 => x"73",
         15168 => x"20",
         15169 => x"58",
         15170 => x"00",
         15171 => x"20",
         15172 => x"61",
         15173 => x"53",
         15174 => x"74",
         15175 => x"64",
         15176 => x"73",
         15177 => x"20",
         15178 => x"20",
         15179 => x"58",
         15180 => x"00",
         15181 => x"73",
         15182 => x"00",
         15183 => x"20",
         15184 => x"55",
         15185 => x"20",
         15186 => x"20",
         15187 => x"20",
         15188 => x"20",
         15189 => x"20",
         15190 => x"20",
         15191 => x"58",
         15192 => x"00",
         15193 => x"20",
         15194 => x"73",
         15195 => x"20",
         15196 => x"63",
         15197 => x"72",
         15198 => x"20",
         15199 => x"20",
         15200 => x"20",
         15201 => x"25",
         15202 => x"4d",
         15203 => x"00",
         15204 => x"20",
         15205 => x"73",
         15206 => x"6e",
         15207 => x"44",
         15208 => x"20",
         15209 => x"63",
         15210 => x"72",
         15211 => x"20",
         15212 => x"25",
         15213 => x"4d",
         15214 => x"00",
         15215 => x"20",
         15216 => x"52",
         15217 => x"43",
         15218 => x"6b",
         15219 => x"65",
         15220 => x"20",
         15221 => x"20",
         15222 => x"20",
         15223 => x"25",
         15224 => x"4d",
         15225 => x"00",
         15226 => x"20",
         15227 => x"49",
         15228 => x"20",
         15229 => x"32",
         15230 => x"20",
         15231 => x"43",
         15232 => x"00",
         15233 => x"20",
         15234 => x"20",
         15235 => x"00",
         15236 => x"20",
         15237 => x"53",
         15238 => x"4e",
         15239 => x"55",
         15240 => x"00",
         15241 => x"20",
         15242 => x"54",
         15243 => x"54",
         15244 => x"28",
         15245 => x"6e",
         15246 => x"73",
         15247 => x"32",
         15248 => x"0a",
         15249 => x"20",
         15250 => x"4d",
         15251 => x"20",
         15252 => x"28",
         15253 => x"65",
         15254 => x"20",
         15255 => x"32",
         15256 => x"0a",
         15257 => x"20",
         15258 => x"20",
         15259 => x"44",
         15260 => x"28",
         15261 => x"69",
         15262 => x"20",
         15263 => x"32",
         15264 => x"0a",
         15265 => x"20",
         15266 => x"4d",
         15267 => x"20",
         15268 => x"28",
         15269 => x"58",
         15270 => x"38",
         15271 => x"0a",
         15272 => x"20",
         15273 => x"41",
         15274 => x"20",
         15275 => x"28",
         15276 => x"58",
         15277 => x"38",
         15278 => x"0a",
         15279 => x"20",
         15280 => x"53",
         15281 => x"52",
         15282 => x"28",
         15283 => x"58",
         15284 => x"38",
         15285 => x"0a",
         15286 => x"20",
         15287 => x"52",
         15288 => x"20",
         15289 => x"28",
         15290 => x"58",
         15291 => x"38",
         15292 => x"0a",
         15293 => x"20",
         15294 => x"20",
         15295 => x"41",
         15296 => x"28",
         15297 => x"58",
         15298 => x"38",
         15299 => x"0a",
         15300 => x"66",
         15301 => x"20",
         15302 => x"20",
         15303 => x"66",
         15304 => x"00",
         15305 => x"6b",
         15306 => x"6e",
         15307 => x"4f",
         15308 => x"00",
         15309 => x"61",
         15310 => x"00",
         15311 => x"64",
         15312 => x"00",
         15313 => x"65",
         15314 => x"00",
         15315 => x"4f",
         15316 => x"f0",
         15317 => x"00",
         15318 => x"00",
         15319 => x"f0",
         15320 => x"00",
         15321 => x"00",
         15322 => x"f0",
         15323 => x"00",
         15324 => x"00",
         15325 => x"f0",
         15326 => x"00",
         15327 => x"00",
         15328 => x"f0",
         15329 => x"00",
         15330 => x"00",
         15331 => x"f0",
         15332 => x"00",
         15333 => x"00",
         15334 => x"f0",
         15335 => x"00",
         15336 => x"00",
         15337 => x"f0",
         15338 => x"00",
         15339 => x"00",
         15340 => x"f0",
         15341 => x"00",
         15342 => x"00",
         15343 => x"f0",
         15344 => x"00",
         15345 => x"00",
         15346 => x"f0",
         15347 => x"00",
         15348 => x"00",
         15349 => x"f0",
         15350 => x"00",
         15351 => x"00",
         15352 => x"f0",
         15353 => x"00",
         15354 => x"00",
         15355 => x"f0",
         15356 => x"00",
         15357 => x"00",
         15358 => x"f0",
         15359 => x"00",
         15360 => x"00",
         15361 => x"f0",
         15362 => x"00",
         15363 => x"00",
         15364 => x"f0",
         15365 => x"00",
         15366 => x"00",
         15367 => x"f0",
         15368 => x"00",
         15369 => x"00",
         15370 => x"f0",
         15371 => x"00",
         15372 => x"00",
         15373 => x"f0",
         15374 => x"00",
         15375 => x"00",
         15376 => x"f0",
         15377 => x"00",
         15378 => x"00",
         15379 => x"f0",
         15380 => x"00",
         15381 => x"00",
         15382 => x"44",
         15383 => x"43",
         15384 => x"42",
         15385 => x"41",
         15386 => x"36",
         15387 => x"35",
         15388 => x"34",
         15389 => x"46",
         15390 => x"33",
         15391 => x"32",
         15392 => x"31",
         15393 => x"00",
         15394 => x"00",
         15395 => x"00",
         15396 => x"00",
         15397 => x"00",
         15398 => x"00",
         15399 => x"00",
         15400 => x"00",
         15401 => x"00",
         15402 => x"00",
         15403 => x"00",
         15404 => x"6e",
         15405 => x"20",
         15406 => x"6e",
         15407 => x"65",
         15408 => x"20",
         15409 => x"74",
         15410 => x"20",
         15411 => x"65",
         15412 => x"69",
         15413 => x"6c",
         15414 => x"2e",
         15415 => x"73",
         15416 => x"79",
         15417 => x"73",
         15418 => x"00",
         15419 => x"00",
         15420 => x"36",
         15421 => x"20",
         15422 => x"00",
         15423 => x"69",
         15424 => x"20",
         15425 => x"72",
         15426 => x"74",
         15427 => x"65",
         15428 => x"73",
         15429 => x"79",
         15430 => x"6c",
         15431 => x"6f",
         15432 => x"46",
         15433 => x"00",
         15434 => x"73",
         15435 => x"00",
         15436 => x"31",
         15437 => x"00",
         15438 => x"41",
         15439 => x"42",
         15440 => x"43",
         15441 => x"44",
         15442 => x"31",
         15443 => x"00",
         15444 => x"31",
         15445 => x"00",
         15446 => x"31",
         15447 => x"00",
         15448 => x"31",
         15449 => x"00",
         15450 => x"31",
         15451 => x"00",
         15452 => x"31",
         15453 => x"00",
         15454 => x"31",
         15455 => x"00",
         15456 => x"31",
         15457 => x"00",
         15458 => x"31",
         15459 => x"00",
         15460 => x"32",
         15461 => x"00",
         15462 => x"32",
         15463 => x"00",
         15464 => x"33",
         15465 => x"00",
         15466 => x"46",
         15467 => x"35",
         15468 => x"00",
         15469 => x"36",
         15470 => x"00",
         15471 => x"25",
         15472 => x"64",
         15473 => x"2c",
         15474 => x"25",
         15475 => x"64",
         15476 => x"32",
         15477 => x"00",
         15478 => x"25",
         15479 => x"64",
         15480 => x"3a",
         15481 => x"25",
         15482 => x"64",
         15483 => x"3a",
         15484 => x"2c",
         15485 => x"25",
         15486 => x"00",
         15487 => x"32",
         15488 => x"00",
         15489 => x"5b",
         15490 => x"25",
         15491 => x"00",
         15492 => x"70",
         15493 => x"20",
         15494 => x"73",
         15495 => x"00",
         15496 => x"3a",
         15497 => x"78",
         15498 => x"32",
         15499 => x"00",
         15500 => x"3a",
         15501 => x"78",
         15502 => x"32",
         15503 => x"00",
         15504 => x"3a",
         15505 => x"78",
         15506 => x"00",
         15507 => x"20",
         15508 => x"74",
         15509 => x"66",
         15510 => x"64",
         15511 => x"00",
         15512 => x"00",
         15513 => x"3a",
         15514 => x"7c",
         15515 => x"00",
         15516 => x"3b",
         15517 => x"00",
         15518 => x"54",
         15519 => x"54",
         15520 => x"00",
         15521 => x"90",
         15522 => x"4f",
         15523 => x"30",
         15524 => x"20",
         15525 => x"45",
         15526 => x"20",
         15527 => x"20",
         15528 => x"20",
         15529 => x"20",
         15530 => x"45",
         15531 => x"20",
         15532 => x"33",
         15533 => x"20",
         15534 => x"f2",
         15535 => x"00",
         15536 => x"00",
         15537 => x"00",
         15538 => x"05",
         15539 => x"10",
         15540 => x"18",
         15541 => x"00",
         15542 => x"45",
         15543 => x"8f",
         15544 => x"45",
         15545 => x"8e",
         15546 => x"92",
         15547 => x"55",
         15548 => x"9a",
         15549 => x"9e",
         15550 => x"4f",
         15551 => x"a6",
         15552 => x"aa",
         15553 => x"ae",
         15554 => x"b2",
         15555 => x"b6",
         15556 => x"ba",
         15557 => x"be",
         15558 => x"c2",
         15559 => x"c6",
         15560 => x"ca",
         15561 => x"ce",
         15562 => x"d2",
         15563 => x"d6",
         15564 => x"da",
         15565 => x"de",
         15566 => x"e2",
         15567 => x"e6",
         15568 => x"ea",
         15569 => x"ee",
         15570 => x"f2",
         15571 => x"f6",
         15572 => x"fa",
         15573 => x"fe",
         15574 => x"2c",
         15575 => x"5d",
         15576 => x"2a",
         15577 => x"3f",
         15578 => x"00",
         15579 => x"00",
         15580 => x"00",
         15581 => x"02",
         15582 => x"00",
         15583 => x"00",
         15584 => x"00",
         15585 => x"00",
         15586 => x"00",
         15587 => x"00",
         15588 => x"00",
         15589 => x"00",
         15590 => x"00",
         15591 => x"00",
         15592 => x"00",
         15593 => x"00",
         15594 => x"00",
         15595 => x"00",
         15596 => x"00",
         15597 => x"00",
         15598 => x"00",
         15599 => x"00",
         15600 => x"00",
         15601 => x"00",
         15602 => x"01",
         15603 => x"00",
         15604 => x"00",
         15605 => x"00",
         15606 => x"00",
         15607 => x"23",
         15608 => x"00",
         15609 => x"00",
         15610 => x"00",
         15611 => x"25",
         15612 => x"25",
         15613 => x"25",
         15614 => x"25",
         15615 => x"25",
         15616 => x"25",
         15617 => x"25",
         15618 => x"25",
         15619 => x"25",
         15620 => x"25",
         15621 => x"25",
         15622 => x"25",
         15623 => x"25",
         15624 => x"25",
         15625 => x"25",
         15626 => x"25",
         15627 => x"25",
         15628 => x"25",
         15629 => x"25",
         15630 => x"25",
         15631 => x"25",
         15632 => x"25",
         15633 => x"25",
         15634 => x"25",
         15635 => x"00",
         15636 => x"03",
         15637 => x"03",
         15638 => x"03",
         15639 => x"03",
         15640 => x"03",
         15641 => x"03",
         15642 => x"22",
         15643 => x"00",
         15644 => x"22",
         15645 => x"23",
         15646 => x"22",
         15647 => x"22",
         15648 => x"22",
         15649 => x"00",
         15650 => x"00",
         15651 => x"03",
         15652 => x"03",
         15653 => x"03",
         15654 => x"00",
         15655 => x"01",
         15656 => x"01",
         15657 => x"01",
         15658 => x"01",
         15659 => x"01",
         15660 => x"01",
         15661 => x"02",
         15662 => x"01",
         15663 => x"01",
         15664 => x"01",
         15665 => x"01",
         15666 => x"01",
         15667 => x"01",
         15668 => x"01",
         15669 => x"01",
         15670 => x"01",
         15671 => x"01",
         15672 => x"01",
         15673 => x"01",
         15674 => x"02",
         15675 => x"01",
         15676 => x"02",
         15677 => x"01",
         15678 => x"01",
         15679 => x"01",
         15680 => x"01",
         15681 => x"01",
         15682 => x"01",
         15683 => x"01",
         15684 => x"01",
         15685 => x"01",
         15686 => x"01",
         15687 => x"01",
         15688 => x"01",
         15689 => x"01",
         15690 => x"01",
         15691 => x"01",
         15692 => x"01",
         15693 => x"01",
         15694 => x"01",
         15695 => x"01",
         15696 => x"01",
         15697 => x"01",
         15698 => x"01",
         15699 => x"01",
         15700 => x"01",
         15701 => x"00",
         15702 => x"01",
         15703 => x"01",
         15704 => x"01",
         15705 => x"01",
         15706 => x"01",
         15707 => x"01",
         15708 => x"00",
         15709 => x"02",
         15710 => x"02",
         15711 => x"02",
         15712 => x"02",
         15713 => x"02",
         15714 => x"02",
         15715 => x"01",
         15716 => x"02",
         15717 => x"01",
         15718 => x"01",
         15719 => x"01",
         15720 => x"02",
         15721 => x"02",
         15722 => x"02",
         15723 => x"01",
         15724 => x"02",
         15725 => x"02",
         15726 => x"01",
         15727 => x"2c",
         15728 => x"02",
         15729 => x"01",
         15730 => x"02",
         15731 => x"02",
         15732 => x"01",
         15733 => x"02",
         15734 => x"02",
         15735 => x"02",
         15736 => x"2c",
         15737 => x"02",
         15738 => x"02",
         15739 => x"01",
         15740 => x"02",
         15741 => x"02",
         15742 => x"02",
         15743 => x"01",
         15744 => x"02",
         15745 => x"02",
         15746 => x"02",
         15747 => x"03",
         15748 => x"03",
         15749 => x"03",
         15750 => x"00",
         15751 => x"03",
         15752 => x"03",
         15753 => x"03",
         15754 => x"00",
         15755 => x"03",
         15756 => x"03",
         15757 => x"00",
         15758 => x"03",
         15759 => x"03",
         15760 => x"03",
         15761 => x"03",
         15762 => x"03",
         15763 => x"03",
         15764 => x"03",
         15765 => x"03",
         15766 => x"04",
         15767 => x"04",
         15768 => x"04",
         15769 => x"04",
         15770 => x"04",
         15771 => x"04",
         15772 => x"04",
         15773 => x"01",
         15774 => x"04",
         15775 => x"00",
         15776 => x"00",
         15777 => x"1e",
         15778 => x"1e",
         15779 => x"1f",
         15780 => x"1f",
         15781 => x"1f",
         15782 => x"1f",
         15783 => x"1f",
         15784 => x"1f",
         15785 => x"1f",
         15786 => x"1f",
         15787 => x"1f",
         15788 => x"1f",
         15789 => x"06",
         15790 => x"00",
         15791 => x"1f",
         15792 => x"1f",
         15793 => x"1f",
         15794 => x"1f",
         15795 => x"1f",
         15796 => x"1f",
         15797 => x"1f",
         15798 => x"06",
         15799 => x"06",
         15800 => x"06",
         15801 => x"00",
         15802 => x"1f",
         15803 => x"1f",
         15804 => x"00",
         15805 => x"1f",
         15806 => x"1f",
         15807 => x"1f",
         15808 => x"1f",
         15809 => x"00",
         15810 => x"21",
         15811 => x"21",
         15812 => x"02",
         15813 => x"00",
         15814 => x"24",
         15815 => x"2c",
         15816 => x"2c",
         15817 => x"2c",
         15818 => x"2c",
         15819 => x"2c",
         15820 => x"2d",
         15821 => x"ff",
         15822 => x"00",
         15823 => x"00",
         15824 => x"e6",
         15825 => x"01",
         15826 => x"00",
         15827 => x"00",
         15828 => x"e6",
         15829 => x"01",
         15830 => x"00",
         15831 => x"00",
         15832 => x"e6",
         15833 => x"03",
         15834 => x"00",
         15835 => x"00",
         15836 => x"e6",
         15837 => x"03",
         15838 => x"00",
         15839 => x"00",
         15840 => x"e6",
         15841 => x"03",
         15842 => x"00",
         15843 => x"00",
         15844 => x"e6",
         15845 => x"04",
         15846 => x"00",
         15847 => x"00",
         15848 => x"e6",
         15849 => x"04",
         15850 => x"00",
         15851 => x"00",
         15852 => x"e6",
         15853 => x"04",
         15854 => x"00",
         15855 => x"00",
         15856 => x"e6",
         15857 => x"04",
         15858 => x"00",
         15859 => x"00",
         15860 => x"e6",
         15861 => x"04",
         15862 => x"00",
         15863 => x"00",
         15864 => x"e6",
         15865 => x"04",
         15866 => x"00",
         15867 => x"00",
         15868 => x"e6",
         15869 => x"04",
         15870 => x"00",
         15871 => x"00",
         15872 => x"e6",
         15873 => x"05",
         15874 => x"00",
         15875 => x"00",
         15876 => x"e6",
         15877 => x"05",
         15878 => x"00",
         15879 => x"00",
         15880 => x"e6",
         15881 => x"05",
         15882 => x"00",
         15883 => x"00",
         15884 => x"e6",
         15885 => x"05",
         15886 => x"00",
         15887 => x"00",
         15888 => x"e6",
         15889 => x"07",
         15890 => x"00",
         15891 => x"00",
         15892 => x"e6",
         15893 => x"07",
         15894 => x"00",
         15895 => x"00",
         15896 => x"e6",
         15897 => x"08",
         15898 => x"00",
         15899 => x"00",
         15900 => x"e6",
         15901 => x"08",
         15902 => x"00",
         15903 => x"00",
         15904 => x"e6",
         15905 => x"08",
         15906 => x"00",
         15907 => x"00",
         15908 => x"e6",
         15909 => x"08",
         15910 => x"00",
         15911 => x"00",
         15912 => x"e6",
         15913 => x"08",
         15914 => x"00",
         15915 => x"00",
         15916 => x"e6",
         15917 => x"08",
         15918 => x"00",
         15919 => x"00",
         15920 => x"e7",
         15921 => x"09",
         15922 => x"00",
         15923 => x"00",
         15924 => x"e7",
         15925 => x"09",
         15926 => x"00",
         15927 => x"00",
         15928 => x"e7",
         15929 => x"09",
         15930 => x"00",
         15931 => x"00",
         15932 => x"e7",
         15933 => x"09",
         15934 => x"00",
         15935 => x"00",
         15936 => x"00",
         15937 => x"00",
         15938 => x"7f",
         15939 => x"00",
         15940 => x"7f",
         15941 => x"00",
         15942 => x"7f",
         15943 => x"00",
         15944 => x"00",
         15945 => x"00",
         15946 => x"ff",
         15947 => x"00",
         15948 => x"00",
         15949 => x"78",
         15950 => x"00",
         15951 => x"e1",
         15952 => x"e1",
         15953 => x"e1",
         15954 => x"00",
         15955 => x"01",
         15956 => x"01",
         15957 => x"10",
         15958 => x"00",
         15959 => x"00",
         15960 => x"00",
         15961 => x"00",
         15962 => x"00",
         15963 => x"00",
         15964 => x"00",
         15965 => x"00",
         15966 => x"00",
         15967 => x"00",
         15968 => x"00",
         15969 => x"00",
         15970 => x"00",
         15971 => x"00",
         15972 => x"00",
         15973 => x"00",
         15974 => x"00",
         15975 => x"00",
         15976 => x"00",
         15977 => x"00",
         15978 => x"00",
         15979 => x"00",
         15980 => x"00",
         15981 => x"00",
         15982 => x"00",
         15983 => x"f0",
         15984 => x"00",
         15985 => x"f0",
         15986 => x"00",
         15987 => x"f0",
         15988 => x"00",
         15989 => x"fd",
         15990 => x"5f",
         15991 => x"3a",
         15992 => x"40",
         15993 => x"f0",
         15994 => x"73",
         15995 => x"77",
         15996 => x"6b",
         15997 => x"6f",
         15998 => x"63",
         15999 => x"67",
         16000 => x"33",
         16001 => x"37",
         16002 => x"2d",
         16003 => x"2c",
         16004 => x"f3",
         16005 => x"3f",
         16006 => x"f0",
         16007 => x"f0",
         16008 => x"82",
         16009 => x"f0",
         16010 => x"58",
         16011 => x"3b",
         16012 => x"40",
         16013 => x"f0",
         16014 => x"53",
         16015 => x"57",
         16016 => x"4b",
         16017 => x"4f",
         16018 => x"43",
         16019 => x"47",
         16020 => x"33",
         16021 => x"37",
         16022 => x"2d",
         16023 => x"2c",
         16024 => x"f3",
         16025 => x"3f",
         16026 => x"f0",
         16027 => x"f0",
         16028 => x"82",
         16029 => x"f0",
         16030 => x"58",
         16031 => x"2a",
         16032 => x"60",
         16033 => x"f0",
         16034 => x"53",
         16035 => x"57",
         16036 => x"4b",
         16037 => x"4f",
         16038 => x"43",
         16039 => x"47",
         16040 => x"23",
         16041 => x"27",
         16042 => x"3d",
         16043 => x"3c",
         16044 => x"e0",
         16045 => x"3f",
         16046 => x"f0",
         16047 => x"f0",
         16048 => x"87",
         16049 => x"f0",
         16050 => x"1e",
         16051 => x"f0",
         16052 => x"00",
         16053 => x"f0",
         16054 => x"13",
         16055 => x"17",
         16056 => x"0b",
         16057 => x"0f",
         16058 => x"03",
         16059 => x"07",
         16060 => x"f0",
         16061 => x"f0",
         16062 => x"f0",
         16063 => x"f0",
         16064 => x"f0",
         16065 => x"f0",
         16066 => x"f0",
         16067 => x"f0",
         16068 => x"82",
         16069 => x"f0",
         16070 => x"cf",
         16071 => x"4d",
         16072 => x"d7",
         16073 => x"f0",
         16074 => x"41",
         16075 => x"78",
         16076 => x"6c",
         16077 => x"d5",
         16078 => x"d9",
         16079 => x"4c",
         16080 => x"7e",
         16081 => x"5f",
         16082 => x"d1",
         16083 => x"d0",
         16084 => x"c2",
         16085 => x"bb",
         16086 => x"f0",
         16087 => x"f0",
         16088 => x"82",
         16089 => x"f0",
         16090 => x"00",
         16091 => x"00",
         16092 => x"00",
         16093 => x"00",
         16094 => x"00",
         16095 => x"00",
         16096 => x"00",
         16097 => x"00",
         16098 => x"00",
         16099 => x"00",
         16100 => x"00",
         16101 => x"00",
         16102 => x"00",
         16103 => x"00",
         16104 => x"00",
         16105 => x"00",
         16106 => x"00",
         16107 => x"00",
         16108 => x"00",
         16109 => x"00",
         16110 => x"00",
         16111 => x"00",
         16112 => x"00",
         16113 => x"00",
         16114 => x"00",
         16115 => x"00",
         16116 => x"00",
         16117 => x"00",
         16118 => x"f1",
         16119 => x"00",
         16120 => x"f1",
         16121 => x"00",
         16122 => x"f1",
         16123 => x"00",
         16124 => x"f1",
         16125 => x"00",
         16126 => x"f1",
         16127 => x"00",
         16128 => x"f1",
         16129 => x"00",
         16130 => x"f1",
         16131 => x"00",
         16132 => x"f1",
         16133 => x"00",
         16134 => x"f1",
         16135 => x"00",
         16136 => x"f1",
         16137 => x"00",
         16138 => x"f1",
         16139 => x"00",
         16140 => x"f1",
         16141 => x"00",
         16142 => x"f1",
         16143 => x"00",
         16144 => x"f1",
         16145 => x"00",
         16146 => x"f1",
         16147 => x"00",
         16148 => x"f1",
         16149 => x"00",
         16150 => x"f1",
         16151 => x"00",
         16152 => x"f1",
         16153 => x"00",
         16154 => x"f1",
         16155 => x"00",
         16156 => x"f1",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"00",
         16166 => x"00",
         16167 => x"00",
         16168 => x"00",
         16169 => x"00",
         16170 => x"00",
         16171 => x"00",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"32",
         18159 => x"01",
         18160 => x"00",
         18161 => x"f2",
         18162 => x"f6",
         18163 => x"fa",
         18164 => x"fe",
         18165 => x"c2",
         18166 => x"c6",
         18167 => x"e5",
         18168 => x"ef",
         18169 => x"62",
         18170 => x"66",
         18171 => x"6b",
         18172 => x"2e",
         18173 => x"22",
         18174 => x"26",
         18175 => x"4f",
         18176 => x"57",
         18177 => x"02",
         18178 => x"06",
         18179 => x"0a",
         18180 => x"0e",
         18181 => x"12",
         18182 => x"16",
         18183 => x"1a",
         18184 => x"be",
         18185 => x"82",
         18186 => x"86",
         18187 => x"8a",
         18188 => x"8e",
         18189 => x"92",
         18190 => x"96",
         18191 => x"9a",
         18192 => x"a5",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"00",
         18199 => x"00",
         18200 => x"00",
         18201 => x"00",
         18202 => x"00",
         18203 => x"00",
         18204 => x"00",
         18205 => x"00",
         18206 => x"00",
         18207 => x"00",
         18208 => x"00",
         18209 => x"00",
         18210 => x"00",
         18211 => x"00",
         18212 => x"00",
         18213 => x"00",
         18214 => x"00",
         18215 => x"00",
         18216 => x"00",
         18217 => x"00",
         18218 => x"00",
         18219 => x"00",
         18220 => x"00",
         18221 => x"00",
         18222 => x"00",
         18223 => x"00",
         18224 => x"01",
         18225 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"b5",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8e",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8f",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"90",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"91",
           324 => x"0b",
           325 => x"04",
           326 => x"91",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"92",
           336 => x"0b",
           337 => x"04",
           338 => x"92",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"84",
           386 => x"80",
           387 => x"84",
           388 => x"80",
           389 => x"04",
           390 => x"0c",
           391 => x"84",
           392 => x"80",
           393 => x"04",
           394 => x"0c",
           395 => x"84",
           396 => x"80",
           397 => x"04",
           398 => x"0c",
           399 => x"84",
           400 => x"80",
           401 => x"04",
           402 => x"0c",
           403 => x"84",
           404 => x"80",
           405 => x"04",
           406 => x"0c",
           407 => x"84",
           408 => x"80",
           409 => x"04",
           410 => x"0c",
           411 => x"84",
           412 => x"80",
           413 => x"04",
           414 => x"0c",
           415 => x"84",
           416 => x"80",
           417 => x"04",
           418 => x"0c",
           419 => x"84",
           420 => x"80",
           421 => x"04",
           422 => x"0c",
           423 => x"84",
           424 => x"80",
           425 => x"04",
           426 => x"0c",
           427 => x"84",
           428 => x"80",
           429 => x"04",
           430 => x"0c",
           431 => x"84",
           432 => x"80",
           433 => x"04",
           434 => x"0c",
           435 => x"2d",
           436 => x"08",
           437 => x"90",
           438 => x"d4",
           439 => x"d1",
           440 => x"d4",
           441 => x"80",
           442 => x"b9",
           443 => x"d2",
           444 => x"b9",
           445 => x"c0",
           446 => x"84",
           447 => x"80",
           448 => x"84",
           449 => x"80",
           450 => x"04",
           451 => x"0c",
           452 => x"2d",
           453 => x"08",
           454 => x"90",
           455 => x"d4",
           456 => x"80",
           457 => x"d4",
           458 => x"80",
           459 => x"b9",
           460 => x"d2",
           461 => x"b9",
           462 => x"c0",
           463 => x"84",
           464 => x"82",
           465 => x"84",
           466 => x"80",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"90",
           472 => x"d4",
           473 => x"a5",
           474 => x"d4",
           475 => x"80",
           476 => x"b9",
           477 => x"df",
           478 => x"b9",
           479 => x"c0",
           480 => x"84",
           481 => x"82",
           482 => x"84",
           483 => x"80",
           484 => x"04",
           485 => x"0c",
           486 => x"2d",
           487 => x"08",
           488 => x"90",
           489 => x"d4",
           490 => x"e0",
           491 => x"d4",
           492 => x"80",
           493 => x"b9",
           494 => x"84",
           495 => x"b9",
           496 => x"c0",
           497 => x"84",
           498 => x"82",
           499 => x"84",
           500 => x"80",
           501 => x"04",
           502 => x"0c",
           503 => x"2d",
           504 => x"08",
           505 => x"90",
           506 => x"d4",
           507 => x"bd",
           508 => x"d4",
           509 => x"80",
           510 => x"b9",
           511 => x"93",
           512 => x"b9",
           513 => x"c0",
           514 => x"84",
           515 => x"83",
           516 => x"84",
           517 => x"80",
           518 => x"04",
           519 => x"0c",
           520 => x"2d",
           521 => x"08",
           522 => x"90",
           523 => x"d4",
           524 => x"e7",
           525 => x"d4",
           526 => x"80",
           527 => x"b9",
           528 => x"e7",
           529 => x"b9",
           530 => x"c0",
           531 => x"84",
           532 => x"82",
           533 => x"84",
           534 => x"80",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"90",
           540 => x"d4",
           541 => x"f7",
           542 => x"d4",
           543 => x"80",
           544 => x"b9",
           545 => x"a0",
           546 => x"b9",
           547 => x"c0",
           548 => x"84",
           549 => x"82",
           550 => x"84",
           551 => x"80",
           552 => x"04",
           553 => x"0c",
           554 => x"2d",
           555 => x"08",
           556 => x"90",
           557 => x"d4",
           558 => x"93",
           559 => x"d4",
           560 => x"80",
           561 => x"b9",
           562 => x"b7",
           563 => x"b9",
           564 => x"c0",
           565 => x"84",
           566 => x"81",
           567 => x"84",
           568 => x"80",
           569 => x"04",
           570 => x"0c",
           571 => x"2d",
           572 => x"08",
           573 => x"90",
           574 => x"d4",
           575 => x"e1",
           576 => x"d4",
           577 => x"80",
           578 => x"b9",
           579 => x"d0",
           580 => x"b9",
           581 => x"c0",
           582 => x"84",
           583 => x"80",
           584 => x"84",
           585 => x"80",
           586 => x"04",
           587 => x"0c",
           588 => x"2d",
           589 => x"08",
           590 => x"90",
           591 => x"d4",
           592 => x"2d",
           593 => x"08",
           594 => x"90",
           595 => x"d4",
           596 => x"81",
           597 => x"d4",
           598 => x"80",
           599 => x"b9",
           600 => x"dc",
           601 => x"b9",
           602 => x"c0",
           603 => x"84",
           604 => x"81",
           605 => x"84",
           606 => x"80",
           607 => x"04",
           608 => x"0c",
           609 => x"2d",
           610 => x"08",
           611 => x"90",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"51",
           621 => x"73",
           622 => x"73",
           623 => x"81",
           624 => x"10",
           625 => x"07",
           626 => x"0c",
           627 => x"72",
           628 => x"81",
           629 => x"09",
           630 => x"71",
           631 => x"0a",
           632 => x"72",
           633 => x"51",
           634 => x"84",
           635 => x"84",
           636 => x"8e",
           637 => x"70",
           638 => x"0c",
           639 => x"93",
           640 => x"81",
           641 => x"ba",
           642 => x"3d",
           643 => x"70",
           644 => x"52",
           645 => x"74",
           646 => x"ac",
           647 => x"c5",
           648 => x"0d",
           649 => x"0d",
           650 => x"85",
           651 => x"32",
           652 => x"73",
           653 => x"58",
           654 => x"52",
           655 => x"09",
           656 => x"d3",
           657 => x"77",
           658 => x"70",
           659 => x"07",
           660 => x"55",
           661 => x"80",
           662 => x"38",
           663 => x"b2",
           664 => x"8e",
           665 => x"b9",
           666 => x"84",
           667 => x"ff",
           668 => x"84",
           669 => x"75",
           670 => x"57",
           671 => x"73",
           672 => x"30",
           673 => x"9f",
           674 => x"54",
           675 => x"24",
           676 => x"75",
           677 => x"71",
           678 => x"0c",
           679 => x"04",
           680 => x"b9",
           681 => x"3d",
           682 => x"3d",
           683 => x"86",
           684 => x"99",
           685 => x"56",
           686 => x"8e",
           687 => x"53",
           688 => x"3d",
           689 => x"9d",
           690 => x"54",
           691 => x"8d",
           692 => x"fd",
           693 => x"3d",
           694 => x"76",
           695 => x"85",
           696 => x"0d",
           697 => x"0d",
           698 => x"42",
           699 => x"70",
           700 => x"85",
           701 => x"81",
           702 => x"81",
           703 => x"5b",
           704 => x"7b",
           705 => x"06",
           706 => x"7b",
           707 => x"7b",
           708 => x"38",
           709 => x"81",
           710 => x"72",
           711 => x"81",
           712 => x"5f",
           713 => x"81",
           714 => x"b0",
           715 => x"70",
           716 => x"54",
           717 => x"38",
           718 => x"a9",
           719 => x"2a",
           720 => x"81",
           721 => x"7e",
           722 => x"38",
           723 => x"07",
           724 => x"57",
           725 => x"38",
           726 => x"54",
           727 => x"c8",
           728 => x"0d",
           729 => x"2a",
           730 => x"10",
           731 => x"05",
           732 => x"70",
           733 => x"70",
           734 => x"29",
           735 => x"70",
           736 => x"5a",
           737 => x"80",
           738 => x"86",
           739 => x"06",
           740 => x"bd",
           741 => x"33",
           742 => x"fe",
           743 => x"b8",
           744 => x"2e",
           745 => x"93",
           746 => x"74",
           747 => x"8a",
           748 => x"5a",
           749 => x"38",
           750 => x"7c",
           751 => x"8b",
           752 => x"33",
           753 => x"cc",
           754 => x"39",
           755 => x"70",
           756 => x"55",
           757 => x"81",
           758 => x"40",
           759 => x"38",
           760 => x"72",
           761 => x"97",
           762 => x"10",
           763 => x"05",
           764 => x"04",
           765 => x"54",
           766 => x"73",
           767 => x"7c",
           768 => x"8a",
           769 => x"7c",
           770 => x"76",
           771 => x"fe",
           772 => x"ff",
           773 => x"39",
           774 => x"60",
           775 => x"08",
           776 => x"cf",
           777 => x"41",
           778 => x"d8",
           779 => x"75",
           780 => x"3f",
           781 => x"08",
           782 => x"84",
           783 => x"18",
           784 => x"53",
           785 => x"88",
           786 => x"c8",
           787 => x"55",
           788 => x"81",
           789 => x"79",
           790 => x"90",
           791 => x"b9",
           792 => x"84",
           793 => x"c5",
           794 => x"b9",
           795 => x"2b",
           796 => x"40",
           797 => x"2e",
           798 => x"84",
           799 => x"fc",
           800 => x"70",
           801 => x"55",
           802 => x"70",
           803 => x"5f",
           804 => x"9e",
           805 => x"80",
           806 => x"80",
           807 => x"79",
           808 => x"38",
           809 => x"80",
           810 => x"80",
           811 => x"90",
           812 => x"83",
           813 => x"06",
           814 => x"80",
           815 => x"75",
           816 => x"81",
           817 => x"54",
           818 => x"86",
           819 => x"83",
           820 => x"70",
           821 => x"86",
           822 => x"5b",
           823 => x"54",
           824 => x"85",
           825 => x"79",
           826 => x"70",
           827 => x"83",
           828 => x"59",
           829 => x"2e",
           830 => x"7a",
           831 => x"06",
           832 => x"eb",
           833 => x"2a",
           834 => x"73",
           835 => x"7a",
           836 => x"06",
           837 => x"97",
           838 => x"06",
           839 => x"8f",
           840 => x"2a",
           841 => x"7e",
           842 => x"38",
           843 => x"80",
           844 => x"80",
           845 => x"90",
           846 => x"54",
           847 => x"9d",
           848 => x"b0",
           849 => x"3f",
           850 => x"80",
           851 => x"80",
           852 => x"90",
           853 => x"54",
           854 => x"e5",
           855 => x"06",
           856 => x"2e",
           857 => x"79",
           858 => x"29",
           859 => x"05",
           860 => x"5b",
           861 => x"75",
           862 => x"7c",
           863 => x"87",
           864 => x"79",
           865 => x"29",
           866 => x"05",
           867 => x"5b",
           868 => x"80",
           869 => x"7a",
           870 => x"81",
           871 => x"7a",
           872 => x"b9",
           873 => x"e3",
           874 => x"38",
           875 => x"2e",
           876 => x"76",
           877 => x"81",
           878 => x"84",
           879 => x"96",
           880 => x"ff",
           881 => x"52",
           882 => x"3f",
           883 => x"d8",
           884 => x"06",
           885 => x"81",
           886 => x"80",
           887 => x"38",
           888 => x"80",
           889 => x"80",
           890 => x"90",
           891 => x"55",
           892 => x"fc",
           893 => x"52",
           894 => x"f4",
           895 => x"7a",
           896 => x"7a",
           897 => x"33",
           898 => x"fa",
           899 => x"c8",
           900 => x"c0",
           901 => x"f8",
           902 => x"61",
           903 => x"08",
           904 => x"cf",
           905 => x"42",
           906 => x"fd",
           907 => x"84",
           908 => x"80",
           909 => x"13",
           910 => x"2b",
           911 => x"84",
           912 => x"fc",
           913 => x"70",
           914 => x"52",
           915 => x"41",
           916 => x"2a",
           917 => x"5c",
           918 => x"c9",
           919 => x"84",
           920 => x"fc",
           921 => x"70",
           922 => x"54",
           923 => x"25",
           924 => x"7c",
           925 => x"85",
           926 => x"39",
           927 => x"83",
           928 => x"5b",
           929 => x"ff",
           930 => x"ca",
           931 => x"75",
           932 => x"57",
           933 => x"d8",
           934 => x"ff",
           935 => x"ff",
           936 => x"54",
           937 => x"ff",
           938 => x"38",
           939 => x"70",
           940 => x"33",
           941 => x"3f",
           942 => x"fc",
           943 => x"fc",
           944 => x"84",
           945 => x"fc",
           946 => x"70",
           947 => x"58",
           948 => x"7b",
           949 => x"81",
           950 => x"57",
           951 => x"38",
           952 => x"7f",
           953 => x"71",
           954 => x"40",
           955 => x"7e",
           956 => x"38",
           957 => x"bf",
           958 => x"b9",
           959 => x"ad",
           960 => x"07",
           961 => x"5b",
           962 => x"38",
           963 => x"7a",
           964 => x"80",
           965 => x"59",
           966 => x"38",
           967 => x"7f",
           968 => x"71",
           969 => x"06",
           970 => x"5f",
           971 => x"38",
           972 => x"f6",
           973 => x"c8",
           974 => x"ff",
           975 => x"31",
           976 => x"5a",
           977 => x"58",
           978 => x"7a",
           979 => x"7c",
           980 => x"76",
           981 => x"f7",
           982 => x"60",
           983 => x"08",
           984 => x"5d",
           985 => x"79",
           986 => x"75",
           987 => x"3f",
           988 => x"08",
           989 => x"06",
           990 => x"90",
           991 => x"c4",
           992 => x"80",
           993 => x"58",
           994 => x"88",
           995 => x"39",
           996 => x"80",
           997 => x"80",
           998 => x"90",
           999 => x"54",
          1000 => x"fa",
          1001 => x"52",
          1002 => x"c4",
          1003 => x"7c",
          1004 => x"83",
          1005 => x"90",
          1006 => x"06",
          1007 => x"7c",
          1008 => x"83",
          1009 => x"88",
          1010 => x"5f",
          1011 => x"fb",
          1012 => x"d8",
          1013 => x"2c",
          1014 => x"90",
          1015 => x"2c",
          1016 => x"06",
          1017 => x"53",
          1018 => x"38",
          1019 => x"7c",
          1020 => x"82",
          1021 => x"81",
          1022 => x"80",
          1023 => x"38",
          1024 => x"7c",
          1025 => x"2a",
          1026 => x"3f",
          1027 => x"5b",
          1028 => x"f7",
          1029 => x"c8",
          1030 => x"31",
          1031 => x"98",
          1032 => x"f9",
          1033 => x"52",
          1034 => x"c4",
          1035 => x"7c",
          1036 => x"82",
          1037 => x"be",
          1038 => x"75",
          1039 => x"3f",
          1040 => x"08",
          1041 => x"06",
          1042 => x"90",
          1043 => x"fd",
          1044 => x"82",
          1045 => x"71",
          1046 => x"06",
          1047 => x"fd",
          1048 => x"3d",
          1049 => x"a8",
          1050 => x"52",
          1051 => x"b5",
          1052 => x"0d",
          1053 => x"0d",
          1054 => x"0b",
          1055 => x"08",
          1056 => x"70",
          1057 => x"32",
          1058 => x"51",
          1059 => x"57",
          1060 => x"77",
          1061 => x"06",
          1062 => x"74",
          1063 => x"56",
          1064 => x"77",
          1065 => x"84",
          1066 => x"52",
          1067 => x"14",
          1068 => x"2d",
          1069 => x"08",
          1070 => x"38",
          1071 => x"70",
          1072 => x"33",
          1073 => x"2e",
          1074 => x"d5",
          1075 => x"d7",
          1076 => x"ac",
          1077 => x"d5",
          1078 => x"8a",
          1079 => x"08",
          1080 => x"84",
          1081 => x"80",
          1082 => x"ff",
          1083 => x"75",
          1084 => x"0c",
          1085 => x"04",
          1086 => x"78",
          1087 => x"80",
          1088 => x"33",
          1089 => x"81",
          1090 => x"06",
          1091 => x"57",
          1092 => x"77",
          1093 => x"06",
          1094 => x"70",
          1095 => x"33",
          1096 => x"2e",
          1097 => x"98",
          1098 => x"75",
          1099 => x"0c",
          1100 => x"04",
          1101 => x"05",
          1102 => x"72",
          1103 => x"38",
          1104 => x"51",
          1105 => x"53",
          1106 => x"b9",
          1107 => x"2e",
          1108 => x"74",
          1109 => x"56",
          1110 => x"72",
          1111 => x"39",
          1112 => x"84",
          1113 => x"52",
          1114 => x"3f",
          1115 => x"04",
          1116 => x"78",
          1117 => x"33",
          1118 => x"81",
          1119 => x"56",
          1120 => x"ff",
          1121 => x"38",
          1122 => x"81",
          1123 => x"80",
          1124 => x"8c",
          1125 => x"72",
          1126 => x"25",
          1127 => x"08",
          1128 => x"34",
          1129 => x"05",
          1130 => x"15",
          1131 => x"13",
          1132 => x"76",
          1133 => x"b9",
          1134 => x"3d",
          1135 => x"52",
          1136 => x"06",
          1137 => x"08",
          1138 => x"ff",
          1139 => x"c8",
          1140 => x"8c",
          1141 => x"05",
          1142 => x"76",
          1143 => x"fb",
          1144 => x"85",
          1145 => x"81",
          1146 => x"81",
          1147 => x"55",
          1148 => x"ff",
          1149 => x"38",
          1150 => x"81",
          1151 => x"b3",
          1152 => x"2a",
          1153 => x"71",
          1154 => x"c3",
          1155 => x"70",
          1156 => x"71",
          1157 => x"f0",
          1158 => x"76",
          1159 => x"08",
          1160 => x"17",
          1161 => x"ff",
          1162 => x"84",
          1163 => x"87",
          1164 => x"74",
          1165 => x"53",
          1166 => x"34",
          1167 => x"81",
          1168 => x"0c",
          1169 => x"84",
          1170 => x"87",
          1171 => x"75",
          1172 => x"08",
          1173 => x"84",
          1174 => x"52",
          1175 => x"08",
          1176 => x"b9",
          1177 => x"33",
          1178 => x"54",
          1179 => x"c8",
          1180 => x"85",
          1181 => x"07",
          1182 => x"17",
          1183 => x"73",
          1184 => x"0c",
          1185 => x"04",
          1186 => x"53",
          1187 => x"34",
          1188 => x"39",
          1189 => x"75",
          1190 => x"54",
          1191 => x"81",
          1192 => x"51",
          1193 => x"ff",
          1194 => x"70",
          1195 => x"33",
          1196 => x"70",
          1197 => x"34",
          1198 => x"73",
          1199 => x"0c",
          1200 => x"04",
          1201 => x"76",
          1202 => x"55",
          1203 => x"70",
          1204 => x"38",
          1205 => x"a1",
          1206 => x"2e",
          1207 => x"70",
          1208 => x"33",
          1209 => x"05",
          1210 => x"11",
          1211 => x"38",
          1212 => x"c8",
          1213 => x"0d",
          1214 => x"55",
          1215 => x"d9",
          1216 => x"75",
          1217 => x"13",
          1218 => x"53",
          1219 => x"34",
          1220 => x"70",
          1221 => x"38",
          1222 => x"13",
          1223 => x"33",
          1224 => x"11",
          1225 => x"38",
          1226 => x"3d",
          1227 => x"53",
          1228 => x"81",
          1229 => x"51",
          1230 => x"ff",
          1231 => x"31",
          1232 => x"0c",
          1233 => x"0d",
          1234 => x"0d",
          1235 => x"54",
          1236 => x"70",
          1237 => x"33",
          1238 => x"70",
          1239 => x"34",
          1240 => x"73",
          1241 => x"0c",
          1242 => x"04",
          1243 => x"75",
          1244 => x"55",
          1245 => x"70",
          1246 => x"38",
          1247 => x"05",
          1248 => x"70",
          1249 => x"34",
          1250 => x"70",
          1251 => x"84",
          1252 => x"85",
          1253 => x"fc",
          1254 => x"78",
          1255 => x"54",
          1256 => x"a1",
          1257 => x"75",
          1258 => x"57",
          1259 => x"71",
          1260 => x"81",
          1261 => x"81",
          1262 => x"80",
          1263 => x"ff",
          1264 => x"e1",
          1265 => x"70",
          1266 => x"0c",
          1267 => x"04",
          1268 => x"f1",
          1269 => x"53",
          1270 => x"80",
          1271 => x"ff",
          1272 => x"81",
          1273 => x"2e",
          1274 => x"72",
          1275 => x"c8",
          1276 => x"0d",
          1277 => x"b9",
          1278 => x"3d",
          1279 => x"3d",
          1280 => x"53",
          1281 => x"80",
          1282 => x"b9",
          1283 => x"b9",
          1284 => x"05",
          1285 => x"b2",
          1286 => x"b9",
          1287 => x"84",
          1288 => x"80",
          1289 => x"84",
          1290 => x"15",
          1291 => x"34",
          1292 => x"52",
          1293 => x"08",
          1294 => x"3f",
          1295 => x"08",
          1296 => x"b9",
          1297 => x"3d",
          1298 => x"3d",
          1299 => x"71",
          1300 => x"53",
          1301 => x"2e",
          1302 => x"70",
          1303 => x"33",
          1304 => x"2e",
          1305 => x"12",
          1306 => x"2e",
          1307 => x"ea",
          1308 => x"70",
          1309 => x"52",
          1310 => x"c8",
          1311 => x"0d",
          1312 => x"0d",
          1313 => x"72",
          1314 => x"54",
          1315 => x"8e",
          1316 => x"70",
          1317 => x"34",
          1318 => x"70",
          1319 => x"84",
          1320 => x"85",
          1321 => x"fa",
          1322 => x"7a",
          1323 => x"52",
          1324 => x"8b",
          1325 => x"80",
          1326 => x"b9",
          1327 => x"e0",
          1328 => x"80",
          1329 => x"73",
          1330 => x"3f",
          1331 => x"c8",
          1332 => x"80",
          1333 => x"26",
          1334 => x"73",
          1335 => x"2e",
          1336 => x"81",
          1337 => x"2a",
          1338 => x"76",
          1339 => x"54",
          1340 => x"56",
          1341 => x"a8",
          1342 => x"74",
          1343 => x"74",
          1344 => x"78",
          1345 => x"11",
          1346 => x"81",
          1347 => x"06",
          1348 => x"ff",
          1349 => x"52",
          1350 => x"55",
          1351 => x"38",
          1352 => x"07",
          1353 => x"b9",
          1354 => x"3d",
          1355 => x"3d",
          1356 => x"fc",
          1357 => x"70",
          1358 => x"07",
          1359 => x"84",
          1360 => x"31",
          1361 => x"70",
          1362 => x"06",
          1363 => x"80",
          1364 => x"88",
          1365 => x"71",
          1366 => x"f0",
          1367 => x"70",
          1368 => x"2b",
          1369 => x"74",
          1370 => x"53",
          1371 => x"73",
          1372 => x"30",
          1373 => x"10",
          1374 => x"77",
          1375 => x"81",
          1376 => x"70",
          1377 => x"30",
          1378 => x"06",
          1379 => x"84",
          1380 => x"51",
          1381 => x"51",
          1382 => x"53",
          1383 => x"51",
          1384 => x"56",
          1385 => x"54",
          1386 => x"0d",
          1387 => x"0d",
          1388 => x"54",
          1389 => x"54",
          1390 => x"84",
          1391 => x"73",
          1392 => x"31",
          1393 => x"0c",
          1394 => x"0d",
          1395 => x"0d",
          1396 => x"54",
          1397 => x"80",
          1398 => x"76",
          1399 => x"3f",
          1400 => x"08",
          1401 => x"52",
          1402 => x"8d",
          1403 => x"fe",
          1404 => x"84",
          1405 => x"31",
          1406 => x"71",
          1407 => x"c5",
          1408 => x"71",
          1409 => x"38",
          1410 => x"71",
          1411 => x"31",
          1412 => x"57",
          1413 => x"80",
          1414 => x"2e",
          1415 => x"10",
          1416 => x"07",
          1417 => x"07",
          1418 => x"ff",
          1419 => x"70",
          1420 => x"72",
          1421 => x"31",
          1422 => x"56",
          1423 => x"58",
          1424 => x"da",
          1425 => x"b9",
          1426 => x"3d",
          1427 => x"3d",
          1428 => x"2c",
          1429 => x"7a",
          1430 => x"32",
          1431 => x"7d",
          1432 => x"32",
          1433 => x"57",
          1434 => x"56",
          1435 => x"55",
          1436 => x"3f",
          1437 => x"08",
          1438 => x"31",
          1439 => x"0c",
          1440 => x"04",
          1441 => x"7b",
          1442 => x"80",
          1443 => x"77",
          1444 => x"56",
          1445 => x"a0",
          1446 => x"06",
          1447 => x"15",
          1448 => x"70",
          1449 => x"73",
          1450 => x"38",
          1451 => x"80",
          1452 => x"b0",
          1453 => x"38",
          1454 => x"80",
          1455 => x"26",
          1456 => x"8a",
          1457 => x"a0",
          1458 => x"c4",
          1459 => x"74",
          1460 => x"e0",
          1461 => x"ff",
          1462 => x"d0",
          1463 => x"ff",
          1464 => x"90",
          1465 => x"38",
          1466 => x"81",
          1467 => x"54",
          1468 => x"81",
          1469 => x"78",
          1470 => x"38",
          1471 => x"13",
          1472 => x"79",
          1473 => x"56",
          1474 => x"a0",
          1475 => x"38",
          1476 => x"84",
          1477 => x"56",
          1478 => x"81",
          1479 => x"b9",
          1480 => x"3d",
          1481 => x"70",
          1482 => x"0c",
          1483 => x"56",
          1484 => x"2e",
          1485 => x"fe",
          1486 => x"15",
          1487 => x"70",
          1488 => x"73",
          1489 => x"a6",
          1490 => x"73",
          1491 => x"a0",
          1492 => x"a0",
          1493 => x"38",
          1494 => x"80",
          1495 => x"89",
          1496 => x"e1",
          1497 => x"b9",
          1498 => x"3d",
          1499 => x"58",
          1500 => x"78",
          1501 => x"55",
          1502 => x"fe",
          1503 => x"0b",
          1504 => x"0c",
          1505 => x"04",
          1506 => x"7b",
          1507 => x"80",
          1508 => x"77",
          1509 => x"56",
          1510 => x"a0",
          1511 => x"06",
          1512 => x"15",
          1513 => x"70",
          1514 => x"73",
          1515 => x"38",
          1516 => x"80",
          1517 => x"b0",
          1518 => x"38",
          1519 => x"80",
          1520 => x"26",
          1521 => x"8a",
          1522 => x"a0",
          1523 => x"c4",
          1524 => x"74",
          1525 => x"e0",
          1526 => x"ff",
          1527 => x"d0",
          1528 => x"ff",
          1529 => x"90",
          1530 => x"38",
          1531 => x"81",
          1532 => x"54",
          1533 => x"81",
          1534 => x"78",
          1535 => x"38",
          1536 => x"13",
          1537 => x"79",
          1538 => x"56",
          1539 => x"a0",
          1540 => x"38",
          1541 => x"84",
          1542 => x"56",
          1543 => x"81",
          1544 => x"b9",
          1545 => x"3d",
          1546 => x"70",
          1547 => x"0c",
          1548 => x"56",
          1549 => x"2e",
          1550 => x"fe",
          1551 => x"15",
          1552 => x"70",
          1553 => x"73",
          1554 => x"a6",
          1555 => x"73",
          1556 => x"a0",
          1557 => x"a0",
          1558 => x"38",
          1559 => x"80",
          1560 => x"89",
          1561 => x"e1",
          1562 => x"b9",
          1563 => x"3d",
          1564 => x"58",
          1565 => x"78",
          1566 => x"55",
          1567 => x"fe",
          1568 => x"0b",
          1569 => x"0c",
          1570 => x"04",
          1571 => x"3f",
          1572 => x"08",
          1573 => x"84",
          1574 => x"04",
          1575 => x"73",
          1576 => x"26",
          1577 => x"10",
          1578 => x"84",
          1579 => x"08",
          1580 => x"9c",
          1581 => x"3f",
          1582 => x"04",
          1583 => x"51",
          1584 => x"83",
          1585 => x"83",
          1586 => x"ef",
          1587 => x"3d",
          1588 => x"ce",
          1589 => x"9d",
          1590 => x"0d",
          1591 => x"f4",
          1592 => x"3f",
          1593 => x"04",
          1594 => x"51",
          1595 => x"83",
          1596 => x"83",
          1597 => x"ee",
          1598 => x"3d",
          1599 => x"cf",
          1600 => x"f1",
          1601 => x"0d",
          1602 => x"dc",
          1603 => x"3f",
          1604 => x"04",
          1605 => x"51",
          1606 => x"83",
          1607 => x"83",
          1608 => x"ee",
          1609 => x"3d",
          1610 => x"d0",
          1611 => x"c5",
          1612 => x"0d",
          1613 => x"bc",
          1614 => x"3f",
          1615 => x"04",
          1616 => x"51",
          1617 => x"83",
          1618 => x"83",
          1619 => x"ee",
          1620 => x"3d",
          1621 => x"d0",
          1622 => x"99",
          1623 => x"0d",
          1624 => x"88",
          1625 => x"3f",
          1626 => x"04",
          1627 => x"51",
          1628 => x"83",
          1629 => x"83",
          1630 => x"ed",
          1631 => x"3d",
          1632 => x"d1",
          1633 => x"ed",
          1634 => x"0d",
          1635 => x"c4",
          1636 => x"3f",
          1637 => x"04",
          1638 => x"66",
          1639 => x"80",
          1640 => x"5b",
          1641 => x"79",
          1642 => x"07",
          1643 => x"57",
          1644 => x"57",
          1645 => x"26",
          1646 => x"57",
          1647 => x"70",
          1648 => x"51",
          1649 => x"74",
          1650 => x"81",
          1651 => x"8c",
          1652 => x"58",
          1653 => x"3f",
          1654 => x"08",
          1655 => x"c8",
          1656 => x"80",
          1657 => x"51",
          1658 => x"3f",
          1659 => x"78",
          1660 => x"7b",
          1661 => x"2a",
          1662 => x"57",
          1663 => x"80",
          1664 => x"87",
          1665 => x"08",
          1666 => x"e7",
          1667 => x"38",
          1668 => x"87",
          1669 => x"f5",
          1670 => x"b9",
          1671 => x"83",
          1672 => x"78",
          1673 => x"d0",
          1674 => x"3f",
          1675 => x"c8",
          1676 => x"0d",
          1677 => x"c8",
          1678 => x"98",
          1679 => x"b9",
          1680 => x"96",
          1681 => x"54",
          1682 => x"75",
          1683 => x"82",
          1684 => x"84",
          1685 => x"57",
          1686 => x"08",
          1687 => x"7a",
          1688 => x"2e",
          1689 => x"74",
          1690 => x"57",
          1691 => x"87",
          1692 => x"51",
          1693 => x"84",
          1694 => x"52",
          1695 => x"a7",
          1696 => x"c8",
          1697 => x"d1",
          1698 => x"52",
          1699 => x"51",
          1700 => x"ff",
          1701 => x"3d",
          1702 => x"84",
          1703 => x"33",
          1704 => x"58",
          1705 => x"52",
          1706 => x"ec",
          1707 => x"c8",
          1708 => x"76",
          1709 => x"38",
          1710 => x"8a",
          1711 => x"b9",
          1712 => x"3d",
          1713 => x"04",
          1714 => x"56",
          1715 => x"54",
          1716 => x"53",
          1717 => x"51",
          1718 => x"b9",
          1719 => x"b9",
          1720 => x"3d",
          1721 => x"3d",
          1722 => x"63",
          1723 => x"80",
          1724 => x"73",
          1725 => x"41",
          1726 => x"5f",
          1727 => x"80",
          1728 => x"38",
          1729 => x"d1",
          1730 => x"fe",
          1731 => x"84",
          1732 => x"3f",
          1733 => x"79",
          1734 => x"7c",
          1735 => x"ed",
          1736 => x"2e",
          1737 => x"73",
          1738 => x"7a",
          1739 => x"38",
          1740 => x"83",
          1741 => x"dd",
          1742 => x"14",
          1743 => x"08",
          1744 => x"51",
          1745 => x"78",
          1746 => x"38",
          1747 => x"51",
          1748 => x"80",
          1749 => x"27",
          1750 => x"75",
          1751 => x"55",
          1752 => x"72",
          1753 => x"38",
          1754 => x"53",
          1755 => x"83",
          1756 => x"74",
          1757 => x"81",
          1758 => x"57",
          1759 => x"88",
          1760 => x"74",
          1761 => x"38",
          1762 => x"08",
          1763 => x"eb",
          1764 => x"16",
          1765 => x"26",
          1766 => x"d2",
          1767 => x"d5",
          1768 => x"79",
          1769 => x"80",
          1770 => x"3f",
          1771 => x"08",
          1772 => x"98",
          1773 => x"76",
          1774 => x"ee",
          1775 => x"2e",
          1776 => x"7b",
          1777 => x"78",
          1778 => x"38",
          1779 => x"b9",
          1780 => x"3d",
          1781 => x"d2",
          1782 => x"ae",
          1783 => x"84",
          1784 => x"53",
          1785 => x"eb",
          1786 => x"74",
          1787 => x"38",
          1788 => x"83",
          1789 => x"dc",
          1790 => x"14",
          1791 => x"08",
          1792 => x"51",
          1793 => x"73",
          1794 => x"c0",
          1795 => x"53",
          1796 => x"df",
          1797 => x"52",
          1798 => x"51",
          1799 => x"82",
          1800 => x"ac",
          1801 => x"a0",
          1802 => x"3f",
          1803 => x"dd",
          1804 => x"39",
          1805 => x"51",
          1806 => x"84",
          1807 => x"ac",
          1808 => x"a0",
          1809 => x"3f",
          1810 => x"fd",
          1811 => x"18",
          1812 => x"27",
          1813 => x"08",
          1814 => x"fc",
          1815 => x"3f",
          1816 => x"d5",
          1817 => x"54",
          1818 => x"84",
          1819 => x"26",
          1820 => x"d8",
          1821 => x"ac",
          1822 => x"51",
          1823 => x"81",
          1824 => x"91",
          1825 => x"e9",
          1826 => x"c8",
          1827 => x"06",
          1828 => x"72",
          1829 => x"ec",
          1830 => x"72",
          1831 => x"09",
          1832 => x"e0",
          1833 => x"fc",
          1834 => x"51",
          1835 => x"84",
          1836 => x"98",
          1837 => x"2c",
          1838 => x"70",
          1839 => x"32",
          1840 => x"72",
          1841 => x"07",
          1842 => x"58",
          1843 => x"53",
          1844 => x"fd",
          1845 => x"51",
          1846 => x"84",
          1847 => x"98",
          1848 => x"2c",
          1849 => x"70",
          1850 => x"32",
          1851 => x"72",
          1852 => x"07",
          1853 => x"58",
          1854 => x"53",
          1855 => x"ff",
          1856 => x"b9",
          1857 => x"84",
          1858 => x"8f",
          1859 => x"fe",
          1860 => x"c0",
          1861 => x"53",
          1862 => x"81",
          1863 => x"3f",
          1864 => x"51",
          1865 => x"80",
          1866 => x"3f",
          1867 => x"70",
          1868 => x"52",
          1869 => x"38",
          1870 => x"70",
          1871 => x"52",
          1872 => x"38",
          1873 => x"70",
          1874 => x"52",
          1875 => x"38",
          1876 => x"70",
          1877 => x"52",
          1878 => x"38",
          1879 => x"70",
          1880 => x"52",
          1881 => x"38",
          1882 => x"70",
          1883 => x"52",
          1884 => x"38",
          1885 => x"70",
          1886 => x"52",
          1887 => x"72",
          1888 => x"06",
          1889 => x"38",
          1890 => x"84",
          1891 => x"81",
          1892 => x"3f",
          1893 => x"51",
          1894 => x"80",
          1895 => x"3f",
          1896 => x"84",
          1897 => x"81",
          1898 => x"3f",
          1899 => x"51",
          1900 => x"80",
          1901 => x"3f",
          1902 => x"81",
          1903 => x"80",
          1904 => x"cb",
          1905 => x"9b",
          1906 => x"d4",
          1907 => x"ef",
          1908 => x"9b",
          1909 => x"87",
          1910 => x"06",
          1911 => x"80",
          1912 => x"38",
          1913 => x"51",
          1914 => x"83",
          1915 => x"9b",
          1916 => x"51",
          1917 => x"72",
          1918 => x"81",
          1919 => x"71",
          1920 => x"f0",
          1921 => x"39",
          1922 => x"9b",
          1923 => x"a8",
          1924 => x"3f",
          1925 => x"8f",
          1926 => x"2a",
          1927 => x"51",
          1928 => x"2e",
          1929 => x"ff",
          1930 => x"51",
          1931 => x"83",
          1932 => x"9b",
          1933 => x"51",
          1934 => x"72",
          1935 => x"81",
          1936 => x"71",
          1937 => x"94",
          1938 => x"39",
          1939 => x"d7",
          1940 => x"d0",
          1941 => x"3f",
          1942 => x"cb",
          1943 => x"2a",
          1944 => x"51",
          1945 => x"2e",
          1946 => x"ff",
          1947 => x"51",
          1948 => x"83",
          1949 => x"9a",
          1950 => x"51",
          1951 => x"72",
          1952 => x"81",
          1953 => x"71",
          1954 => x"b8",
          1955 => x"39",
          1956 => x"80",
          1957 => x"ff",
          1958 => x"d4",
          1959 => x"52",
          1960 => x"b6",
          1961 => x"b9",
          1962 => x"ff",
          1963 => x"40",
          1964 => x"2e",
          1965 => x"83",
          1966 => x"e3",
          1967 => x"3d",
          1968 => x"ec",
          1969 => x"3f",
          1970 => x"f8",
          1971 => x"7e",
          1972 => x"3f",
          1973 => x"ee",
          1974 => x"81",
          1975 => x"59",
          1976 => x"82",
          1977 => x"81",
          1978 => x"38",
          1979 => x"06",
          1980 => x"2e",
          1981 => x"67",
          1982 => x"79",
          1983 => x"dc",
          1984 => x"5c",
          1985 => x"09",
          1986 => x"38",
          1987 => x"33",
          1988 => x"a0",
          1989 => x"80",
          1990 => x"26",
          1991 => x"90",
          1992 => x"c0",
          1993 => x"52",
          1994 => x"3f",
          1995 => x"08",
          1996 => x"08",
          1997 => x"7b",
          1998 => x"e8",
          1999 => x"b9",
          2000 => x"38",
          2001 => x"5e",
          2002 => x"83",
          2003 => x"1c",
          2004 => x"06",
          2005 => x"7c",
          2006 => x"9a",
          2007 => x"7b",
          2008 => x"dd",
          2009 => x"52",
          2010 => x"92",
          2011 => x"c8",
          2012 => x"b9",
          2013 => x"2e",
          2014 => x"84",
          2015 => x"48",
          2016 => x"80",
          2017 => x"a4",
          2018 => x"c8",
          2019 => x"06",
          2020 => x"80",
          2021 => x"38",
          2022 => x"08",
          2023 => x"3f",
          2024 => x"08",
          2025 => x"f3",
          2026 => x"a5",
          2027 => x"7a",
          2028 => x"85",
          2029 => x"24",
          2030 => x"7a",
          2031 => x"e4",
          2032 => x"80",
          2033 => x"f0",
          2034 => x"d5",
          2035 => x"f2",
          2036 => x"b9",
          2037 => x"56",
          2038 => x"54",
          2039 => x"53",
          2040 => x"52",
          2041 => x"ae",
          2042 => x"c8",
          2043 => x"c8",
          2044 => x"30",
          2045 => x"80",
          2046 => x"5b",
          2047 => x"7a",
          2048 => x"38",
          2049 => x"7a",
          2050 => x"80",
          2051 => x"81",
          2052 => x"ff",
          2053 => x"7a",
          2054 => x"7f",
          2055 => x"81",
          2056 => x"7c",
          2057 => x"61",
          2058 => x"e8",
          2059 => x"81",
          2060 => x"83",
          2061 => x"d3",
          2062 => x"48",
          2063 => x"80",
          2064 => x"e8",
          2065 => x"0b",
          2066 => x"33",
          2067 => x"06",
          2068 => x"fd",
          2069 => x"53",
          2070 => x"52",
          2071 => x"51",
          2072 => x"3f",
          2073 => x"08",
          2074 => x"81",
          2075 => x"83",
          2076 => x"84",
          2077 => x"80",
          2078 => x"51",
          2079 => x"3f",
          2080 => x"08",
          2081 => x"38",
          2082 => x"08",
          2083 => x"3f",
          2084 => x"ee",
          2085 => x"81",
          2086 => x"59",
          2087 => x"09",
          2088 => x"d3",
          2089 => x"84",
          2090 => x"82",
          2091 => x"82",
          2092 => x"83",
          2093 => x"83",
          2094 => x"80",
          2095 => x"51",
          2096 => x"67",
          2097 => x"79",
          2098 => x"90",
          2099 => x"63",
          2100 => x"33",
          2101 => x"89",
          2102 => x"38",
          2103 => x"83",
          2104 => x"5a",
          2105 => x"83",
          2106 => x"f8",
          2107 => x"e4",
          2108 => x"53",
          2109 => x"ba",
          2110 => x"85",
          2111 => x"b9",
          2112 => x"2e",
          2113 => x"fb",
          2114 => x"70",
          2115 => x"41",
          2116 => x"39",
          2117 => x"51",
          2118 => x"7d",
          2119 => x"f3",
          2120 => x"39",
          2121 => x"56",
          2122 => x"d6",
          2123 => x"53",
          2124 => x"52",
          2125 => x"f2",
          2126 => x"39",
          2127 => x"3f",
          2128 => x"9a",
          2129 => x"f9",
          2130 => x"83",
          2131 => x"3f",
          2132 => x"81",
          2133 => x"fa",
          2134 => x"d6",
          2135 => x"95",
          2136 => x"78",
          2137 => x"b8",
          2138 => x"3f",
          2139 => x"fa",
          2140 => x"3d",
          2141 => x"53",
          2142 => x"51",
          2143 => x"84",
          2144 => x"80",
          2145 => x"38",
          2146 => x"d6",
          2147 => x"fa",
          2148 => x"79",
          2149 => x"c8",
          2150 => x"fa",
          2151 => x"b9",
          2152 => x"83",
          2153 => x"d0",
          2154 => x"95",
          2155 => x"ff",
          2156 => x"ff",
          2157 => x"eb",
          2158 => x"b9",
          2159 => x"2e",
          2160 => x"68",
          2161 => x"8c",
          2162 => x"3f",
          2163 => x"04",
          2164 => x"f4",
          2165 => x"80",
          2166 => x"a8",
          2167 => x"c8",
          2168 => x"f9",
          2169 => x"3d",
          2170 => x"53",
          2171 => x"51",
          2172 => x"84",
          2173 => x"86",
          2174 => x"59",
          2175 => x"78",
          2176 => x"a8",
          2177 => x"3f",
          2178 => x"08",
          2179 => x"52",
          2180 => x"91",
          2181 => x"7e",
          2182 => x"ae",
          2183 => x"38",
          2184 => x"87",
          2185 => x"84",
          2186 => x"59",
          2187 => x"3d",
          2188 => x"53",
          2189 => x"51",
          2190 => x"84",
          2191 => x"80",
          2192 => x"38",
          2193 => x"f0",
          2194 => x"80",
          2195 => x"b4",
          2196 => x"c8",
          2197 => x"38",
          2198 => x"22",
          2199 => x"83",
          2200 => x"cf",
          2201 => x"d5",
          2202 => x"80",
          2203 => x"51",
          2204 => x"7e",
          2205 => x"59",
          2206 => x"f8",
          2207 => x"9f",
          2208 => x"38",
          2209 => x"70",
          2210 => x"39",
          2211 => x"84",
          2212 => x"80",
          2213 => x"f0",
          2214 => x"c8",
          2215 => x"f8",
          2216 => x"3d",
          2217 => x"53",
          2218 => x"51",
          2219 => x"84",
          2220 => x"80",
          2221 => x"38",
          2222 => x"f8",
          2223 => x"80",
          2224 => x"c4",
          2225 => x"c8",
          2226 => x"f7",
          2227 => x"d7",
          2228 => x"b6",
          2229 => x"5d",
          2230 => x"27",
          2231 => x"65",
          2232 => x"33",
          2233 => x"7a",
          2234 => x"38",
          2235 => x"54",
          2236 => x"78",
          2237 => x"d4",
          2238 => x"3f",
          2239 => x"5c",
          2240 => x"1b",
          2241 => x"39",
          2242 => x"84",
          2243 => x"80",
          2244 => x"f4",
          2245 => x"c8",
          2246 => x"f7",
          2247 => x"3d",
          2248 => x"53",
          2249 => x"51",
          2250 => x"84",
          2251 => x"80",
          2252 => x"38",
          2253 => x"f8",
          2254 => x"80",
          2255 => x"c8",
          2256 => x"c8",
          2257 => x"f6",
          2258 => x"d7",
          2259 => x"ba",
          2260 => x"79",
          2261 => x"93",
          2262 => x"79",
          2263 => x"5b",
          2264 => x"65",
          2265 => x"eb",
          2266 => x"ff",
          2267 => x"ff",
          2268 => x"e8",
          2269 => x"b9",
          2270 => x"2e",
          2271 => x"b8",
          2272 => x"11",
          2273 => x"05",
          2274 => x"3f",
          2275 => x"08",
          2276 => x"70",
          2277 => x"83",
          2278 => x"cc",
          2279 => x"d5",
          2280 => x"80",
          2281 => x"51",
          2282 => x"7e",
          2283 => x"59",
          2284 => x"f6",
          2285 => x"9f",
          2286 => x"38",
          2287 => x"49",
          2288 => x"59",
          2289 => x"05",
          2290 => x"68",
          2291 => x"b8",
          2292 => x"11",
          2293 => x"05",
          2294 => x"3f",
          2295 => x"08",
          2296 => x"dd",
          2297 => x"02",
          2298 => x"33",
          2299 => x"81",
          2300 => x"3d",
          2301 => x"53",
          2302 => x"51",
          2303 => x"84",
          2304 => x"ff",
          2305 => x"b9",
          2306 => x"ff",
          2307 => x"ff",
          2308 => x"e6",
          2309 => x"b9",
          2310 => x"2e",
          2311 => x"b8",
          2312 => x"11",
          2313 => x"05",
          2314 => x"3f",
          2315 => x"08",
          2316 => x"8d",
          2317 => x"fe",
          2318 => x"ff",
          2319 => x"e6",
          2320 => x"b9",
          2321 => x"38",
          2322 => x"08",
          2323 => x"88",
          2324 => x"3f",
          2325 => x"59",
          2326 => x"8f",
          2327 => x"7a",
          2328 => x"05",
          2329 => x"79",
          2330 => x"8a",
          2331 => x"3f",
          2332 => x"b8",
          2333 => x"05",
          2334 => x"3f",
          2335 => x"08",
          2336 => x"80",
          2337 => x"88",
          2338 => x"53",
          2339 => x"08",
          2340 => x"ea",
          2341 => x"b9",
          2342 => x"2e",
          2343 => x"84",
          2344 => x"51",
          2345 => x"f4",
          2346 => x"3d",
          2347 => x"53",
          2348 => x"51",
          2349 => x"84",
          2350 => x"91",
          2351 => x"cc",
          2352 => x"80",
          2353 => x"38",
          2354 => x"08",
          2355 => x"fe",
          2356 => x"ff",
          2357 => x"e5",
          2358 => x"b9",
          2359 => x"38",
          2360 => x"33",
          2361 => x"2e",
          2362 => x"83",
          2363 => x"47",
          2364 => x"f8",
          2365 => x"80",
          2366 => x"8c",
          2367 => x"c8",
          2368 => x"a5",
          2369 => x"5c",
          2370 => x"2e",
          2371 => x"5c",
          2372 => x"70",
          2373 => x"07",
          2374 => x"06",
          2375 => x"79",
          2376 => x"38",
          2377 => x"83",
          2378 => x"83",
          2379 => x"d6",
          2380 => x"55",
          2381 => x"53",
          2382 => x"51",
          2383 => x"83",
          2384 => x"d6",
          2385 => x"f9",
          2386 => x"71",
          2387 => x"84",
          2388 => x"3d",
          2389 => x"53",
          2390 => x"51",
          2391 => x"84",
          2392 => x"80",
          2393 => x"38",
          2394 => x"0c",
          2395 => x"05",
          2396 => x"fe",
          2397 => x"ff",
          2398 => x"e2",
          2399 => x"b9",
          2400 => x"38",
          2401 => x"64",
          2402 => x"ce",
          2403 => x"70",
          2404 => x"23",
          2405 => x"3d",
          2406 => x"53",
          2407 => x"51",
          2408 => x"84",
          2409 => x"80",
          2410 => x"38",
          2411 => x"80",
          2412 => x"7e",
          2413 => x"40",
          2414 => x"b8",
          2415 => x"11",
          2416 => x"05",
          2417 => x"3f",
          2418 => x"08",
          2419 => x"f1",
          2420 => x"3d",
          2421 => x"53",
          2422 => x"51",
          2423 => x"84",
          2424 => x"80",
          2425 => x"38",
          2426 => x"80",
          2427 => x"7c",
          2428 => x"05",
          2429 => x"39",
          2430 => x"f0",
          2431 => x"80",
          2432 => x"80",
          2433 => x"c8",
          2434 => x"81",
          2435 => x"64",
          2436 => x"64",
          2437 => x"46",
          2438 => x"39",
          2439 => x"09",
          2440 => x"9d",
          2441 => x"83",
          2442 => x"80",
          2443 => x"b0",
          2444 => x"c8",
          2445 => x"96",
          2446 => x"7c",
          2447 => x"3f",
          2448 => x"83",
          2449 => x"d4",
          2450 => x"f5",
          2451 => x"fe",
          2452 => x"ff",
          2453 => x"e0",
          2454 => x"b9",
          2455 => x"2e",
          2456 => x"59",
          2457 => x"05",
          2458 => x"82",
          2459 => x"78",
          2460 => x"39",
          2461 => x"33",
          2462 => x"2e",
          2463 => x"83",
          2464 => x"47",
          2465 => x"83",
          2466 => x"5c",
          2467 => x"a1",
          2468 => x"8c",
          2469 => x"b5",
          2470 => x"e8",
          2471 => x"3f",
          2472 => x"b6",
          2473 => x"e8",
          2474 => x"3f",
          2475 => x"cc",
          2476 => x"ce",
          2477 => x"80",
          2478 => x"83",
          2479 => x"49",
          2480 => x"83",
          2481 => x"d3",
          2482 => x"c6",
          2483 => x"ce",
          2484 => x"80",
          2485 => x"83",
          2486 => x"47",
          2487 => x"83",
          2488 => x"5e",
          2489 => x"9b",
          2490 => x"9c",
          2491 => x"dd",
          2492 => x"cf",
          2493 => x"80",
          2494 => x"83",
          2495 => x"47",
          2496 => x"83",
          2497 => x"5d",
          2498 => x"9b",
          2499 => x"a4",
          2500 => x"b9",
          2501 => x"ca",
          2502 => x"80",
          2503 => x"83",
          2504 => x"47",
          2505 => x"83",
          2506 => x"fc",
          2507 => x"fb",
          2508 => x"f2",
          2509 => x"05",
          2510 => x"39",
          2511 => x"80",
          2512 => x"f8",
          2513 => x"94",
          2514 => x"56",
          2515 => x"80",
          2516 => x"da",
          2517 => x"b9",
          2518 => x"2b",
          2519 => x"55",
          2520 => x"52",
          2521 => x"bf",
          2522 => x"b9",
          2523 => x"77",
          2524 => x"94",
          2525 => x"56",
          2526 => x"80",
          2527 => x"da",
          2528 => x"b9",
          2529 => x"2b",
          2530 => x"55",
          2531 => x"52",
          2532 => x"93",
          2533 => x"b9",
          2534 => x"77",
          2535 => x"83",
          2536 => x"94",
          2537 => x"80",
          2538 => x"c0",
          2539 => x"81",
          2540 => x"81",
          2541 => x"83",
          2542 => x"a1",
          2543 => x"5e",
          2544 => x"0b",
          2545 => x"88",
          2546 => x"72",
          2547 => x"ac",
          2548 => x"85",
          2549 => x"3f",
          2550 => x"ba",
          2551 => x"8c",
          2552 => x"b0",
          2553 => x"b4",
          2554 => x"3f",
          2555 => x"70",
          2556 => x"94",
          2557 => x"d2",
          2558 => x"d2",
          2559 => x"15",
          2560 => x"d2",
          2561 => x"82",
          2562 => x"3f",
          2563 => x"51",
          2564 => x"80",
          2565 => x"f0",
          2566 => x"3f",
          2567 => x"52",
          2568 => x"51",
          2569 => x"ec",
          2570 => x"04",
          2571 => x"77",
          2572 => x"56",
          2573 => x"53",
          2574 => x"81",
          2575 => x"33",
          2576 => x"06",
          2577 => x"a0",
          2578 => x"06",
          2579 => x"15",
          2580 => x"81",
          2581 => x"53",
          2582 => x"2e",
          2583 => x"81",
          2584 => x"73",
          2585 => x"82",
          2586 => x"72",
          2587 => x"e7",
          2588 => x"33",
          2589 => x"06",
          2590 => x"70",
          2591 => x"38",
          2592 => x"80",
          2593 => x"73",
          2594 => x"38",
          2595 => x"e1",
          2596 => x"81",
          2597 => x"54",
          2598 => x"09",
          2599 => x"38",
          2600 => x"a2",
          2601 => x"70",
          2602 => x"07",
          2603 => x"72",
          2604 => x"38",
          2605 => x"81",
          2606 => x"71",
          2607 => x"51",
          2608 => x"c8",
          2609 => x"0d",
          2610 => x"2e",
          2611 => x"80",
          2612 => x"38",
          2613 => x"80",
          2614 => x"81",
          2615 => x"54",
          2616 => x"2e",
          2617 => x"54",
          2618 => x"15",
          2619 => x"53",
          2620 => x"2e",
          2621 => x"fe",
          2622 => x"39",
          2623 => x"76",
          2624 => x"8b",
          2625 => x"84",
          2626 => x"86",
          2627 => x"86",
          2628 => x"52",
          2629 => x"ec",
          2630 => x"c8",
          2631 => x"e5",
          2632 => x"b9",
          2633 => x"3d",
          2634 => x"3d",
          2635 => x"11",
          2636 => x"52",
          2637 => x"70",
          2638 => x"98",
          2639 => x"33",
          2640 => x"82",
          2641 => x"26",
          2642 => x"84",
          2643 => x"83",
          2644 => x"26",
          2645 => x"85",
          2646 => x"84",
          2647 => x"26",
          2648 => x"86",
          2649 => x"85",
          2650 => x"26",
          2651 => x"88",
          2652 => x"86",
          2653 => x"e7",
          2654 => x"38",
          2655 => x"54",
          2656 => x"87",
          2657 => x"cc",
          2658 => x"87",
          2659 => x"0c",
          2660 => x"c0",
          2661 => x"82",
          2662 => x"c0",
          2663 => x"83",
          2664 => x"c0",
          2665 => x"84",
          2666 => x"c0",
          2667 => x"85",
          2668 => x"c0",
          2669 => x"86",
          2670 => x"c0",
          2671 => x"74",
          2672 => x"a4",
          2673 => x"c0",
          2674 => x"80",
          2675 => x"98",
          2676 => x"52",
          2677 => x"c8",
          2678 => x"0d",
          2679 => x"0d",
          2680 => x"c0",
          2681 => x"81",
          2682 => x"c0",
          2683 => x"5e",
          2684 => x"87",
          2685 => x"08",
          2686 => x"1c",
          2687 => x"98",
          2688 => x"79",
          2689 => x"87",
          2690 => x"08",
          2691 => x"1c",
          2692 => x"98",
          2693 => x"79",
          2694 => x"87",
          2695 => x"08",
          2696 => x"1c",
          2697 => x"98",
          2698 => x"7b",
          2699 => x"87",
          2700 => x"08",
          2701 => x"1c",
          2702 => x"0c",
          2703 => x"ff",
          2704 => x"83",
          2705 => x"58",
          2706 => x"57",
          2707 => x"56",
          2708 => x"55",
          2709 => x"54",
          2710 => x"53",
          2711 => x"ff",
          2712 => x"d8",
          2713 => x"bf",
          2714 => x"3d",
          2715 => x"3d",
          2716 => x"05",
          2717 => x"81",
          2718 => x"72",
          2719 => x"a6",
          2720 => x"c8",
          2721 => x"70",
          2722 => x"52",
          2723 => x"09",
          2724 => x"38",
          2725 => x"e3",
          2726 => x"b9",
          2727 => x"3d",
          2728 => x"51",
          2729 => x"3f",
          2730 => x"08",
          2731 => x"98",
          2732 => x"71",
          2733 => x"81",
          2734 => x"72",
          2735 => x"e6",
          2736 => x"c8",
          2737 => x"70",
          2738 => x"52",
          2739 => x"d2",
          2740 => x"fd",
          2741 => x"70",
          2742 => x"88",
          2743 => x"51",
          2744 => x"3f",
          2745 => x"08",
          2746 => x"98",
          2747 => x"71",
          2748 => x"38",
          2749 => x"81",
          2750 => x"83",
          2751 => x"38",
          2752 => x"c8",
          2753 => x"0d",
          2754 => x"0d",
          2755 => x"33",
          2756 => x"33",
          2757 => x"06",
          2758 => x"70",
          2759 => x"f4",
          2760 => x"94",
          2761 => x"96",
          2762 => x"06",
          2763 => x"70",
          2764 => x"38",
          2765 => x"70",
          2766 => x"51",
          2767 => x"72",
          2768 => x"06",
          2769 => x"2e",
          2770 => x"93",
          2771 => x"52",
          2772 => x"73",
          2773 => x"51",
          2774 => x"80",
          2775 => x"2e",
          2776 => x"c0",
          2777 => x"74",
          2778 => x"84",
          2779 => x"86",
          2780 => x"71",
          2781 => x"81",
          2782 => x"70",
          2783 => x"81",
          2784 => x"53",
          2785 => x"cb",
          2786 => x"2a",
          2787 => x"71",
          2788 => x"38",
          2789 => x"84",
          2790 => x"2a",
          2791 => x"53",
          2792 => x"cf",
          2793 => x"ff",
          2794 => x"8f",
          2795 => x"30",
          2796 => x"51",
          2797 => x"83",
          2798 => x"83",
          2799 => x"fa",
          2800 => x"55",
          2801 => x"70",
          2802 => x"70",
          2803 => x"e7",
          2804 => x"83",
          2805 => x"70",
          2806 => x"54",
          2807 => x"80",
          2808 => x"38",
          2809 => x"94",
          2810 => x"2a",
          2811 => x"53",
          2812 => x"80",
          2813 => x"71",
          2814 => x"81",
          2815 => x"70",
          2816 => x"81",
          2817 => x"53",
          2818 => x"8a",
          2819 => x"2a",
          2820 => x"71",
          2821 => x"81",
          2822 => x"87",
          2823 => x"52",
          2824 => x"86",
          2825 => x"94",
          2826 => x"72",
          2827 => x"75",
          2828 => x"73",
          2829 => x"76",
          2830 => x"0c",
          2831 => x"04",
          2832 => x"70",
          2833 => x"51",
          2834 => x"72",
          2835 => x"06",
          2836 => x"2e",
          2837 => x"93",
          2838 => x"52",
          2839 => x"ff",
          2840 => x"c0",
          2841 => x"70",
          2842 => x"81",
          2843 => x"52",
          2844 => x"d7",
          2845 => x"0d",
          2846 => x"80",
          2847 => x"2a",
          2848 => x"52",
          2849 => x"84",
          2850 => x"c0",
          2851 => x"83",
          2852 => x"87",
          2853 => x"08",
          2854 => x"0c",
          2855 => x"94",
          2856 => x"8c",
          2857 => x"9e",
          2858 => x"f2",
          2859 => x"c0",
          2860 => x"83",
          2861 => x"87",
          2862 => x"08",
          2863 => x"0c",
          2864 => x"ac",
          2865 => x"9c",
          2866 => x"9e",
          2867 => x"f2",
          2868 => x"c0",
          2869 => x"83",
          2870 => x"87",
          2871 => x"08",
          2872 => x"0c",
          2873 => x"bc",
          2874 => x"ac",
          2875 => x"9e",
          2876 => x"f2",
          2877 => x"c0",
          2878 => x"83",
          2879 => x"87",
          2880 => x"08",
          2881 => x"f2",
          2882 => x"c0",
          2883 => x"83",
          2884 => x"87",
          2885 => x"08",
          2886 => x"0c",
          2887 => x"8c",
          2888 => x"c4",
          2889 => x"83",
          2890 => x"80",
          2891 => x"9e",
          2892 => x"84",
          2893 => x"51",
          2894 => x"82",
          2895 => x"83",
          2896 => x"80",
          2897 => x"9e",
          2898 => x"88",
          2899 => x"51",
          2900 => x"80",
          2901 => x"81",
          2902 => x"f2",
          2903 => x"0b",
          2904 => x"90",
          2905 => x"80",
          2906 => x"52",
          2907 => x"2e",
          2908 => x"52",
          2909 => x"cb",
          2910 => x"87",
          2911 => x"08",
          2912 => x"80",
          2913 => x"52",
          2914 => x"83",
          2915 => x"71",
          2916 => x"34",
          2917 => x"c0",
          2918 => x"70",
          2919 => x"06",
          2920 => x"70",
          2921 => x"38",
          2922 => x"83",
          2923 => x"80",
          2924 => x"9e",
          2925 => x"90",
          2926 => x"51",
          2927 => x"80",
          2928 => x"81",
          2929 => x"f2",
          2930 => x"0b",
          2931 => x"90",
          2932 => x"80",
          2933 => x"52",
          2934 => x"2e",
          2935 => x"52",
          2936 => x"cf",
          2937 => x"87",
          2938 => x"08",
          2939 => x"80",
          2940 => x"52",
          2941 => x"83",
          2942 => x"71",
          2943 => x"34",
          2944 => x"c0",
          2945 => x"70",
          2946 => x"06",
          2947 => x"70",
          2948 => x"38",
          2949 => x"83",
          2950 => x"80",
          2951 => x"9e",
          2952 => x"80",
          2953 => x"51",
          2954 => x"80",
          2955 => x"81",
          2956 => x"f2",
          2957 => x"0b",
          2958 => x"90",
          2959 => x"80",
          2960 => x"52",
          2961 => x"83",
          2962 => x"71",
          2963 => x"34",
          2964 => x"90",
          2965 => x"06",
          2966 => x"53",
          2967 => x"f2",
          2968 => x"0b",
          2969 => x"90",
          2970 => x"80",
          2971 => x"52",
          2972 => x"83",
          2973 => x"71",
          2974 => x"34",
          2975 => x"90",
          2976 => x"06",
          2977 => x"53",
          2978 => x"f2",
          2979 => x"0b",
          2980 => x"90",
          2981 => x"06",
          2982 => x"70",
          2983 => x"38",
          2984 => x"83",
          2985 => x"87",
          2986 => x"08",
          2987 => x"70",
          2988 => x"34",
          2989 => x"04",
          2990 => x"82",
          2991 => x"0d",
          2992 => x"51",
          2993 => x"3f",
          2994 => x"33",
          2995 => x"9f",
          2996 => x"98",
          2997 => x"3f",
          2998 => x"33",
          2999 => x"ef",
          3000 => x"cf",
          3001 => x"85",
          3002 => x"f2",
          3003 => x"75",
          3004 => x"83",
          3005 => x"55",
          3006 => x"38",
          3007 => x"33",
          3008 => x"cb",
          3009 => x"d3",
          3010 => x"84",
          3011 => x"f2",
          3012 => x"73",
          3013 => x"83",
          3014 => x"55",
          3015 => x"38",
          3016 => x"33",
          3017 => x"c4",
          3018 => x"cb",
          3019 => x"83",
          3020 => x"f2",
          3021 => x"74",
          3022 => x"83",
          3023 => x"56",
          3024 => x"38",
          3025 => x"33",
          3026 => x"e1",
          3027 => x"b0",
          3028 => x"3f",
          3029 => x"08",
          3030 => x"bc",
          3031 => x"aa",
          3032 => x"b0",
          3033 => x"d9",
          3034 => x"b5",
          3035 => x"f2",
          3036 => x"83",
          3037 => x"ff",
          3038 => x"83",
          3039 => x"c1",
          3040 => x"f2",
          3041 => x"83",
          3042 => x"ff",
          3043 => x"83",
          3044 => x"56",
          3045 => x"52",
          3046 => x"8b",
          3047 => x"c8",
          3048 => x"c0",
          3049 => x"31",
          3050 => x"b9",
          3051 => x"83",
          3052 => x"ff",
          3053 => x"83",
          3054 => x"55",
          3055 => x"83",
          3056 => x"55",
          3057 => x"87",
          3058 => x"83",
          3059 => x"56",
          3060 => x"52",
          3061 => x"cf",
          3062 => x"c8",
          3063 => x"c0",
          3064 => x"31",
          3065 => x"b9",
          3066 => x"83",
          3067 => x"ff",
          3068 => x"87",
          3069 => x"83",
          3070 => x"56",
          3071 => x"52",
          3072 => x"a3",
          3073 => x"c8",
          3074 => x"c0",
          3075 => x"31",
          3076 => x"b9",
          3077 => x"83",
          3078 => x"ff",
          3079 => x"83",
          3080 => x"55",
          3081 => x"ff",
          3082 => x"9f",
          3083 => x"e8",
          3084 => x"3f",
          3085 => x"51",
          3086 => x"83",
          3087 => x"52",
          3088 => x"51",
          3089 => x"3f",
          3090 => x"08",
          3091 => x"e4",
          3092 => x"b6",
          3093 => x"b4",
          3094 => x"da",
          3095 => x"b3",
          3096 => x"da",
          3097 => x"8d",
          3098 => x"b8",
          3099 => x"da",
          3100 => x"b3",
          3101 => x"f2",
          3102 => x"bd",
          3103 => x"75",
          3104 => x"3f",
          3105 => x"08",
          3106 => x"29",
          3107 => x"54",
          3108 => x"c8",
          3109 => x"da",
          3110 => x"b2",
          3111 => x"f2",
          3112 => x"74",
          3113 => x"97",
          3114 => x"39",
          3115 => x"51",
          3116 => x"3f",
          3117 => x"33",
          3118 => x"2e",
          3119 => x"fe",
          3120 => x"db",
          3121 => x"bf",
          3122 => x"f2",
          3123 => x"75",
          3124 => x"f0",
          3125 => x"83",
          3126 => x"ff",
          3127 => x"83",
          3128 => x"55",
          3129 => x"fc",
          3130 => x"39",
          3131 => x"51",
          3132 => x"3f",
          3133 => x"33",
          3134 => x"2e",
          3135 => x"d7",
          3136 => x"d6",
          3137 => x"dc",
          3138 => x"b1",
          3139 => x"f2",
          3140 => x"75",
          3141 => x"91",
          3142 => x"83",
          3143 => x"52",
          3144 => x"51",
          3145 => x"3f",
          3146 => x"33",
          3147 => x"2e",
          3148 => x"cd",
          3149 => x"d4",
          3150 => x"dc",
          3151 => x"b1",
          3152 => x"f2",
          3153 => x"73",
          3154 => x"cb",
          3155 => x"83",
          3156 => x"83",
          3157 => x"11",
          3158 => x"dd",
          3159 => x"b1",
          3160 => x"f2",
          3161 => x"75",
          3162 => x"a2",
          3163 => x"83",
          3164 => x"83",
          3165 => x"11",
          3166 => x"dd",
          3167 => x"b1",
          3168 => x"f2",
          3169 => x"73",
          3170 => x"f9",
          3171 => x"83",
          3172 => x"83",
          3173 => x"11",
          3174 => x"dd",
          3175 => x"b0",
          3176 => x"f2",
          3177 => x"74",
          3178 => x"d0",
          3179 => x"83",
          3180 => x"83",
          3181 => x"11",
          3182 => x"dd",
          3183 => x"b0",
          3184 => x"f2",
          3185 => x"75",
          3186 => x"a7",
          3187 => x"83",
          3188 => x"83",
          3189 => x"11",
          3190 => x"dd",
          3191 => x"b0",
          3192 => x"f2",
          3193 => x"73",
          3194 => x"fe",
          3195 => x"83",
          3196 => x"ff",
          3197 => x"83",
          3198 => x"ff",
          3199 => x"83",
          3200 => x"55",
          3201 => x"f9",
          3202 => x"39",
          3203 => x"02",
          3204 => x"52",
          3205 => x"8c",
          3206 => x"10",
          3207 => x"05",
          3208 => x"04",
          3209 => x"51",
          3210 => x"3f",
          3211 => x"04",
          3212 => x"51",
          3213 => x"3f",
          3214 => x"04",
          3215 => x"51",
          3216 => x"3f",
          3217 => x"04",
          3218 => x"51",
          3219 => x"3f",
          3220 => x"04",
          3221 => x"51",
          3222 => x"3f",
          3223 => x"04",
          3224 => x"51",
          3225 => x"3f",
          3226 => x"04",
          3227 => x"0c",
          3228 => x"87",
          3229 => x"0c",
          3230 => x"dc",
          3231 => x"96",
          3232 => x"d9",
          3233 => x"3d",
          3234 => x"08",
          3235 => x"70",
          3236 => x"52",
          3237 => x"08",
          3238 => x"83",
          3239 => x"c8",
          3240 => x"38",
          3241 => x"ff",
          3242 => x"b4",
          3243 => x"80",
          3244 => x"51",
          3245 => x"3f",
          3246 => x"08",
          3247 => x"38",
          3248 => x"e6",
          3249 => x"c8",
          3250 => x"57",
          3251 => x"84",
          3252 => x"25",
          3253 => x"b9",
          3254 => x"05",
          3255 => x"55",
          3256 => x"74",
          3257 => x"70",
          3258 => x"2a",
          3259 => x"78",
          3260 => x"38",
          3261 => x"38",
          3262 => x"08",
          3263 => x"53",
          3264 => x"9b",
          3265 => x"c8",
          3266 => x"78",
          3267 => x"38",
          3268 => x"c8",
          3269 => x"0d",
          3270 => x"fc",
          3271 => x"ea",
          3272 => x"2e",
          3273 => x"e8",
          3274 => x"79",
          3275 => x"3f",
          3276 => x"bf",
          3277 => x"3d",
          3278 => x"b9",
          3279 => x"34",
          3280 => x"e2",
          3281 => x"ad",
          3282 => x"0b",
          3283 => x"0c",
          3284 => x"04",
          3285 => x"ab",
          3286 => x"3d",
          3287 => x"5d",
          3288 => x"57",
          3289 => x"a0",
          3290 => x"38",
          3291 => x"3d",
          3292 => x"10",
          3293 => x"f3",
          3294 => x"08",
          3295 => x"bf",
          3296 => x"b9",
          3297 => x"79",
          3298 => x"51",
          3299 => x"84",
          3300 => x"90",
          3301 => x"33",
          3302 => x"2e",
          3303 => x"73",
          3304 => x"38",
          3305 => x"81",
          3306 => x"54",
          3307 => x"c2",
          3308 => x"73",
          3309 => x"0c",
          3310 => x"04",
          3311 => x"aa",
          3312 => x"11",
          3313 => x"05",
          3314 => x"3f",
          3315 => x"08",
          3316 => x"38",
          3317 => x"78",
          3318 => x"fd",
          3319 => x"b9",
          3320 => x"ff",
          3321 => x"80",
          3322 => x"81",
          3323 => x"ff",
          3324 => x"82",
          3325 => x"fa",
          3326 => x"39",
          3327 => x"05",
          3328 => x"27",
          3329 => x"81",
          3330 => x"70",
          3331 => x"73",
          3332 => x"81",
          3333 => x"38",
          3334 => x"eb",
          3335 => x"8d",
          3336 => x"fe",
          3337 => x"84",
          3338 => x"53",
          3339 => x"08",
          3340 => x"84",
          3341 => x"b9",
          3342 => x"d0",
          3343 => x"b4",
          3344 => x"f8",
          3345 => x"82",
          3346 => x"84",
          3347 => x"80",
          3348 => x"77",
          3349 => x"d2",
          3350 => x"c8",
          3351 => x"0b",
          3352 => x"08",
          3353 => x"84",
          3354 => x"ff",
          3355 => x"58",
          3356 => x"34",
          3357 => x"52",
          3358 => x"e1",
          3359 => x"ff",
          3360 => x"74",
          3361 => x"81",
          3362 => x"38",
          3363 => x"b9",
          3364 => x"3d",
          3365 => x"3d",
          3366 => x"08",
          3367 => x"b9",
          3368 => x"41",
          3369 => x"b4",
          3370 => x"f3",
          3371 => x"f3",
          3372 => x"5d",
          3373 => x"74",
          3374 => x"33",
          3375 => x"80",
          3376 => x"38",
          3377 => x"91",
          3378 => x"70",
          3379 => x"57",
          3380 => x"38",
          3381 => x"90",
          3382 => x"3d",
          3383 => x"5f",
          3384 => x"8a",
          3385 => x"c8",
          3386 => x"70",
          3387 => x"56",
          3388 => x"ec",
          3389 => x"ff",
          3390 => x"84",
          3391 => x"2b",
          3392 => x"84",
          3393 => x"70",
          3394 => x"97",
          3395 => x"2c",
          3396 => x"10",
          3397 => x"05",
          3398 => x"70",
          3399 => x"5c",
          3400 => x"5b",
          3401 => x"81",
          3402 => x"2e",
          3403 => x"78",
          3404 => x"87",
          3405 => x"80",
          3406 => x"ff",
          3407 => x"98",
          3408 => x"80",
          3409 => x"cb",
          3410 => x"16",
          3411 => x"56",
          3412 => x"83",
          3413 => x"33",
          3414 => x"61",
          3415 => x"83",
          3416 => x"08",
          3417 => x"56",
          3418 => x"2e",
          3419 => x"76",
          3420 => x"38",
          3421 => x"80",
          3422 => x"76",
          3423 => x"99",
          3424 => x"70",
          3425 => x"98",
          3426 => x"80",
          3427 => x"2b",
          3428 => x"71",
          3429 => x"70",
          3430 => x"de",
          3431 => x"5f",
          3432 => x"58",
          3433 => x"7a",
          3434 => x"90",
          3435 => x"d1",
          3436 => x"ac",
          3437 => x"76",
          3438 => x"75",
          3439 => x"29",
          3440 => x"05",
          3441 => x"70",
          3442 => x"59",
          3443 => x"95",
          3444 => x"38",
          3445 => x"70",
          3446 => x"55",
          3447 => x"de",
          3448 => x"42",
          3449 => x"25",
          3450 => x"de",
          3451 => x"18",
          3452 => x"55",
          3453 => x"ff",
          3454 => x"80",
          3455 => x"38",
          3456 => x"81",
          3457 => x"2e",
          3458 => x"fe",
          3459 => x"56",
          3460 => x"80",
          3461 => x"e9",
          3462 => x"d1",
          3463 => x"84",
          3464 => x"79",
          3465 => x"7f",
          3466 => x"74",
          3467 => x"b0",
          3468 => x"10",
          3469 => x"05",
          3470 => x"04",
          3471 => x"15",
          3472 => x"80",
          3473 => x"84",
          3474 => x"84",
          3475 => x"d9",
          3476 => x"8c",
          3477 => x"80",
          3478 => x"38",
          3479 => x"08",
          3480 => x"ff",
          3481 => x"84",
          3482 => x"ff",
          3483 => x"84",
          3484 => x"fc",
          3485 => x"d1",
          3486 => x"81",
          3487 => x"d1",
          3488 => x"57",
          3489 => x"27",
          3490 => x"84",
          3491 => x"52",
          3492 => x"77",
          3493 => x"34",
          3494 => x"33",
          3495 => x"b5",
          3496 => x"bc",
          3497 => x"2e",
          3498 => x"7c",
          3499 => x"f2",
          3500 => x"08",
          3501 => x"8f",
          3502 => x"84",
          3503 => x"75",
          3504 => x"d1",
          3505 => x"d1",
          3506 => x"56",
          3507 => x"b6",
          3508 => x"ac",
          3509 => x"51",
          3510 => x"3f",
          3511 => x"08",
          3512 => x"ff",
          3513 => x"84",
          3514 => x"52",
          3515 => x"b4",
          3516 => x"d1",
          3517 => x"05",
          3518 => x"d1",
          3519 => x"81",
          3520 => x"74",
          3521 => x"51",
          3522 => x"3f",
          3523 => x"8c",
          3524 => x"39",
          3525 => x"83",
          3526 => x"56",
          3527 => x"38",
          3528 => x"83",
          3529 => x"fc",
          3530 => x"55",
          3531 => x"38",
          3532 => x"75",
          3533 => x"a8",
          3534 => x"ff",
          3535 => x"84",
          3536 => x"84",
          3537 => x"84",
          3538 => x"81",
          3539 => x"05",
          3540 => x"7b",
          3541 => x"94",
          3542 => x"88",
          3543 => x"8c",
          3544 => x"74",
          3545 => x"9e",
          3546 => x"ac",
          3547 => x"51",
          3548 => x"3f",
          3549 => x"08",
          3550 => x"ff",
          3551 => x"84",
          3552 => x"52",
          3553 => x"b3",
          3554 => x"d1",
          3555 => x"05",
          3556 => x"d1",
          3557 => x"81",
          3558 => x"c7",
          3559 => x"8c",
          3560 => x"ff",
          3561 => x"88",
          3562 => x"55",
          3563 => x"fa",
          3564 => x"d5",
          3565 => x"81",
          3566 => x"84",
          3567 => x"7b",
          3568 => x"52",
          3569 => x"a8",
          3570 => x"8c",
          3571 => x"ff",
          3572 => x"88",
          3573 => x"55",
          3574 => x"fa",
          3575 => x"d5",
          3576 => x"81",
          3577 => x"84",
          3578 => x"7b",
          3579 => x"52",
          3580 => x"fc",
          3581 => x"8c",
          3582 => x"ff",
          3583 => x"88",
          3584 => x"55",
          3585 => x"ff",
          3586 => x"d4",
          3587 => x"8c",
          3588 => x"88",
          3589 => x"74",
          3590 => x"c4",
          3591 => x"5b",
          3592 => x"88",
          3593 => x"2b",
          3594 => x"7c",
          3595 => x"43",
          3596 => x"76",
          3597 => x"38",
          3598 => x"08",
          3599 => x"ff",
          3600 => x"84",
          3601 => x"70",
          3602 => x"98",
          3603 => x"88",
          3604 => x"57",
          3605 => x"24",
          3606 => x"84",
          3607 => x"52",
          3608 => x"b2",
          3609 => x"81",
          3610 => x"81",
          3611 => x"70",
          3612 => x"d1",
          3613 => x"56",
          3614 => x"24",
          3615 => x"84",
          3616 => x"52",
          3617 => x"b1",
          3618 => x"81",
          3619 => x"81",
          3620 => x"70",
          3621 => x"d1",
          3622 => x"56",
          3623 => x"25",
          3624 => x"f8",
          3625 => x"16",
          3626 => x"33",
          3627 => x"d5",
          3628 => x"77",
          3629 => x"b1",
          3630 => x"81",
          3631 => x"81",
          3632 => x"70",
          3633 => x"d1",
          3634 => x"57",
          3635 => x"25",
          3636 => x"7b",
          3637 => x"18",
          3638 => x"84",
          3639 => x"52",
          3640 => x"ff",
          3641 => x"75",
          3642 => x"29",
          3643 => x"05",
          3644 => x"84",
          3645 => x"5b",
          3646 => x"76",
          3647 => x"38",
          3648 => x"84",
          3649 => x"55",
          3650 => x"f7",
          3651 => x"d5",
          3652 => x"88",
          3653 => x"d8",
          3654 => x"8c",
          3655 => x"57",
          3656 => x"8c",
          3657 => x"ff",
          3658 => x"39",
          3659 => x"33",
          3660 => x"80",
          3661 => x"d5",
          3662 => x"8a",
          3663 => x"b0",
          3664 => x"88",
          3665 => x"f4",
          3666 => x"b9",
          3667 => x"ff",
          3668 => x"89",
          3669 => x"d1",
          3670 => x"76",
          3671 => x"d8",
          3672 => x"b8",
          3673 => x"10",
          3674 => x"05",
          3675 => x"5e",
          3676 => x"a0",
          3677 => x"2b",
          3678 => x"83",
          3679 => x"81",
          3680 => x"57",
          3681 => x"fb",
          3682 => x"c8",
          3683 => x"83",
          3684 => x"70",
          3685 => x"f2",
          3686 => x"08",
          3687 => x"74",
          3688 => x"83",
          3689 => x"56",
          3690 => x"8c",
          3691 => x"b0",
          3692 => x"80",
          3693 => x"38",
          3694 => x"d1",
          3695 => x"0b",
          3696 => x"34",
          3697 => x"c8",
          3698 => x"0d",
          3699 => x"8c",
          3700 => x"80",
          3701 => x"84",
          3702 => x"52",
          3703 => x"af",
          3704 => x"d5",
          3705 => x"a0",
          3706 => x"84",
          3707 => x"ac",
          3708 => x"51",
          3709 => x"3f",
          3710 => x"33",
          3711 => x"75",
          3712 => x"34",
          3713 => x"06",
          3714 => x"38",
          3715 => x"51",
          3716 => x"3f",
          3717 => x"d1",
          3718 => x"0b",
          3719 => x"34",
          3720 => x"83",
          3721 => x"0b",
          3722 => x"84",
          3723 => x"55",
          3724 => x"b6",
          3725 => x"ac",
          3726 => x"51",
          3727 => x"3f",
          3728 => x"08",
          3729 => x"ff",
          3730 => x"84",
          3731 => x"52",
          3732 => x"ae",
          3733 => x"d1",
          3734 => x"05",
          3735 => x"d1",
          3736 => x"81",
          3737 => x"74",
          3738 => x"d1",
          3739 => x"9f",
          3740 => x"0b",
          3741 => x"34",
          3742 => x"d1",
          3743 => x"84",
          3744 => x"b4",
          3745 => x"84",
          3746 => x"70",
          3747 => x"5c",
          3748 => x"2e",
          3749 => x"84",
          3750 => x"ff",
          3751 => x"84",
          3752 => x"ff",
          3753 => x"84",
          3754 => x"84",
          3755 => x"52",
          3756 => x"ad",
          3757 => x"d1",
          3758 => x"98",
          3759 => x"2c",
          3760 => x"33",
          3761 => x"56",
          3762 => x"80",
          3763 => x"d5",
          3764 => x"a0",
          3765 => x"98",
          3766 => x"8c",
          3767 => x"2b",
          3768 => x"84",
          3769 => x"5d",
          3770 => x"74",
          3771 => x"f0",
          3772 => x"ac",
          3773 => x"51",
          3774 => x"3f",
          3775 => x"0a",
          3776 => x"0a",
          3777 => x"2c",
          3778 => x"33",
          3779 => x"74",
          3780 => x"cc",
          3781 => x"ac",
          3782 => x"51",
          3783 => x"3f",
          3784 => x"0a",
          3785 => x"0a",
          3786 => x"2c",
          3787 => x"33",
          3788 => x"78",
          3789 => x"b9",
          3790 => x"39",
          3791 => x"81",
          3792 => x"34",
          3793 => x"08",
          3794 => x"51",
          3795 => x"3f",
          3796 => x"0a",
          3797 => x"0a",
          3798 => x"2c",
          3799 => x"33",
          3800 => x"75",
          3801 => x"e6",
          3802 => x"57",
          3803 => x"77",
          3804 => x"ac",
          3805 => x"33",
          3806 => x"f4",
          3807 => x"80",
          3808 => x"80",
          3809 => x"98",
          3810 => x"88",
          3811 => x"5b",
          3812 => x"ff",
          3813 => x"b6",
          3814 => x"8c",
          3815 => x"ff",
          3816 => x"76",
          3817 => x"b8",
          3818 => x"88",
          3819 => x"75",
          3820 => x"74",
          3821 => x"98",
          3822 => x"76",
          3823 => x"38",
          3824 => x"7a",
          3825 => x"34",
          3826 => x"0a",
          3827 => x"0a",
          3828 => x"2c",
          3829 => x"33",
          3830 => x"75",
          3831 => x"38",
          3832 => x"74",
          3833 => x"34",
          3834 => x"06",
          3835 => x"b3",
          3836 => x"34",
          3837 => x"33",
          3838 => x"25",
          3839 => x"17",
          3840 => x"d1",
          3841 => x"57",
          3842 => x"33",
          3843 => x"0a",
          3844 => x"0a",
          3845 => x"2c",
          3846 => x"06",
          3847 => x"58",
          3848 => x"81",
          3849 => x"98",
          3850 => x"2c",
          3851 => x"06",
          3852 => x"75",
          3853 => x"a8",
          3854 => x"ac",
          3855 => x"51",
          3856 => x"3f",
          3857 => x"0a",
          3858 => x"0a",
          3859 => x"2c",
          3860 => x"33",
          3861 => x"75",
          3862 => x"84",
          3863 => x"ac",
          3864 => x"51",
          3865 => x"3f",
          3866 => x"0a",
          3867 => x"0a",
          3868 => x"2c",
          3869 => x"33",
          3870 => x"74",
          3871 => x"b9",
          3872 => x"39",
          3873 => x"08",
          3874 => x"2e",
          3875 => x"75",
          3876 => x"96",
          3877 => x"c8",
          3878 => x"88",
          3879 => x"c8",
          3880 => x"06",
          3881 => x"75",
          3882 => x"ff",
          3883 => x"84",
          3884 => x"84",
          3885 => x"56",
          3886 => x"2e",
          3887 => x"84",
          3888 => x"52",
          3889 => x"a9",
          3890 => x"d5",
          3891 => x"a0",
          3892 => x"9c",
          3893 => x"ac",
          3894 => x"51",
          3895 => x"3f",
          3896 => x"33",
          3897 => x"7a",
          3898 => x"34",
          3899 => x"06",
          3900 => x"a8",
          3901 => x"8b",
          3902 => x"c8",
          3903 => x"b4",
          3904 => x"c8",
          3905 => x"38",
          3906 => x"b0",
          3907 => x"ca",
          3908 => x"39",
          3909 => x"08",
          3910 => x"70",
          3911 => x"ff",
          3912 => x"75",
          3913 => x"29",
          3914 => x"05",
          3915 => x"84",
          3916 => x"52",
          3917 => x"76",
          3918 => x"84",
          3919 => x"70",
          3920 => x"98",
          3921 => x"ff",
          3922 => x"5a",
          3923 => x"25",
          3924 => x"fd",
          3925 => x"f3",
          3926 => x"2e",
          3927 => x"83",
          3928 => x"93",
          3929 => x"55",
          3930 => x"ff",
          3931 => x"58",
          3932 => x"25",
          3933 => x"0b",
          3934 => x"34",
          3935 => x"08",
          3936 => x"2e",
          3937 => x"74",
          3938 => x"f6",
          3939 => x"b4",
          3940 => x"d9",
          3941 => x"0b",
          3942 => x"0c",
          3943 => x"3d",
          3944 => x"bc",
          3945 => x"80",
          3946 => x"80",
          3947 => x"16",
          3948 => x"56",
          3949 => x"ff",
          3950 => x"ba",
          3951 => x"ff",
          3952 => x"84",
          3953 => x"84",
          3954 => x"84",
          3955 => x"81",
          3956 => x"05",
          3957 => x"7b",
          3958 => x"90",
          3959 => x"84",
          3960 => x"84",
          3961 => x"57",
          3962 => x"80",
          3963 => x"38",
          3964 => x"08",
          3965 => x"ff",
          3966 => x"84",
          3967 => x"52",
          3968 => x"a6",
          3969 => x"d5",
          3970 => x"88",
          3971 => x"e0",
          3972 => x"8c",
          3973 => x"5a",
          3974 => x"8c",
          3975 => x"ff",
          3976 => x"39",
          3977 => x"80",
          3978 => x"8c",
          3979 => x"84",
          3980 => x"7b",
          3981 => x"0c",
          3982 => x"04",
          3983 => x"a9",
          3984 => x"b9",
          3985 => x"d1",
          3986 => x"b9",
          3987 => x"ff",
          3988 => x"53",
          3989 => x"51",
          3990 => x"3f",
          3991 => x"81",
          3992 => x"d1",
          3993 => x"d1",
          3994 => x"52",
          3995 => x"80",
          3996 => x"38",
          3997 => x"08",
          3998 => x"ff",
          3999 => x"84",
          4000 => x"52",
          4001 => x"a5",
          4002 => x"d5",
          4003 => x"88",
          4004 => x"dc",
          4005 => x"8c",
          4006 => x"57",
          4007 => x"8c",
          4008 => x"ff",
          4009 => x"39",
          4010 => x"a8",
          4011 => x"b9",
          4012 => x"d1",
          4013 => x"b9",
          4014 => x"ff",
          4015 => x"53",
          4016 => x"51",
          4017 => x"3f",
          4018 => x"81",
          4019 => x"d1",
          4020 => x"d1",
          4021 => x"58",
          4022 => x"80",
          4023 => x"38",
          4024 => x"08",
          4025 => x"ff",
          4026 => x"84",
          4027 => x"52",
          4028 => x"a4",
          4029 => x"d5",
          4030 => x"88",
          4031 => x"f0",
          4032 => x"8c",
          4033 => x"41",
          4034 => x"8c",
          4035 => x"ff",
          4036 => x"39",
          4037 => x"d6",
          4038 => x"f3",
          4039 => x"82",
          4040 => x"06",
          4041 => x"05",
          4042 => x"54",
          4043 => x"80",
          4044 => x"84",
          4045 => x"7b",
          4046 => x"b8",
          4047 => x"10",
          4048 => x"05",
          4049 => x"41",
          4050 => x"2e",
          4051 => x"75",
          4052 => x"74",
          4053 => x"94",
          4054 => x"b8",
          4055 => x"70",
          4056 => x"5a",
          4057 => x"27",
          4058 => x"77",
          4059 => x"34",
          4060 => x"b4",
          4061 => x"05",
          4062 => x"7b",
          4063 => x"81",
          4064 => x"83",
          4065 => x"52",
          4066 => x"ba",
          4067 => x"f3",
          4068 => x"81",
          4069 => x"80",
          4070 => x"8c",
          4071 => x"84",
          4072 => x"7b",
          4073 => x"0c",
          4074 => x"04",
          4075 => x"52",
          4076 => x"08",
          4077 => x"f8",
          4078 => x"c8",
          4079 => x"38",
          4080 => x"08",
          4081 => x"5d",
          4082 => x"08",
          4083 => x"52",
          4084 => x"b7",
          4085 => x"b9",
          4086 => x"84",
          4087 => x"7b",
          4088 => x"06",
          4089 => x"84",
          4090 => x"51",
          4091 => x"3f",
          4092 => x"08",
          4093 => x"84",
          4094 => x"25",
          4095 => x"84",
          4096 => x"ff",
          4097 => x"58",
          4098 => x"34",
          4099 => x"06",
          4100 => x"33",
          4101 => x"83",
          4102 => x"70",
          4103 => x"58",
          4104 => x"f2",
          4105 => x"2b",
          4106 => x"83",
          4107 => x"81",
          4108 => x"58",
          4109 => x"cb",
          4110 => x"c8",
          4111 => x"83",
          4112 => x"70",
          4113 => x"f2",
          4114 => x"08",
          4115 => x"74",
          4116 => x"1d",
          4117 => x"06",
          4118 => x"7d",
          4119 => x"80",
          4120 => x"2e",
          4121 => x"fe",
          4122 => x"e8",
          4123 => x"e6",
          4124 => x"79",
          4125 => x"ff",
          4126 => x"83",
          4127 => x"81",
          4128 => x"ff",
          4129 => x"93",
          4130 => x"c8",
          4131 => x"83",
          4132 => x"ff",
          4133 => x"51",
          4134 => x"3f",
          4135 => x"33",
          4136 => x"87",
          4137 => x"f2",
          4138 => x"1b",
          4139 => x"56",
          4140 => x"cf",
          4141 => x"c8",
          4142 => x"83",
          4143 => x"70",
          4144 => x"f2",
          4145 => x"08",
          4146 => x"74",
          4147 => x"82",
          4148 => x"39",
          4149 => x"b8",
          4150 => x"39",
          4151 => x"b8",
          4152 => x"39",
          4153 => x"51",
          4154 => x"3f",
          4155 => x"38",
          4156 => x"f2",
          4157 => x"80",
          4158 => x"02",
          4159 => x"c7",
          4160 => x"53",
          4161 => x"81",
          4162 => x"81",
          4163 => x"38",
          4164 => x"83",
          4165 => x"82",
          4166 => x"38",
          4167 => x"80",
          4168 => x"b0",
          4169 => x"57",
          4170 => x"a0",
          4171 => x"2e",
          4172 => x"83",
          4173 => x"75",
          4174 => x"34",
          4175 => x"f6",
          4176 => x"f4",
          4177 => x"2b",
          4178 => x"07",
          4179 => x"07",
          4180 => x"7f",
          4181 => x"5b",
          4182 => x"94",
          4183 => x"70",
          4184 => x"0c",
          4185 => x"84",
          4186 => x"76",
          4187 => x"38",
          4188 => x"a2",
          4189 => x"f4",
          4190 => x"9a",
          4191 => x"31",
          4192 => x"a0",
          4193 => x"15",
          4194 => x"70",
          4195 => x"34",
          4196 => x"72",
          4197 => x"3d",
          4198 => x"a7",
          4199 => x"83",
          4200 => x"70",
          4201 => x"83",
          4202 => x"71",
          4203 => x"74",
          4204 => x"58",
          4205 => x"a7",
          4206 => x"84",
          4207 => x"70",
          4208 => x"84",
          4209 => x"70",
          4210 => x"83",
          4211 => x"70",
          4212 => x"06",
          4213 => x"5d",
          4214 => x"5e",
          4215 => x"73",
          4216 => x"38",
          4217 => x"75",
          4218 => x"81",
          4219 => x"81",
          4220 => x"81",
          4221 => x"83",
          4222 => x"62",
          4223 => x"70",
          4224 => x"5d",
          4225 => x"5b",
          4226 => x"26",
          4227 => x"f8",
          4228 => x"76",
          4229 => x"7d",
          4230 => x"5f",
          4231 => x"5c",
          4232 => x"fe",
          4233 => x"7d",
          4234 => x"77",
          4235 => x"38",
          4236 => x"81",
          4237 => x"83",
          4238 => x"74",
          4239 => x"56",
          4240 => x"86",
          4241 => x"59",
          4242 => x"80",
          4243 => x"bc",
          4244 => x"ff",
          4245 => x"bb",
          4246 => x"ff",
          4247 => x"f6",
          4248 => x"29",
          4249 => x"57",
          4250 => x"57",
          4251 => x"81",
          4252 => x"81",
          4253 => x"81",
          4254 => x"71",
          4255 => x"54",
          4256 => x"2e",
          4257 => x"80",
          4258 => x"f8",
          4259 => x"83",
          4260 => x"83",
          4261 => x"70",
          4262 => x"90",
          4263 => x"88",
          4264 => x"07",
          4265 => x"56",
          4266 => x"79",
          4267 => x"38",
          4268 => x"72",
          4269 => x"83",
          4270 => x"70",
          4271 => x"70",
          4272 => x"83",
          4273 => x"71",
          4274 => x"86",
          4275 => x"11",
          4276 => x"56",
          4277 => x"a7",
          4278 => x"14",
          4279 => x"33",
          4280 => x"06",
          4281 => x"33",
          4282 => x"06",
          4283 => x"22",
          4284 => x"ff",
          4285 => x"29",
          4286 => x"5a",
          4287 => x"5f",
          4288 => x"79",
          4289 => x"38",
          4290 => x"15",
          4291 => x"19",
          4292 => x"81",
          4293 => x"81",
          4294 => x"71",
          4295 => x"ff",
          4296 => x"81",
          4297 => x"75",
          4298 => x"5b",
          4299 => x"7b",
          4300 => x"38",
          4301 => x"53",
          4302 => x"16",
          4303 => x"5b",
          4304 => x"e2",
          4305 => x"06",
          4306 => x"da",
          4307 => x"39",
          4308 => x"7b",
          4309 => x"9a",
          4310 => x"0d",
          4311 => x"8c",
          4312 => x"73",
          4313 => x"34",
          4314 => x"81",
          4315 => x"8e",
          4316 => x"80",
          4317 => x"ff",
          4318 => x"87",
          4319 => x"56",
          4320 => x"80",
          4321 => x"8e",
          4322 => x"8a",
          4323 => x"74",
          4324 => x"75",
          4325 => x"83",
          4326 => x"3f",
          4327 => x"e0",
          4328 => x"54",
          4329 => x"86",
          4330 => x"73",
          4331 => x"07",
          4332 => x"75",
          4333 => x"70",
          4334 => x"80",
          4335 => x"53",
          4336 => x"86",
          4337 => x"08",
          4338 => x"81",
          4339 => x"72",
          4340 => x"f3",
          4341 => x"81",
          4342 => x"07",
          4343 => x"34",
          4344 => x"84",
          4345 => x"80",
          4346 => x"c8",
          4347 => x"0d",
          4348 => x"bc",
          4349 => x"c8",
          4350 => x"3d",
          4351 => x"05",
          4352 => x"05",
          4353 => x"84",
          4354 => x"5b",
          4355 => x"53",
          4356 => x"82",
          4357 => x"b7",
          4358 => x"f8",
          4359 => x"f8",
          4360 => x"71",
          4361 => x"a7",
          4362 => x"83",
          4363 => x"5f",
          4364 => x"71",
          4365 => x"70",
          4366 => x"06",
          4367 => x"33",
          4368 => x"53",
          4369 => x"83",
          4370 => x"f8",
          4371 => x"05",
          4372 => x"f8",
          4373 => x"f8",
          4374 => x"05",
          4375 => x"06",
          4376 => x"06",
          4377 => x"72",
          4378 => x"8c",
          4379 => x"53",
          4380 => x"f8",
          4381 => x"f6",
          4382 => x"ff",
          4383 => x"b7",
          4384 => x"55",
          4385 => x"26",
          4386 => x"84",
          4387 => x"76",
          4388 => x"58",
          4389 => x"9f",
          4390 => x"38",
          4391 => x"70",
          4392 => x"e0",
          4393 => x"e0",
          4394 => x"72",
          4395 => x"54",
          4396 => x"81",
          4397 => x"81",
          4398 => x"b7",
          4399 => x"e3",
          4400 => x"9f",
          4401 => x"83",
          4402 => x"84",
          4403 => x"54",
          4404 => x"e0",
          4405 => x"74",
          4406 => x"05",
          4407 => x"14",
          4408 => x"74",
          4409 => x"84",
          4410 => x"ff",
          4411 => x"83",
          4412 => x"75",
          4413 => x"ff",
          4414 => x"ff",
          4415 => x"54",
          4416 => x"81",
          4417 => x"74",
          4418 => x"84",
          4419 => x"71",
          4420 => x"55",
          4421 => x"86",
          4422 => x"58",
          4423 => x"80",
          4424 => x"06",
          4425 => x"06",
          4426 => x"19",
          4427 => x"57",
          4428 => x"b9",
          4429 => x"9a",
          4430 => x"e0",
          4431 => x"84",
          4432 => x"33",
          4433 => x"05",
          4434 => x"70",
          4435 => x"33",
          4436 => x"05",
          4437 => x"15",
          4438 => x"33",
          4439 => x"33",
          4440 => x"19",
          4441 => x"55",
          4442 => x"ce",
          4443 => x"72",
          4444 => x"0c",
          4445 => x"04",
          4446 => x"f8",
          4447 => x"f6",
          4448 => x"ff",
          4449 => x"b7",
          4450 => x"55",
          4451 => x"27",
          4452 => x"77",
          4453 => x"dd",
          4454 => x"ff",
          4455 => x"83",
          4456 => x"56",
          4457 => x"2e",
          4458 => x"fe",
          4459 => x"76",
          4460 => x"84",
          4461 => x"71",
          4462 => x"72",
          4463 => x"52",
          4464 => x"73",
          4465 => x"38",
          4466 => x"33",
          4467 => x"15",
          4468 => x"55",
          4469 => x"0b",
          4470 => x"34",
          4471 => x"81",
          4472 => x"ff",
          4473 => x"80",
          4474 => x"38",
          4475 => x"e0",
          4476 => x"75",
          4477 => x"57",
          4478 => x"53",
          4479 => x"fd",
          4480 => x"0b",
          4481 => x"33",
          4482 => x"89",
          4483 => x"fa",
          4484 => x"84",
          4485 => x"33",
          4486 => x"b7",
          4487 => x"fc",
          4488 => x"3d",
          4489 => x"84",
          4490 => x"33",
          4491 => x"86",
          4492 => x"70",
          4493 => x"c3",
          4494 => x"70",
          4495 => x"b7",
          4496 => x"71",
          4497 => x"38",
          4498 => x"f9",
          4499 => x"84",
          4500 => x"86",
          4501 => x"80",
          4502 => x"f9",
          4503 => x"f8",
          4504 => x"ff",
          4505 => x"72",
          4506 => x"38",
          4507 => x"70",
          4508 => x"34",
          4509 => x"b9",
          4510 => x"3d",
          4511 => x"f8",
          4512 => x"73",
          4513 => x"70",
          4514 => x"06",
          4515 => x"54",
          4516 => x"f8",
          4517 => x"83",
          4518 => x"72",
          4519 => x"bb",
          4520 => x"55",
          4521 => x"75",
          4522 => x"70",
          4523 => x"f8",
          4524 => x"0b",
          4525 => x"0c",
          4526 => x"04",
          4527 => x"33",
          4528 => x"70",
          4529 => x"2c",
          4530 => x"56",
          4531 => x"83",
          4532 => x"80",
          4533 => x"c8",
          4534 => x"0d",
          4535 => x"f9",
          4536 => x"84",
          4537 => x"ff",
          4538 => x"51",
          4539 => x"83",
          4540 => x"72",
          4541 => x"34",
          4542 => x"b9",
          4543 => x"3d",
          4544 => x"0b",
          4545 => x"34",
          4546 => x"33",
          4547 => x"33",
          4548 => x"52",
          4549 => x"fe",
          4550 => x"12",
          4551 => x"f8",
          4552 => x"d0",
          4553 => x"0d",
          4554 => x"33",
          4555 => x"26",
          4556 => x"10",
          4557 => x"88",
          4558 => x"08",
          4559 => x"f4",
          4560 => x"f0",
          4561 => x"2b",
          4562 => x"70",
          4563 => x"07",
          4564 => x"51",
          4565 => x"2e",
          4566 => x"9c",
          4567 => x"0b",
          4568 => x"34",
          4569 => x"b9",
          4570 => x"3d",
          4571 => x"f8",
          4572 => x"9f",
          4573 => x"51",
          4574 => x"f4",
          4575 => x"84",
          4576 => x"83",
          4577 => x"83",
          4578 => x"80",
          4579 => x"70",
          4580 => x"34",
          4581 => x"f8",
          4582 => x"fe",
          4583 => x"51",
          4584 => x"f4",
          4585 => x"80",
          4586 => x"f8",
          4587 => x"0b",
          4588 => x"0c",
          4589 => x"04",
          4590 => x"33",
          4591 => x"84",
          4592 => x"83",
          4593 => x"ff",
          4594 => x"f8",
          4595 => x"07",
          4596 => x"f8",
          4597 => x"a5",
          4598 => x"f4",
          4599 => x"06",
          4600 => x"70",
          4601 => x"34",
          4602 => x"83",
          4603 => x"81",
          4604 => x"07",
          4605 => x"f8",
          4606 => x"81",
          4607 => x"f4",
          4608 => x"06",
          4609 => x"70",
          4610 => x"34",
          4611 => x"83",
          4612 => x"81",
          4613 => x"70",
          4614 => x"34",
          4615 => x"83",
          4616 => x"81",
          4617 => x"d0",
          4618 => x"83",
          4619 => x"fe",
          4620 => x"f8",
          4621 => x"bf",
          4622 => x"51",
          4623 => x"f4",
          4624 => x"39",
          4625 => x"33",
          4626 => x"80",
          4627 => x"70",
          4628 => x"34",
          4629 => x"83",
          4630 => x"81",
          4631 => x"c0",
          4632 => x"83",
          4633 => x"fe",
          4634 => x"f8",
          4635 => x"af",
          4636 => x"51",
          4637 => x"f4",
          4638 => x"39",
          4639 => x"33",
          4640 => x"51",
          4641 => x"f4",
          4642 => x"39",
          4643 => x"33",
          4644 => x"82",
          4645 => x"83",
          4646 => x"fd",
          4647 => x"3d",
          4648 => x"05",
          4649 => x"05",
          4650 => x"33",
          4651 => x"33",
          4652 => x"33",
          4653 => x"33",
          4654 => x"33",
          4655 => x"5d",
          4656 => x"82",
          4657 => x"38",
          4658 => x"a5",
          4659 => x"2e",
          4660 => x"7d",
          4661 => x"34",
          4662 => x"b7",
          4663 => x"83",
          4664 => x"7b",
          4665 => x"23",
          4666 => x"f9",
          4667 => x"0d",
          4668 => x"2e",
          4669 => x"db",
          4670 => x"84",
          4671 => x"81",
          4672 => x"c0",
          4673 => x"83",
          4674 => x"a8",
          4675 => x"f9",
          4676 => x"83",
          4677 => x"79",
          4678 => x"bc",
          4679 => x"b7",
          4680 => x"84",
          4681 => x"55",
          4682 => x"53",
          4683 => x"e3",
          4684 => x"81",
          4685 => x"84",
          4686 => x"80",
          4687 => x"c0",
          4688 => x"f8",
          4689 => x"83",
          4690 => x"7c",
          4691 => x"34",
          4692 => x"04",
          4693 => x"b7",
          4694 => x"0b",
          4695 => x"34",
          4696 => x"f8",
          4697 => x"0b",
          4698 => x"34",
          4699 => x"f8",
          4700 => x"b8",
          4701 => x"84",
          4702 => x"57",
          4703 => x"33",
          4704 => x"7b",
          4705 => x"7a",
          4706 => x"d8",
          4707 => x"fa",
          4708 => x"84",
          4709 => x"5a",
          4710 => x"27",
          4711 => x"10",
          4712 => x"05",
          4713 => x"59",
          4714 => x"51",
          4715 => x"3f",
          4716 => x"81",
          4717 => x"b8",
          4718 => x"5b",
          4719 => x"26",
          4720 => x"d2",
          4721 => x"80",
          4722 => x"84",
          4723 => x"80",
          4724 => x"c0",
          4725 => x"f8",
          4726 => x"83",
          4727 => x"7c",
          4728 => x"34",
          4729 => x"04",
          4730 => x"b7",
          4731 => x"0b",
          4732 => x"34",
          4733 => x"f8",
          4734 => x"0b",
          4735 => x"34",
          4736 => x"f8",
          4737 => x"f7",
          4738 => x"92",
          4739 => x"b9",
          4740 => x"83",
          4741 => x"fe",
          4742 => x"80",
          4743 => x"ac",
          4744 => x"86",
          4745 => x"b9",
          4746 => x"fd",
          4747 => x"f7",
          4748 => x"52",
          4749 => x"51",
          4750 => x"3f",
          4751 => x"81",
          4752 => x"5a",
          4753 => x"3d",
          4754 => x"84",
          4755 => x"33",
          4756 => x"33",
          4757 => x"33",
          4758 => x"33",
          4759 => x"12",
          4760 => x"80",
          4761 => x"f6",
          4762 => x"59",
          4763 => x"29",
          4764 => x"ff",
          4765 => x"f7",
          4766 => x"59",
          4767 => x"57",
          4768 => x"81",
          4769 => x"89",
          4770 => x"38",
          4771 => x"81",
          4772 => x"81",
          4773 => x"38",
          4774 => x"82",
          4775 => x"b7",
          4776 => x"f8",
          4777 => x"f8",
          4778 => x"72",
          4779 => x"56",
          4780 => x"c4",
          4781 => x"a7",
          4782 => x"34",
          4783 => x"33",
          4784 => x"33",
          4785 => x"22",
          4786 => x"12",
          4787 => x"53",
          4788 => x"fa",
          4789 => x"f8",
          4790 => x"71",
          4791 => x"54",
          4792 => x"33",
          4793 => x"80",
          4794 => x"b7",
          4795 => x"81",
          4796 => x"f8",
          4797 => x"f8",
          4798 => x"72",
          4799 => x"5b",
          4800 => x"83",
          4801 => x"84",
          4802 => x"34",
          4803 => x"81",
          4804 => x"55",
          4805 => x"81",
          4806 => x"b7",
          4807 => x"77",
          4808 => x"ff",
          4809 => x"83",
          4810 => x"84",
          4811 => x"53",
          4812 => x"8c",
          4813 => x"c0",
          4814 => x"80",
          4815 => x"38",
          4816 => x"b9",
          4817 => x"3d",
          4818 => x"8d",
          4819 => x"75",
          4820 => x"f7",
          4821 => x"2e",
          4822 => x"fe",
          4823 => x"52",
          4824 => x"96",
          4825 => x"83",
          4826 => x"ff",
          4827 => x"f8",
          4828 => x"53",
          4829 => x"13",
          4830 => x"75",
          4831 => x"81",
          4832 => x"38",
          4833 => x"52",
          4834 => x"ba",
          4835 => x"70",
          4836 => x"54",
          4837 => x"26",
          4838 => x"76",
          4839 => x"fd",
          4840 => x"13",
          4841 => x"06",
          4842 => x"73",
          4843 => x"fe",
          4844 => x"83",
          4845 => x"fe",
          4846 => x"52",
          4847 => x"de",
          4848 => x"84",
          4849 => x"89",
          4850 => x"75",
          4851 => x"09",
          4852 => x"ca",
          4853 => x"f9",
          4854 => x"ff",
          4855 => x"05",
          4856 => x"38",
          4857 => x"83",
          4858 => x"76",
          4859 => x"fc",
          4860 => x"f8",
          4861 => x"81",
          4862 => x"ff",
          4863 => x"fe",
          4864 => x"53",
          4865 => x"f9",
          4866 => x"39",
          4867 => x"f8",
          4868 => x"52",
          4869 => x"e2",
          4870 => x"39",
          4871 => x"51",
          4872 => x"fe",
          4873 => x"3d",
          4874 => x"f3",
          4875 => x"b8",
          4876 => x"59",
          4877 => x"81",
          4878 => x"82",
          4879 => x"38",
          4880 => x"84",
          4881 => x"8a",
          4882 => x"38",
          4883 => x"84",
          4884 => x"89",
          4885 => x"38",
          4886 => x"33",
          4887 => x"33",
          4888 => x"33",
          4889 => x"05",
          4890 => x"84",
          4891 => x"33",
          4892 => x"80",
          4893 => x"b7",
          4894 => x"f8",
          4895 => x"f8",
          4896 => x"71",
          4897 => x"5a",
          4898 => x"83",
          4899 => x"34",
          4900 => x"33",
          4901 => x"62",
          4902 => x"83",
          4903 => x"7f",
          4904 => x"80",
          4905 => x"b7",
          4906 => x"81",
          4907 => x"f8",
          4908 => x"f8",
          4909 => x"72",
          4910 => x"40",
          4911 => x"83",
          4912 => x"84",
          4913 => x"34",
          4914 => x"81",
          4915 => x"58",
          4916 => x"81",
          4917 => x"b7",
          4918 => x"79",
          4919 => x"ff",
          4920 => x"83",
          4921 => x"80",
          4922 => x"c8",
          4923 => x"0d",
          4924 => x"2e",
          4925 => x"b7",
          4926 => x"fd",
          4927 => x"2e",
          4928 => x"78",
          4929 => x"89",
          4930 => x"0b",
          4931 => x"0c",
          4932 => x"33",
          4933 => x"33",
          4934 => x"33",
          4935 => x"05",
          4936 => x"84",
          4937 => x"33",
          4938 => x"80",
          4939 => x"b7",
          4940 => x"f8",
          4941 => x"f8",
          4942 => x"71",
          4943 => x"5f",
          4944 => x"83",
          4945 => x"34",
          4946 => x"33",
          4947 => x"19",
          4948 => x"f8",
          4949 => x"a7",
          4950 => x"34",
          4951 => x"33",
          4952 => x"06",
          4953 => x"22",
          4954 => x"33",
          4955 => x"11",
          4956 => x"58",
          4957 => x"f4",
          4958 => x"98",
          4959 => x"81",
          4960 => x"81",
          4961 => x"60",
          4962 => x"ca",
          4963 => x"f8",
          4964 => x"0b",
          4965 => x"0c",
          4966 => x"04",
          4967 => x"82",
          4968 => x"9b",
          4969 => x"38",
          4970 => x"09",
          4971 => x"a8",
          4972 => x"83",
          4973 => x"80",
          4974 => x"c8",
          4975 => x"0d",
          4976 => x"2e",
          4977 => x"d0",
          4978 => x"89",
          4979 => x"38",
          4980 => x"33",
          4981 => x"57",
          4982 => x"c8",
          4983 => x"b8",
          4984 => x"77",
          4985 => x"59",
          4986 => x"b8",
          4987 => x"80",
          4988 => x"c8",
          4989 => x"0d",
          4990 => x"2e",
          4991 => x"80",
          4992 => x"c4",
          4993 => x"bc",
          4994 => x"f8",
          4995 => x"f9",
          4996 => x"29",
          4997 => x"40",
          4998 => x"19",
          4999 => x"a0",
          5000 => x"84",
          5001 => x"83",
          5002 => x"83",
          5003 => x"72",
          5004 => x"41",
          5005 => x"78",
          5006 => x"1f",
          5007 => x"f8",
          5008 => x"29",
          5009 => x"83",
          5010 => x"86",
          5011 => x"1b",
          5012 => x"bc",
          5013 => x"ff",
          5014 => x"f6",
          5015 => x"f9",
          5016 => x"29",
          5017 => x"43",
          5018 => x"f8",
          5019 => x"84",
          5020 => x"34",
          5021 => x"fe",
          5022 => x"52",
          5023 => x"fa",
          5024 => x"83",
          5025 => x"fe",
          5026 => x"b7",
          5027 => x"f8",
          5028 => x"81",
          5029 => x"f8",
          5030 => x"71",
          5031 => x"a7",
          5032 => x"83",
          5033 => x"40",
          5034 => x"7e",
          5035 => x"83",
          5036 => x"83",
          5037 => x"5a",
          5038 => x"5c",
          5039 => x"86",
          5040 => x"81",
          5041 => x"1a",
          5042 => x"fc",
          5043 => x"56",
          5044 => x"f9",
          5045 => x"39",
          5046 => x"b8",
          5047 => x"0b",
          5048 => x"34",
          5049 => x"b8",
          5050 => x"0b",
          5051 => x"34",
          5052 => x"b8",
          5053 => x"0b",
          5054 => x"0c",
          5055 => x"04",
          5056 => x"33",
          5057 => x"34",
          5058 => x"33",
          5059 => x"34",
          5060 => x"33",
          5061 => x"34",
          5062 => x"b8",
          5063 => x"0b",
          5064 => x"0c",
          5065 => x"04",
          5066 => x"2e",
          5067 => x"fa",
          5068 => x"f8",
          5069 => x"b7",
          5070 => x"81",
          5071 => x"f8",
          5072 => x"81",
          5073 => x"75",
          5074 => x"a7",
          5075 => x"83",
          5076 => x"5c",
          5077 => x"29",
          5078 => x"ff",
          5079 => x"f7",
          5080 => x"5c",
          5081 => x"5b",
          5082 => x"2e",
          5083 => x"78",
          5084 => x"ff",
          5085 => x"75",
          5086 => x"57",
          5087 => x"f9",
          5088 => x"ff",
          5089 => x"ff",
          5090 => x"ff",
          5091 => x"29",
          5092 => x"5b",
          5093 => x"33",
          5094 => x"80",
          5095 => x"b7",
          5096 => x"f8",
          5097 => x"f8",
          5098 => x"71",
          5099 => x"5e",
          5100 => x"0b",
          5101 => x"18",
          5102 => x"f8",
          5103 => x"29",
          5104 => x"56",
          5105 => x"33",
          5106 => x"80",
          5107 => x"b7",
          5108 => x"81",
          5109 => x"f8",
          5110 => x"f8",
          5111 => x"72",
          5112 => x"5d",
          5113 => x"83",
          5114 => x"7f",
          5115 => x"05",
          5116 => x"70",
          5117 => x"5c",
          5118 => x"26",
          5119 => x"84",
          5120 => x"5a",
          5121 => x"38",
          5122 => x"77",
          5123 => x"34",
          5124 => x"33",
          5125 => x"06",
          5126 => x"56",
          5127 => x"78",
          5128 => x"d8",
          5129 => x"2e",
          5130 => x"78",
          5131 => x"a8",
          5132 => x"c8",
          5133 => x"83",
          5134 => x"bf",
          5135 => x"b4",
          5136 => x"38",
          5137 => x"83",
          5138 => x"58",
          5139 => x"80",
          5140 => x"f9",
          5141 => x"81",
          5142 => x"3f",
          5143 => x"b9",
          5144 => x"3d",
          5145 => x"f8",
          5146 => x"b7",
          5147 => x"81",
          5148 => x"f8",
          5149 => x"81",
          5150 => x"75",
          5151 => x"a7",
          5152 => x"83",
          5153 => x"5c",
          5154 => x"29",
          5155 => x"ff",
          5156 => x"f7",
          5157 => x"53",
          5158 => x"5b",
          5159 => x"2e",
          5160 => x"80",
          5161 => x"ff",
          5162 => x"ff",
          5163 => x"ff",
          5164 => x"29",
          5165 => x"40",
          5166 => x"33",
          5167 => x"80",
          5168 => x"b7",
          5169 => x"f8",
          5170 => x"f8",
          5171 => x"71",
          5172 => x"41",
          5173 => x"0b",
          5174 => x"1c",
          5175 => x"f8",
          5176 => x"29",
          5177 => x"83",
          5178 => x"86",
          5179 => x"1a",
          5180 => x"bc",
          5181 => x"ff",
          5182 => x"f6",
          5183 => x"f9",
          5184 => x"29",
          5185 => x"5a",
          5186 => x"f8",
          5187 => x"98",
          5188 => x"60",
          5189 => x"81",
          5190 => x"58",
          5191 => x"81",
          5192 => x"b7",
          5193 => x"77",
          5194 => x"ff",
          5195 => x"83",
          5196 => x"81",
          5197 => x"ff",
          5198 => x"7b",
          5199 => x"a7",
          5200 => x"f8",
          5201 => x"bc",
          5202 => x"f9",
          5203 => x"ff",
          5204 => x"ff",
          5205 => x"ff",
          5206 => x"29",
          5207 => x"43",
          5208 => x"84",
          5209 => x"86",
          5210 => x"1b",
          5211 => x"bc",
          5212 => x"f9",
          5213 => x"f6",
          5214 => x"29",
          5215 => x"5e",
          5216 => x"83",
          5217 => x"34",
          5218 => x"33",
          5219 => x"1e",
          5220 => x"f8",
          5221 => x"a7",
          5222 => x"34",
          5223 => x"33",
          5224 => x"06",
          5225 => x"22",
          5226 => x"33",
          5227 => x"11",
          5228 => x"40",
          5229 => x"f4",
          5230 => x"9a",
          5231 => x"81",
          5232 => x"ff",
          5233 => x"79",
          5234 => x"d6",
          5235 => x"f8",
          5236 => x"df",
          5237 => x"84",
          5238 => x"80",
          5239 => x"c8",
          5240 => x"0d",
          5241 => x"fa",
          5242 => x"84",
          5243 => x"33",
          5244 => x"f8",
          5245 => x"81",
          5246 => x"ff",
          5247 => x"ca",
          5248 => x"84",
          5249 => x"80",
          5250 => x"c8",
          5251 => x"0d",
          5252 => x"fa",
          5253 => x"84",
          5254 => x"33",
          5255 => x"f8",
          5256 => x"b7",
          5257 => x"f8",
          5258 => x"5b",
          5259 => x"fc",
          5260 => x"b8",
          5261 => x"3d",
          5262 => x"d8",
          5263 => x"8a",
          5264 => x"b9",
          5265 => x"2e",
          5266 => x"84",
          5267 => x"81",
          5268 => x"75",
          5269 => x"34",
          5270 => x"fe",
          5271 => x"80",
          5272 => x"61",
          5273 => x"05",
          5274 => x"39",
          5275 => x"17",
          5276 => x"b7",
          5277 => x"7b",
          5278 => x"f8",
          5279 => x"bc",
          5280 => x"f9",
          5281 => x"5c",
          5282 => x"84",
          5283 => x"83",
          5284 => x"83",
          5285 => x"72",
          5286 => x"41",
          5287 => x"b7",
          5288 => x"7f",
          5289 => x"80",
          5290 => x"b7",
          5291 => x"f8",
          5292 => x"f8",
          5293 => x"71",
          5294 => x"43",
          5295 => x"83",
          5296 => x"34",
          5297 => x"33",
          5298 => x"1b",
          5299 => x"f8",
          5300 => x"86",
          5301 => x"05",
          5302 => x"bc",
          5303 => x"ff",
          5304 => x"f6",
          5305 => x"f9",
          5306 => x"29",
          5307 => x"5a",
          5308 => x"f8",
          5309 => x"98",
          5310 => x"81",
          5311 => x"ff",
          5312 => x"60",
          5313 => x"a2",
          5314 => x"bd",
          5315 => x"90",
          5316 => x"1a",
          5317 => x"f8",
          5318 => x"0b",
          5319 => x"0c",
          5320 => x"33",
          5321 => x"2e",
          5322 => x"84",
          5323 => x"56",
          5324 => x"38",
          5325 => x"51",
          5326 => x"80",
          5327 => x"c8",
          5328 => x"0d",
          5329 => x"b0",
          5330 => x"f8",
          5331 => x"b1",
          5332 => x"f9",
          5333 => x"b2",
          5334 => x"83",
          5335 => x"ff",
          5336 => x"f8",
          5337 => x"b9",
          5338 => x"f8",
          5339 => x"b9",
          5340 => x"f8",
          5341 => x"b9",
          5342 => x"9e",
          5343 => x"c9",
          5344 => x"80",
          5345 => x"38",
          5346 => x"22",
          5347 => x"2e",
          5348 => x"ff",
          5349 => x"f8",
          5350 => x"05",
          5351 => x"f8",
          5352 => x"54",
          5353 => x"e4",
          5354 => x"3d",
          5355 => x"fe",
          5356 => x"76",
          5357 => x"f2",
          5358 => x"c8",
          5359 => x"06",
          5360 => x"33",
          5361 => x"41",
          5362 => x"fe",
          5363 => x"52",
          5364 => x"51",
          5365 => x"3f",
          5366 => x"80",
          5367 => x"c9",
          5368 => x"79",
          5369 => x"5b",
          5370 => x"fe",
          5371 => x"10",
          5372 => x"05",
          5373 => x"57",
          5374 => x"26",
          5375 => x"75",
          5376 => x"c7",
          5377 => x"7e",
          5378 => x"b8",
          5379 => x"7d",
          5380 => x"a4",
          5381 => x"f8",
          5382 => x"9d",
          5383 => x"31",
          5384 => x"9f",
          5385 => x"5a",
          5386 => x"5c",
          5387 => x"f8",
          5388 => x"39",
          5389 => x"33",
          5390 => x"2e",
          5391 => x"84",
          5392 => x"ff",
          5393 => x"ff",
          5394 => x"bc",
          5395 => x"5f",
          5396 => x"fd",
          5397 => x"83",
          5398 => x"fd",
          5399 => x"0b",
          5400 => x"34",
          5401 => x"33",
          5402 => x"06",
          5403 => x"80",
          5404 => x"38",
          5405 => x"75",
          5406 => x"34",
          5407 => x"80",
          5408 => x"f9",
          5409 => x"f8",
          5410 => x"bb",
          5411 => x"57",
          5412 => x"25",
          5413 => x"81",
          5414 => x"83",
          5415 => x"fc",
          5416 => x"b8",
          5417 => x"7f",
          5418 => x"e0",
          5419 => x"f9",
          5420 => x"9d",
          5421 => x"31",
          5422 => x"9f",
          5423 => x"5a",
          5424 => x"5a",
          5425 => x"f9",
          5426 => x"39",
          5427 => x"33",
          5428 => x"2e",
          5429 => x"84",
          5430 => x"41",
          5431 => x"09",
          5432 => x"b6",
          5433 => x"bc",
          5434 => x"f9",
          5435 => x"f8",
          5436 => x"29",
          5437 => x"a0",
          5438 => x"f8",
          5439 => x"51",
          5440 => x"60",
          5441 => x"83",
          5442 => x"83",
          5443 => x"87",
          5444 => x"06",
          5445 => x"5d",
          5446 => x"80",
          5447 => x"38",
          5448 => x"f7",
          5449 => x"f2",
          5450 => x"c9",
          5451 => x"80",
          5452 => x"38",
          5453 => x"22",
          5454 => x"2e",
          5455 => x"fb",
          5456 => x"0b",
          5457 => x"34",
          5458 => x"84",
          5459 => x"56",
          5460 => x"90",
          5461 => x"b9",
          5462 => x"f8",
          5463 => x"7c",
          5464 => x"bc",
          5465 => x"59",
          5466 => x"7d",
          5467 => x"75",
          5468 => x"f8",
          5469 => x"a2",
          5470 => x"c9",
          5471 => x"80",
          5472 => x"38",
          5473 => x"33",
          5474 => x"33",
          5475 => x"84",
          5476 => x"ff",
          5477 => x"56",
          5478 => x"83",
          5479 => x"76",
          5480 => x"34",
          5481 => x"83",
          5482 => x"fe",
          5483 => x"80",
          5484 => x"c9",
          5485 => x"76",
          5486 => x"c7",
          5487 => x"84",
          5488 => x"70",
          5489 => x"83",
          5490 => x"fe",
          5491 => x"81",
          5492 => x"ff",
          5493 => x"c9",
          5494 => x"58",
          5495 => x"0b",
          5496 => x"33",
          5497 => x"80",
          5498 => x"84",
          5499 => x"56",
          5500 => x"83",
          5501 => x"81",
          5502 => x"ff",
          5503 => x"f3",
          5504 => x"39",
          5505 => x"33",
          5506 => x"27",
          5507 => x"84",
          5508 => x"ff",
          5509 => x"ff",
          5510 => x"9d",
          5511 => x"70",
          5512 => x"84",
          5513 => x"70",
          5514 => x"ff",
          5515 => x"52",
          5516 => x"5c",
          5517 => x"83",
          5518 => x"79",
          5519 => x"23",
          5520 => x"06",
          5521 => x"5f",
          5522 => x"83",
          5523 => x"76",
          5524 => x"34",
          5525 => x"33",
          5526 => x"40",
          5527 => x"f9",
          5528 => x"56",
          5529 => x"f9",
          5530 => x"39",
          5531 => x"33",
          5532 => x"2e",
          5533 => x"84",
          5534 => x"84",
          5535 => x"40",
          5536 => x"26",
          5537 => x"83",
          5538 => x"84",
          5539 => x"70",
          5540 => x"83",
          5541 => x"71",
          5542 => x"86",
          5543 => x"05",
          5544 => x"22",
          5545 => x"7e",
          5546 => x"83",
          5547 => x"83",
          5548 => x"46",
          5549 => x"5f",
          5550 => x"2e",
          5551 => x"79",
          5552 => x"06",
          5553 => x"5d",
          5554 => x"24",
          5555 => x"84",
          5556 => x"56",
          5557 => x"8e",
          5558 => x"16",
          5559 => x"f8",
          5560 => x"81",
          5561 => x"7c",
          5562 => x"80",
          5563 => x"e5",
          5564 => x"bb",
          5565 => x"76",
          5566 => x"38",
          5567 => x"75",
          5568 => x"34",
          5569 => x"06",
          5570 => x"22",
          5571 => x"5a",
          5572 => x"90",
          5573 => x"31",
          5574 => x"81",
          5575 => x"71",
          5576 => x"5b",
          5577 => x"a7",
          5578 => x"86",
          5579 => x"7f",
          5580 => x"7f",
          5581 => x"71",
          5582 => x"42",
          5583 => x"79",
          5584 => x"d6",
          5585 => x"9a",
          5586 => x"e0",
          5587 => x"84",
          5588 => x"33",
          5589 => x"05",
          5590 => x"70",
          5591 => x"33",
          5592 => x"05",
          5593 => x"18",
          5594 => x"33",
          5595 => x"33",
          5596 => x"1d",
          5597 => x"58",
          5598 => x"f7",
          5599 => x"e0",
          5600 => x"84",
          5601 => x"33",
          5602 => x"05",
          5603 => x"70",
          5604 => x"33",
          5605 => x"05",
          5606 => x"18",
          5607 => x"33",
          5608 => x"33",
          5609 => x"1d",
          5610 => x"58",
          5611 => x"ff",
          5612 => x"e6",
          5613 => x"c9",
          5614 => x"80",
          5615 => x"38",
          5616 => x"b9",
          5617 => x"d8",
          5618 => x"ce",
          5619 => x"84",
          5620 => x"ff",
          5621 => x"c9",
          5622 => x"40",
          5623 => x"2e",
          5624 => x"b9",
          5625 => x"75",
          5626 => x"81",
          5627 => x"38",
          5628 => x"33",
          5629 => x"ff",
          5630 => x"f8",
          5631 => x"5c",
          5632 => x"2e",
          5633 => x"84",
          5634 => x"40",
          5635 => x"f6",
          5636 => x"81",
          5637 => x"60",
          5638 => x"fe",
          5639 => x"26",
          5640 => x"07",
          5641 => x"f2",
          5642 => x"10",
          5643 => x"29",
          5644 => x"a7",
          5645 => x"70",
          5646 => x"86",
          5647 => x"05",
          5648 => x"58",
          5649 => x"8b",
          5650 => x"83",
          5651 => x"8b",
          5652 => x"f8",
          5653 => x"98",
          5654 => x"2b",
          5655 => x"2b",
          5656 => x"79",
          5657 => x"5f",
          5658 => x"27",
          5659 => x"77",
          5660 => x"59",
          5661 => x"70",
          5662 => x"0c",
          5663 => x"ee",
          5664 => x"bc",
          5665 => x"bb",
          5666 => x"7e",
          5667 => x"60",
          5668 => x"83",
          5669 => x"7d",
          5670 => x"05",
          5671 => x"5a",
          5672 => x"8c",
          5673 => x"31",
          5674 => x"29",
          5675 => x"40",
          5676 => x"57",
          5677 => x"26",
          5678 => x"83",
          5679 => x"84",
          5680 => x"59",
          5681 => x"e0",
          5682 => x"79",
          5683 => x"05",
          5684 => x"17",
          5685 => x"26",
          5686 => x"a0",
          5687 => x"19",
          5688 => x"70",
          5689 => x"34",
          5690 => x"75",
          5691 => x"38",
          5692 => x"ff",
          5693 => x"ff",
          5694 => x"fe",
          5695 => x"f8",
          5696 => x"80",
          5697 => x"84",
          5698 => x"06",
          5699 => x"07",
          5700 => x"7b",
          5701 => x"09",
          5702 => x"38",
          5703 => x"83",
          5704 => x"81",
          5705 => x"ff",
          5706 => x"f5",
          5707 => x"f8",
          5708 => x"5e",
          5709 => x"1e",
          5710 => x"83",
          5711 => x"84",
          5712 => x"83",
          5713 => x"84",
          5714 => x"42",
          5715 => x"fa",
          5716 => x"f8",
          5717 => x"07",
          5718 => x"f8",
          5719 => x"18",
          5720 => x"06",
          5721 => x"fb",
          5722 => x"f4",
          5723 => x"06",
          5724 => x"75",
          5725 => x"34",
          5726 => x"f8",
          5727 => x"fb",
          5728 => x"56",
          5729 => x"f4",
          5730 => x"83",
          5731 => x"81",
          5732 => x"07",
          5733 => x"f8",
          5734 => x"39",
          5735 => x"33",
          5736 => x"90",
          5737 => x"83",
          5738 => x"ff",
          5739 => x"f1",
          5740 => x"f4",
          5741 => x"70",
          5742 => x"59",
          5743 => x"39",
          5744 => x"33",
          5745 => x"56",
          5746 => x"f4",
          5747 => x"39",
          5748 => x"33",
          5749 => x"90",
          5750 => x"83",
          5751 => x"fe",
          5752 => x"f8",
          5753 => x"ef",
          5754 => x"07",
          5755 => x"f8",
          5756 => x"ea",
          5757 => x"f4",
          5758 => x"06",
          5759 => x"56",
          5760 => x"f4",
          5761 => x"39",
          5762 => x"33",
          5763 => x"a0",
          5764 => x"83",
          5765 => x"fe",
          5766 => x"f8",
          5767 => x"fe",
          5768 => x"56",
          5769 => x"f4",
          5770 => x"39",
          5771 => x"33",
          5772 => x"84",
          5773 => x"83",
          5774 => x"fe",
          5775 => x"f8",
          5776 => x"fa",
          5777 => x"56",
          5778 => x"f4",
          5779 => x"39",
          5780 => x"33",
          5781 => x"56",
          5782 => x"f4",
          5783 => x"39",
          5784 => x"33",
          5785 => x"56",
          5786 => x"f4",
          5787 => x"39",
          5788 => x"33",
          5789 => x"56",
          5790 => x"f4",
          5791 => x"39",
          5792 => x"33",
          5793 => x"80",
          5794 => x"75",
          5795 => x"34",
          5796 => x"83",
          5797 => x"81",
          5798 => x"07",
          5799 => x"f8",
          5800 => x"ba",
          5801 => x"83",
          5802 => x"80",
          5803 => x"d2",
          5804 => x"ff",
          5805 => x"b0",
          5806 => x"f8",
          5807 => x"b1",
          5808 => x"f9",
          5809 => x"b2",
          5810 => x"83",
          5811 => x"80",
          5812 => x"c4",
          5813 => x"39",
          5814 => x"b8",
          5815 => x"0b",
          5816 => x"0c",
          5817 => x"04",
          5818 => x"f9",
          5819 => x"f9",
          5820 => x"ff",
          5821 => x"05",
          5822 => x"39",
          5823 => x"42",
          5824 => x"11",
          5825 => x"51",
          5826 => x"3f",
          5827 => x"08",
          5828 => x"b9",
          5829 => x"b8",
          5830 => x"0b",
          5831 => x"34",
          5832 => x"b9",
          5833 => x"3d",
          5834 => x"83",
          5835 => x"ef",
          5836 => x"b8",
          5837 => x"11",
          5838 => x"84",
          5839 => x"7b",
          5840 => x"06",
          5841 => x"ca",
          5842 => x"b9",
          5843 => x"80",
          5844 => x"c8",
          5845 => x"80",
          5846 => x"f9",
          5847 => x"81",
          5848 => x"3f",
          5849 => x"33",
          5850 => x"06",
          5851 => x"56",
          5852 => x"80",
          5853 => x"f9",
          5854 => x"81",
          5855 => x"3f",
          5856 => x"8a",
          5857 => x"d8",
          5858 => x"39",
          5859 => x"33",
          5860 => x"09",
          5861 => x"72",
          5862 => x"57",
          5863 => x"75",
          5864 => x"d9",
          5865 => x"bc",
          5866 => x"60",
          5867 => x"38",
          5868 => x"f9",
          5869 => x"39",
          5870 => x"33",
          5871 => x"09",
          5872 => x"72",
          5873 => x"57",
          5874 => x"83",
          5875 => x"81",
          5876 => x"bb",
          5877 => x"59",
          5878 => x"78",
          5879 => x"38",
          5880 => x"bb",
          5881 => x"bb",
          5882 => x"ff",
          5883 => x"81",
          5884 => x"a6",
          5885 => x"f8",
          5886 => x"bc",
          5887 => x"ff",
          5888 => x"f9",
          5889 => x"29",
          5890 => x"a0",
          5891 => x"f8",
          5892 => x"5f",
          5893 => x"05",
          5894 => x"ff",
          5895 => x"ce",
          5896 => x"44",
          5897 => x"77",
          5898 => x"f5",
          5899 => x"ff",
          5900 => x"11",
          5901 => x"7b",
          5902 => x"38",
          5903 => x"33",
          5904 => x"27",
          5905 => x"ff",
          5906 => x"83",
          5907 => x"7c",
          5908 => x"ff",
          5909 => x"80",
          5910 => x"df",
          5911 => x"bb",
          5912 => x"76",
          5913 => x"38",
          5914 => x"75",
          5915 => x"34",
          5916 => x"06",
          5917 => x"22",
          5918 => x"5a",
          5919 => x"90",
          5920 => x"31",
          5921 => x"81",
          5922 => x"71",
          5923 => x"5f",
          5924 => x"a7",
          5925 => x"86",
          5926 => x"7c",
          5927 => x"7f",
          5928 => x"71",
          5929 => x"41",
          5930 => x"79",
          5931 => x"ea",
          5932 => x"9a",
          5933 => x"e0",
          5934 => x"84",
          5935 => x"33",
          5936 => x"05",
          5937 => x"70",
          5938 => x"33",
          5939 => x"05",
          5940 => x"18",
          5941 => x"33",
          5942 => x"33",
          5943 => x"1d",
          5944 => x"58",
          5945 => x"ec",
          5946 => x"e0",
          5947 => x"84",
          5948 => x"33",
          5949 => x"05",
          5950 => x"70",
          5951 => x"33",
          5952 => x"05",
          5953 => x"18",
          5954 => x"33",
          5955 => x"33",
          5956 => x"1d",
          5957 => x"58",
          5958 => x"ff",
          5959 => x"fa",
          5960 => x"fa",
          5961 => x"84",
          5962 => x"33",
          5963 => x"f8",
          5964 => x"b7",
          5965 => x"f8",
          5966 => x"b7",
          5967 => x"5c",
          5968 => x"e9",
          5969 => x"d2",
          5970 => x"bb",
          5971 => x"ff",
          5972 => x"5c",
          5973 => x"61",
          5974 => x"76",
          5975 => x"f8",
          5976 => x"81",
          5977 => x"19",
          5978 => x"7a",
          5979 => x"80",
          5980 => x"f8",
          5981 => x"b7",
          5982 => x"81",
          5983 => x"12",
          5984 => x"80",
          5985 => x"8d",
          5986 => x"75",
          5987 => x"34",
          5988 => x"83",
          5989 => x"81",
          5990 => x"bc",
          5991 => x"59",
          5992 => x"7f",
          5993 => x"38",
          5994 => x"c5",
          5995 => x"2e",
          5996 => x"f4",
          5997 => x"f8",
          5998 => x"81",
          5999 => x"f8",
          6000 => x"44",
          6001 => x"76",
          6002 => x"81",
          6003 => x"38",
          6004 => x"ff",
          6005 => x"83",
          6006 => x"fd",
          6007 => x"1a",
          6008 => x"f8",
          6009 => x"e7",
          6010 => x"31",
          6011 => x"f8",
          6012 => x"90",
          6013 => x"58",
          6014 => x"26",
          6015 => x"80",
          6016 => x"05",
          6017 => x"f8",
          6018 => x"70",
          6019 => x"34",
          6020 => x"f4",
          6021 => x"76",
          6022 => x"58",
          6023 => x"f4",
          6024 => x"81",
          6025 => x"79",
          6026 => x"38",
          6027 => x"79",
          6028 => x"75",
          6029 => x"23",
          6030 => x"80",
          6031 => x"f8",
          6032 => x"39",
          6033 => x"f6",
          6034 => x"39",
          6035 => x"f8",
          6036 => x"8e",
          6037 => x"83",
          6038 => x"f1",
          6039 => x"f8",
          6040 => x"5a",
          6041 => x"1a",
          6042 => x"80",
          6043 => x"cd",
          6044 => x"39",
          6045 => x"02",
          6046 => x"84",
          6047 => x"54",
          6048 => x"2e",
          6049 => x"51",
          6050 => x"80",
          6051 => x"c8",
          6052 => x"0d",
          6053 => x"73",
          6054 => x"3f",
          6055 => x"b9",
          6056 => x"3d",
          6057 => x"3d",
          6058 => x"05",
          6059 => x"0b",
          6060 => x"33",
          6061 => x"06",
          6062 => x"11",
          6063 => x"55",
          6064 => x"2e",
          6065 => x"81",
          6066 => x"83",
          6067 => x"74",
          6068 => x"b9",
          6069 => x"3d",
          6070 => x"f7",
          6071 => x"82",
          6072 => x"2e",
          6073 => x"73",
          6074 => x"71",
          6075 => x"70",
          6076 => x"5d",
          6077 => x"83",
          6078 => x"ff",
          6079 => x"7b",
          6080 => x"81",
          6081 => x"7b",
          6082 => x"32",
          6083 => x"80",
          6084 => x"5c",
          6085 => x"80",
          6086 => x"38",
          6087 => x"33",
          6088 => x"33",
          6089 => x"33",
          6090 => x"12",
          6091 => x"80",
          6092 => x"f6",
          6093 => x"5d",
          6094 => x"05",
          6095 => x"ff",
          6096 => x"cd",
          6097 => x"55",
          6098 => x"2e",
          6099 => x"81",
          6100 => x"87",
          6101 => x"34",
          6102 => x"c0",
          6103 => x"87",
          6104 => x"08",
          6105 => x"2e",
          6106 => x"8e",
          6107 => x"57",
          6108 => x"f8",
          6109 => x"14",
          6110 => x"06",
          6111 => x"f9",
          6112 => x"38",
          6113 => x"f6",
          6114 => x"70",
          6115 => x"83",
          6116 => x"33",
          6117 => x"72",
          6118 => x"c1",
          6119 => x"ff",
          6120 => x"38",
          6121 => x"fc",
          6122 => x"81",
          6123 => x"79",
          6124 => x"85",
          6125 => x"83",
          6126 => x"34",
          6127 => x"14",
          6128 => x"f2",
          6129 => x"14",
          6130 => x"06",
          6131 => x"74",
          6132 => x"38",
          6133 => x"33",
          6134 => x"70",
          6135 => x"56",
          6136 => x"f7",
          6137 => x"81",
          6138 => x"86",
          6139 => x"70",
          6140 => x"54",
          6141 => x"2e",
          6142 => x"81",
          6143 => x"a1",
          6144 => x"81",
          6145 => x"80",
          6146 => x"38",
          6147 => x"f7",
          6148 => x"0b",
          6149 => x"33",
          6150 => x"08",
          6151 => x"33",
          6152 => x"a4",
          6153 => x"a3",
          6154 => x"42",
          6155 => x"56",
          6156 => x"16",
          6157 => x"81",
          6158 => x"38",
          6159 => x"16",
          6160 => x"80",
          6161 => x"38",
          6162 => x"16",
          6163 => x"81",
          6164 => x"38",
          6165 => x"16",
          6166 => x"81",
          6167 => x"81",
          6168 => x"73",
          6169 => x"8d",
          6170 => x"90",
          6171 => x"72",
          6172 => x"da",
          6173 => x"ff",
          6174 => x"81",
          6175 => x"8c",
          6176 => x"90",
          6177 => x"81",
          6178 => x"80",
          6179 => x"9c",
          6180 => x"05",
          6181 => x"9c",
          6182 => x"73",
          6183 => x"ec",
          6184 => x"87",
          6185 => x"08",
          6186 => x"0c",
          6187 => x"70",
          6188 => x"57",
          6189 => x"27",
          6190 => x"76",
          6191 => x"34",
          6192 => x"a4",
          6193 => x"19",
          6194 => x"26",
          6195 => x"72",
          6196 => x"c8",
          6197 => x"79",
          6198 => x"f7",
          6199 => x"73",
          6200 => x"38",
          6201 => x"87",
          6202 => x"08",
          6203 => x"7d",
          6204 => x"38",
          6205 => x"f7",
          6206 => x"54",
          6207 => x"83",
          6208 => x"73",
          6209 => x"34",
          6210 => x"9c",
          6211 => x"d0",
          6212 => x"ff",
          6213 => x"81",
          6214 => x"83",
          6215 => x"33",
          6216 => x"c4",
          6217 => x"34",
          6218 => x"fc",
          6219 => x"f7",
          6220 => x"72",
          6221 => x"9c",
          6222 => x"2e",
          6223 => x"80",
          6224 => x"81",
          6225 => x"8a",
          6226 => x"fe",
          6227 => x"74",
          6228 => x"59",
          6229 => x"9b",
          6230 => x"2e",
          6231 => x"83",
          6232 => x"81",
          6233 => x"38",
          6234 => x"80",
          6235 => x"81",
          6236 => x"87",
          6237 => x"98",
          6238 => x"72",
          6239 => x"38",
          6240 => x"9c",
          6241 => x"70",
          6242 => x"76",
          6243 => x"06",
          6244 => x"71",
          6245 => x"53",
          6246 => x"80",
          6247 => x"38",
          6248 => x"10",
          6249 => x"76",
          6250 => x"78",
          6251 => x"d8",
          6252 => x"5b",
          6253 => x"87",
          6254 => x"08",
          6255 => x"0c",
          6256 => x"39",
          6257 => x"81",
          6258 => x"38",
          6259 => x"06",
          6260 => x"39",
          6261 => x"9b",
          6262 => x"2e",
          6263 => x"80",
          6264 => x"be",
          6265 => x"72",
          6266 => x"e8",
          6267 => x"32",
          6268 => x"80",
          6269 => x"40",
          6270 => x"8a",
          6271 => x"2e",
          6272 => x"f9",
          6273 => x"ff",
          6274 => x"38",
          6275 => x"10",
          6276 => x"f7",
          6277 => x"33",
          6278 => x"7c",
          6279 => x"38",
          6280 => x"81",
          6281 => x"57",
          6282 => x"e2",
          6283 => x"bf",
          6284 => x"80",
          6285 => x"38",
          6286 => x"33",
          6287 => x"91",
          6288 => x"ff",
          6289 => x"51",
          6290 => x"78",
          6291 => x"0c",
          6292 => x"04",
          6293 => x"81",
          6294 => x"f6",
          6295 => x"ff",
          6296 => x"83",
          6297 => x"33",
          6298 => x"7a",
          6299 => x"15",
          6300 => x"39",
          6301 => x"f7",
          6302 => x"ff",
          6303 => x"fc",
          6304 => x"0b",
          6305 => x"15",
          6306 => x"39",
          6307 => x"06",
          6308 => x"ff",
          6309 => x"38",
          6310 => x"16",
          6311 => x"75",
          6312 => x"38",
          6313 => x"06",
          6314 => x"2e",
          6315 => x"fb",
          6316 => x"f7",
          6317 => x"fa",
          6318 => x"98",
          6319 => x"55",
          6320 => x"fb",
          6321 => x"c0",
          6322 => x"83",
          6323 => x"76",
          6324 => x"59",
          6325 => x"ff",
          6326 => x"fc",
          6327 => x"ca",
          6328 => x"f7",
          6329 => x"09",
          6330 => x"72",
          6331 => x"72",
          6332 => x"34",
          6333 => x"f7",
          6334 => x"f7",
          6335 => x"f7",
          6336 => x"83",
          6337 => x"83",
          6338 => x"5d",
          6339 => x"5c",
          6340 => x"9c",
          6341 => x"2e",
          6342 => x"fc",
          6343 => x"59",
          6344 => x"fc",
          6345 => x"81",
          6346 => x"06",
          6347 => x"fd",
          6348 => x"76",
          6349 => x"54",
          6350 => x"80",
          6351 => x"bf",
          6352 => x"75",
          6353 => x"54",
          6354 => x"bf",
          6355 => x"f7",
          6356 => x"0b",
          6357 => x"33",
          6358 => x"83",
          6359 => x"73",
          6360 => x"34",
          6361 => x"95",
          6362 => x"83",
          6363 => x"84",
          6364 => x"38",
          6365 => x"f7",
          6366 => x"ff",
          6367 => x"bb",
          6368 => x"ff",
          6369 => x"57",
          6370 => x"79",
          6371 => x"80",
          6372 => x"f8",
          6373 => x"81",
          6374 => x"15",
          6375 => x"73",
          6376 => x"80",
          6377 => x"f8",
          6378 => x"b7",
          6379 => x"81",
          6380 => x"ff",
          6381 => x"75",
          6382 => x"80",
          6383 => x"f8",
          6384 => x"59",
          6385 => x"81",
          6386 => x"ff",
          6387 => x"ff",
          6388 => x"39",
          6389 => x"95",
          6390 => x"08",
          6391 => x"ac",
          6392 => x"e5",
          6393 => x"83",
          6394 => x"83",
          6395 => x"59",
          6396 => x"80",
          6397 => x"51",
          6398 => x"82",
          6399 => x"fa",
          6400 => x"0b",
          6401 => x"08",
          6402 => x"a3",
          6403 => x"13",
          6404 => x"d4",
          6405 => x"e0",
          6406 => x"0b",
          6407 => x"08",
          6408 => x"0b",
          6409 => x"80",
          6410 => x"80",
          6411 => x"c0",
          6412 => x"83",
          6413 => x"55",
          6414 => x"05",
          6415 => x"98",
          6416 => x"87",
          6417 => x"08",
          6418 => x"2e",
          6419 => x"14",
          6420 => x"98",
          6421 => x"52",
          6422 => x"87",
          6423 => x"fe",
          6424 => x"87",
          6425 => x"08",
          6426 => x"70",
          6427 => x"c8",
          6428 => x"71",
          6429 => x"c0",
          6430 => x"98",
          6431 => x"ce",
          6432 => x"87",
          6433 => x"08",
          6434 => x"98",
          6435 => x"74",
          6436 => x"38",
          6437 => x"87",
          6438 => x"08",
          6439 => x"73",
          6440 => x"71",
          6441 => x"db",
          6442 => x"98",
          6443 => x"72",
          6444 => x"38",
          6445 => x"55",
          6446 => x"81",
          6447 => x"53",
          6448 => x"98",
          6449 => x"ff",
          6450 => x"fe",
          6451 => x"ff",
          6452 => x"76",
          6453 => x"0c",
          6454 => x"04",
          6455 => x"b9",
          6456 => x"3d",
          6457 => x"3d",
          6458 => x"84",
          6459 => x"33",
          6460 => x"0b",
          6461 => x"08",
          6462 => x"87",
          6463 => x"06",
          6464 => x"2a",
          6465 => x"55",
          6466 => x"15",
          6467 => x"2a",
          6468 => x"15",
          6469 => x"2a",
          6470 => x"15",
          6471 => x"15",
          6472 => x"d4",
          6473 => x"82",
          6474 => x"f3",
          6475 => x"80",
          6476 => x"85",
          6477 => x"d4",
          6478 => x"fe",
          6479 => x"34",
          6480 => x"90",
          6481 => x"87",
          6482 => x"08",
          6483 => x"08",
          6484 => x"90",
          6485 => x"c0",
          6486 => x"52",
          6487 => x"9c",
          6488 => x"72",
          6489 => x"81",
          6490 => x"c0",
          6491 => x"56",
          6492 => x"27",
          6493 => x"81",
          6494 => x"38",
          6495 => x"a4",
          6496 => x"55",
          6497 => x"80",
          6498 => x"55",
          6499 => x"80",
          6500 => x"c0",
          6501 => x"80",
          6502 => x"53",
          6503 => x"9c",
          6504 => x"c0",
          6505 => x"55",
          6506 => x"f6",
          6507 => x"33",
          6508 => x"9c",
          6509 => x"70",
          6510 => x"38",
          6511 => x"2e",
          6512 => x"c0",
          6513 => x"55",
          6514 => x"83",
          6515 => x"71",
          6516 => x"70",
          6517 => x"57",
          6518 => x"2e",
          6519 => x"74",
          6520 => x"52",
          6521 => x"38",
          6522 => x"81",
          6523 => x"75",
          6524 => x"c6",
          6525 => x"80",
          6526 => x"52",
          6527 => x"92",
          6528 => x"81",
          6529 => x"71",
          6530 => x"53",
          6531 => x"26",
          6532 => x"84",
          6533 => x"88",
          6534 => x"81",
          6535 => x"c8",
          6536 => x"0d",
          6537 => x"c2",
          6538 => x"0d",
          6539 => x"05",
          6540 => x"56",
          6541 => x"83",
          6542 => x"77",
          6543 => x"fc",
          6544 => x"70",
          6545 => x"07",
          6546 => x"57",
          6547 => x"34",
          6548 => x"51",
          6549 => x"34",
          6550 => x"52",
          6551 => x"34",
          6552 => x"34",
          6553 => x"d4",
          6554 => x"11",
          6555 => x"56",
          6556 => x"70",
          6557 => x"38",
          6558 => x"05",
          6559 => x"70",
          6560 => x"34",
          6561 => x"f0",
          6562 => x"d4",
          6563 => x"82",
          6564 => x"f3",
          6565 => x"80",
          6566 => x"85",
          6567 => x"d4",
          6568 => x"fe",
          6569 => x"34",
          6570 => x"90",
          6571 => x"87",
          6572 => x"08",
          6573 => x"08",
          6574 => x"90",
          6575 => x"c0",
          6576 => x"52",
          6577 => x"9c",
          6578 => x"72",
          6579 => x"81",
          6580 => x"c0",
          6581 => x"56",
          6582 => x"27",
          6583 => x"81",
          6584 => x"38",
          6585 => x"a4",
          6586 => x"55",
          6587 => x"80",
          6588 => x"55",
          6589 => x"80",
          6590 => x"c0",
          6591 => x"80",
          6592 => x"53",
          6593 => x"9c",
          6594 => x"c0",
          6595 => x"55",
          6596 => x"f6",
          6597 => x"33",
          6598 => x"9c",
          6599 => x"70",
          6600 => x"38",
          6601 => x"2e",
          6602 => x"c0",
          6603 => x"55",
          6604 => x"83",
          6605 => x"71",
          6606 => x"70",
          6607 => x"57",
          6608 => x"2e",
          6609 => x"81",
          6610 => x"71",
          6611 => x"74",
          6612 => x"ff",
          6613 => x"80",
          6614 => x"81",
          6615 => x"b9",
          6616 => x"3d",
          6617 => x"51",
          6618 => x"3d",
          6619 => x"d4",
          6620 => x"d0",
          6621 => x"0b",
          6622 => x"08",
          6623 => x"0b",
          6624 => x"80",
          6625 => x"80",
          6626 => x"c0",
          6627 => x"83",
          6628 => x"56",
          6629 => x"05",
          6630 => x"98",
          6631 => x"87",
          6632 => x"08",
          6633 => x"2e",
          6634 => x"15",
          6635 => x"98",
          6636 => x"52",
          6637 => x"87",
          6638 => x"fe",
          6639 => x"87",
          6640 => x"08",
          6641 => x"70",
          6642 => x"c8",
          6643 => x"71",
          6644 => x"c0",
          6645 => x"98",
          6646 => x"ce",
          6647 => x"87",
          6648 => x"08",
          6649 => x"98",
          6650 => x"70",
          6651 => x"38",
          6652 => x"87",
          6653 => x"08",
          6654 => x"73",
          6655 => x"71",
          6656 => x"db",
          6657 => x"98",
          6658 => x"72",
          6659 => x"38",
          6660 => x"53",
          6661 => x"81",
          6662 => x"52",
          6663 => x"8a",
          6664 => x"ff",
          6665 => x"fe",
          6666 => x"39",
          6667 => x"83",
          6668 => x"fe",
          6669 => x"82",
          6670 => x"f9",
          6671 => x"b9",
          6672 => x"71",
          6673 => x"70",
          6674 => x"06",
          6675 => x"73",
          6676 => x"81",
          6677 => x"8b",
          6678 => x"2b",
          6679 => x"70",
          6680 => x"33",
          6681 => x"71",
          6682 => x"5c",
          6683 => x"53",
          6684 => x"52",
          6685 => x"80",
          6686 => x"af",
          6687 => x"82",
          6688 => x"12",
          6689 => x"2b",
          6690 => x"07",
          6691 => x"33",
          6692 => x"71",
          6693 => x"90",
          6694 => x"53",
          6695 => x"56",
          6696 => x"24",
          6697 => x"84",
          6698 => x"14",
          6699 => x"2b",
          6700 => x"07",
          6701 => x"88",
          6702 => x"56",
          6703 => x"13",
          6704 => x"ff",
          6705 => x"87",
          6706 => x"b9",
          6707 => x"17",
          6708 => x"85",
          6709 => x"88",
          6710 => x"88",
          6711 => x"59",
          6712 => x"84",
          6713 => x"85",
          6714 => x"b9",
          6715 => x"52",
          6716 => x"13",
          6717 => x"87",
          6718 => x"b9",
          6719 => x"74",
          6720 => x"73",
          6721 => x"84",
          6722 => x"16",
          6723 => x"12",
          6724 => x"2b",
          6725 => x"80",
          6726 => x"2a",
          6727 => x"52",
          6728 => x"75",
          6729 => x"89",
          6730 => x"86",
          6731 => x"13",
          6732 => x"2b",
          6733 => x"07",
          6734 => x"16",
          6735 => x"33",
          6736 => x"07",
          6737 => x"58",
          6738 => x"53",
          6739 => x"84",
          6740 => x"85",
          6741 => x"b9",
          6742 => x"16",
          6743 => x"85",
          6744 => x"8b",
          6745 => x"2b",
          6746 => x"5a",
          6747 => x"86",
          6748 => x"13",
          6749 => x"2b",
          6750 => x"2a",
          6751 => x"52",
          6752 => x"34",
          6753 => x"34",
          6754 => x"08",
          6755 => x"81",
          6756 => x"88",
          6757 => x"ff",
          6758 => x"88",
          6759 => x"54",
          6760 => x"34",
          6761 => x"34",
          6762 => x"08",
          6763 => x"33",
          6764 => x"71",
          6765 => x"83",
          6766 => x"05",
          6767 => x"12",
          6768 => x"2b",
          6769 => x"2b",
          6770 => x"06",
          6771 => x"88",
          6772 => x"53",
          6773 => x"57",
          6774 => x"82",
          6775 => x"83",
          6776 => x"b9",
          6777 => x"17",
          6778 => x"12",
          6779 => x"2b",
          6780 => x"07",
          6781 => x"33",
          6782 => x"71",
          6783 => x"81",
          6784 => x"70",
          6785 => x"52",
          6786 => x"57",
          6787 => x"73",
          6788 => x"14",
          6789 => x"b8",
          6790 => x"82",
          6791 => x"12",
          6792 => x"2b",
          6793 => x"07",
          6794 => x"33",
          6795 => x"71",
          6796 => x"90",
          6797 => x"53",
          6798 => x"57",
          6799 => x"80",
          6800 => x"38",
          6801 => x"13",
          6802 => x"2b",
          6803 => x"80",
          6804 => x"2a",
          6805 => x"76",
          6806 => x"81",
          6807 => x"b9",
          6808 => x"17",
          6809 => x"12",
          6810 => x"2b",
          6811 => x"07",
          6812 => x"14",
          6813 => x"33",
          6814 => x"07",
          6815 => x"57",
          6816 => x"58",
          6817 => x"72",
          6818 => x"75",
          6819 => x"89",
          6820 => x"f9",
          6821 => x"84",
          6822 => x"58",
          6823 => x"2e",
          6824 => x"80",
          6825 => x"77",
          6826 => x"3f",
          6827 => x"04",
          6828 => x"0b",
          6829 => x"0c",
          6830 => x"84",
          6831 => x"82",
          6832 => x"76",
          6833 => x"f4",
          6834 => x"b5",
          6835 => x"b8",
          6836 => x"75",
          6837 => x"81",
          6838 => x"b9",
          6839 => x"76",
          6840 => x"81",
          6841 => x"34",
          6842 => x"08",
          6843 => x"17",
          6844 => x"87",
          6845 => x"b9",
          6846 => x"b9",
          6847 => x"05",
          6848 => x"07",
          6849 => x"ff",
          6850 => x"2a",
          6851 => x"56",
          6852 => x"34",
          6853 => x"34",
          6854 => x"22",
          6855 => x"10",
          6856 => x"08",
          6857 => x"55",
          6858 => x"15",
          6859 => x"83",
          6860 => x"ee",
          6861 => x"0d",
          6862 => x"53",
          6863 => x"72",
          6864 => x"fb",
          6865 => x"82",
          6866 => x"ff",
          6867 => x"51",
          6868 => x"ff",
          6869 => x"b8",
          6870 => x"33",
          6871 => x"71",
          6872 => x"70",
          6873 => x"58",
          6874 => x"ff",
          6875 => x"2e",
          6876 => x"75",
          6877 => x"17",
          6878 => x"12",
          6879 => x"2b",
          6880 => x"ff",
          6881 => x"31",
          6882 => x"ff",
          6883 => x"27",
          6884 => x"5c",
          6885 => x"74",
          6886 => x"70",
          6887 => x"38",
          6888 => x"58",
          6889 => x"85",
          6890 => x"88",
          6891 => x"5a",
          6892 => x"73",
          6893 => x"2e",
          6894 => x"74",
          6895 => x"76",
          6896 => x"11",
          6897 => x"12",
          6898 => x"2b",
          6899 => x"ff",
          6900 => x"56",
          6901 => x"59",
          6902 => x"83",
          6903 => x"80",
          6904 => x"26",
          6905 => x"78",
          6906 => x"2e",
          6907 => x"72",
          6908 => x"88",
          6909 => x"70",
          6910 => x"11",
          6911 => x"80",
          6912 => x"2a",
          6913 => x"56",
          6914 => x"34",
          6915 => x"34",
          6916 => x"08",
          6917 => x"2a",
          6918 => x"82",
          6919 => x"83",
          6920 => x"b9",
          6921 => x"19",
          6922 => x"12",
          6923 => x"2b",
          6924 => x"2b",
          6925 => x"06",
          6926 => x"83",
          6927 => x"70",
          6928 => x"58",
          6929 => x"52",
          6930 => x"12",
          6931 => x"ff",
          6932 => x"83",
          6933 => x"b9",
          6934 => x"54",
          6935 => x"72",
          6936 => x"84",
          6937 => x"70",
          6938 => x"33",
          6939 => x"71",
          6940 => x"83",
          6941 => x"05",
          6942 => x"53",
          6943 => x"15",
          6944 => x"15",
          6945 => x"b8",
          6946 => x"55",
          6947 => x"11",
          6948 => x"33",
          6949 => x"07",
          6950 => x"54",
          6951 => x"70",
          6952 => x"71",
          6953 => x"84",
          6954 => x"70",
          6955 => x"33",
          6956 => x"71",
          6957 => x"83",
          6958 => x"05",
          6959 => x"5a",
          6960 => x"15",
          6961 => x"15",
          6962 => x"b8",
          6963 => x"55",
          6964 => x"11",
          6965 => x"33",
          6966 => x"07",
          6967 => x"54",
          6968 => x"70",
          6969 => x"79",
          6970 => x"84",
          6971 => x"18",
          6972 => x"70",
          6973 => x"0c",
          6974 => x"04",
          6975 => x"87",
          6976 => x"8b",
          6977 => x"2b",
          6978 => x"84",
          6979 => x"18",
          6980 => x"2b",
          6981 => x"2a",
          6982 => x"53",
          6983 => x"84",
          6984 => x"85",
          6985 => x"b9",
          6986 => x"19",
          6987 => x"85",
          6988 => x"8b",
          6989 => x"2b",
          6990 => x"86",
          6991 => x"15",
          6992 => x"2b",
          6993 => x"2a",
          6994 => x"52",
          6995 => x"52",
          6996 => x"34",
          6997 => x"34",
          6998 => x"08",
          6999 => x"81",
          7000 => x"88",
          7001 => x"ff",
          7002 => x"88",
          7003 => x"54",
          7004 => x"34",
          7005 => x"34",
          7006 => x"08",
          7007 => x"51",
          7008 => x"f9",
          7009 => x"84",
          7010 => x"58",
          7011 => x"2e",
          7012 => x"54",
          7013 => x"73",
          7014 => x"0c",
          7015 => x"04",
          7016 => x"91",
          7017 => x"c8",
          7018 => x"c8",
          7019 => x"0d",
          7020 => x"f4",
          7021 => x"b8",
          7022 => x"0b",
          7023 => x"23",
          7024 => x"53",
          7025 => x"ff",
          7026 => x"cd",
          7027 => x"b9",
          7028 => x"76",
          7029 => x"0b",
          7030 => x"84",
          7031 => x"54",
          7032 => x"34",
          7033 => x"15",
          7034 => x"b8",
          7035 => x"86",
          7036 => x"0b",
          7037 => x"84",
          7038 => x"84",
          7039 => x"ff",
          7040 => x"80",
          7041 => x"ff",
          7042 => x"88",
          7043 => x"55",
          7044 => x"17",
          7045 => x"17",
          7046 => x"b4",
          7047 => x"10",
          7048 => x"b8",
          7049 => x"05",
          7050 => x"82",
          7051 => x"0b",
          7052 => x"77",
          7053 => x"2e",
          7054 => x"fe",
          7055 => x"3d",
          7056 => x"41",
          7057 => x"84",
          7058 => x"59",
          7059 => x"61",
          7060 => x"38",
          7061 => x"85",
          7062 => x"80",
          7063 => x"38",
          7064 => x"60",
          7065 => x"7f",
          7066 => x"2a",
          7067 => x"83",
          7068 => x"55",
          7069 => x"ff",
          7070 => x"78",
          7071 => x"70",
          7072 => x"06",
          7073 => x"7a",
          7074 => x"81",
          7075 => x"88",
          7076 => x"75",
          7077 => x"ff",
          7078 => x"10",
          7079 => x"05",
          7080 => x"61",
          7081 => x"81",
          7082 => x"88",
          7083 => x"90",
          7084 => x"2c",
          7085 => x"46",
          7086 => x"43",
          7087 => x"59",
          7088 => x"42",
          7089 => x"85",
          7090 => x"15",
          7091 => x"33",
          7092 => x"07",
          7093 => x"10",
          7094 => x"81",
          7095 => x"98",
          7096 => x"2b",
          7097 => x"53",
          7098 => x"80",
          7099 => x"c9",
          7100 => x"27",
          7101 => x"63",
          7102 => x"62",
          7103 => x"38",
          7104 => x"85",
          7105 => x"1b",
          7106 => x"25",
          7107 => x"63",
          7108 => x"79",
          7109 => x"38",
          7110 => x"33",
          7111 => x"71",
          7112 => x"83",
          7113 => x"11",
          7114 => x"12",
          7115 => x"2b",
          7116 => x"07",
          7117 => x"52",
          7118 => x"58",
          7119 => x"8c",
          7120 => x"1e",
          7121 => x"83",
          7122 => x"8b",
          7123 => x"2b",
          7124 => x"86",
          7125 => x"12",
          7126 => x"2b",
          7127 => x"07",
          7128 => x"14",
          7129 => x"33",
          7130 => x"07",
          7131 => x"59",
          7132 => x"5b",
          7133 => x"5c",
          7134 => x"84",
          7135 => x"85",
          7136 => x"b9",
          7137 => x"17",
          7138 => x"85",
          7139 => x"8b",
          7140 => x"2b",
          7141 => x"86",
          7142 => x"15",
          7143 => x"2b",
          7144 => x"2a",
          7145 => x"52",
          7146 => x"57",
          7147 => x"34",
          7148 => x"34",
          7149 => x"08",
          7150 => x"81",
          7151 => x"88",
          7152 => x"ff",
          7153 => x"88",
          7154 => x"5e",
          7155 => x"34",
          7156 => x"34",
          7157 => x"08",
          7158 => x"11",
          7159 => x"33",
          7160 => x"71",
          7161 => x"74",
          7162 => x"81",
          7163 => x"88",
          7164 => x"88",
          7165 => x"45",
          7166 => x"55",
          7167 => x"34",
          7168 => x"34",
          7169 => x"08",
          7170 => x"33",
          7171 => x"71",
          7172 => x"83",
          7173 => x"05",
          7174 => x"83",
          7175 => x"88",
          7176 => x"88",
          7177 => x"45",
          7178 => x"55",
          7179 => x"1a",
          7180 => x"1a",
          7181 => x"b8",
          7182 => x"82",
          7183 => x"12",
          7184 => x"2b",
          7185 => x"62",
          7186 => x"2b",
          7187 => x"5d",
          7188 => x"05",
          7189 => x"ec",
          7190 => x"b8",
          7191 => x"05",
          7192 => x"1c",
          7193 => x"ff",
          7194 => x"5f",
          7195 => x"81",
          7196 => x"54",
          7197 => x"c8",
          7198 => x"0d",
          7199 => x"f4",
          7200 => x"b8",
          7201 => x"0b",
          7202 => x"23",
          7203 => x"53",
          7204 => x"ff",
          7205 => x"c7",
          7206 => x"b9",
          7207 => x"60",
          7208 => x"0b",
          7209 => x"84",
          7210 => x"5d",
          7211 => x"34",
          7212 => x"1e",
          7213 => x"b8",
          7214 => x"86",
          7215 => x"0b",
          7216 => x"84",
          7217 => x"84",
          7218 => x"ff",
          7219 => x"80",
          7220 => x"ff",
          7221 => x"88",
          7222 => x"5b",
          7223 => x"18",
          7224 => x"18",
          7225 => x"b4",
          7226 => x"10",
          7227 => x"b8",
          7228 => x"05",
          7229 => x"82",
          7230 => x"0b",
          7231 => x"84",
          7232 => x"57",
          7233 => x"38",
          7234 => x"82",
          7235 => x"54",
          7236 => x"fe",
          7237 => x"51",
          7238 => x"84",
          7239 => x"84",
          7240 => x"95",
          7241 => x"61",
          7242 => x"b8",
          7243 => x"2b",
          7244 => x"44",
          7245 => x"33",
          7246 => x"71",
          7247 => x"81",
          7248 => x"70",
          7249 => x"44",
          7250 => x"63",
          7251 => x"81",
          7252 => x"84",
          7253 => x"05",
          7254 => x"57",
          7255 => x"19",
          7256 => x"19",
          7257 => x"b8",
          7258 => x"70",
          7259 => x"33",
          7260 => x"07",
          7261 => x"8f",
          7262 => x"74",
          7263 => x"ff",
          7264 => x"88",
          7265 => x"47",
          7266 => x"5d",
          7267 => x"05",
          7268 => x"ff",
          7269 => x"63",
          7270 => x"84",
          7271 => x"1e",
          7272 => x"34",
          7273 => x"34",
          7274 => x"b8",
          7275 => x"05",
          7276 => x"3f",
          7277 => x"bc",
          7278 => x"31",
          7279 => x"ff",
          7280 => x"fa",
          7281 => x"81",
          7282 => x"76",
          7283 => x"ff",
          7284 => x"17",
          7285 => x"33",
          7286 => x"07",
          7287 => x"10",
          7288 => x"81",
          7289 => x"98",
          7290 => x"2b",
          7291 => x"53",
          7292 => x"45",
          7293 => x"25",
          7294 => x"ff",
          7295 => x"78",
          7296 => x"38",
          7297 => x"8b",
          7298 => x"83",
          7299 => x"5b",
          7300 => x"fc",
          7301 => x"8f",
          7302 => x"f4",
          7303 => x"b8",
          7304 => x"0b",
          7305 => x"23",
          7306 => x"53",
          7307 => x"ff",
          7308 => x"c4",
          7309 => x"b9",
          7310 => x"7e",
          7311 => x"0b",
          7312 => x"84",
          7313 => x"59",
          7314 => x"34",
          7315 => x"1a",
          7316 => x"b8",
          7317 => x"86",
          7318 => x"0b",
          7319 => x"84",
          7320 => x"84",
          7321 => x"ff",
          7322 => x"80",
          7323 => x"ff",
          7324 => x"88",
          7325 => x"57",
          7326 => x"88",
          7327 => x"64",
          7328 => x"84",
          7329 => x"70",
          7330 => x"84",
          7331 => x"05",
          7332 => x"43",
          7333 => x"05",
          7334 => x"83",
          7335 => x"ee",
          7336 => x"24",
          7337 => x"61",
          7338 => x"06",
          7339 => x"27",
          7340 => x"fc",
          7341 => x"80",
          7342 => x"38",
          7343 => x"fb",
          7344 => x"73",
          7345 => x"0c",
          7346 => x"04",
          7347 => x"11",
          7348 => x"33",
          7349 => x"71",
          7350 => x"7a",
          7351 => x"33",
          7352 => x"71",
          7353 => x"83",
          7354 => x"05",
          7355 => x"85",
          7356 => x"88",
          7357 => x"88",
          7358 => x"45",
          7359 => x"58",
          7360 => x"56",
          7361 => x"05",
          7362 => x"85",
          7363 => x"b9",
          7364 => x"17",
          7365 => x"85",
          7366 => x"8b",
          7367 => x"2b",
          7368 => x"86",
          7369 => x"15",
          7370 => x"2b",
          7371 => x"2a",
          7372 => x"48",
          7373 => x"41",
          7374 => x"05",
          7375 => x"87",
          7376 => x"b9",
          7377 => x"70",
          7378 => x"33",
          7379 => x"07",
          7380 => x"06",
          7381 => x"5f",
          7382 => x"7b",
          7383 => x"81",
          7384 => x"b9",
          7385 => x"1f",
          7386 => x"83",
          7387 => x"8b",
          7388 => x"2b",
          7389 => x"73",
          7390 => x"33",
          7391 => x"07",
          7392 => x"5e",
          7393 => x"43",
          7394 => x"76",
          7395 => x"81",
          7396 => x"b9",
          7397 => x"1f",
          7398 => x"12",
          7399 => x"2b",
          7400 => x"07",
          7401 => x"14",
          7402 => x"33",
          7403 => x"07",
          7404 => x"40",
          7405 => x"40",
          7406 => x"78",
          7407 => x"60",
          7408 => x"84",
          7409 => x"70",
          7410 => x"33",
          7411 => x"71",
          7412 => x"66",
          7413 => x"70",
          7414 => x"52",
          7415 => x"05",
          7416 => x"fe",
          7417 => x"84",
          7418 => x"1e",
          7419 => x"83",
          7420 => x"5c",
          7421 => x"39",
          7422 => x"0b",
          7423 => x"0c",
          7424 => x"84",
          7425 => x"82",
          7426 => x"7f",
          7427 => x"f4",
          7428 => x"ed",
          7429 => x"b8",
          7430 => x"76",
          7431 => x"81",
          7432 => x"b9",
          7433 => x"7f",
          7434 => x"81",
          7435 => x"34",
          7436 => x"08",
          7437 => x"15",
          7438 => x"87",
          7439 => x"b9",
          7440 => x"b9",
          7441 => x"05",
          7442 => x"07",
          7443 => x"ff",
          7444 => x"2a",
          7445 => x"5e",
          7446 => x"34",
          7447 => x"34",
          7448 => x"22",
          7449 => x"10",
          7450 => x"08",
          7451 => x"5c",
          7452 => x"1c",
          7453 => x"83",
          7454 => x"51",
          7455 => x"7f",
          7456 => x"39",
          7457 => x"87",
          7458 => x"8b",
          7459 => x"2b",
          7460 => x"84",
          7461 => x"1d",
          7462 => x"2b",
          7463 => x"2a",
          7464 => x"43",
          7465 => x"61",
          7466 => x"63",
          7467 => x"34",
          7468 => x"08",
          7469 => x"11",
          7470 => x"33",
          7471 => x"71",
          7472 => x"74",
          7473 => x"33",
          7474 => x"71",
          7475 => x"70",
          7476 => x"5f",
          7477 => x"56",
          7478 => x"64",
          7479 => x"78",
          7480 => x"34",
          7481 => x"08",
          7482 => x"81",
          7483 => x"88",
          7484 => x"ff",
          7485 => x"88",
          7486 => x"58",
          7487 => x"34",
          7488 => x"34",
          7489 => x"08",
          7490 => x"33",
          7491 => x"71",
          7492 => x"83",
          7493 => x"05",
          7494 => x"12",
          7495 => x"2b",
          7496 => x"2b",
          7497 => x"06",
          7498 => x"88",
          7499 => x"5d",
          7500 => x"5d",
          7501 => x"82",
          7502 => x"83",
          7503 => x"b9",
          7504 => x"1f",
          7505 => x"12",
          7506 => x"2b",
          7507 => x"07",
          7508 => x"33",
          7509 => x"71",
          7510 => x"81",
          7511 => x"70",
          7512 => x"5d",
          7513 => x"5a",
          7514 => x"60",
          7515 => x"81",
          7516 => x"83",
          7517 => x"5b",
          7518 => x"86",
          7519 => x"16",
          7520 => x"2b",
          7521 => x"07",
          7522 => x"18",
          7523 => x"33",
          7524 => x"07",
          7525 => x"5e",
          7526 => x"41",
          7527 => x"1e",
          7528 => x"1e",
          7529 => x"b8",
          7530 => x"84",
          7531 => x"12",
          7532 => x"2b",
          7533 => x"07",
          7534 => x"14",
          7535 => x"33",
          7536 => x"07",
          7537 => x"44",
          7538 => x"5a",
          7539 => x"7c",
          7540 => x"34",
          7541 => x"05",
          7542 => x"b8",
          7543 => x"33",
          7544 => x"71",
          7545 => x"81",
          7546 => x"70",
          7547 => x"5b",
          7548 => x"75",
          7549 => x"16",
          7550 => x"b8",
          7551 => x"70",
          7552 => x"33",
          7553 => x"71",
          7554 => x"74",
          7555 => x"81",
          7556 => x"88",
          7557 => x"83",
          7558 => x"f8",
          7559 => x"63",
          7560 => x"54",
          7561 => x"59",
          7562 => x"7f",
          7563 => x"7b",
          7564 => x"84",
          7565 => x"70",
          7566 => x"81",
          7567 => x"8b",
          7568 => x"2b",
          7569 => x"70",
          7570 => x"33",
          7571 => x"07",
          7572 => x"06",
          7573 => x"5d",
          7574 => x"5b",
          7575 => x"75",
          7576 => x"81",
          7577 => x"b9",
          7578 => x"1f",
          7579 => x"83",
          7580 => x"8b",
          7581 => x"2b",
          7582 => x"86",
          7583 => x"12",
          7584 => x"2b",
          7585 => x"07",
          7586 => x"14",
          7587 => x"33",
          7588 => x"07",
          7589 => x"59",
          7590 => x"5c",
          7591 => x"5d",
          7592 => x"77",
          7593 => x"79",
          7594 => x"84",
          7595 => x"70",
          7596 => x"33",
          7597 => x"71",
          7598 => x"83",
          7599 => x"05",
          7600 => x"87",
          7601 => x"88",
          7602 => x"88",
          7603 => x"5e",
          7604 => x"41",
          7605 => x"16",
          7606 => x"16",
          7607 => x"b8",
          7608 => x"33",
          7609 => x"71",
          7610 => x"81",
          7611 => x"70",
          7612 => x"5c",
          7613 => x"79",
          7614 => x"1a",
          7615 => x"b8",
          7616 => x"82",
          7617 => x"12",
          7618 => x"2b",
          7619 => x"07",
          7620 => x"33",
          7621 => x"71",
          7622 => x"70",
          7623 => x"5c",
          7624 => x"5a",
          7625 => x"79",
          7626 => x"1a",
          7627 => x"b8",
          7628 => x"70",
          7629 => x"33",
          7630 => x"71",
          7631 => x"74",
          7632 => x"33",
          7633 => x"71",
          7634 => x"70",
          7635 => x"5c",
          7636 => x"5a",
          7637 => x"82",
          7638 => x"83",
          7639 => x"b9",
          7640 => x"1f",
          7641 => x"83",
          7642 => x"88",
          7643 => x"57",
          7644 => x"83",
          7645 => x"5a",
          7646 => x"84",
          7647 => x"b6",
          7648 => x"b9",
          7649 => x"84",
          7650 => x"05",
          7651 => x"ff",
          7652 => x"44",
          7653 => x"39",
          7654 => x"87",
          7655 => x"8b",
          7656 => x"2b",
          7657 => x"84",
          7658 => x"1d",
          7659 => x"2b",
          7660 => x"2a",
          7661 => x"43",
          7662 => x"61",
          7663 => x"63",
          7664 => x"34",
          7665 => x"08",
          7666 => x"11",
          7667 => x"33",
          7668 => x"71",
          7669 => x"74",
          7670 => x"33",
          7671 => x"71",
          7672 => x"70",
          7673 => x"41",
          7674 => x"59",
          7675 => x"64",
          7676 => x"7a",
          7677 => x"34",
          7678 => x"08",
          7679 => x"81",
          7680 => x"88",
          7681 => x"ff",
          7682 => x"88",
          7683 => x"42",
          7684 => x"34",
          7685 => x"34",
          7686 => x"08",
          7687 => x"33",
          7688 => x"71",
          7689 => x"83",
          7690 => x"05",
          7691 => x"12",
          7692 => x"2b",
          7693 => x"2b",
          7694 => x"06",
          7695 => x"88",
          7696 => x"5c",
          7697 => x"45",
          7698 => x"82",
          7699 => x"83",
          7700 => x"b9",
          7701 => x"1f",
          7702 => x"12",
          7703 => x"2b",
          7704 => x"07",
          7705 => x"33",
          7706 => x"71",
          7707 => x"81",
          7708 => x"70",
          7709 => x"5f",
          7710 => x"59",
          7711 => x"7d",
          7712 => x"1e",
          7713 => x"ff",
          7714 => x"f3",
          7715 => x"60",
          7716 => x"a1",
          7717 => x"c8",
          7718 => x"b9",
          7719 => x"2e",
          7720 => x"53",
          7721 => x"b9",
          7722 => x"fe",
          7723 => x"73",
          7724 => x"3f",
          7725 => x"7b",
          7726 => x"38",
          7727 => x"f9",
          7728 => x"7a",
          7729 => x"b8",
          7730 => x"76",
          7731 => x"38",
          7732 => x"8a",
          7733 => x"b9",
          7734 => x"3d",
          7735 => x"51",
          7736 => x"84",
          7737 => x"54",
          7738 => x"08",
          7739 => x"38",
          7740 => x"52",
          7741 => x"08",
          7742 => x"85",
          7743 => x"b9",
          7744 => x"3d",
          7745 => x"ff",
          7746 => x"b9",
          7747 => x"80",
          7748 => x"b4",
          7749 => x"80",
          7750 => x"84",
          7751 => x"fe",
          7752 => x"84",
          7753 => x"55",
          7754 => x"81",
          7755 => x"34",
          7756 => x"08",
          7757 => x"15",
          7758 => x"85",
          7759 => x"b9",
          7760 => x"76",
          7761 => x"81",
          7762 => x"34",
          7763 => x"08",
          7764 => x"22",
          7765 => x"80",
          7766 => x"83",
          7767 => x"70",
          7768 => x"51",
          7769 => x"88",
          7770 => x"89",
          7771 => x"b9",
          7772 => x"10",
          7773 => x"b9",
          7774 => x"f8",
          7775 => x"76",
          7776 => x"81",
          7777 => x"34",
          7778 => x"80",
          7779 => x"38",
          7780 => x"ff",
          7781 => x"8f",
          7782 => x"81",
          7783 => x"26",
          7784 => x"b9",
          7785 => x"52",
          7786 => x"c8",
          7787 => x"0d",
          7788 => x"0d",
          7789 => x"33",
          7790 => x"71",
          7791 => x"38",
          7792 => x"bb",
          7793 => x"c8",
          7794 => x"06",
          7795 => x"38",
          7796 => x"c4",
          7797 => x"b9",
          7798 => x"53",
          7799 => x"c8",
          7800 => x"0d",
          7801 => x"0d",
          7802 => x"02",
          7803 => x"05",
          7804 => x"57",
          7805 => x"76",
          7806 => x"38",
          7807 => x"17",
          7808 => x"81",
          7809 => x"55",
          7810 => x"73",
          7811 => x"87",
          7812 => x"0c",
          7813 => x"52",
          7814 => x"ca",
          7815 => x"c8",
          7816 => x"06",
          7817 => x"2e",
          7818 => x"c0",
          7819 => x"54",
          7820 => x"79",
          7821 => x"38",
          7822 => x"80",
          7823 => x"80",
          7824 => x"81",
          7825 => x"74",
          7826 => x"0c",
          7827 => x"04",
          7828 => x"81",
          7829 => x"ff",
          7830 => x"56",
          7831 => x"ff",
          7832 => x"39",
          7833 => x"7c",
          7834 => x"8c",
          7835 => x"33",
          7836 => x"59",
          7837 => x"74",
          7838 => x"84",
          7839 => x"33",
          7840 => x"06",
          7841 => x"73",
          7842 => x"58",
          7843 => x"c0",
          7844 => x"78",
          7845 => x"76",
          7846 => x"3f",
          7847 => x"08",
          7848 => x"55",
          7849 => x"a7",
          7850 => x"98",
          7851 => x"73",
          7852 => x"78",
          7853 => x"74",
          7854 => x"06",
          7855 => x"2e",
          7856 => x"54",
          7857 => x"84",
          7858 => x"8b",
          7859 => x"84",
          7860 => x"19",
          7861 => x"06",
          7862 => x"79",
          7863 => x"ac",
          7864 => x"fc",
          7865 => x"02",
          7866 => x"05",
          7867 => x"05",
          7868 => x"53",
          7869 => x"53",
          7870 => x"87",
          7871 => x"c4",
          7872 => x"72",
          7873 => x"83",
          7874 => x"38",
          7875 => x"c0",
          7876 => x"81",
          7877 => x"2e",
          7878 => x"71",
          7879 => x"70",
          7880 => x"38",
          7881 => x"84",
          7882 => x"86",
          7883 => x"88",
          7884 => x"0c",
          7885 => x"c8",
          7886 => x"0d",
          7887 => x"75",
          7888 => x"84",
          7889 => x"86",
          7890 => x"71",
          7891 => x"c0",
          7892 => x"53",
          7893 => x"38",
          7894 => x"81",
          7895 => x"51",
          7896 => x"2e",
          7897 => x"c0",
          7898 => x"55",
          7899 => x"87",
          7900 => x"08",
          7901 => x"38",
          7902 => x"87",
          7903 => x"14",
          7904 => x"82",
          7905 => x"80",
          7906 => x"38",
          7907 => x"06",
          7908 => x"38",
          7909 => x"f6",
          7910 => x"58",
          7911 => x"19",
          7912 => x"56",
          7913 => x"2e",
          7914 => x"a8",
          7915 => x"56",
          7916 => x"81",
          7917 => x"53",
          7918 => x"18",
          7919 => x"a3",
          7920 => x"c8",
          7921 => x"83",
          7922 => x"78",
          7923 => x"0c",
          7924 => x"04",
          7925 => x"18",
          7926 => x"18",
          7927 => x"19",
          7928 => x"fc",
          7929 => x"59",
          7930 => x"08",
          7931 => x"81",
          7932 => x"84",
          7933 => x"83",
          7934 => x"18",
          7935 => x"1a",
          7936 => x"1a",
          7937 => x"c8",
          7938 => x"56",
          7939 => x"27",
          7940 => x"82",
          7941 => x"74",
          7942 => x"81",
          7943 => x"38",
          7944 => x"1b",
          7945 => x"81",
          7946 => x"fc",
          7947 => x"78",
          7948 => x"75",
          7949 => x"81",
          7950 => x"38",
          7951 => x"57",
          7952 => x"09",
          7953 => x"ee",
          7954 => x"5a",
          7955 => x"56",
          7956 => x"70",
          7957 => x"34",
          7958 => x"76",
          7959 => x"d5",
          7960 => x"19",
          7961 => x"0b",
          7962 => x"34",
          7963 => x"34",
          7964 => x"b9",
          7965 => x"e1",
          7966 => x"34",
          7967 => x"bb",
          7968 => x"f2",
          7969 => x"19",
          7970 => x"0b",
          7971 => x"34",
          7972 => x"84",
          7973 => x"80",
          7974 => x"9f",
          7975 => x"18",
          7976 => x"84",
          7977 => x"74",
          7978 => x"7a",
          7979 => x"34",
          7980 => x"56",
          7981 => x"19",
          7982 => x"2a",
          7983 => x"a3",
          7984 => x"18",
          7985 => x"84",
          7986 => x"7a",
          7987 => x"74",
          7988 => x"34",
          7989 => x"56",
          7990 => x"19",
          7991 => x"2a",
          7992 => x"a7",
          7993 => x"18",
          7994 => x"70",
          7995 => x"5b",
          7996 => x"53",
          7997 => x"18",
          7998 => x"e8",
          7999 => x"19",
          8000 => x"80",
          8001 => x"33",
          8002 => x"3f",
          8003 => x"08",
          8004 => x"b7",
          8005 => x"39",
          8006 => x"60",
          8007 => x"59",
          8008 => x"76",
          8009 => x"9c",
          8010 => x"26",
          8011 => x"58",
          8012 => x"c8",
          8013 => x"0d",
          8014 => x"33",
          8015 => x"82",
          8016 => x"38",
          8017 => x"82",
          8018 => x"81",
          8019 => x"06",
          8020 => x"81",
          8021 => x"89",
          8022 => x"08",
          8023 => x"80",
          8024 => x"08",
          8025 => x"38",
          8026 => x"5c",
          8027 => x"09",
          8028 => x"de",
          8029 => x"78",
          8030 => x"52",
          8031 => x"51",
          8032 => x"84",
          8033 => x"80",
          8034 => x"ff",
          8035 => x"78",
          8036 => x"7a",
          8037 => x"79",
          8038 => x"17",
          8039 => x"81",
          8040 => x"2a",
          8041 => x"05",
          8042 => x"59",
          8043 => x"79",
          8044 => x"80",
          8045 => x"33",
          8046 => x"5d",
          8047 => x"09",
          8048 => x"b5",
          8049 => x"78",
          8050 => x"52",
          8051 => x"51",
          8052 => x"84",
          8053 => x"80",
          8054 => x"ff",
          8055 => x"78",
          8056 => x"79",
          8057 => x"7a",
          8058 => x"17",
          8059 => x"70",
          8060 => x"07",
          8061 => x"71",
          8062 => x"5d",
          8063 => x"79",
          8064 => x"76",
          8065 => x"84",
          8066 => x"8f",
          8067 => x"75",
          8068 => x"18",
          8069 => x"b4",
          8070 => x"2e",
          8071 => x"0b",
          8072 => x"71",
          8073 => x"7b",
          8074 => x"81",
          8075 => x"38",
          8076 => x"53",
          8077 => x"81",
          8078 => x"f7",
          8079 => x"b9",
          8080 => x"2e",
          8081 => x"59",
          8082 => x"b4",
          8083 => x"fd",
          8084 => x"10",
          8085 => x"77",
          8086 => x"81",
          8087 => x"33",
          8088 => x"07",
          8089 => x"0c",
          8090 => x"3d",
          8091 => x"83",
          8092 => x"06",
          8093 => x"75",
          8094 => x"18",
          8095 => x"b4",
          8096 => x"2e",
          8097 => x"0b",
          8098 => x"71",
          8099 => x"7c",
          8100 => x"81",
          8101 => x"38",
          8102 => x"53",
          8103 => x"81",
          8104 => x"f6",
          8105 => x"b9",
          8106 => x"2e",
          8107 => x"59",
          8108 => x"b4",
          8109 => x"fc",
          8110 => x"82",
          8111 => x"06",
          8112 => x"05",
          8113 => x"82",
          8114 => x"90",
          8115 => x"2b",
          8116 => x"33",
          8117 => x"88",
          8118 => x"71",
          8119 => x"fe",
          8120 => x"84",
          8121 => x"41",
          8122 => x"5a",
          8123 => x"0d",
          8124 => x"b4",
          8125 => x"b8",
          8126 => x"81",
          8127 => x"5c",
          8128 => x"81",
          8129 => x"c8",
          8130 => x"09",
          8131 => x"be",
          8132 => x"c8",
          8133 => x"34",
          8134 => x"a8",
          8135 => x"84",
          8136 => x"5b",
          8137 => x"18",
          8138 => x"84",
          8139 => x"33",
          8140 => x"2e",
          8141 => x"fd",
          8142 => x"54",
          8143 => x"a0",
          8144 => x"53",
          8145 => x"17",
          8146 => x"98",
          8147 => x"fd",
          8148 => x"54",
          8149 => x"53",
          8150 => x"53",
          8151 => x"52",
          8152 => x"3f",
          8153 => x"08",
          8154 => x"81",
          8155 => x"38",
          8156 => x"08",
          8157 => x"b4",
          8158 => x"18",
          8159 => x"7c",
          8160 => x"27",
          8161 => x"17",
          8162 => x"82",
          8163 => x"38",
          8164 => x"08",
          8165 => x"39",
          8166 => x"17",
          8167 => x"17",
          8168 => x"18",
          8169 => x"f5",
          8170 => x"5a",
          8171 => x"08",
          8172 => x"81",
          8173 => x"38",
          8174 => x"08",
          8175 => x"b4",
          8176 => x"18",
          8177 => x"b9",
          8178 => x"5e",
          8179 => x"08",
          8180 => x"38",
          8181 => x"55",
          8182 => x"09",
          8183 => x"b8",
          8184 => x"b4",
          8185 => x"18",
          8186 => x"7b",
          8187 => x"33",
          8188 => x"3f",
          8189 => x"a0",
          8190 => x"b4",
          8191 => x"b8",
          8192 => x"81",
          8193 => x"5e",
          8194 => x"81",
          8195 => x"c8",
          8196 => x"09",
          8197 => x"cb",
          8198 => x"c8",
          8199 => x"34",
          8200 => x"a8",
          8201 => x"84",
          8202 => x"5b",
          8203 => x"18",
          8204 => x"91",
          8205 => x"33",
          8206 => x"2e",
          8207 => x"fb",
          8208 => x"54",
          8209 => x"a0",
          8210 => x"53",
          8211 => x"17",
          8212 => x"90",
          8213 => x"fa",
          8214 => x"54",
          8215 => x"a0",
          8216 => x"53",
          8217 => x"17",
          8218 => x"f8",
          8219 => x"39",
          8220 => x"f9",
          8221 => x"9f",
          8222 => x"0d",
          8223 => x"5d",
          8224 => x"58",
          8225 => x"9c",
          8226 => x"1a",
          8227 => x"38",
          8228 => x"74",
          8229 => x"38",
          8230 => x"81",
          8231 => x"81",
          8232 => x"38",
          8233 => x"c8",
          8234 => x"0d",
          8235 => x"2a",
          8236 => x"05",
          8237 => x"b4",
          8238 => x"5c",
          8239 => x"86",
          8240 => x"19",
          8241 => x"5d",
          8242 => x"09",
          8243 => x"fa",
          8244 => x"77",
          8245 => x"52",
          8246 => x"51",
          8247 => x"84",
          8248 => x"80",
          8249 => x"ff",
          8250 => x"77",
          8251 => x"79",
          8252 => x"b0",
          8253 => x"83",
          8254 => x"05",
          8255 => x"ff",
          8256 => x"76",
          8257 => x"76",
          8258 => x"79",
          8259 => x"81",
          8260 => x"34",
          8261 => x"c8",
          8262 => x"0d",
          8263 => x"2e",
          8264 => x"fe",
          8265 => x"87",
          8266 => x"08",
          8267 => x"0b",
          8268 => x"58",
          8269 => x"2e",
          8270 => x"83",
          8271 => x"5b",
          8272 => x"2e",
          8273 => x"84",
          8274 => x"54",
          8275 => x"19",
          8276 => x"33",
          8277 => x"3f",
          8278 => x"08",
          8279 => x"38",
          8280 => x"5a",
          8281 => x"0c",
          8282 => x"fe",
          8283 => x"82",
          8284 => x"06",
          8285 => x"11",
          8286 => x"70",
          8287 => x"0a",
          8288 => x"0a",
          8289 => x"57",
          8290 => x"7d",
          8291 => x"2a",
          8292 => x"1d",
          8293 => x"2a",
          8294 => x"1d",
          8295 => x"2a",
          8296 => x"1d",
          8297 => x"83",
          8298 => x"e8",
          8299 => x"2a",
          8300 => x"2a",
          8301 => x"05",
          8302 => x"59",
          8303 => x"78",
          8304 => x"80",
          8305 => x"33",
          8306 => x"5d",
          8307 => x"09",
          8308 => x"d4",
          8309 => x"77",
          8310 => x"52",
          8311 => x"51",
          8312 => x"84",
          8313 => x"80",
          8314 => x"ff",
          8315 => x"77",
          8316 => x"7b",
          8317 => x"ac",
          8318 => x"ff",
          8319 => x"05",
          8320 => x"81",
          8321 => x"57",
          8322 => x"80",
          8323 => x"7a",
          8324 => x"f0",
          8325 => x"8f",
          8326 => x"56",
          8327 => x"34",
          8328 => x"1a",
          8329 => x"2a",
          8330 => x"05",
          8331 => x"b4",
          8332 => x"5f",
          8333 => x"83",
          8334 => x"54",
          8335 => x"19",
          8336 => x"1a",
          8337 => x"f0",
          8338 => x"58",
          8339 => x"08",
          8340 => x"81",
          8341 => x"38",
          8342 => x"08",
          8343 => x"b4",
          8344 => x"a8",
          8345 => x"a0",
          8346 => x"b9",
          8347 => x"5c",
          8348 => x"7a",
          8349 => x"82",
          8350 => x"74",
          8351 => x"e4",
          8352 => x"75",
          8353 => x"81",
          8354 => x"ee",
          8355 => x"b9",
          8356 => x"2e",
          8357 => x"56",
          8358 => x"b4",
          8359 => x"fc",
          8360 => x"83",
          8361 => x"b8",
          8362 => x"2a",
          8363 => x"8f",
          8364 => x"2a",
          8365 => x"f0",
          8366 => x"06",
          8367 => x"74",
          8368 => x"0b",
          8369 => x"fc",
          8370 => x"54",
          8371 => x"19",
          8372 => x"1a",
          8373 => x"ef",
          8374 => x"5a",
          8375 => x"08",
          8376 => x"81",
          8377 => x"38",
          8378 => x"08",
          8379 => x"b4",
          8380 => x"a8",
          8381 => x"a0",
          8382 => x"b9",
          8383 => x"59",
          8384 => x"77",
          8385 => x"38",
          8386 => x"55",
          8387 => x"09",
          8388 => x"bd",
          8389 => x"76",
          8390 => x"52",
          8391 => x"51",
          8392 => x"7b",
          8393 => x"39",
          8394 => x"53",
          8395 => x"53",
          8396 => x"52",
          8397 => x"3f",
          8398 => x"b9",
          8399 => x"2e",
          8400 => x"fd",
          8401 => x"b9",
          8402 => x"1a",
          8403 => x"08",
          8404 => x"08",
          8405 => x"08",
          8406 => x"08",
          8407 => x"5f",
          8408 => x"fc",
          8409 => x"19",
          8410 => x"82",
          8411 => x"06",
          8412 => x"81",
          8413 => x"53",
          8414 => x"19",
          8415 => x"e4",
          8416 => x"fc",
          8417 => x"54",
          8418 => x"19",
          8419 => x"1a",
          8420 => x"ed",
          8421 => x"5a",
          8422 => x"08",
          8423 => x"81",
          8424 => x"38",
          8425 => x"08",
          8426 => x"b4",
          8427 => x"a8",
          8428 => x"a0",
          8429 => x"b9",
          8430 => x"5f",
          8431 => x"7d",
          8432 => x"38",
          8433 => x"55",
          8434 => x"09",
          8435 => x"fa",
          8436 => x"7c",
          8437 => x"52",
          8438 => x"51",
          8439 => x"7b",
          8440 => x"39",
          8441 => x"1c",
          8442 => x"81",
          8443 => x"ec",
          8444 => x"58",
          8445 => x"7b",
          8446 => x"fe",
          8447 => x"7c",
          8448 => x"06",
          8449 => x"76",
          8450 => x"76",
          8451 => x"79",
          8452 => x"f9",
          8453 => x"58",
          8454 => x"7b",
          8455 => x"83",
          8456 => x"05",
          8457 => x"11",
          8458 => x"2b",
          8459 => x"7f",
          8460 => x"07",
          8461 => x"5d",
          8462 => x"34",
          8463 => x"56",
          8464 => x"34",
          8465 => x"5a",
          8466 => x"34",
          8467 => x"5b",
          8468 => x"34",
          8469 => x"f6",
          8470 => x"7e",
          8471 => x"5c",
          8472 => x"8a",
          8473 => x"08",
          8474 => x"2e",
          8475 => x"76",
          8476 => x"27",
          8477 => x"94",
          8478 => x"56",
          8479 => x"2e",
          8480 => x"76",
          8481 => x"93",
          8482 => x"81",
          8483 => x"19",
          8484 => x"89",
          8485 => x"75",
          8486 => x"b2",
          8487 => x"79",
          8488 => x"3f",
          8489 => x"08",
          8490 => x"d0",
          8491 => x"84",
          8492 => x"81",
          8493 => x"84",
          8494 => x"09",
          8495 => x"72",
          8496 => x"70",
          8497 => x"51",
          8498 => x"82",
          8499 => x"77",
          8500 => x"06",
          8501 => x"73",
          8502 => x"b9",
          8503 => x"3d",
          8504 => x"57",
          8505 => x"84",
          8506 => x"58",
          8507 => x"52",
          8508 => x"a4",
          8509 => x"74",
          8510 => x"08",
          8511 => x"84",
          8512 => x"55",
          8513 => x"08",
          8514 => x"38",
          8515 => x"84",
          8516 => x"26",
          8517 => x"57",
          8518 => x"81",
          8519 => x"19",
          8520 => x"83",
          8521 => x"75",
          8522 => x"ef",
          8523 => x"58",
          8524 => x"08",
          8525 => x"a0",
          8526 => x"c8",
          8527 => x"30",
          8528 => x"80",
          8529 => x"07",
          8530 => x"08",
          8531 => x"55",
          8532 => x"85",
          8533 => x"c8",
          8534 => x"9a",
          8535 => x"08",
          8536 => x"27",
          8537 => x"73",
          8538 => x"27",
          8539 => x"73",
          8540 => x"fe",
          8541 => x"80",
          8542 => x"38",
          8543 => x"52",
          8544 => x"f5",
          8545 => x"c8",
          8546 => x"c8",
          8547 => x"84",
          8548 => x"07",
          8549 => x"58",
          8550 => x"c4",
          8551 => x"e3",
          8552 => x"1a",
          8553 => x"08",
          8554 => x"1a",
          8555 => x"74",
          8556 => x"38",
          8557 => x"1a",
          8558 => x"33",
          8559 => x"79",
          8560 => x"75",
          8561 => x"b9",
          8562 => x"3d",
          8563 => x"0b",
          8564 => x"0c",
          8565 => x"04",
          8566 => x"08",
          8567 => x"39",
          8568 => x"ff",
          8569 => x"53",
          8570 => x"51",
          8571 => x"84",
          8572 => x"55",
          8573 => x"84",
          8574 => x"84",
          8575 => x"8c",
          8576 => x"ff",
          8577 => x"2e",
          8578 => x"81",
          8579 => x"39",
          8580 => x"7a",
          8581 => x"59",
          8582 => x"f0",
          8583 => x"80",
          8584 => x"9f",
          8585 => x"80",
          8586 => x"90",
          8587 => x"18",
          8588 => x"80",
          8589 => x"33",
          8590 => x"26",
          8591 => x"73",
          8592 => x"82",
          8593 => x"22",
          8594 => x"79",
          8595 => x"ac",
          8596 => x"19",
          8597 => x"19",
          8598 => x"08",
          8599 => x"72",
          8600 => x"38",
          8601 => x"13",
          8602 => x"73",
          8603 => x"17",
          8604 => x"19",
          8605 => x"75",
          8606 => x"0c",
          8607 => x"04",
          8608 => x"b9",
          8609 => x"3d",
          8610 => x"17",
          8611 => x"80",
          8612 => x"38",
          8613 => x"70",
          8614 => x"59",
          8615 => x"a5",
          8616 => x"08",
          8617 => x"fe",
          8618 => x"80",
          8619 => x"27",
          8620 => x"17",
          8621 => x"29",
          8622 => x"05",
          8623 => x"98",
          8624 => x"91",
          8625 => x"77",
          8626 => x"3f",
          8627 => x"08",
          8628 => x"c8",
          8629 => x"a4",
          8630 => x"84",
          8631 => x"27",
          8632 => x"9c",
          8633 => x"84",
          8634 => x"73",
          8635 => x"38",
          8636 => x"54",
          8637 => x"cd",
          8638 => x"39",
          8639 => x"b9",
          8640 => x"3d",
          8641 => x"3d",
          8642 => x"08",
          8643 => x"a0",
          8644 => x"57",
          8645 => x"7a",
          8646 => x"80",
          8647 => x"0c",
          8648 => x"55",
          8649 => x"80",
          8650 => x"79",
          8651 => x"5b",
          8652 => x"81",
          8653 => x"08",
          8654 => x"a9",
          8655 => x"2a",
          8656 => x"57",
          8657 => x"27",
          8658 => x"77",
          8659 => x"79",
          8660 => x"78",
          8661 => x"9c",
          8662 => x"56",
          8663 => x"c8",
          8664 => x"0d",
          8665 => x"18",
          8666 => x"22",
          8667 => x"89",
          8668 => x"7b",
          8669 => x"52",
          8670 => x"9c",
          8671 => x"c8",
          8672 => x"56",
          8673 => x"b9",
          8674 => x"d0",
          8675 => x"84",
          8676 => x"ff",
          8677 => x"9c",
          8678 => x"b9",
          8679 => x"82",
          8680 => x"80",
          8681 => x"38",
          8682 => x"52",
          8683 => x"a7",
          8684 => x"c8",
          8685 => x"56",
          8686 => x"08",
          8687 => x"9c",
          8688 => x"84",
          8689 => x"81",
          8690 => x"38",
          8691 => x"b9",
          8692 => x"2e",
          8693 => x"84",
          8694 => x"83",
          8695 => x"58",
          8696 => x"38",
          8697 => x"1a",
          8698 => x"59",
          8699 => x"75",
          8700 => x"38",
          8701 => x"76",
          8702 => x"1b",
          8703 => x"5e",
          8704 => x"0c",
          8705 => x"84",
          8706 => x"55",
          8707 => x"81",
          8708 => x"ff",
          8709 => x"f4",
          8710 => x"8a",
          8711 => x"75",
          8712 => x"80",
          8713 => x"75",
          8714 => x"52",
          8715 => x"51",
          8716 => x"84",
          8717 => x"80",
          8718 => x"16",
          8719 => x"7a",
          8720 => x"84",
          8721 => x"c8",
          8722 => x"0d",
          8723 => x"b4",
          8724 => x"b8",
          8725 => x"81",
          8726 => x"56",
          8727 => x"84",
          8728 => x"80",
          8729 => x"b9",
          8730 => x"1a",
          8731 => x"08",
          8732 => x"31",
          8733 => x"1a",
          8734 => x"e8",
          8735 => x"33",
          8736 => x"2e",
          8737 => x"fe",
          8738 => x"54",
          8739 => x"a0",
          8740 => x"53",
          8741 => x"19",
          8742 => x"c8",
          8743 => x"39",
          8744 => x"55",
          8745 => x"ff",
          8746 => x"76",
          8747 => x"06",
          8748 => x"94",
          8749 => x"1d",
          8750 => x"fe",
          8751 => x"80",
          8752 => x"27",
          8753 => x"8a",
          8754 => x"71",
          8755 => x"08",
          8756 => x"0c",
          8757 => x"39",
          8758 => x"b9",
          8759 => x"3d",
          8760 => x"3d",
          8761 => x"41",
          8762 => x"08",
          8763 => x"ff",
          8764 => x"08",
          8765 => x"75",
          8766 => x"d2",
          8767 => x"5f",
          8768 => x"58",
          8769 => x"76",
          8770 => x"38",
          8771 => x"78",
          8772 => x"78",
          8773 => x"06",
          8774 => x"81",
          8775 => x"b8",
          8776 => x"19",
          8777 => x"bd",
          8778 => x"c8",
          8779 => x"85",
          8780 => x"81",
          8781 => x"1a",
          8782 => x"76",
          8783 => x"9c",
          8784 => x"33",
          8785 => x"80",
          8786 => x"38",
          8787 => x"bf",
          8788 => x"ff",
          8789 => x"60",
          8790 => x"76",
          8791 => x"70",
          8792 => x"32",
          8793 => x"80",
          8794 => x"25",
          8795 => x"45",
          8796 => x"93",
          8797 => x"df",
          8798 => x"61",
          8799 => x"bf",
          8800 => x"2e",
          8801 => x"81",
          8802 => x"52",
          8803 => x"f6",
          8804 => x"c8",
          8805 => x"b9",
          8806 => x"b2",
          8807 => x"08",
          8808 => x"dc",
          8809 => x"b9",
          8810 => x"3d",
          8811 => x"54",
          8812 => x"53",
          8813 => x"19",
          8814 => x"a8",
          8815 => x"84",
          8816 => x"78",
          8817 => x"06",
          8818 => x"84",
          8819 => x"83",
          8820 => x"19",
          8821 => x"08",
          8822 => x"c8",
          8823 => x"7a",
          8824 => x"27",
          8825 => x"82",
          8826 => x"60",
          8827 => x"81",
          8828 => x"38",
          8829 => x"19",
          8830 => x"08",
          8831 => x"52",
          8832 => x"51",
          8833 => x"77",
          8834 => x"39",
          8835 => x"09",
          8836 => x"e7",
          8837 => x"2a",
          8838 => x"7a",
          8839 => x"38",
          8840 => x"77",
          8841 => x"70",
          8842 => x"7f",
          8843 => x"59",
          8844 => x"7d",
          8845 => x"81",
          8846 => x"5d",
          8847 => x"81",
          8848 => x"2e",
          8849 => x"fe",
          8850 => x"39",
          8851 => x"0b",
          8852 => x"7a",
          8853 => x"0c",
          8854 => x"04",
          8855 => x"df",
          8856 => x"33",
          8857 => x"2e",
          8858 => x"cb",
          8859 => x"08",
          8860 => x"9a",
          8861 => x"88",
          8862 => x"56",
          8863 => x"b7",
          8864 => x"70",
          8865 => x"8d",
          8866 => x"51",
          8867 => x"58",
          8868 => x"c8",
          8869 => x"05",
          8870 => x"71",
          8871 => x"2b",
          8872 => x"56",
          8873 => x"80",
          8874 => x"81",
          8875 => x"87",
          8876 => x"61",
          8877 => x"42",
          8878 => x"81",
          8879 => x"17",
          8880 => x"27",
          8881 => x"33",
          8882 => x"81",
          8883 => x"77",
          8884 => x"38",
          8885 => x"26",
          8886 => x"79",
          8887 => x"43",
          8888 => x"ff",
          8889 => x"ff",
          8890 => x"fd",
          8891 => x"83",
          8892 => x"ca",
          8893 => x"55",
          8894 => x"7c",
          8895 => x"55",
          8896 => x"81",
          8897 => x"80",
          8898 => x"70",
          8899 => x"33",
          8900 => x"70",
          8901 => x"ff",
          8902 => x"59",
          8903 => x"74",
          8904 => x"81",
          8905 => x"ac",
          8906 => x"84",
          8907 => x"94",
          8908 => x"ef",
          8909 => x"70",
          8910 => x"80",
          8911 => x"f5",
          8912 => x"b9",
          8913 => x"84",
          8914 => x"82",
          8915 => x"ff",
          8916 => x"ff",
          8917 => x"0c",
          8918 => x"98",
          8919 => x"80",
          8920 => x"08",
          8921 => x"cc",
          8922 => x"33",
          8923 => x"74",
          8924 => x"81",
          8925 => x"38",
          8926 => x"53",
          8927 => x"81",
          8928 => x"dc",
          8929 => x"b9",
          8930 => x"2e",
          8931 => x"56",
          8932 => x"b4",
          8933 => x"5a",
          8934 => x"38",
          8935 => x"70",
          8936 => x"76",
          8937 => x"99",
          8938 => x"33",
          8939 => x"81",
          8940 => x"58",
          8941 => x"34",
          8942 => x"2e",
          8943 => x"75",
          8944 => x"06",
          8945 => x"2e",
          8946 => x"74",
          8947 => x"75",
          8948 => x"e5",
          8949 => x"38",
          8950 => x"58",
          8951 => x"81",
          8952 => x"80",
          8953 => x"70",
          8954 => x"33",
          8955 => x"70",
          8956 => x"ff",
          8957 => x"5d",
          8958 => x"74",
          8959 => x"cd",
          8960 => x"33",
          8961 => x"76",
          8962 => x"0b",
          8963 => x"57",
          8964 => x"05",
          8965 => x"70",
          8966 => x"33",
          8967 => x"ff",
          8968 => x"42",
          8969 => x"2e",
          8970 => x"75",
          8971 => x"38",
          8972 => x"ff",
          8973 => x"0c",
          8974 => x"51",
          8975 => x"84",
          8976 => x"5a",
          8977 => x"08",
          8978 => x"8f",
          8979 => x"b9",
          8980 => x"3d",
          8981 => x"54",
          8982 => x"53",
          8983 => x"1b",
          8984 => x"80",
          8985 => x"84",
          8986 => x"78",
          8987 => x"06",
          8988 => x"84",
          8989 => x"83",
          8990 => x"1b",
          8991 => x"08",
          8992 => x"c8",
          8993 => x"78",
          8994 => x"27",
          8995 => x"82",
          8996 => x"79",
          8997 => x"81",
          8998 => x"38",
          8999 => x"1b",
          9000 => x"08",
          9001 => x"52",
          9002 => x"51",
          9003 => x"77",
          9004 => x"39",
          9005 => x"e4",
          9006 => x"33",
          9007 => x"81",
          9008 => x"60",
          9009 => x"76",
          9010 => x"06",
          9011 => x"2e",
          9012 => x"19",
          9013 => x"bf",
          9014 => x"1f",
          9015 => x"05",
          9016 => x"5f",
          9017 => x"af",
          9018 => x"55",
          9019 => x"52",
          9020 => x"92",
          9021 => x"c8",
          9022 => x"b9",
          9023 => x"2e",
          9024 => x"fe",
          9025 => x"80",
          9026 => x"38",
          9027 => x"ff",
          9028 => x"0c",
          9029 => x"8d",
          9030 => x"7e",
          9031 => x"81",
          9032 => x"8c",
          9033 => x"1a",
          9034 => x"33",
          9035 => x"07",
          9036 => x"76",
          9037 => x"78",
          9038 => x"06",
          9039 => x"05",
          9040 => x"77",
          9041 => x"e5",
          9042 => x"79",
          9043 => x"33",
          9044 => x"88",
          9045 => x"42",
          9046 => x"2e",
          9047 => x"79",
          9048 => x"ff",
          9049 => x"51",
          9050 => x"3f",
          9051 => x"08",
          9052 => x"05",
          9053 => x"43",
          9054 => x"56",
          9055 => x"3f",
          9056 => x"c8",
          9057 => x"81",
          9058 => x"38",
          9059 => x"18",
          9060 => x"27",
          9061 => x"78",
          9062 => x"2a",
          9063 => x"59",
          9064 => x"92",
          9065 => x"2e",
          9066 => x"10",
          9067 => x"22",
          9068 => x"fe",
          9069 => x"1d",
          9070 => x"06",
          9071 => x"ae",
          9072 => x"84",
          9073 => x"93",
          9074 => x"76",
          9075 => x"2e",
          9076 => x"81",
          9077 => x"94",
          9078 => x"0d",
          9079 => x"70",
          9080 => x"81",
          9081 => x"5a",
          9082 => x"56",
          9083 => x"38",
          9084 => x"08",
          9085 => x"57",
          9086 => x"2e",
          9087 => x"1d",
          9088 => x"70",
          9089 => x"5d",
          9090 => x"95",
          9091 => x"5b",
          9092 => x"7b",
          9093 => x"75",
          9094 => x"57",
          9095 => x"81",
          9096 => x"ff",
          9097 => x"ef",
          9098 => x"db",
          9099 => x"81",
          9100 => x"76",
          9101 => x"aa",
          9102 => x"0b",
          9103 => x"81",
          9104 => x"40",
          9105 => x"08",
          9106 => x"8b",
          9107 => x"57",
          9108 => x"81",
          9109 => x"76",
          9110 => x"58",
          9111 => x"55",
          9112 => x"85",
          9113 => x"c2",
          9114 => x"22",
          9115 => x"80",
          9116 => x"74",
          9117 => x"56",
          9118 => x"81",
          9119 => x"07",
          9120 => x"70",
          9121 => x"06",
          9122 => x"81",
          9123 => x"56",
          9124 => x"2e",
          9125 => x"84",
          9126 => x"57",
          9127 => x"77",
          9128 => x"38",
          9129 => x"74",
          9130 => x"02",
          9131 => x"cf",
          9132 => x"76",
          9133 => x"06",
          9134 => x"27",
          9135 => x"15",
          9136 => x"34",
          9137 => x"19",
          9138 => x"59",
          9139 => x"e3",
          9140 => x"59",
          9141 => x"34",
          9142 => x"56",
          9143 => x"a0",
          9144 => x"55",
          9145 => x"98",
          9146 => x"56",
          9147 => x"88",
          9148 => x"1a",
          9149 => x"57",
          9150 => x"09",
          9151 => x"38",
          9152 => x"a0",
          9153 => x"26",
          9154 => x"3d",
          9155 => x"05",
          9156 => x"33",
          9157 => x"74",
          9158 => x"76",
          9159 => x"38",
          9160 => x"8f",
          9161 => x"c8",
          9162 => x"81",
          9163 => x"e3",
          9164 => x"91",
          9165 => x"7a",
          9166 => x"82",
          9167 => x"b9",
          9168 => x"84",
          9169 => x"84",
          9170 => x"06",
          9171 => x"02",
          9172 => x"33",
          9173 => x"7d",
          9174 => x"05",
          9175 => x"33",
          9176 => x"81",
          9177 => x"5f",
          9178 => x"80",
          9179 => x"8d",
          9180 => x"51",
          9181 => x"3f",
          9182 => x"08",
          9183 => x"52",
          9184 => x"8c",
          9185 => x"c8",
          9186 => x"b9",
          9187 => x"82",
          9188 => x"c8",
          9189 => x"5e",
          9190 => x"08",
          9191 => x"b4",
          9192 => x"2e",
          9193 => x"83",
          9194 => x"7f",
          9195 => x"81",
          9196 => x"38",
          9197 => x"53",
          9198 => x"81",
          9199 => x"d4",
          9200 => x"b9",
          9201 => x"2e",
          9202 => x"56",
          9203 => x"b4",
          9204 => x"56",
          9205 => x"9c",
          9206 => x"33",
          9207 => x"81",
          9208 => x"c9",
          9209 => x"70",
          9210 => x"07",
          9211 => x"80",
          9212 => x"38",
          9213 => x"78",
          9214 => x"89",
          9215 => x"7d",
          9216 => x"3f",
          9217 => x"08",
          9218 => x"c8",
          9219 => x"ff",
          9220 => x"58",
          9221 => x"81",
          9222 => x"58",
          9223 => x"38",
          9224 => x"7f",
          9225 => x"98",
          9226 => x"b4",
          9227 => x"2e",
          9228 => x"1c",
          9229 => x"40",
          9230 => x"38",
          9231 => x"53",
          9232 => x"81",
          9233 => x"d3",
          9234 => x"b9",
          9235 => x"2e",
          9236 => x"57",
          9237 => x"b4",
          9238 => x"58",
          9239 => x"38",
          9240 => x"1f",
          9241 => x"80",
          9242 => x"05",
          9243 => x"15",
          9244 => x"38",
          9245 => x"1f",
          9246 => x"58",
          9247 => x"81",
          9248 => x"77",
          9249 => x"59",
          9250 => x"55",
          9251 => x"9c",
          9252 => x"1f",
          9253 => x"5e",
          9254 => x"1b",
          9255 => x"83",
          9256 => x"56",
          9257 => x"c8",
          9258 => x"0d",
          9259 => x"30",
          9260 => x"72",
          9261 => x"57",
          9262 => x"38",
          9263 => x"52",
          9264 => x"c2",
          9265 => x"c8",
          9266 => x"b9",
          9267 => x"2e",
          9268 => x"fe",
          9269 => x"54",
          9270 => x"53",
          9271 => x"18",
          9272 => x"80",
          9273 => x"c8",
          9274 => x"09",
          9275 => x"bf",
          9276 => x"c8",
          9277 => x"34",
          9278 => x"a8",
          9279 => x"55",
          9280 => x"08",
          9281 => x"82",
          9282 => x"60",
          9283 => x"ac",
          9284 => x"c8",
          9285 => x"9c",
          9286 => x"2b",
          9287 => x"71",
          9288 => x"7d",
          9289 => x"3f",
          9290 => x"08",
          9291 => x"c8",
          9292 => x"38",
          9293 => x"c8",
          9294 => x"8b",
          9295 => x"2a",
          9296 => x"29",
          9297 => x"81",
          9298 => x"57",
          9299 => x"81",
          9300 => x"19",
          9301 => x"76",
          9302 => x"81",
          9303 => x"1d",
          9304 => x"1e",
          9305 => x"56",
          9306 => x"77",
          9307 => x"83",
          9308 => x"7a",
          9309 => x"81",
          9310 => x"38",
          9311 => x"53",
          9312 => x"81",
          9313 => x"d0",
          9314 => x"b9",
          9315 => x"2e",
          9316 => x"57",
          9317 => x"b4",
          9318 => x"58",
          9319 => x"38",
          9320 => x"9c",
          9321 => x"81",
          9322 => x"5c",
          9323 => x"1c",
          9324 => x"8b",
          9325 => x"8c",
          9326 => x"9a",
          9327 => x"9b",
          9328 => x"8d",
          9329 => x"76",
          9330 => x"59",
          9331 => x"ff",
          9332 => x"78",
          9333 => x"22",
          9334 => x"58",
          9335 => x"c8",
          9336 => x"05",
          9337 => x"70",
          9338 => x"34",
          9339 => x"56",
          9340 => x"76",
          9341 => x"ff",
          9342 => x"18",
          9343 => x"27",
          9344 => x"83",
          9345 => x"81",
          9346 => x"10",
          9347 => x"58",
          9348 => x"2e",
          9349 => x"7c",
          9350 => x"0b",
          9351 => x"80",
          9352 => x"e9",
          9353 => x"b9",
          9354 => x"84",
          9355 => x"fc",
          9356 => x"ff",
          9357 => x"fe",
          9358 => x"eb",
          9359 => x"b4",
          9360 => x"b8",
          9361 => x"81",
          9362 => x"59",
          9363 => x"81",
          9364 => x"c8",
          9365 => x"38",
          9366 => x"08",
          9367 => x"b4",
          9368 => x"1d",
          9369 => x"b9",
          9370 => x"41",
          9371 => x"08",
          9372 => x"38",
          9373 => x"42",
          9374 => x"09",
          9375 => x"bc",
          9376 => x"b4",
          9377 => x"1d",
          9378 => x"78",
          9379 => x"33",
          9380 => x"3f",
          9381 => x"a4",
          9382 => x"1f",
          9383 => x"57",
          9384 => x"81",
          9385 => x"81",
          9386 => x"38",
          9387 => x"81",
          9388 => x"76",
          9389 => x"9f",
          9390 => x"39",
          9391 => x"07",
          9392 => x"39",
          9393 => x"1c",
          9394 => x"52",
          9395 => x"51",
          9396 => x"84",
          9397 => x"76",
          9398 => x"06",
          9399 => x"b9",
          9400 => x"1d",
          9401 => x"08",
          9402 => x"31",
          9403 => x"1d",
          9404 => x"38",
          9405 => x"5f",
          9406 => x"aa",
          9407 => x"c8",
          9408 => x"f8",
          9409 => x"1c",
          9410 => x"80",
          9411 => x"38",
          9412 => x"75",
          9413 => x"e8",
          9414 => x"59",
          9415 => x"2e",
          9416 => x"fa",
          9417 => x"54",
          9418 => x"a0",
          9419 => x"53",
          9420 => x"1c",
          9421 => x"ac",
          9422 => x"39",
          9423 => x"18",
          9424 => x"08",
          9425 => x"52",
          9426 => x"51",
          9427 => x"f8",
          9428 => x"3d",
          9429 => x"71",
          9430 => x"5c",
          9431 => x"1e",
          9432 => x"08",
          9433 => x"b5",
          9434 => x"08",
          9435 => x"d9",
          9436 => x"71",
          9437 => x"08",
          9438 => x"58",
          9439 => x"72",
          9440 => x"38",
          9441 => x"14",
          9442 => x"1b",
          9443 => x"7a",
          9444 => x"80",
          9445 => x"70",
          9446 => x"06",
          9447 => x"8f",
          9448 => x"83",
          9449 => x"1a",
          9450 => x"22",
          9451 => x"5b",
          9452 => x"7a",
          9453 => x"25",
          9454 => x"06",
          9455 => x"7c",
          9456 => x"57",
          9457 => x"18",
          9458 => x"89",
          9459 => x"58",
          9460 => x"16",
          9461 => x"18",
          9462 => x"74",
          9463 => x"38",
          9464 => x"81",
          9465 => x"89",
          9466 => x"70",
          9467 => x"25",
          9468 => x"77",
          9469 => x"38",
          9470 => x"8b",
          9471 => x"70",
          9472 => x"34",
          9473 => x"74",
          9474 => x"05",
          9475 => x"18",
          9476 => x"27",
          9477 => x"7c",
          9478 => x"55",
          9479 => x"16",
          9480 => x"33",
          9481 => x"38",
          9482 => x"38",
          9483 => x"1e",
          9484 => x"7c",
          9485 => x"56",
          9486 => x"17",
          9487 => x"08",
          9488 => x"55",
          9489 => x"38",
          9490 => x"34",
          9491 => x"53",
          9492 => x"88",
          9493 => x"1c",
          9494 => x"83",
          9495 => x"12",
          9496 => x"2b",
          9497 => x"07",
          9498 => x"70",
          9499 => x"2b",
          9500 => x"07",
          9501 => x"97",
          9502 => x"17",
          9503 => x"2b",
          9504 => x"5b",
          9505 => x"5b",
          9506 => x"1e",
          9507 => x"33",
          9508 => x"71",
          9509 => x"5d",
          9510 => x"1e",
          9511 => x"0d",
          9512 => x"55",
          9513 => x"77",
          9514 => x"81",
          9515 => x"58",
          9516 => x"b5",
          9517 => x"2b",
          9518 => x"81",
          9519 => x"84",
          9520 => x"83",
          9521 => x"55",
          9522 => x"27",
          9523 => x"76",
          9524 => x"38",
          9525 => x"54",
          9526 => x"74",
          9527 => x"82",
          9528 => x"80",
          9529 => x"08",
          9530 => x"19",
          9531 => x"22",
          9532 => x"79",
          9533 => x"fd",
          9534 => x"30",
          9535 => x"78",
          9536 => x"72",
          9537 => x"58",
          9538 => x"80",
          9539 => x"7a",
          9540 => x"05",
          9541 => x"8c",
          9542 => x"5b",
          9543 => x"73",
          9544 => x"5a",
          9545 => x"80",
          9546 => x"38",
          9547 => x"7e",
          9548 => x"89",
          9549 => x"bf",
          9550 => x"78",
          9551 => x"38",
          9552 => x"8c",
          9553 => x"5b",
          9554 => x"b4",
          9555 => x"2a",
          9556 => x"06",
          9557 => x"2e",
          9558 => x"14",
          9559 => x"ff",
          9560 => x"73",
          9561 => x"05",
          9562 => x"16",
          9563 => x"19",
          9564 => x"33",
          9565 => x"56",
          9566 => x"b7",
          9567 => x"39",
          9568 => x"53",
          9569 => x"7b",
          9570 => x"25",
          9571 => x"06",
          9572 => x"58",
          9573 => x"ef",
          9574 => x"70",
          9575 => x"57",
          9576 => x"70",
          9577 => x"53",
          9578 => x"83",
          9579 => x"74",
          9580 => x"81",
          9581 => x"80",
          9582 => x"38",
          9583 => x"88",
          9584 => x"33",
          9585 => x"3d",
          9586 => x"9f",
          9587 => x"a7",
          9588 => x"8c",
          9589 => x"80",
          9590 => x"70",
          9591 => x"33",
          9592 => x"81",
          9593 => x"7f",
          9594 => x"2e",
          9595 => x"83",
          9596 => x"27",
          9597 => x"10",
          9598 => x"76",
          9599 => x"57",
          9600 => x"ff",
          9601 => x"32",
          9602 => x"73",
          9603 => x"25",
          9604 => x"5b",
          9605 => x"90",
          9606 => x"dc",
          9607 => x"38",
          9608 => x"26",
          9609 => x"e4",
          9610 => x"e4",
          9611 => x"81",
          9612 => x"54",
          9613 => x"2e",
          9614 => x"73",
          9615 => x"38",
          9616 => x"33",
          9617 => x"06",
          9618 => x"73",
          9619 => x"81",
          9620 => x"7a",
          9621 => x"76",
          9622 => x"80",
          9623 => x"10",
          9624 => x"7d",
          9625 => x"62",
          9626 => x"05",
          9627 => x"54",
          9628 => x"2e",
          9629 => x"80",
          9630 => x"73",
          9631 => x"70",
          9632 => x"25",
          9633 => x"55",
          9634 => x"80",
          9635 => x"81",
          9636 => x"54",
          9637 => x"54",
          9638 => x"2e",
          9639 => x"80",
          9640 => x"30",
          9641 => x"77",
          9642 => x"57",
          9643 => x"72",
          9644 => x"73",
          9645 => x"94",
          9646 => x"55",
          9647 => x"fe",
          9648 => x"39",
          9649 => x"73",
          9650 => x"e7",
          9651 => x"c8",
          9652 => x"ff",
          9653 => x"fe",
          9654 => x"54",
          9655 => x"c8",
          9656 => x"0d",
          9657 => x"e4",
          9658 => x"ff",
          9659 => x"7a",
          9660 => x"e3",
          9661 => x"ff",
          9662 => x"1d",
          9663 => x"7b",
          9664 => x"3f",
          9665 => x"08",
          9666 => x"0c",
          9667 => x"04",
          9668 => x"dc",
          9669 => x"70",
          9670 => x"07",
          9671 => x"56",
          9672 => x"a1",
          9673 => x"42",
          9674 => x"33",
          9675 => x"72",
          9676 => x"38",
          9677 => x"32",
          9678 => x"80",
          9679 => x"40",
          9680 => x"e1",
          9681 => x"0c",
          9682 => x"82",
          9683 => x"81",
          9684 => x"38",
          9685 => x"83",
          9686 => x"17",
          9687 => x"2e",
          9688 => x"17",
          9689 => x"05",
          9690 => x"a0",
          9691 => x"70",
          9692 => x"42",
          9693 => x"59",
          9694 => x"84",
          9695 => x"38",
          9696 => x"76",
          9697 => x"59",
          9698 => x"80",
          9699 => x"80",
          9700 => x"38",
          9701 => x"70",
          9702 => x"06",
          9703 => x"55",
          9704 => x"2e",
          9705 => x"73",
          9706 => x"06",
          9707 => x"2e",
          9708 => x"76",
          9709 => x"38",
          9710 => x"05",
          9711 => x"54",
          9712 => x"9d",
          9713 => x"18",
          9714 => x"ff",
          9715 => x"80",
          9716 => x"fe",
          9717 => x"5e",
          9718 => x"2e",
          9719 => x"eb",
          9720 => x"a0",
          9721 => x"a0",
          9722 => x"05",
          9723 => x"13",
          9724 => x"38",
          9725 => x"5e",
          9726 => x"70",
          9727 => x"59",
          9728 => x"74",
          9729 => x"ed",
          9730 => x"2e",
          9731 => x"74",
          9732 => x"30",
          9733 => x"55",
          9734 => x"77",
          9735 => x"38",
          9736 => x"38",
          9737 => x"7b",
          9738 => x"81",
          9739 => x"32",
          9740 => x"72",
          9741 => x"70",
          9742 => x"51",
          9743 => x"80",
          9744 => x"38",
          9745 => x"86",
          9746 => x"77",
          9747 => x"79",
          9748 => x"75",
          9749 => x"38",
          9750 => x"5b",
          9751 => x"2b",
          9752 => x"77",
          9753 => x"5d",
          9754 => x"22",
          9755 => x"56",
          9756 => x"95",
          9757 => x"33",
          9758 => x"e5",
          9759 => x"38",
          9760 => x"82",
          9761 => x"8c",
          9762 => x"8c",
          9763 => x"38",
          9764 => x"55",
          9765 => x"82",
          9766 => x"81",
          9767 => x"56",
          9768 => x"7d",
          9769 => x"7c",
          9770 => x"38",
          9771 => x"5a",
          9772 => x"81",
          9773 => x"80",
          9774 => x"79",
          9775 => x"79",
          9776 => x"7b",
          9777 => x"3f",
          9778 => x"08",
          9779 => x"56",
          9780 => x"c8",
          9781 => x"81",
          9782 => x"b9",
          9783 => x"2e",
          9784 => x"fb",
          9785 => x"85",
          9786 => x"5a",
          9787 => x"84",
          9788 => x"82",
          9789 => x"59",
          9790 => x"38",
          9791 => x"55",
          9792 => x"8c",
          9793 => x"80",
          9794 => x"39",
          9795 => x"11",
          9796 => x"22",
          9797 => x"56",
          9798 => x"f0",
          9799 => x"2e",
          9800 => x"79",
          9801 => x"fd",
          9802 => x"18",
          9803 => x"ae",
          9804 => x"06",
          9805 => x"77",
          9806 => x"ae",
          9807 => x"06",
          9808 => x"76",
          9809 => x"80",
          9810 => x"0b",
          9811 => x"53",
          9812 => x"73",
          9813 => x"a0",
          9814 => x"70",
          9815 => x"34",
          9816 => x"8a",
          9817 => x"38",
          9818 => x"58",
          9819 => x"34",
          9820 => x"bf",
          9821 => x"c8",
          9822 => x"33",
          9823 => x"b9",
          9824 => x"d6",
          9825 => x"2a",
          9826 => x"77",
          9827 => x"86",
          9828 => x"84",
          9829 => x"56",
          9830 => x"2e",
          9831 => x"90",
          9832 => x"ff",
          9833 => x"80",
          9834 => x"80",
          9835 => x"71",
          9836 => x"62",
          9837 => x"54",
          9838 => x"2e",
          9839 => x"74",
          9840 => x"7b",
          9841 => x"56",
          9842 => x"77",
          9843 => x"ae",
          9844 => x"38",
          9845 => x"76",
          9846 => x"fb",
          9847 => x"83",
          9848 => x"56",
          9849 => x"39",
          9850 => x"81",
          9851 => x"8c",
          9852 => x"77",
          9853 => x"81",
          9854 => x"38",
          9855 => x"5a",
          9856 => x"85",
          9857 => x"34",
          9858 => x"09",
          9859 => x"f6",
          9860 => x"ff",
          9861 => x"1d",
          9862 => x"84",
          9863 => x"93",
          9864 => x"74",
          9865 => x"9d",
          9866 => x"75",
          9867 => x"38",
          9868 => x"78",
          9869 => x"f7",
          9870 => x"07",
          9871 => x"57",
          9872 => x"a4",
          9873 => x"07",
          9874 => x"52",
          9875 => x"85",
          9876 => x"b9",
          9877 => x"ff",
          9878 => x"87",
          9879 => x"5a",
          9880 => x"2e",
          9881 => x"80",
          9882 => x"e5",
          9883 => x"56",
          9884 => x"ff",
          9885 => x"38",
          9886 => x"81",
          9887 => x"e4",
          9888 => x"e4",
          9889 => x"81",
          9890 => x"54",
          9891 => x"2e",
          9892 => x"73",
          9893 => x"38",
          9894 => x"33",
          9895 => x"06",
          9896 => x"73",
          9897 => x"81",
          9898 => x"78",
          9899 => x"ff",
          9900 => x"73",
          9901 => x"38",
          9902 => x"70",
          9903 => x"5f",
          9904 => x"15",
          9905 => x"26",
          9906 => x"81",
          9907 => x"ff",
          9908 => x"70",
          9909 => x"06",
          9910 => x"53",
          9911 => x"05",
          9912 => x"34",
          9913 => x"75",
          9914 => x"fc",
          9915 => x"fa",
          9916 => x"e4",
          9917 => x"81",
          9918 => x"53",
          9919 => x"ff",
          9920 => x"df",
          9921 => x"7d",
          9922 => x"5b",
          9923 => x"79",
          9924 => x"5b",
          9925 => x"cd",
          9926 => x"cc",
          9927 => x"98",
          9928 => x"2b",
          9929 => x"88",
          9930 => x"57",
          9931 => x"7b",
          9932 => x"75",
          9933 => x"54",
          9934 => x"81",
          9935 => x"a0",
          9936 => x"74",
          9937 => x"1b",
          9938 => x"39",
          9939 => x"a0",
          9940 => x"5a",
          9941 => x"2e",
          9942 => x"fa",
          9943 => x"a3",
          9944 => x"2a",
          9945 => x"7b",
          9946 => x"85",
          9947 => x"c8",
          9948 => x"0d",
          9949 => x"0d",
          9950 => x"88",
          9951 => x"05",
          9952 => x"5e",
          9953 => x"ff",
          9954 => x"59",
          9955 => x"80",
          9956 => x"38",
          9957 => x"05",
          9958 => x"9f",
          9959 => x"75",
          9960 => x"d0",
          9961 => x"38",
          9962 => x"85",
          9963 => x"d1",
          9964 => x"80",
          9965 => x"b2",
          9966 => x"10",
          9967 => x"05",
          9968 => x"5a",
          9969 => x"80",
          9970 => x"38",
          9971 => x"7f",
          9972 => x"77",
          9973 => x"7b",
          9974 => x"38",
          9975 => x"51",
          9976 => x"3f",
          9977 => x"08",
          9978 => x"70",
          9979 => x"58",
          9980 => x"86",
          9981 => x"77",
          9982 => x"5d",
          9983 => x"1d",
          9984 => x"34",
          9985 => x"17",
          9986 => x"bb",
          9987 => x"b9",
          9988 => x"ff",
          9989 => x"06",
          9990 => x"58",
          9991 => x"38",
          9992 => x"8d",
          9993 => x"2a",
          9994 => x"8a",
          9995 => x"b1",
          9996 => x"7a",
          9997 => x"ff",
          9998 => x"0c",
          9999 => x"55",
         10000 => x"53",
         10001 => x"53",
         10002 => x"52",
         10003 => x"95",
         10004 => x"c8",
         10005 => x"85",
         10006 => x"81",
         10007 => x"18",
         10008 => x"78",
         10009 => x"b7",
         10010 => x"b6",
         10011 => x"88",
         10012 => x"56",
         10013 => x"82",
         10014 => x"85",
         10015 => x"81",
         10016 => x"84",
         10017 => x"33",
         10018 => x"bf",
         10019 => x"75",
         10020 => x"cd",
         10021 => x"75",
         10022 => x"c5",
         10023 => x"17",
         10024 => x"18",
         10025 => x"2b",
         10026 => x"7c",
         10027 => x"09",
         10028 => x"ad",
         10029 => x"17",
         10030 => x"18",
         10031 => x"2b",
         10032 => x"75",
         10033 => x"dc",
         10034 => x"33",
         10035 => x"71",
         10036 => x"88",
         10037 => x"14",
         10038 => x"07",
         10039 => x"33",
         10040 => x"5a",
         10041 => x"5f",
         10042 => x"18",
         10043 => x"17",
         10044 => x"34",
         10045 => x"33",
         10046 => x"81",
         10047 => x"40",
         10048 => x"7c",
         10049 => x"d9",
         10050 => x"ff",
         10051 => x"29",
         10052 => x"33",
         10053 => x"77",
         10054 => x"77",
         10055 => x"2e",
         10056 => x"ff",
         10057 => x"42",
         10058 => x"38",
         10059 => x"33",
         10060 => x"33",
         10061 => x"07",
         10062 => x"88",
         10063 => x"75",
         10064 => x"5a",
         10065 => x"82",
         10066 => x"cc",
         10067 => x"cb",
         10068 => x"88",
         10069 => x"5c",
         10070 => x"80",
         10071 => x"11",
         10072 => x"33",
         10073 => x"71",
         10074 => x"81",
         10075 => x"72",
         10076 => x"75",
         10077 => x"53",
         10078 => x"42",
         10079 => x"c7",
         10080 => x"c6",
         10081 => x"88",
         10082 => x"58",
         10083 => x"80",
         10084 => x"38",
         10085 => x"84",
         10086 => x"79",
         10087 => x"c1",
         10088 => x"74",
         10089 => x"fd",
         10090 => x"84",
         10091 => x"56",
         10092 => x"08",
         10093 => x"a9",
         10094 => x"c8",
         10095 => x"ff",
         10096 => x"83",
         10097 => x"75",
         10098 => x"26",
         10099 => x"5d",
         10100 => x"26",
         10101 => x"81",
         10102 => x"70",
         10103 => x"7b",
         10104 => x"7b",
         10105 => x"1a",
         10106 => x"b0",
         10107 => x"59",
         10108 => x"8a",
         10109 => x"17",
         10110 => x"58",
         10111 => x"80",
         10112 => x"16",
         10113 => x"78",
         10114 => x"82",
         10115 => x"78",
         10116 => x"81",
         10117 => x"06",
         10118 => x"83",
         10119 => x"2a",
         10120 => x"78",
         10121 => x"26",
         10122 => x"0b",
         10123 => x"ff",
         10124 => x"0c",
         10125 => x"84",
         10126 => x"83",
         10127 => x"38",
         10128 => x"84",
         10129 => x"81",
         10130 => x"84",
         10131 => x"7c",
         10132 => x"84",
         10133 => x"8c",
         10134 => x"0b",
         10135 => x"80",
         10136 => x"b9",
         10137 => x"3d",
         10138 => x"0b",
         10139 => x"0c",
         10140 => x"04",
         10141 => x"11",
         10142 => x"06",
         10143 => x"74",
         10144 => x"38",
         10145 => x"81",
         10146 => x"05",
         10147 => x"7a",
         10148 => x"38",
         10149 => x"83",
         10150 => x"40",
         10151 => x"7f",
         10152 => x"70",
         10153 => x"33",
         10154 => x"05",
         10155 => x"9f",
         10156 => x"56",
         10157 => x"89",
         10158 => x"70",
         10159 => x"57",
         10160 => x"17",
         10161 => x"26",
         10162 => x"17",
         10163 => x"06",
         10164 => x"30",
         10165 => x"59",
         10166 => x"2e",
         10167 => x"85",
         10168 => x"be",
         10169 => x"32",
         10170 => x"72",
         10171 => x"7a",
         10172 => x"55",
         10173 => x"87",
         10174 => x"1c",
         10175 => x"5c",
         10176 => x"ff",
         10177 => x"56",
         10178 => x"78",
         10179 => x"cf",
         10180 => x"2a",
         10181 => x"8a",
         10182 => x"c5",
         10183 => x"fe",
         10184 => x"78",
         10185 => x"75",
         10186 => x"09",
         10187 => x"38",
         10188 => x"81",
         10189 => x"30",
         10190 => x"7b",
         10191 => x"5c",
         10192 => x"38",
         10193 => x"2e",
         10194 => x"93",
         10195 => x"5a",
         10196 => x"fa",
         10197 => x"59",
         10198 => x"2e",
         10199 => x"81",
         10200 => x"80",
         10201 => x"90",
         10202 => x"2b",
         10203 => x"19",
         10204 => x"07",
         10205 => x"fe",
         10206 => x"07",
         10207 => x"40",
         10208 => x"7a",
         10209 => x"5c",
         10210 => x"90",
         10211 => x"78",
         10212 => x"be",
         10213 => x"bd",
         10214 => x"30",
         10215 => x"72",
         10216 => x"3d",
         10217 => x"05",
         10218 => x"b6",
         10219 => x"52",
         10220 => x"78",
         10221 => x"56",
         10222 => x"80",
         10223 => x"0b",
         10224 => x"ff",
         10225 => x"0c",
         10226 => x"56",
         10227 => x"a5",
         10228 => x"7a",
         10229 => x"52",
         10230 => x"51",
         10231 => x"3f",
         10232 => x"08",
         10233 => x"38",
         10234 => x"56",
         10235 => x"0c",
         10236 => x"bf",
         10237 => x"33",
         10238 => x"88",
         10239 => x"5e",
         10240 => x"82",
         10241 => x"09",
         10242 => x"38",
         10243 => x"18",
         10244 => x"75",
         10245 => x"82",
         10246 => x"81",
         10247 => x"30",
         10248 => x"7a",
         10249 => x"42",
         10250 => x"75",
         10251 => x"b6",
         10252 => x"77",
         10253 => x"56",
         10254 => x"b9",
         10255 => x"5d",
         10256 => x"2e",
         10257 => x"83",
         10258 => x"81",
         10259 => x"bd",
         10260 => x"2e",
         10261 => x"81",
         10262 => x"5a",
         10263 => x"27",
         10264 => x"f8",
         10265 => x"0b",
         10266 => x"83",
         10267 => x"5d",
         10268 => x"81",
         10269 => x"7e",
         10270 => x"40",
         10271 => x"31",
         10272 => x"52",
         10273 => x"80",
         10274 => x"38",
         10275 => x"e1",
         10276 => x"81",
         10277 => x"e4",
         10278 => x"58",
         10279 => x"05",
         10280 => x"70",
         10281 => x"33",
         10282 => x"ff",
         10283 => x"42",
         10284 => x"2e",
         10285 => x"75",
         10286 => x"38",
         10287 => x"f3",
         10288 => x"7c",
         10289 => x"77",
         10290 => x"0c",
         10291 => x"04",
         10292 => x"80",
         10293 => x"38",
         10294 => x"8a",
         10295 => x"fc",
         10296 => x"ff",
         10297 => x"0b",
         10298 => x"0c",
         10299 => x"04",
         10300 => x"ee",
         10301 => x"f8",
         10302 => x"78",
         10303 => x"5a",
         10304 => x"81",
         10305 => x"71",
         10306 => x"1b",
         10307 => x"5f",
         10308 => x"83",
         10309 => x"80",
         10310 => x"85",
         10311 => x"18",
         10312 => x"5c",
         10313 => x"70",
         10314 => x"33",
         10315 => x"05",
         10316 => x"71",
         10317 => x"5b",
         10318 => x"77",
         10319 => x"91",
         10320 => x"2e",
         10321 => x"3d",
         10322 => x"83",
         10323 => x"39",
         10324 => x"c6",
         10325 => x"17",
         10326 => x"18",
         10327 => x"2b",
         10328 => x"75",
         10329 => x"81",
         10330 => x"38",
         10331 => x"80",
         10332 => x"08",
         10333 => x"38",
         10334 => x"5b",
         10335 => x"09",
         10336 => x"9b",
         10337 => x"77",
         10338 => x"52",
         10339 => x"51",
         10340 => x"3f",
         10341 => x"08",
         10342 => x"38",
         10343 => x"5a",
         10344 => x"0c",
         10345 => x"38",
         10346 => x"34",
         10347 => x"33",
         10348 => x"33",
         10349 => x"07",
         10350 => x"82",
         10351 => x"09",
         10352 => x"fc",
         10353 => x"83",
         10354 => x"12",
         10355 => x"2b",
         10356 => x"07",
         10357 => x"70",
         10358 => x"2b",
         10359 => x"07",
         10360 => x"45",
         10361 => x"77",
         10362 => x"a4",
         10363 => x"81",
         10364 => x"38",
         10365 => x"83",
         10366 => x"12",
         10367 => x"2b",
         10368 => x"07",
         10369 => x"70",
         10370 => x"2b",
         10371 => x"07",
         10372 => x"5b",
         10373 => x"60",
         10374 => x"e4",
         10375 => x"81",
         10376 => x"38",
         10377 => x"83",
         10378 => x"12",
         10379 => x"2b",
         10380 => x"07",
         10381 => x"70",
         10382 => x"2b",
         10383 => x"07",
         10384 => x"5d",
         10385 => x"83",
         10386 => x"12",
         10387 => x"2b",
         10388 => x"07",
         10389 => x"70",
         10390 => x"2b",
         10391 => x"07",
         10392 => x"0c",
         10393 => x"46",
         10394 => x"45",
         10395 => x"7c",
         10396 => x"d1",
         10397 => x"05",
         10398 => x"d1",
         10399 => x"86",
         10400 => x"d1",
         10401 => x"18",
         10402 => x"98",
         10403 => x"cf",
         10404 => x"24",
         10405 => x"7b",
         10406 => x"56",
         10407 => x"75",
         10408 => x"08",
         10409 => x"70",
         10410 => x"33",
         10411 => x"af",
         10412 => x"b9",
         10413 => x"2e",
         10414 => x"81",
         10415 => x"b9",
         10416 => x"18",
         10417 => x"08",
         10418 => x"31",
         10419 => x"18",
         10420 => x"38",
         10421 => x"41",
         10422 => x"81",
         10423 => x"b9",
         10424 => x"fd",
         10425 => x"56",
         10426 => x"f3",
         10427 => x"0b",
         10428 => x"83",
         10429 => x"5a",
         10430 => x"39",
         10431 => x"33",
         10432 => x"33",
         10433 => x"07",
         10434 => x"58",
         10435 => x"38",
         10436 => x"42",
         10437 => x"38",
         10438 => x"83",
         10439 => x"12",
         10440 => x"2b",
         10441 => x"07",
         10442 => x"70",
         10443 => x"2b",
         10444 => x"07",
         10445 => x"5a",
         10446 => x"5a",
         10447 => x"59",
         10448 => x"39",
         10449 => x"80",
         10450 => x"38",
         10451 => x"e3",
         10452 => x"2e",
         10453 => x"93",
         10454 => x"5a",
         10455 => x"f2",
         10456 => x"79",
         10457 => x"fc",
         10458 => x"54",
         10459 => x"a0",
         10460 => x"53",
         10461 => x"17",
         10462 => x"ad",
         10463 => x"85",
         10464 => x"0d",
         10465 => x"05",
         10466 => x"43",
         10467 => x"57",
         10468 => x"5a",
         10469 => x"2e",
         10470 => x"78",
         10471 => x"5a",
         10472 => x"26",
         10473 => x"ba",
         10474 => x"38",
         10475 => x"74",
         10476 => x"d9",
         10477 => x"a4",
         10478 => x"74",
         10479 => x"38",
         10480 => x"84",
         10481 => x"70",
         10482 => x"73",
         10483 => x"38",
         10484 => x"62",
         10485 => x"2e",
         10486 => x"74",
         10487 => x"73",
         10488 => x"54",
         10489 => x"92",
         10490 => x"93",
         10491 => x"84",
         10492 => x"81",
         10493 => x"c8",
         10494 => x"84",
         10495 => x"92",
         10496 => x"8b",
         10497 => x"c8",
         10498 => x"0d",
         10499 => x"d0",
         10500 => x"ff",
         10501 => x"57",
         10502 => x"91",
         10503 => x"77",
         10504 => x"d0",
         10505 => x"77",
         10506 => x"f7",
         10507 => x"08",
         10508 => x"5e",
         10509 => x"08",
         10510 => x"79",
         10511 => x"5b",
         10512 => x"81",
         10513 => x"ff",
         10514 => x"57",
         10515 => x"26",
         10516 => x"15",
         10517 => x"06",
         10518 => x"9f",
         10519 => x"99",
         10520 => x"e0",
         10521 => x"ff",
         10522 => x"74",
         10523 => x"2a",
         10524 => x"76",
         10525 => x"06",
         10526 => x"ff",
         10527 => x"79",
         10528 => x"70",
         10529 => x"2a",
         10530 => x"57",
         10531 => x"2e",
         10532 => x"1b",
         10533 => x"5b",
         10534 => x"ff",
         10535 => x"54",
         10536 => x"7a",
         10537 => x"38",
         10538 => x"0c",
         10539 => x"39",
         10540 => x"6c",
         10541 => x"80",
         10542 => x"56",
         10543 => x"78",
         10544 => x"38",
         10545 => x"70",
         10546 => x"cc",
         10547 => x"3d",
         10548 => x"58",
         10549 => x"84",
         10550 => x"57",
         10551 => x"08",
         10552 => x"38",
         10553 => x"76",
         10554 => x"b9",
         10555 => x"3d",
         10556 => x"40",
         10557 => x"3d",
         10558 => x"e1",
         10559 => x"b9",
         10560 => x"84",
         10561 => x"80",
         10562 => x"38",
         10563 => x"5d",
         10564 => x"81",
         10565 => x"80",
         10566 => x"38",
         10567 => x"83",
         10568 => x"88",
         10569 => x"ff",
         10570 => x"83",
         10571 => x"5b",
         10572 => x"81",
         10573 => x"9b",
         10574 => x"12",
         10575 => x"2b",
         10576 => x"33",
         10577 => x"5e",
         10578 => x"2e",
         10579 => x"80",
         10580 => x"34",
         10581 => x"17",
         10582 => x"90",
         10583 => x"cc",
         10584 => x"34",
         10585 => x"0b",
         10586 => x"7e",
         10587 => x"80",
         10588 => x"34",
         10589 => x"17",
         10590 => x"5d",
         10591 => x"84",
         10592 => x"5b",
         10593 => x"1c",
         10594 => x"9d",
         10595 => x"0b",
         10596 => x"80",
         10597 => x"34",
         10598 => x"0b",
         10599 => x"7b",
         10600 => x"e2",
         10601 => x"11",
         10602 => x"08",
         10603 => x"57",
         10604 => x"89",
         10605 => x"08",
         10606 => x"8a",
         10607 => x"80",
         10608 => x"a3",
         10609 => x"e7",
         10610 => x"98",
         10611 => x"7b",
         10612 => x"b8",
         10613 => x"9c",
         10614 => x"7c",
         10615 => x"76",
         10616 => x"02",
         10617 => x"33",
         10618 => x"81",
         10619 => x"7b",
         10620 => x"77",
         10621 => x"06",
         10622 => x"2e",
         10623 => x"81",
         10624 => x"81",
         10625 => x"83",
         10626 => x"56",
         10627 => x"86",
         10628 => x"c0",
         10629 => x"b4",
         10630 => x"1b",
         10631 => x"1b",
         10632 => x"11",
         10633 => x"33",
         10634 => x"07",
         10635 => x"5e",
         10636 => x"7b",
         10637 => x"f1",
         10638 => x"1a",
         10639 => x"83",
         10640 => x"12",
         10641 => x"2b",
         10642 => x"07",
         10643 => x"70",
         10644 => x"2b",
         10645 => x"07",
         10646 => x"05",
         10647 => x"0c",
         10648 => x"59",
         10649 => x"86",
         10650 => x"1a",
         10651 => x"1a",
         10652 => x"91",
         10653 => x"0b",
         10654 => x"77",
         10655 => x"06",
         10656 => x"2e",
         10657 => x"75",
         10658 => x"f1",
         10659 => x"1a",
         10660 => x"22",
         10661 => x"7c",
         10662 => x"76",
         10663 => x"07",
         10664 => x"5b",
         10665 => x"84",
         10666 => x"70",
         10667 => x"5b",
         10668 => x"84",
         10669 => x"52",
         10670 => x"ac",
         10671 => x"b9",
         10672 => x"84",
         10673 => x"81",
         10674 => x"82",
         10675 => x"c8",
         10676 => x"80",
         10677 => x"7a",
         10678 => x"39",
         10679 => x"05",
         10680 => x"5e",
         10681 => x"77",
         10682 => x"06",
         10683 => x"2e",
         10684 => x"88",
         10685 => x"0c",
         10686 => x"87",
         10687 => x"0c",
         10688 => x"84",
         10689 => x"0c",
         10690 => x"79",
         10691 => x"3f",
         10692 => x"08",
         10693 => x"59",
         10694 => x"c8",
         10695 => x"39",
         10696 => x"31",
         10697 => x"f3",
         10698 => x"33",
         10699 => x"71",
         10700 => x"90",
         10701 => x"07",
         10702 => x"fd",
         10703 => x"55",
         10704 => x"81",
         10705 => x"52",
         10706 => x"ab",
         10707 => x"b9",
         10708 => x"84",
         10709 => x"80",
         10710 => x"38",
         10711 => x"08",
         10712 => x"d9",
         10713 => x"c8",
         10714 => x"83",
         10715 => x"53",
         10716 => x"51",
         10717 => x"3f",
         10718 => x"08",
         10719 => x"9c",
         10720 => x"11",
         10721 => x"58",
         10722 => x"75",
         10723 => x"38",
         10724 => x"18",
         10725 => x"33",
         10726 => x"74",
         10727 => x"7c",
         10728 => x"26",
         10729 => x"80",
         10730 => x"0b",
         10731 => x"80",
         10732 => x"34",
         10733 => x"95",
         10734 => x"17",
         10735 => x"2b",
         10736 => x"07",
         10737 => x"56",
         10738 => x"8e",
         10739 => x"0b",
         10740 => x"a1",
         10741 => x"34",
         10742 => x"91",
         10743 => x"56",
         10744 => x"17",
         10745 => x"57",
         10746 => x"9a",
         10747 => x"0b",
         10748 => x"7d",
         10749 => x"83",
         10750 => x"06",
         10751 => x"ff",
         10752 => x"7f",
         10753 => x"59",
         10754 => x"16",
         10755 => x"ae",
         10756 => x"33",
         10757 => x"2e",
         10758 => x"b5",
         10759 => x"7d",
         10760 => x"52",
         10761 => x"51",
         10762 => x"3f",
         10763 => x"08",
         10764 => x"38",
         10765 => x"5b",
         10766 => x"0c",
         10767 => x"ff",
         10768 => x"0c",
         10769 => x"2e",
         10770 => x"80",
         10771 => x"97",
         10772 => x"b4",
         10773 => x"b8",
         10774 => x"81",
         10775 => x"5a",
         10776 => x"3f",
         10777 => x"08",
         10778 => x"81",
         10779 => x"38",
         10780 => x"08",
         10781 => x"b4",
         10782 => x"17",
         10783 => x"b9",
         10784 => x"55",
         10785 => x"08",
         10786 => x"38",
         10787 => x"55",
         10788 => x"09",
         10789 => x"85",
         10790 => x"b4",
         10791 => x"17",
         10792 => x"79",
         10793 => x"33",
         10794 => x"b8",
         10795 => x"fe",
         10796 => x"94",
         10797 => x"56",
         10798 => x"77",
         10799 => x"76",
         10800 => x"75",
         10801 => x"5a",
         10802 => x"f8",
         10803 => x"fe",
         10804 => x"08",
         10805 => x"59",
         10806 => x"27",
         10807 => x"8a",
         10808 => x"71",
         10809 => x"08",
         10810 => x"74",
         10811 => x"cd",
         10812 => x"2a",
         10813 => x"0c",
         10814 => x"ed",
         10815 => x"1a",
         10816 => x"f7",
         10817 => x"57",
         10818 => x"f7",
         10819 => x"b9",
         10820 => x"80",
         10821 => x"cf",
         10822 => x"57",
         10823 => x"39",
         10824 => x"62",
         10825 => x"40",
         10826 => x"80",
         10827 => x"57",
         10828 => x"9f",
         10829 => x"56",
         10830 => x"97",
         10831 => x"55",
         10832 => x"8f",
         10833 => x"22",
         10834 => x"59",
         10835 => x"2e",
         10836 => x"80",
         10837 => x"76",
         10838 => x"8c",
         10839 => x"33",
         10840 => x"84",
         10841 => x"33",
         10842 => x"87",
         10843 => x"2e",
         10844 => x"94",
         10845 => x"1b",
         10846 => x"56",
         10847 => x"26",
         10848 => x"7b",
         10849 => x"d5",
         10850 => x"75",
         10851 => x"5b",
         10852 => x"38",
         10853 => x"ff",
         10854 => x"2a",
         10855 => x"9b",
         10856 => x"d3",
         10857 => x"08",
         10858 => x"27",
         10859 => x"74",
         10860 => x"f0",
         10861 => x"1b",
         10862 => x"98",
         10863 => x"05",
         10864 => x"fe",
         10865 => x"76",
         10866 => x"e7",
         10867 => x"22",
         10868 => x"b0",
         10869 => x"56",
         10870 => x"2e",
         10871 => x"7a",
         10872 => x"2a",
         10873 => x"80",
         10874 => x"38",
         10875 => x"75",
         10876 => x"38",
         10877 => x"58",
         10878 => x"53",
         10879 => x"19",
         10880 => x"9f",
         10881 => x"b9",
         10882 => x"98",
         10883 => x"11",
         10884 => x"75",
         10885 => x"38",
         10886 => x"77",
         10887 => x"78",
         10888 => x"84",
         10889 => x"29",
         10890 => x"58",
         10891 => x"70",
         10892 => x"33",
         10893 => x"05",
         10894 => x"15",
         10895 => x"38",
         10896 => x"58",
         10897 => x"7e",
         10898 => x"0c",
         10899 => x"1c",
         10900 => x"59",
         10901 => x"5e",
         10902 => x"af",
         10903 => x"75",
         10904 => x"0c",
         10905 => x"04",
         10906 => x"c8",
         10907 => x"0d",
         10908 => x"fe",
         10909 => x"1a",
         10910 => x"83",
         10911 => x"80",
         10912 => x"5b",
         10913 => x"83",
         10914 => x"76",
         10915 => x"08",
         10916 => x"38",
         10917 => x"1a",
         10918 => x"41",
         10919 => x"2e",
         10920 => x"80",
         10921 => x"54",
         10922 => x"19",
         10923 => x"33",
         10924 => x"b1",
         10925 => x"c8",
         10926 => x"85",
         10927 => x"81",
         10928 => x"1a",
         10929 => x"dc",
         10930 => x"1b",
         10931 => x"06",
         10932 => x"5a",
         10933 => x"56",
         10934 => x"2e",
         10935 => x"74",
         10936 => x"56",
         10937 => x"81",
         10938 => x"ff",
         10939 => x"80",
         10940 => x"38",
         10941 => x"05",
         10942 => x"70",
         10943 => x"34",
         10944 => x"75",
         10945 => x"bc",
         10946 => x"b4",
         10947 => x"b8",
         10948 => x"81",
         10949 => x"40",
         10950 => x"3f",
         10951 => x"b9",
         10952 => x"2e",
         10953 => x"ff",
         10954 => x"b9",
         10955 => x"1a",
         10956 => x"08",
         10957 => x"31",
         10958 => x"08",
         10959 => x"a0",
         10960 => x"fe",
         10961 => x"19",
         10962 => x"82",
         10963 => x"06",
         10964 => x"81",
         10965 => x"08",
         10966 => x"05",
         10967 => x"81",
         10968 => x"ff",
         10969 => x"7e",
         10970 => x"39",
         10971 => x"0c",
         10972 => x"56",
         10973 => x"98",
         10974 => x"79",
         10975 => x"98",
         10976 => x"c8",
         10977 => x"a1",
         10978 => x"33",
         10979 => x"83",
         10980 => x"c8",
         10981 => x"55",
         10982 => x"38",
         10983 => x"56",
         10984 => x"39",
         10985 => x"1b",
         10986 => x"84",
         10987 => x"92",
         10988 => x"82",
         10989 => x"34",
         10990 => x"b9",
         10991 => x"3d",
         10992 => x"3d",
         10993 => x"67",
         10994 => x"5c",
         10995 => x"0c",
         10996 => x"80",
         10997 => x"79",
         10998 => x"80",
         10999 => x"75",
         11000 => x"80",
         11001 => x"86",
         11002 => x"1b",
         11003 => x"78",
         11004 => x"fd",
         11005 => x"74",
         11006 => x"76",
         11007 => x"91",
         11008 => x"74",
         11009 => x"90",
         11010 => x"81",
         11011 => x"58",
         11012 => x"76",
         11013 => x"a1",
         11014 => x"08",
         11015 => x"57",
         11016 => x"84",
         11017 => x"5b",
         11018 => x"82",
         11019 => x"83",
         11020 => x"7e",
         11021 => x"60",
         11022 => x"ff",
         11023 => x"2a",
         11024 => x"78",
         11025 => x"84",
         11026 => x"1a",
         11027 => x"80",
         11028 => x"38",
         11029 => x"86",
         11030 => x"ff",
         11031 => x"38",
         11032 => x"0c",
         11033 => x"85",
         11034 => x"1b",
         11035 => x"b4",
         11036 => x"1b",
         11037 => x"d3",
         11038 => x"08",
         11039 => x"17",
         11040 => x"58",
         11041 => x"27",
         11042 => x"8a",
         11043 => x"79",
         11044 => x"08",
         11045 => x"74",
         11046 => x"de",
         11047 => x"7b",
         11048 => x"5c",
         11049 => x"83",
         11050 => x"19",
         11051 => x"27",
         11052 => x"79",
         11053 => x"54",
         11054 => x"52",
         11055 => x"51",
         11056 => x"3f",
         11057 => x"08",
         11058 => x"60",
         11059 => x"7d",
         11060 => x"74",
         11061 => x"38",
         11062 => x"b8",
         11063 => x"29",
         11064 => x"56",
         11065 => x"05",
         11066 => x"70",
         11067 => x"34",
         11068 => x"75",
         11069 => x"59",
         11070 => x"34",
         11071 => x"59",
         11072 => x"7e",
         11073 => x"0c",
         11074 => x"1c",
         11075 => x"71",
         11076 => x"8c",
         11077 => x"5a",
         11078 => x"75",
         11079 => x"38",
         11080 => x"8c",
         11081 => x"fe",
         11082 => x"1a",
         11083 => x"80",
         11084 => x"7a",
         11085 => x"80",
         11086 => x"b9",
         11087 => x"3d",
         11088 => x"84",
         11089 => x"92",
         11090 => x"83",
         11091 => x"74",
         11092 => x"60",
         11093 => x"39",
         11094 => x"08",
         11095 => x"83",
         11096 => x"80",
         11097 => x"5c",
         11098 => x"83",
         11099 => x"77",
         11100 => x"08",
         11101 => x"38",
         11102 => x"17",
         11103 => x"41",
         11104 => x"2e",
         11105 => x"80",
         11106 => x"54",
         11107 => x"16",
         11108 => x"33",
         11109 => x"cd",
         11110 => x"c8",
         11111 => x"85",
         11112 => x"81",
         11113 => x"17",
         11114 => x"bf",
         11115 => x"1b",
         11116 => x"06",
         11117 => x"b8",
         11118 => x"56",
         11119 => x"2e",
         11120 => x"70",
         11121 => x"33",
         11122 => x"05",
         11123 => x"16",
         11124 => x"38",
         11125 => x"0b",
         11126 => x"fe",
         11127 => x"54",
         11128 => x"53",
         11129 => x"53",
         11130 => x"52",
         11131 => x"f4",
         11132 => x"84",
         11133 => x"7f",
         11134 => x"06",
         11135 => x"84",
         11136 => x"83",
         11137 => x"16",
         11138 => x"08",
         11139 => x"c8",
         11140 => x"74",
         11141 => x"27",
         11142 => x"82",
         11143 => x"74",
         11144 => x"81",
         11145 => x"38",
         11146 => x"16",
         11147 => x"08",
         11148 => x"52",
         11149 => x"51",
         11150 => x"3f",
         11151 => x"ca",
         11152 => x"08",
         11153 => x"08",
         11154 => x"38",
         11155 => x"40",
         11156 => x"38",
         11157 => x"12",
         11158 => x"08",
         11159 => x"7c",
         11160 => x"58",
         11161 => x"98",
         11162 => x"79",
         11163 => x"e7",
         11164 => x"c8",
         11165 => x"b9",
         11166 => x"d8",
         11167 => x"33",
         11168 => x"39",
         11169 => x"51",
         11170 => x"3f",
         11171 => x"08",
         11172 => x"c8",
         11173 => x"38",
         11174 => x"54",
         11175 => x"53",
         11176 => x"53",
         11177 => x"52",
         11178 => x"b8",
         11179 => x"c8",
         11180 => x"38",
         11181 => x"08",
         11182 => x"b4",
         11183 => x"17",
         11184 => x"77",
         11185 => x"27",
         11186 => x"82",
         11187 => x"7b",
         11188 => x"81",
         11189 => x"38",
         11190 => x"16",
         11191 => x"08",
         11192 => x"52",
         11193 => x"51",
         11194 => x"3f",
         11195 => x"89",
         11196 => x"33",
         11197 => x"9b",
         11198 => x"c8",
         11199 => x"55",
         11200 => x"38",
         11201 => x"56",
         11202 => x"39",
         11203 => x"16",
         11204 => x"16",
         11205 => x"17",
         11206 => x"ff",
         11207 => x"84",
         11208 => x"80",
         11209 => x"b9",
         11210 => x"17",
         11211 => x"08",
         11212 => x"31",
         11213 => x"17",
         11214 => x"98",
         11215 => x"33",
         11216 => x"2e",
         11217 => x"fe",
         11218 => x"54",
         11219 => x"a0",
         11220 => x"53",
         11221 => x"16",
         11222 => x"96",
         11223 => x"7c",
         11224 => x"94",
         11225 => x"56",
         11226 => x"81",
         11227 => x"34",
         11228 => x"b9",
         11229 => x"3d",
         11230 => x"0b",
         11231 => x"82",
         11232 => x"c8",
         11233 => x"0d",
         11234 => x"0d",
         11235 => x"5a",
         11236 => x"9f",
         11237 => x"56",
         11238 => x"97",
         11239 => x"55",
         11240 => x"8f",
         11241 => x"22",
         11242 => x"58",
         11243 => x"2e",
         11244 => x"80",
         11245 => x"79",
         11246 => x"d8",
         11247 => x"33",
         11248 => x"81",
         11249 => x"7a",
         11250 => x"c8",
         11251 => x"19",
         11252 => x"b4",
         11253 => x"2e",
         11254 => x"17",
         11255 => x"81",
         11256 => x"54",
         11257 => x"17",
         11258 => x"33",
         11259 => x"f5",
         11260 => x"c8",
         11261 => x"85",
         11262 => x"81",
         11263 => x"18",
         11264 => x"90",
         11265 => x"08",
         11266 => x"a0",
         11267 => x"78",
         11268 => x"77",
         11269 => x"08",
         11270 => x"ff",
         11271 => x"56",
         11272 => x"34",
         11273 => x"5a",
         11274 => x"34",
         11275 => x"33",
         11276 => x"56",
         11277 => x"2e",
         11278 => x"8c",
         11279 => x"74",
         11280 => x"88",
         11281 => x"9d",
         11282 => x"90",
         11283 => x"9e",
         11284 => x"98",
         11285 => x"9f",
         11286 => x"7a",
         11287 => x"97",
         11288 => x"0b",
         11289 => x"80",
         11290 => x"18",
         11291 => x"92",
         11292 => x"0b",
         11293 => x"7b",
         11294 => x"83",
         11295 => x"51",
         11296 => x"3f",
         11297 => x"08",
         11298 => x"81",
         11299 => x"56",
         11300 => x"34",
         11301 => x"c8",
         11302 => x"0d",
         11303 => x"b4",
         11304 => x"b8",
         11305 => x"81",
         11306 => x"5b",
         11307 => x"3f",
         11308 => x"b9",
         11309 => x"c9",
         11310 => x"c8",
         11311 => x"34",
         11312 => x"a8",
         11313 => x"84",
         11314 => x"57",
         11315 => x"18",
         11316 => x"8e",
         11317 => x"33",
         11318 => x"2e",
         11319 => x"fe",
         11320 => x"54",
         11321 => x"a0",
         11322 => x"53",
         11323 => x"17",
         11324 => x"92",
         11325 => x"56",
         11326 => x"78",
         11327 => x"74",
         11328 => x"74",
         11329 => x"75",
         11330 => x"8c",
         11331 => x"74",
         11332 => x"88",
         11333 => x"9d",
         11334 => x"90",
         11335 => x"9e",
         11336 => x"98",
         11337 => x"9f",
         11338 => x"7a",
         11339 => x"97",
         11340 => x"0b",
         11341 => x"80",
         11342 => x"18",
         11343 => x"92",
         11344 => x"0b",
         11345 => x"7b",
         11346 => x"83",
         11347 => x"51",
         11348 => x"3f",
         11349 => x"08",
         11350 => x"81",
         11351 => x"56",
         11352 => x"34",
         11353 => x"81",
         11354 => x"ff",
         11355 => x"84",
         11356 => x"81",
         11357 => x"fc",
         11358 => x"78",
         11359 => x"fc",
         11360 => x"3d",
         11361 => x"52",
         11362 => x"3f",
         11363 => x"08",
         11364 => x"c8",
         11365 => x"89",
         11366 => x"2e",
         11367 => x"08",
         11368 => x"2e",
         11369 => x"33",
         11370 => x"2e",
         11371 => x"13",
         11372 => x"22",
         11373 => x"77",
         11374 => x"80",
         11375 => x"75",
         11376 => x"38",
         11377 => x"73",
         11378 => x"0c",
         11379 => x"04",
         11380 => x"51",
         11381 => x"3f",
         11382 => x"08",
         11383 => x"72",
         11384 => x"75",
         11385 => x"d5",
         11386 => x"0d",
         11387 => x"5b",
         11388 => x"80",
         11389 => x"75",
         11390 => x"57",
         11391 => x"26",
         11392 => x"ba",
         11393 => x"70",
         11394 => x"ba",
         11395 => x"84",
         11396 => x"51",
         11397 => x"90",
         11398 => x"d1",
         11399 => x"0b",
         11400 => x"0c",
         11401 => x"04",
         11402 => x"b9",
         11403 => x"3d",
         11404 => x"33",
         11405 => x"81",
         11406 => x"53",
         11407 => x"26",
         11408 => x"19",
         11409 => x"06",
         11410 => x"54",
         11411 => x"80",
         11412 => x"0b",
         11413 => x"5b",
         11414 => x"79",
         11415 => x"70",
         11416 => x"33",
         11417 => x"05",
         11418 => x"9f",
         11419 => x"52",
         11420 => x"89",
         11421 => x"70",
         11422 => x"53",
         11423 => x"13",
         11424 => x"26",
         11425 => x"13",
         11426 => x"06",
         11427 => x"30",
         11428 => x"55",
         11429 => x"2e",
         11430 => x"85",
         11431 => x"be",
         11432 => x"32",
         11433 => x"72",
         11434 => x"76",
         11435 => x"52",
         11436 => x"92",
         11437 => x"84",
         11438 => x"83",
         11439 => x"99",
         11440 => x"fe",
         11441 => x"83",
         11442 => x"77",
         11443 => x"fe",
         11444 => x"3d",
         11445 => x"98",
         11446 => x"52",
         11447 => x"d1",
         11448 => x"b9",
         11449 => x"84",
         11450 => x"80",
         11451 => x"74",
         11452 => x"0c",
         11453 => x"04",
         11454 => x"52",
         11455 => x"05",
         11456 => x"3f",
         11457 => x"08",
         11458 => x"c8",
         11459 => x"38",
         11460 => x"05",
         11461 => x"2b",
         11462 => x"77",
         11463 => x"38",
         11464 => x"33",
         11465 => x"81",
         11466 => x"75",
         11467 => x"38",
         11468 => x"11",
         11469 => x"33",
         11470 => x"07",
         11471 => x"5a",
         11472 => x"79",
         11473 => x"38",
         11474 => x"0c",
         11475 => x"c8",
         11476 => x"0d",
         11477 => x"c8",
         11478 => x"09",
         11479 => x"8f",
         11480 => x"84",
         11481 => x"98",
         11482 => x"95",
         11483 => x"17",
         11484 => x"2b",
         11485 => x"07",
         11486 => x"1b",
         11487 => x"cc",
         11488 => x"98",
         11489 => x"74",
         11490 => x"0c",
         11491 => x"04",
         11492 => x"0d",
         11493 => x"08",
         11494 => x"08",
         11495 => x"7c",
         11496 => x"80",
         11497 => x"b4",
         11498 => x"e5",
         11499 => x"c5",
         11500 => x"c8",
         11501 => x"b9",
         11502 => x"c8",
         11503 => x"d9",
         11504 => x"61",
         11505 => x"80",
         11506 => x"58",
         11507 => x"08",
         11508 => x"80",
         11509 => x"38",
         11510 => x"98",
         11511 => x"a0",
         11512 => x"ff",
         11513 => x"84",
         11514 => x"59",
         11515 => x"08",
         11516 => x"60",
         11517 => x"08",
         11518 => x"16",
         11519 => x"b1",
         11520 => x"c8",
         11521 => x"33",
         11522 => x"83",
         11523 => x"54",
         11524 => x"16",
         11525 => x"33",
         11526 => x"c9",
         11527 => x"c8",
         11528 => x"85",
         11529 => x"81",
         11530 => x"17",
         11531 => x"d4",
         11532 => x"3d",
         11533 => x"33",
         11534 => x"71",
         11535 => x"63",
         11536 => x"40",
         11537 => x"78",
         11538 => x"da",
         11539 => x"db",
         11540 => x"52",
         11541 => x"a3",
         11542 => x"b9",
         11543 => x"84",
         11544 => x"82",
         11545 => x"52",
         11546 => x"a8",
         11547 => x"b9",
         11548 => x"84",
         11549 => x"bb",
         11550 => x"3d",
         11551 => x"33",
         11552 => x"71",
         11553 => x"63",
         11554 => x"58",
         11555 => x"7d",
         11556 => x"fd",
         11557 => x"2e",
         11558 => x"b9",
         11559 => x"7a",
         11560 => x"e2",
         11561 => x"c8",
         11562 => x"b9",
         11563 => x"2e",
         11564 => x"78",
         11565 => x"d8",
         11566 => x"c8",
         11567 => x"3d",
         11568 => x"52",
         11569 => x"bd",
         11570 => x"7f",
         11571 => x"5b",
         11572 => x"2e",
         11573 => x"1f",
         11574 => x"81",
         11575 => x"5f",
         11576 => x"f5",
         11577 => x"56",
         11578 => x"81",
         11579 => x"80",
         11580 => x"7e",
         11581 => x"56",
         11582 => x"e6",
         11583 => x"ff",
         11584 => x"59",
         11585 => x"75",
         11586 => x"76",
         11587 => x"18",
         11588 => x"08",
         11589 => x"af",
         11590 => x"da",
         11591 => x"79",
         11592 => x"77",
         11593 => x"8a",
         11594 => x"84",
         11595 => x"70",
         11596 => x"e5",
         11597 => x"08",
         11598 => x"59",
         11599 => x"7e",
         11600 => x"38",
         11601 => x"17",
         11602 => x"5f",
         11603 => x"38",
         11604 => x"7a",
         11605 => x"38",
         11606 => x"7a",
         11607 => x"76",
         11608 => x"33",
         11609 => x"05",
         11610 => x"17",
         11611 => x"26",
         11612 => x"7c",
         11613 => x"5e",
         11614 => x"2e",
         11615 => x"81",
         11616 => x"59",
         11617 => x"78",
         11618 => x"0c",
         11619 => x"0d",
         11620 => x"33",
         11621 => x"71",
         11622 => x"90",
         11623 => x"07",
         11624 => x"fd",
         11625 => x"16",
         11626 => x"33",
         11627 => x"71",
         11628 => x"79",
         11629 => x"3d",
         11630 => x"80",
         11631 => x"ff",
         11632 => x"84",
         11633 => x"59",
         11634 => x"08",
         11635 => x"96",
         11636 => x"39",
         11637 => x"16",
         11638 => x"16",
         11639 => x"17",
         11640 => x"ff",
         11641 => x"81",
         11642 => x"c8",
         11643 => x"38",
         11644 => x"08",
         11645 => x"b4",
         11646 => x"17",
         11647 => x"b9",
         11648 => x"55",
         11649 => x"08",
         11650 => x"38",
         11651 => x"55",
         11652 => x"09",
         11653 => x"f6",
         11654 => x"b4",
         11655 => x"17",
         11656 => x"7d",
         11657 => x"33",
         11658 => x"b8",
         11659 => x"fb",
         11660 => x"18",
         11661 => x"08",
         11662 => x"af",
         11663 => x"0b",
         11664 => x"33",
         11665 => x"83",
         11666 => x"70",
         11667 => x"43",
         11668 => x"5a",
         11669 => x"09",
         11670 => x"e8",
         11671 => x"39",
         11672 => x"08",
         11673 => x"59",
         11674 => x"7c",
         11675 => x"5e",
         11676 => x"27",
         11677 => x"80",
         11678 => x"18",
         11679 => x"5a",
         11680 => x"70",
         11681 => x"34",
         11682 => x"d4",
         11683 => x"39",
         11684 => x"7c",
         11685 => x"b9",
         11686 => x"e4",
         11687 => x"f7",
         11688 => x"7d",
         11689 => x"56",
         11690 => x"9f",
         11691 => x"54",
         11692 => x"97",
         11693 => x"53",
         11694 => x"8f",
         11695 => x"22",
         11696 => x"59",
         11697 => x"2e",
         11698 => x"80",
         11699 => x"75",
         11700 => x"c2",
         11701 => x"33",
         11702 => x"ba",
         11703 => x"08",
         11704 => x"26",
         11705 => x"94",
         11706 => x"80",
         11707 => x"2e",
         11708 => x"79",
         11709 => x"70",
         11710 => x"5a",
         11711 => x"2e",
         11712 => x"75",
         11713 => x"51",
         11714 => x"3f",
         11715 => x"08",
         11716 => x"54",
         11717 => x"53",
         11718 => x"3f",
         11719 => x"08",
         11720 => x"d5",
         11721 => x"74",
         11722 => x"17",
         11723 => x"31",
         11724 => x"56",
         11725 => x"80",
         11726 => x"38",
         11727 => x"81",
         11728 => x"76",
         11729 => x"08",
         11730 => x"0c",
         11731 => x"70",
         11732 => x"06",
         11733 => x"78",
         11734 => x"fe",
         11735 => x"74",
         11736 => x"f3",
         11737 => x"c8",
         11738 => x"b9",
         11739 => x"2e",
         11740 => x"73",
         11741 => x"38",
         11742 => x"82",
         11743 => x"53",
         11744 => x"08",
         11745 => x"38",
         11746 => x"0c",
         11747 => x"81",
         11748 => x"34",
         11749 => x"84",
         11750 => x"8b",
         11751 => x"90",
         11752 => x"81",
         11753 => x"55",
         11754 => x"bb",
         11755 => x"16",
         11756 => x"80",
         11757 => x"2e",
         11758 => x"fe",
         11759 => x"94",
         11760 => x"15",
         11761 => x"74",
         11762 => x"73",
         11763 => x"90",
         11764 => x"c0",
         11765 => x"90",
         11766 => x"83",
         11767 => x"78",
         11768 => x"38",
         11769 => x"78",
         11770 => x"77",
         11771 => x"80",
         11772 => x"c8",
         11773 => x"0d",
         11774 => x"94",
         11775 => x"15",
         11776 => x"80",
         11777 => x"38",
         11778 => x"0c",
         11779 => x"80",
         11780 => x"a8",
         11781 => x"c8",
         11782 => x"15",
         11783 => x"16",
         11784 => x"ff",
         11785 => x"80",
         11786 => x"79",
         11787 => x"12",
         11788 => x"5a",
         11789 => x"78",
         11790 => x"38",
         11791 => x"74",
         11792 => x"18",
         11793 => x"89",
         11794 => x"5a",
         11795 => x"2e",
         11796 => x"8c",
         11797 => x"fe",
         11798 => x"52",
         11799 => x"89",
         11800 => x"b9",
         11801 => x"fe",
         11802 => x"14",
         11803 => x"82",
         11804 => x"b9",
         11805 => x"06",
         11806 => x"cf",
         11807 => x"08",
         11808 => x"c9",
         11809 => x"74",
         11810 => x"cb",
         11811 => x"c8",
         11812 => x"b9",
         11813 => x"2e",
         11814 => x"b9",
         11815 => x"2e",
         11816 => x"84",
         11817 => x"88",
         11818 => x"98",
         11819 => x"dc",
         11820 => x"91",
         11821 => x"0b",
         11822 => x"0c",
         11823 => x"04",
         11824 => x"7c",
         11825 => x"75",
         11826 => x"38",
         11827 => x"3d",
         11828 => x"8d",
         11829 => x"51",
         11830 => x"84",
         11831 => x"55",
         11832 => x"08",
         11833 => x"38",
         11834 => x"74",
         11835 => x"b9",
         11836 => x"3d",
         11837 => x"76",
         11838 => x"75",
         11839 => x"97",
         11840 => x"c8",
         11841 => x"b9",
         11842 => x"d1",
         11843 => x"33",
         11844 => x"59",
         11845 => x"24",
         11846 => x"16",
         11847 => x"2a",
         11848 => x"54",
         11849 => x"80",
         11850 => x"16",
         11851 => x"33",
         11852 => x"71",
         11853 => x"7d",
         11854 => x"5d",
         11855 => x"78",
         11856 => x"38",
         11857 => x"0c",
         11858 => x"18",
         11859 => x"23",
         11860 => x"51",
         11861 => x"3f",
         11862 => x"08",
         11863 => x"2e",
         11864 => x"80",
         11865 => x"38",
         11866 => x"fe",
         11867 => x"55",
         11868 => x"fe",
         11869 => x"17",
         11870 => x"33",
         11871 => x"71",
         11872 => x"7a",
         11873 => x"0c",
         11874 => x"bc",
         11875 => x"0d",
         11876 => x"54",
         11877 => x"9e",
         11878 => x"53",
         11879 => x"96",
         11880 => x"52",
         11881 => x"8e",
         11882 => x"22",
         11883 => x"57",
         11884 => x"2e",
         11885 => x"52",
         11886 => x"84",
         11887 => x"0c",
         11888 => x"c8",
         11889 => x"0d",
         11890 => x"33",
         11891 => x"c3",
         11892 => x"c8",
         11893 => x"52",
         11894 => x"71",
         11895 => x"54",
         11896 => x"3d",
         11897 => x"58",
         11898 => x"74",
         11899 => x"38",
         11900 => x"73",
         11901 => x"38",
         11902 => x"72",
         11903 => x"38",
         11904 => x"84",
         11905 => x"53",
         11906 => x"81",
         11907 => x"53",
         11908 => x"53",
         11909 => x"38",
         11910 => x"80",
         11911 => x"52",
         11912 => x"9d",
         11913 => x"b9",
         11914 => x"84",
         11915 => x"84",
         11916 => x"84",
         11917 => x"a6",
         11918 => x"74",
         11919 => x"92",
         11920 => x"74",
         11921 => x"be",
         11922 => x"c8",
         11923 => x"70",
         11924 => x"07",
         11925 => x"b9",
         11926 => x"55",
         11927 => x"84",
         11928 => x"8a",
         11929 => x"75",
         11930 => x"52",
         11931 => x"e2",
         11932 => x"74",
         11933 => x"8e",
         11934 => x"c8",
         11935 => x"70",
         11936 => x"07",
         11937 => x"b9",
         11938 => x"55",
         11939 => x"39",
         11940 => x"51",
         11941 => x"3f",
         11942 => x"08",
         11943 => x"0c",
         11944 => x"04",
         11945 => x"51",
         11946 => x"3f",
         11947 => x"08",
         11948 => x"72",
         11949 => x"72",
         11950 => x"56",
         11951 => x"ed",
         11952 => x"57",
         11953 => x"3d",
         11954 => x"3d",
         11955 => x"a5",
         11956 => x"c8",
         11957 => x"b9",
         11958 => x"2e",
         11959 => x"84",
         11960 => x"95",
         11961 => x"65",
         11962 => x"ff",
         11963 => x"84",
         11964 => x"55",
         11965 => x"08",
         11966 => x"80",
         11967 => x"70",
         11968 => x"58",
         11969 => x"97",
         11970 => x"2e",
         11971 => x"52",
         11972 => x"b0",
         11973 => x"84",
         11974 => x"95",
         11975 => x"86",
         11976 => x"c8",
         11977 => x"0d",
         11978 => x"0d",
         11979 => x"5f",
         11980 => x"3d",
         11981 => x"96",
         11982 => x"b9",
         11983 => x"c8",
         11984 => x"b9",
         11985 => x"38",
         11986 => x"74",
         11987 => x"08",
         11988 => x"13",
         11989 => x"59",
         11990 => x"26",
         11991 => x"7f",
         11992 => x"b9",
         11993 => x"3d",
         11994 => x"b9",
         11995 => x"33",
         11996 => x"81",
         11997 => x"38",
         11998 => x"08",
         11999 => x"08",
         12000 => x"77",
         12001 => x"7b",
         12002 => x"5c",
         12003 => x"17",
         12004 => x"82",
         12005 => x"17",
         12006 => x"5d",
         12007 => x"38",
         12008 => x"53",
         12009 => x"81",
         12010 => x"fe",
         12011 => x"84",
         12012 => x"80",
         12013 => x"ff",
         12014 => x"79",
         12015 => x"7f",
         12016 => x"7d",
         12017 => x"76",
         12018 => x"82",
         12019 => x"38",
         12020 => x"05",
         12021 => x"82",
         12022 => x"90",
         12023 => x"2b",
         12024 => x"33",
         12025 => x"88",
         12026 => x"71",
         12027 => x"fe",
         12028 => x"70",
         12029 => x"25",
         12030 => x"84",
         12031 => x"06",
         12032 => x"43",
         12033 => x"54",
         12034 => x"40",
         12035 => x"fe",
         12036 => x"7f",
         12037 => x"18",
         12038 => x"33",
         12039 => x"77",
         12040 => x"79",
         12041 => x"0c",
         12042 => x"04",
         12043 => x"17",
         12044 => x"17",
         12045 => x"18",
         12046 => x"fe",
         12047 => x"81",
         12048 => x"c8",
         12049 => x"38",
         12050 => x"08",
         12051 => x"b4",
         12052 => x"18",
         12053 => x"b9",
         12054 => x"55",
         12055 => x"08",
         12056 => x"38",
         12057 => x"55",
         12058 => x"09",
         12059 => x"b0",
         12060 => x"b4",
         12061 => x"18",
         12062 => x"7c",
         12063 => x"33",
         12064 => x"e0",
         12065 => x"fe",
         12066 => x"77",
         12067 => x"59",
         12068 => x"77",
         12069 => x"80",
         12070 => x"c8",
         12071 => x"80",
         12072 => x"b9",
         12073 => x"2e",
         12074 => x"84",
         12075 => x"30",
         12076 => x"c8",
         12077 => x"25",
         12078 => x"18",
         12079 => x"5c",
         12080 => x"08",
         12081 => x"38",
         12082 => x"7a",
         12083 => x"84",
         12084 => x"07",
         12085 => x"18",
         12086 => x"39",
         12087 => x"05",
         12088 => x"71",
         12089 => x"2b",
         12090 => x"70",
         12091 => x"82",
         12092 => x"06",
         12093 => x"5d",
         12094 => x"5f",
         12095 => x"83",
         12096 => x"39",
         12097 => x"bf",
         12098 => x"58",
         12099 => x"0c",
         12100 => x"0c",
         12101 => x"81",
         12102 => x"84",
         12103 => x"83",
         12104 => x"58",
         12105 => x"f7",
         12106 => x"57",
         12107 => x"80",
         12108 => x"76",
         12109 => x"80",
         12110 => x"74",
         12111 => x"80",
         12112 => x"86",
         12113 => x"18",
         12114 => x"78",
         12115 => x"da",
         12116 => x"73",
         12117 => x"dc",
         12118 => x"33",
         12119 => x"d4",
         12120 => x"33",
         12121 => x"81",
         12122 => x"87",
         12123 => x"2e",
         12124 => x"94",
         12125 => x"73",
         12126 => x"27",
         12127 => x"81",
         12128 => x"17",
         12129 => x"57",
         12130 => x"27",
         12131 => x"16",
         12132 => x"b3",
         12133 => x"80",
         12134 => x"0c",
         12135 => x"8c",
         12136 => x"80",
         12137 => x"78",
         12138 => x"75",
         12139 => x"38",
         12140 => x"34",
         12141 => x"84",
         12142 => x"8b",
         12143 => x"78",
         12144 => x"27",
         12145 => x"73",
         12146 => x"fe",
         12147 => x"84",
         12148 => x"59",
         12149 => x"08",
         12150 => x"e9",
         12151 => x"c8",
         12152 => x"82",
         12153 => x"b9",
         12154 => x"2e",
         12155 => x"80",
         12156 => x"75",
         12157 => x"81",
         12158 => x"c8",
         12159 => x"38",
         12160 => x"fe",
         12161 => x"08",
         12162 => x"74",
         12163 => x"af",
         12164 => x"94",
         12165 => x"16",
         12166 => x"54",
         12167 => x"34",
         12168 => x"79",
         12169 => x"38",
         12170 => x"15",
         12171 => x"f6",
         12172 => x"b9",
         12173 => x"06",
         12174 => x"95",
         12175 => x"08",
         12176 => x"8f",
         12177 => x"90",
         12178 => x"54",
         12179 => x"0b",
         12180 => x"fe",
         12181 => x"17",
         12182 => x"51",
         12183 => x"3f",
         12184 => x"08",
         12185 => x"c2",
         12186 => x"c8",
         12187 => x"81",
         12188 => x"81",
         12189 => x"58",
         12190 => x"08",
         12191 => x"27",
         12192 => x"84",
         12193 => x"98",
         12194 => x"08",
         12195 => x"81",
         12196 => x"c8",
         12197 => x"a1",
         12198 => x"c8",
         12199 => x"08",
         12200 => x"38",
         12201 => x"97",
         12202 => x"74",
         12203 => x"ff",
         12204 => x"84",
         12205 => x"55",
         12206 => x"08",
         12207 => x"73",
         12208 => x"fe",
         12209 => x"84",
         12210 => x"59",
         12211 => x"08",
         12212 => x"cb",
         12213 => x"c8",
         12214 => x"80",
         12215 => x"b9",
         12216 => x"2e",
         12217 => x"80",
         12218 => x"75",
         12219 => x"89",
         12220 => x"c8",
         12221 => x"38",
         12222 => x"fe",
         12223 => x"08",
         12224 => x"74",
         12225 => x"38",
         12226 => x"17",
         12227 => x"33",
         12228 => x"73",
         12229 => x"78",
         12230 => x"26",
         12231 => x"80",
         12232 => x"90",
         12233 => x"fc",
         12234 => x"56",
         12235 => x"82",
         12236 => x"33",
         12237 => x"e4",
         12238 => x"e7",
         12239 => x"90",
         12240 => x"54",
         12241 => x"84",
         12242 => x"90",
         12243 => x"54",
         12244 => x"81",
         12245 => x"33",
         12246 => x"f0",
         12247 => x"c8",
         12248 => x"39",
         12249 => x"bb",
         12250 => x"0d",
         12251 => x"3d",
         12252 => x"52",
         12253 => x"ff",
         12254 => x"84",
         12255 => x"56",
         12256 => x"08",
         12257 => x"38",
         12258 => x"c8",
         12259 => x"0d",
         12260 => x"a8",
         12261 => x"9b",
         12262 => x"59",
         12263 => x"3f",
         12264 => x"08",
         12265 => x"c8",
         12266 => x"02",
         12267 => x"33",
         12268 => x"81",
         12269 => x"86",
         12270 => x"38",
         12271 => x"5b",
         12272 => x"c4",
         12273 => x"ee",
         12274 => x"81",
         12275 => x"87",
         12276 => x"b4",
         12277 => x"3d",
         12278 => x"33",
         12279 => x"71",
         12280 => x"73",
         12281 => x"5c",
         12282 => x"83",
         12283 => x"38",
         12284 => x"81",
         12285 => x"80",
         12286 => x"38",
         12287 => x"18",
         12288 => x"ff",
         12289 => x"5f",
         12290 => x"b9",
         12291 => x"8f",
         12292 => x"55",
         12293 => x"3f",
         12294 => x"08",
         12295 => x"c8",
         12296 => x"38",
         12297 => x"08",
         12298 => x"ff",
         12299 => x"84",
         12300 => x"56",
         12301 => x"08",
         12302 => x"0b",
         12303 => x"0c",
         12304 => x"04",
         12305 => x"94",
         12306 => x"98",
         12307 => x"2b",
         12308 => x"5d",
         12309 => x"98",
         12310 => x"c8",
         12311 => x"88",
         12312 => x"c8",
         12313 => x"38",
         12314 => x"a8",
         12315 => x"5d",
         12316 => x"2e",
         12317 => x"74",
         12318 => x"ff",
         12319 => x"84",
         12320 => x"56",
         12321 => x"08",
         12322 => x"38",
         12323 => x"77",
         12324 => x"56",
         12325 => x"2e",
         12326 => x"80",
         12327 => x"7a",
         12328 => x"55",
         12329 => x"89",
         12330 => x"08",
         12331 => x"fd",
         12332 => x"75",
         12333 => x"7d",
         12334 => x"db",
         12335 => x"c8",
         12336 => x"c8",
         12337 => x"0d",
         12338 => x"5d",
         12339 => x"56",
         12340 => x"17",
         12341 => x"82",
         12342 => x"17",
         12343 => x"55",
         12344 => x"09",
         12345 => x"dd",
         12346 => x"75",
         12347 => x"52",
         12348 => x"51",
         12349 => x"3f",
         12350 => x"08",
         12351 => x"38",
         12352 => x"58",
         12353 => x"0c",
         12354 => x"ab",
         12355 => x"08",
         12356 => x"34",
         12357 => x"18",
         12358 => x"08",
         12359 => x"ec",
         12360 => x"78",
         12361 => x"de",
         12362 => x"c8",
         12363 => x"b9",
         12364 => x"2e",
         12365 => x"75",
         12366 => x"81",
         12367 => x"38",
         12368 => x"c8",
         12369 => x"b4",
         12370 => x"7c",
         12371 => x"33",
         12372 => x"90",
         12373 => x"84",
         12374 => x"7a",
         12375 => x"06",
         12376 => x"84",
         12377 => x"83",
         12378 => x"17",
         12379 => x"08",
         12380 => x"c8",
         12381 => x"74",
         12382 => x"27",
         12383 => x"82",
         12384 => x"74",
         12385 => x"81",
         12386 => x"38",
         12387 => x"17",
         12388 => x"08",
         12389 => x"52",
         12390 => x"51",
         12391 => x"3f",
         12392 => x"c5",
         12393 => x"79",
         12394 => x"e1",
         12395 => x"78",
         12396 => x"e4",
         12397 => x"c8",
         12398 => x"b9",
         12399 => x"2e",
         12400 => x"84",
         12401 => x"81",
         12402 => x"38",
         12403 => x"08",
         12404 => x"cb",
         12405 => x"74",
         12406 => x"fe",
         12407 => x"84",
         12408 => x"b3",
         12409 => x"08",
         12410 => x"19",
         12411 => x"58",
         12412 => x"ff",
         12413 => x"16",
         12414 => x"84",
         12415 => x"07",
         12416 => x"18",
         12417 => x"77",
         12418 => x"a1",
         12419 => x"fd",
         12420 => x"56",
         12421 => x"84",
         12422 => x"56",
         12423 => x"81",
         12424 => x"39",
         12425 => x"82",
         12426 => x"ff",
         12427 => x"a0",
         12428 => x"b2",
         12429 => x"b9",
         12430 => x"84",
         12431 => x"80",
         12432 => x"75",
         12433 => x"0c",
         12434 => x"04",
         12435 => x"52",
         12436 => x"52",
         12437 => x"bf",
         12438 => x"c8",
         12439 => x"b9",
         12440 => x"38",
         12441 => x"b9",
         12442 => x"3d",
         12443 => x"b9",
         12444 => x"2e",
         12445 => x"cb",
         12446 => x"f3",
         12447 => x"85",
         12448 => x"56",
         12449 => x"74",
         12450 => x"7d",
         12451 => x"8f",
         12452 => x"5d",
         12453 => x"3f",
         12454 => x"08",
         12455 => x"84",
         12456 => x"83",
         12457 => x"84",
         12458 => x"81",
         12459 => x"38",
         12460 => x"08",
         12461 => x"cb",
         12462 => x"c9",
         12463 => x"b9",
         12464 => x"12",
         12465 => x"57",
         12466 => x"38",
         12467 => x"18",
         12468 => x"5a",
         12469 => x"75",
         12470 => x"38",
         12471 => x"76",
         12472 => x"19",
         12473 => x"58",
         12474 => x"0c",
         12475 => x"84",
         12476 => x"55",
         12477 => x"81",
         12478 => x"ff",
         12479 => x"f4",
         12480 => x"8a",
         12481 => x"77",
         12482 => x"f9",
         12483 => x"77",
         12484 => x"52",
         12485 => x"51",
         12486 => x"3f",
         12487 => x"08",
         12488 => x"81",
         12489 => x"39",
         12490 => x"84",
         12491 => x"b4",
         12492 => x"b8",
         12493 => x"81",
         12494 => x"58",
         12495 => x"3f",
         12496 => x"b9",
         12497 => x"38",
         12498 => x"08",
         12499 => x"b4",
         12500 => x"18",
         12501 => x"74",
         12502 => x"27",
         12503 => x"82",
         12504 => x"7a",
         12505 => x"81",
         12506 => x"38",
         12507 => x"17",
         12508 => x"08",
         12509 => x"52",
         12510 => x"51",
         12511 => x"3f",
         12512 => x"81",
         12513 => x"08",
         12514 => x"7c",
         12515 => x"38",
         12516 => x"08",
         12517 => x"38",
         12518 => x"51",
         12519 => x"3f",
         12520 => x"08",
         12521 => x"c8",
         12522 => x"fd",
         12523 => x"b9",
         12524 => x"2e",
         12525 => x"84",
         12526 => x"ff",
         12527 => x"38",
         12528 => x"52",
         12529 => x"f9",
         12530 => x"b9",
         12531 => x"f3",
         12532 => x"08",
         12533 => x"19",
         12534 => x"59",
         12535 => x"90",
         12536 => x"94",
         12537 => x"17",
         12538 => x"5c",
         12539 => x"34",
         12540 => x"7a",
         12541 => x"38",
         12542 => x"c8",
         12543 => x"0d",
         12544 => x"22",
         12545 => x"ff",
         12546 => x"81",
         12547 => x"2e",
         12548 => x"fe",
         12549 => x"0b",
         12550 => x"56",
         12551 => x"81",
         12552 => x"ff",
         12553 => x"f4",
         12554 => x"ae",
         12555 => x"34",
         12556 => x"0b",
         12557 => x"34",
         12558 => x"80",
         12559 => x"75",
         12560 => x"34",
         12561 => x"d0",
         12562 => x"cc",
         12563 => x"1a",
         12564 => x"83",
         12565 => x"59",
         12566 => x"d2",
         12567 => x"88",
         12568 => x"80",
         12569 => x"75",
         12570 => x"83",
         12571 => x"38",
         12572 => x"0b",
         12573 => x"b8",
         12574 => x"56",
         12575 => x"05",
         12576 => x"70",
         12577 => x"34",
         12578 => x"75",
         12579 => x"56",
         12580 => x"d9",
         12581 => x"7e",
         12582 => x"ff",
         12583 => x"57",
         12584 => x"17",
         12585 => x"2a",
         12586 => x"f3",
         12587 => x"33",
         12588 => x"2e",
         12589 => x"7d",
         12590 => x"83",
         12591 => x"51",
         12592 => x"3f",
         12593 => x"08",
         12594 => x"c8",
         12595 => x"38",
         12596 => x"b9",
         12597 => x"17",
         12598 => x"c8",
         12599 => x"34",
         12600 => x"17",
         12601 => x"0b",
         12602 => x"7d",
         12603 => x"77",
         12604 => x"77",
         12605 => x"78",
         12606 => x"7c",
         12607 => x"83",
         12608 => x"38",
         12609 => x"0b",
         12610 => x"7d",
         12611 => x"83",
         12612 => x"51",
         12613 => x"3f",
         12614 => x"08",
         12615 => x"b9",
         12616 => x"3d",
         12617 => x"90",
         12618 => x"80",
         12619 => x"74",
         12620 => x"76",
         12621 => x"34",
         12622 => x"7b",
         12623 => x"7a",
         12624 => x"34",
         12625 => x"55",
         12626 => x"17",
         12627 => x"a0",
         12628 => x"1a",
         12629 => x"58",
         12630 => x"39",
         12631 => x"58",
         12632 => x"34",
         12633 => x"5c",
         12634 => x"34",
         12635 => x"0b",
         12636 => x"7d",
         12637 => x"83",
         12638 => x"51",
         12639 => x"3f",
         12640 => x"08",
         12641 => x"39",
         12642 => x"b3",
         12643 => x"08",
         12644 => x"5f",
         12645 => x"9b",
         12646 => x"81",
         12647 => x"70",
         12648 => x"56",
         12649 => x"81",
         12650 => x"ed",
         12651 => x"2e",
         12652 => x"82",
         12653 => x"fe",
         12654 => x"b2",
         12655 => x"ab",
         12656 => x"b9",
         12657 => x"84",
         12658 => x"80",
         12659 => x"75",
         12660 => x"0c",
         12661 => x"04",
         12662 => x"0c",
         12663 => x"52",
         12664 => x"52",
         12665 => x"af",
         12666 => x"c8",
         12667 => x"b9",
         12668 => x"38",
         12669 => x"05",
         12670 => x"06",
         12671 => x"7c",
         12672 => x"0b",
         12673 => x"3d",
         12674 => x"55",
         12675 => x"05",
         12676 => x"70",
         12677 => x"34",
         12678 => x"74",
         12679 => x"3d",
         12680 => x"7a",
         12681 => x"75",
         12682 => x"57",
         12683 => x"81",
         12684 => x"ff",
         12685 => x"ef",
         12686 => x"08",
         12687 => x"ff",
         12688 => x"84",
         12689 => x"56",
         12690 => x"08",
         12691 => x"6a",
         12692 => x"2e",
         12693 => x"88",
         12694 => x"c8",
         12695 => x"0d",
         12696 => x"d0",
         12697 => x"ff",
         12698 => x"58",
         12699 => x"91",
         12700 => x"78",
         12701 => x"d0",
         12702 => x"78",
         12703 => x"fa",
         12704 => x"08",
         12705 => x"70",
         12706 => x"5e",
         12707 => x"7a",
         12708 => x"5c",
         12709 => x"81",
         12710 => x"ff",
         12711 => x"58",
         12712 => x"26",
         12713 => x"16",
         12714 => x"06",
         12715 => x"9f",
         12716 => x"99",
         12717 => x"e0",
         12718 => x"ff",
         12719 => x"75",
         12720 => x"2a",
         12721 => x"77",
         12722 => x"06",
         12723 => x"ff",
         12724 => x"7a",
         12725 => x"70",
         12726 => x"2a",
         12727 => x"58",
         12728 => x"2e",
         12729 => x"1c",
         12730 => x"5c",
         12731 => x"fd",
         12732 => x"08",
         12733 => x"ff",
         12734 => x"83",
         12735 => x"38",
         12736 => x"82",
         12737 => x"fe",
         12738 => x"b2",
         12739 => x"a8",
         12740 => x"b9",
         12741 => x"84",
         12742 => x"fd",
         12743 => x"b8",
         12744 => x"3d",
         12745 => x"81",
         12746 => x"38",
         12747 => x"8d",
         12748 => x"b9",
         12749 => x"84",
         12750 => x"fd",
         12751 => x"58",
         12752 => x"19",
         12753 => x"80",
         12754 => x"56",
         12755 => x"81",
         12756 => x"75",
         12757 => x"57",
         12758 => x"5a",
         12759 => x"02",
         12760 => x"33",
         12761 => x"8b",
         12762 => x"84",
         12763 => x"40",
         12764 => x"38",
         12765 => x"57",
         12766 => x"34",
         12767 => x"0b",
         12768 => x"8b",
         12769 => x"84",
         12770 => x"57",
         12771 => x"2e",
         12772 => x"a7",
         12773 => x"2e",
         12774 => x"7f",
         12775 => x"9a",
         12776 => x"88",
         12777 => x"33",
         12778 => x"57",
         12779 => x"82",
         12780 => x"16",
         12781 => x"fe",
         12782 => x"75",
         12783 => x"c7",
         12784 => x"22",
         12785 => x"b0",
         12786 => x"57",
         12787 => x"2e",
         12788 => x"75",
         12789 => x"b4",
         12790 => x"2e",
         12791 => x"17",
         12792 => x"83",
         12793 => x"54",
         12794 => x"17",
         12795 => x"33",
         12796 => x"f1",
         12797 => x"c8",
         12798 => x"85",
         12799 => x"81",
         12800 => x"18",
         12801 => x"7b",
         12802 => x"56",
         12803 => x"bf",
         12804 => x"33",
         12805 => x"2e",
         12806 => x"bb",
         12807 => x"83",
         12808 => x"5d",
         12809 => x"f2",
         12810 => x"88",
         12811 => x"80",
         12812 => x"76",
         12813 => x"83",
         12814 => x"06",
         12815 => x"90",
         12816 => x"80",
         12817 => x"7d",
         12818 => x"75",
         12819 => x"34",
         12820 => x"0b",
         12821 => x"78",
         12822 => x"08",
         12823 => x"57",
         12824 => x"ff",
         12825 => x"74",
         12826 => x"fe",
         12827 => x"84",
         12828 => x"55",
         12829 => x"08",
         12830 => x"b8",
         12831 => x"19",
         12832 => x"5a",
         12833 => x"77",
         12834 => x"83",
         12835 => x"59",
         12836 => x"2e",
         12837 => x"81",
         12838 => x"54",
         12839 => x"16",
         12840 => x"33",
         12841 => x"bd",
         12842 => x"c8",
         12843 => x"85",
         12844 => x"81",
         12845 => x"17",
         12846 => x"77",
         12847 => x"19",
         12848 => x"7a",
         12849 => x"83",
         12850 => x"19",
         12851 => x"a5",
         12852 => x"78",
         12853 => x"ae",
         12854 => x"c8",
         12855 => x"b9",
         12856 => x"2e",
         12857 => x"82",
         12858 => x"2e",
         12859 => x"74",
         12860 => x"db",
         12861 => x"fe",
         12862 => x"84",
         12863 => x"84",
         12864 => x"b1",
         12865 => x"82",
         12866 => x"c8",
         12867 => x"0d",
         12868 => x"33",
         12869 => x"71",
         12870 => x"90",
         12871 => x"07",
         12872 => x"fd",
         12873 => x"b9",
         12874 => x"2e",
         12875 => x"84",
         12876 => x"80",
         12877 => x"38",
         12878 => x"c8",
         12879 => x"0d",
         12880 => x"b4",
         12881 => x"7b",
         12882 => x"33",
         12883 => x"94",
         12884 => x"84",
         12885 => x"7a",
         12886 => x"06",
         12887 => x"84",
         12888 => x"83",
         12889 => x"16",
         12890 => x"08",
         12891 => x"c8",
         12892 => x"74",
         12893 => x"27",
         12894 => x"82",
         12895 => x"7c",
         12896 => x"81",
         12897 => x"38",
         12898 => x"16",
         12899 => x"08",
         12900 => x"52",
         12901 => x"51",
         12902 => x"3f",
         12903 => x"fa",
         12904 => x"b4",
         12905 => x"b8",
         12906 => x"81",
         12907 => x"5b",
         12908 => x"3f",
         12909 => x"b9",
         12910 => x"c9",
         12911 => x"c8",
         12912 => x"34",
         12913 => x"a8",
         12914 => x"84",
         12915 => x"5d",
         12916 => x"18",
         12917 => x"8e",
         12918 => x"33",
         12919 => x"2e",
         12920 => x"fc",
         12921 => x"54",
         12922 => x"a0",
         12923 => x"53",
         12924 => x"17",
         12925 => x"e0",
         12926 => x"5c",
         12927 => x"ec",
         12928 => x"80",
         12929 => x"02",
         12930 => x"e3",
         12931 => x"57",
         12932 => x"3d",
         12933 => x"97",
         12934 => x"a2",
         12935 => x"b9",
         12936 => x"84",
         12937 => x"80",
         12938 => x"75",
         12939 => x"0c",
         12940 => x"04",
         12941 => x"52",
         12942 => x"05",
         12943 => x"d7",
         12944 => x"c8",
         12945 => x"b9",
         12946 => x"38",
         12947 => x"05",
         12948 => x"06",
         12949 => x"73",
         12950 => x"a7",
         12951 => x"09",
         12952 => x"71",
         12953 => x"06",
         12954 => x"57",
         12955 => x"17",
         12956 => x"81",
         12957 => x"34",
         12958 => x"e2",
         12959 => x"b9",
         12960 => x"b9",
         12961 => x"3d",
         12962 => x"3d",
         12963 => x"82",
         12964 => x"cc",
         12965 => x"3d",
         12966 => x"d9",
         12967 => x"c8",
         12968 => x"b9",
         12969 => x"2e",
         12970 => x"84",
         12971 => x"96",
         12972 => x"78",
         12973 => x"96",
         12974 => x"51",
         12975 => x"3f",
         12976 => x"08",
         12977 => x"c8",
         12978 => x"02",
         12979 => x"33",
         12980 => x"56",
         12981 => x"d2",
         12982 => x"18",
         12983 => x"22",
         12984 => x"07",
         12985 => x"76",
         12986 => x"76",
         12987 => x"74",
         12988 => x"76",
         12989 => x"77",
         12990 => x"76",
         12991 => x"73",
         12992 => x"78",
         12993 => x"83",
         12994 => x"51",
         12995 => x"3f",
         12996 => x"08",
         12997 => x"0c",
         12998 => x"04",
         12999 => x"6b",
         13000 => x"80",
         13001 => x"cc",
         13002 => x"3d",
         13003 => x"c5",
         13004 => x"c8",
         13005 => x"c8",
         13006 => x"84",
         13007 => x"07",
         13008 => x"56",
         13009 => x"2e",
         13010 => x"70",
         13011 => x"56",
         13012 => x"38",
         13013 => x"78",
         13014 => x"56",
         13015 => x"2e",
         13016 => x"81",
         13017 => x"5a",
         13018 => x"2e",
         13019 => x"7c",
         13020 => x"58",
         13021 => x"b4",
         13022 => x"2e",
         13023 => x"83",
         13024 => x"5a",
         13025 => x"2e",
         13026 => x"81",
         13027 => x"54",
         13028 => x"16",
         13029 => x"33",
         13030 => x"c9",
         13031 => x"c8",
         13032 => x"85",
         13033 => x"81",
         13034 => x"17",
         13035 => x"78",
         13036 => x"70",
         13037 => x"80",
         13038 => x"83",
         13039 => x"80",
         13040 => x"84",
         13041 => x"a7",
         13042 => x"b8",
         13043 => x"33",
         13044 => x"71",
         13045 => x"88",
         13046 => x"14",
         13047 => x"07",
         13048 => x"33",
         13049 => x"0c",
         13050 => x"57",
         13051 => x"84",
         13052 => x"9a",
         13053 => x"7c",
         13054 => x"80",
         13055 => x"70",
         13056 => x"f4",
         13057 => x"b9",
         13058 => x"84",
         13059 => x"80",
         13060 => x"38",
         13061 => x"09",
         13062 => x"b8",
         13063 => x"34",
         13064 => x"b0",
         13065 => x"b4",
         13066 => x"b8",
         13067 => x"81",
         13068 => x"5b",
         13069 => x"3f",
         13070 => x"b9",
         13071 => x"2e",
         13072 => x"fe",
         13073 => x"b9",
         13074 => x"17",
         13075 => x"08",
         13076 => x"31",
         13077 => x"08",
         13078 => x"a0",
         13079 => x"fe",
         13080 => x"16",
         13081 => x"82",
         13082 => x"06",
         13083 => x"77",
         13084 => x"08",
         13085 => x"05",
         13086 => x"81",
         13087 => x"fe",
         13088 => x"79",
         13089 => x"76",
         13090 => x"52",
         13091 => x"51",
         13092 => x"3f",
         13093 => x"08",
         13094 => x"8d",
         13095 => x"39",
         13096 => x"51",
         13097 => x"3f",
         13098 => x"08",
         13099 => x"c8",
         13100 => x"38",
         13101 => x"08",
         13102 => x"08",
         13103 => x"59",
         13104 => x"19",
         13105 => x"59",
         13106 => x"75",
         13107 => x"59",
         13108 => x"ec",
         13109 => x"1c",
         13110 => x"76",
         13111 => x"2e",
         13112 => x"ff",
         13113 => x"70",
         13114 => x"58",
         13115 => x"ea",
         13116 => x"39",
         13117 => x"ba",
         13118 => x"0d",
         13119 => x"3d",
         13120 => x"52",
         13121 => x"ff",
         13122 => x"84",
         13123 => x"56",
         13124 => x"08",
         13125 => x"8f",
         13126 => x"7d",
         13127 => x"76",
         13128 => x"58",
         13129 => x"55",
         13130 => x"74",
         13131 => x"70",
         13132 => x"ff",
         13133 => x"58",
         13134 => x"27",
         13135 => x"a2",
         13136 => x"5c",
         13137 => x"ff",
         13138 => x"57",
         13139 => x"f5",
         13140 => x"0c",
         13141 => x"ff",
         13142 => x"38",
         13143 => x"95",
         13144 => x"52",
         13145 => x"08",
         13146 => x"3f",
         13147 => x"08",
         13148 => x"06",
         13149 => x"2e",
         13150 => x"83",
         13151 => x"83",
         13152 => x"70",
         13153 => x"5b",
         13154 => x"80",
         13155 => x"38",
         13156 => x"77",
         13157 => x"81",
         13158 => x"70",
         13159 => x"57",
         13160 => x"80",
         13161 => x"74",
         13162 => x"81",
         13163 => x"75",
         13164 => x"59",
         13165 => x"38",
         13166 => x"27",
         13167 => x"79",
         13168 => x"96",
         13169 => x"77",
         13170 => x"76",
         13171 => x"74",
         13172 => x"05",
         13173 => x"1a",
         13174 => x"70",
         13175 => x"34",
         13176 => x"3d",
         13177 => x"70",
         13178 => x"5b",
         13179 => x"77",
         13180 => x"d1",
         13181 => x"33",
         13182 => x"76",
         13183 => x"bc",
         13184 => x"2e",
         13185 => x"b7",
         13186 => x"16",
         13187 => x"5c",
         13188 => x"09",
         13189 => x"38",
         13190 => x"79",
         13191 => x"45",
         13192 => x"52",
         13193 => x"52",
         13194 => x"e4",
         13195 => x"c8",
         13196 => x"b9",
         13197 => x"2e",
         13198 => x"56",
         13199 => x"c8",
         13200 => x"0d",
         13201 => x"52",
         13202 => x"e7",
         13203 => x"c8",
         13204 => x"ff",
         13205 => x"fd",
         13206 => x"56",
         13207 => x"c8",
         13208 => x"0d",
         13209 => x"d8",
         13210 => x"c3",
         13211 => x"75",
         13212 => x"ee",
         13213 => x"c8",
         13214 => x"b9",
         13215 => x"c1",
         13216 => x"2e",
         13217 => x"8b",
         13218 => x"57",
         13219 => x"81",
         13220 => x"76",
         13221 => x"58",
         13222 => x"55",
         13223 => x"7d",
         13224 => x"83",
         13225 => x"51",
         13226 => x"3f",
         13227 => x"08",
         13228 => x"ff",
         13229 => x"7a",
         13230 => x"38",
         13231 => x"9c",
         13232 => x"c8",
         13233 => x"09",
         13234 => x"ee",
         13235 => x"79",
         13236 => x"e6",
         13237 => x"75",
         13238 => x"58",
         13239 => x"3f",
         13240 => x"08",
         13241 => x"c8",
         13242 => x"09",
         13243 => x"84",
         13244 => x"c8",
         13245 => x"5c",
         13246 => x"08",
         13247 => x"b4",
         13248 => x"2e",
         13249 => x"18",
         13250 => x"79",
         13251 => x"06",
         13252 => x"81",
         13253 => x"b8",
         13254 => x"18",
         13255 => x"d5",
         13256 => x"b9",
         13257 => x"2e",
         13258 => x"57",
         13259 => x"b4",
         13260 => x"57",
         13261 => x"78",
         13262 => x"70",
         13263 => x"57",
         13264 => x"2e",
         13265 => x"74",
         13266 => x"25",
         13267 => x"5c",
         13268 => x"81",
         13269 => x"1a",
         13270 => x"2e",
         13271 => x"52",
         13272 => x"ef",
         13273 => x"b9",
         13274 => x"84",
         13275 => x"80",
         13276 => x"38",
         13277 => x"84",
         13278 => x"38",
         13279 => x"fd",
         13280 => x"6c",
         13281 => x"76",
         13282 => x"58",
         13283 => x"55",
         13284 => x"6b",
         13285 => x"8b",
         13286 => x"6c",
         13287 => x"55",
         13288 => x"05",
         13289 => x"70",
         13290 => x"34",
         13291 => x"74",
         13292 => x"eb",
         13293 => x"81",
         13294 => x"76",
         13295 => x"58",
         13296 => x"55",
         13297 => x"fd",
         13298 => x"5a",
         13299 => x"7d",
         13300 => x"83",
         13301 => x"51",
         13302 => x"3f",
         13303 => x"08",
         13304 => x"39",
         13305 => x"df",
         13306 => x"b4",
         13307 => x"7a",
         13308 => x"33",
         13309 => x"ec",
         13310 => x"c8",
         13311 => x"09",
         13312 => x"c3",
         13313 => x"c8",
         13314 => x"34",
         13315 => x"a8",
         13316 => x"5c",
         13317 => x"08",
         13318 => x"82",
         13319 => x"74",
         13320 => x"38",
         13321 => x"08",
         13322 => x"39",
         13323 => x"52",
         13324 => x"ed",
         13325 => x"b9",
         13326 => x"84",
         13327 => x"80",
         13328 => x"38",
         13329 => x"81",
         13330 => x"78",
         13331 => x"e7",
         13332 => x"39",
         13333 => x"18",
         13334 => x"08",
         13335 => x"52",
         13336 => x"51",
         13337 => x"3f",
         13338 => x"f2",
         13339 => x"62",
         13340 => x"80",
         13341 => x"5e",
         13342 => x"56",
         13343 => x"9f",
         13344 => x"55",
         13345 => x"97",
         13346 => x"54",
         13347 => x"8f",
         13348 => x"22",
         13349 => x"59",
         13350 => x"2e",
         13351 => x"80",
         13352 => x"75",
         13353 => x"91",
         13354 => x"75",
         13355 => x"79",
         13356 => x"a2",
         13357 => x"08",
         13358 => x"90",
         13359 => x"81",
         13360 => x"56",
         13361 => x"2e",
         13362 => x"7e",
         13363 => x"70",
         13364 => x"55",
         13365 => x"5c",
         13366 => x"cb",
         13367 => x"7a",
         13368 => x"70",
         13369 => x"2a",
         13370 => x"08",
         13371 => x"08",
         13372 => x"5f",
         13373 => x"78",
         13374 => x"9c",
         13375 => x"26",
         13376 => x"58",
         13377 => x"5b",
         13378 => x"52",
         13379 => x"d8",
         13380 => x"15",
         13381 => x"9c",
         13382 => x"26",
         13383 => x"55",
         13384 => x"08",
         13385 => x"dc",
         13386 => x"c8",
         13387 => x"81",
         13388 => x"b9",
         13389 => x"c5",
         13390 => x"59",
         13391 => x"bb",
         13392 => x"2e",
         13393 => x"c2",
         13394 => x"75",
         13395 => x"b9",
         13396 => x"3d",
         13397 => x"0b",
         13398 => x"0c",
         13399 => x"04",
         13400 => x"51",
         13401 => x"3f",
         13402 => x"08",
         13403 => x"73",
         13404 => x"73",
         13405 => x"56",
         13406 => x"7b",
         13407 => x"8e",
         13408 => x"56",
         13409 => x"2e",
         13410 => x"18",
         13411 => x"2e",
         13412 => x"73",
         13413 => x"7e",
         13414 => x"dd",
         13415 => x"c8",
         13416 => x"b9",
         13417 => x"a3",
         13418 => x"19",
         13419 => x"59",
         13420 => x"38",
         13421 => x"12",
         13422 => x"80",
         13423 => x"38",
         13424 => x"0c",
         13425 => x"0c",
         13426 => x"80",
         13427 => x"7b",
         13428 => x"9c",
         13429 => x"05",
         13430 => x"58",
         13431 => x"26",
         13432 => x"76",
         13433 => x"16",
         13434 => x"33",
         13435 => x"7c",
         13436 => x"75",
         13437 => x"39",
         13438 => x"97",
         13439 => x"80",
         13440 => x"39",
         13441 => x"c5",
         13442 => x"fe",
         13443 => x"1b",
         13444 => x"39",
         13445 => x"08",
         13446 => x"a3",
         13447 => x"3d",
         13448 => x"05",
         13449 => x"33",
         13450 => x"ff",
         13451 => x"08",
         13452 => x"40",
         13453 => x"85",
         13454 => x"70",
         13455 => x"33",
         13456 => x"56",
         13457 => x"2e",
         13458 => x"74",
         13459 => x"ba",
         13460 => x"38",
         13461 => x"33",
         13462 => x"24",
         13463 => x"75",
         13464 => x"d1",
         13465 => x"08",
         13466 => x"80",
         13467 => x"80",
         13468 => x"16",
         13469 => x"11",
         13470 => x"bd",
         13471 => x"5b",
         13472 => x"79",
         13473 => x"a9",
         13474 => x"c8",
         13475 => x"06",
         13476 => x"5d",
         13477 => x"7b",
         13478 => x"75",
         13479 => x"06",
         13480 => x"7f",
         13481 => x"9f",
         13482 => x"53",
         13483 => x"51",
         13484 => x"3f",
         13485 => x"08",
         13486 => x"6d",
         13487 => x"2e",
         13488 => x"74",
         13489 => x"26",
         13490 => x"ff",
         13491 => x"55",
         13492 => x"38",
         13493 => x"88",
         13494 => x"7f",
         13495 => x"38",
         13496 => x"0a",
         13497 => x"38",
         13498 => x"06",
         13499 => x"e7",
         13500 => x"2a",
         13501 => x"89",
         13502 => x"2b",
         13503 => x"47",
         13504 => x"2e",
         13505 => x"65",
         13506 => x"25",
         13507 => x"5f",
         13508 => x"83",
         13509 => x"80",
         13510 => x"38",
         13511 => x"53",
         13512 => x"51",
         13513 => x"3f",
         13514 => x"b9",
         13515 => x"95",
         13516 => x"ff",
         13517 => x"83",
         13518 => x"71",
         13519 => x"59",
         13520 => x"77",
         13521 => x"2e",
         13522 => x"82",
         13523 => x"90",
         13524 => x"83",
         13525 => x"44",
         13526 => x"2e",
         13527 => x"83",
         13528 => x"11",
         13529 => x"33",
         13530 => x"71",
         13531 => x"81",
         13532 => x"72",
         13533 => x"75",
         13534 => x"83",
         13535 => x"11",
         13536 => x"33",
         13537 => x"71",
         13538 => x"81",
         13539 => x"72",
         13540 => x"75",
         13541 => x"5c",
         13542 => x"42",
         13543 => x"a3",
         13544 => x"4e",
         13545 => x"4f",
         13546 => x"78",
         13547 => x"80",
         13548 => x"82",
         13549 => x"57",
         13550 => x"26",
         13551 => x"61",
         13552 => x"81",
         13553 => x"63",
         13554 => x"f9",
         13555 => x"06",
         13556 => x"2e",
         13557 => x"81",
         13558 => x"83",
         13559 => x"6e",
         13560 => x"46",
         13561 => x"62",
         13562 => x"c2",
         13563 => x"38",
         13564 => x"57",
         13565 => x"e6",
         13566 => x"58",
         13567 => x"9d",
         13568 => x"26",
         13569 => x"e6",
         13570 => x"10",
         13571 => x"22",
         13572 => x"74",
         13573 => x"38",
         13574 => x"ee",
         13575 => x"78",
         13576 => x"83",
         13577 => x"c8",
         13578 => x"05",
         13579 => x"c8",
         13580 => x"26",
         13581 => x"0b",
         13582 => x"08",
         13583 => x"c8",
         13584 => x"11",
         13585 => x"05",
         13586 => x"83",
         13587 => x"2a",
         13588 => x"a0",
         13589 => x"7d",
         13590 => x"66",
         13591 => x"70",
         13592 => x"31",
         13593 => x"44",
         13594 => x"89",
         13595 => x"1d",
         13596 => x"29",
         13597 => x"31",
         13598 => x"79",
         13599 => x"38",
         13600 => x"7d",
         13601 => x"70",
         13602 => x"56",
         13603 => x"3f",
         13604 => x"08",
         13605 => x"2e",
         13606 => x"62",
         13607 => x"81",
         13608 => x"38",
         13609 => x"0b",
         13610 => x"08",
         13611 => x"38",
         13612 => x"38",
         13613 => x"74",
         13614 => x"89",
         13615 => x"5b",
         13616 => x"8b",
         13617 => x"b9",
         13618 => x"3d",
         13619 => x"d4",
         13620 => x"4e",
         13621 => x"93",
         13622 => x"c8",
         13623 => x"0d",
         13624 => x"0c",
         13625 => x"d0",
         13626 => x"ff",
         13627 => x"57",
         13628 => x"91",
         13629 => x"77",
         13630 => x"d0",
         13631 => x"77",
         13632 => x"b2",
         13633 => x"83",
         13634 => x"5c",
         13635 => x"57",
         13636 => x"81",
         13637 => x"76",
         13638 => x"58",
         13639 => x"12",
         13640 => x"62",
         13641 => x"38",
         13642 => x"81",
         13643 => x"44",
         13644 => x"45",
         13645 => x"89",
         13646 => x"70",
         13647 => x"59",
         13648 => x"70",
         13649 => x"47",
         13650 => x"09",
         13651 => x"38",
         13652 => x"38",
         13653 => x"70",
         13654 => x"07",
         13655 => x"07",
         13656 => x"7a",
         13657 => x"ce",
         13658 => x"84",
         13659 => x"83",
         13660 => x"98",
         13661 => x"f9",
         13662 => x"3d",
         13663 => x"81",
         13664 => x"fe",
         13665 => x"81",
         13666 => x"c8",
         13667 => x"38",
         13668 => x"77",
         13669 => x"c8",
         13670 => x"75",
         13671 => x"5f",
         13672 => x"57",
         13673 => x"fe",
         13674 => x"7f",
         13675 => x"fb",
         13676 => x"fa",
         13677 => x"83",
         13678 => x"38",
         13679 => x"3d",
         13680 => x"95",
         13681 => x"06",
         13682 => x"67",
         13683 => x"f5",
         13684 => x"70",
         13685 => x"43",
         13686 => x"84",
         13687 => x"9f",
         13688 => x"38",
         13689 => x"77",
         13690 => x"80",
         13691 => x"f5",
         13692 => x"76",
         13693 => x"0c",
         13694 => x"84",
         13695 => x"04",
         13696 => x"81",
         13697 => x"38",
         13698 => x"27",
         13699 => x"81",
         13700 => x"57",
         13701 => x"38",
         13702 => x"57",
         13703 => x"70",
         13704 => x"34",
         13705 => x"74",
         13706 => x"61",
         13707 => x"59",
         13708 => x"70",
         13709 => x"33",
         13710 => x"05",
         13711 => x"15",
         13712 => x"38",
         13713 => x"45",
         13714 => x"82",
         13715 => x"34",
         13716 => x"05",
         13717 => x"ff",
         13718 => x"6a",
         13719 => x"34",
         13720 => x"5c",
         13721 => x"05",
         13722 => x"90",
         13723 => x"83",
         13724 => x"5a",
         13725 => x"91",
         13726 => x"9e",
         13727 => x"49",
         13728 => x"05",
         13729 => x"75",
         13730 => x"26",
         13731 => x"75",
         13732 => x"06",
         13733 => x"93",
         13734 => x"88",
         13735 => x"61",
         13736 => x"f8",
         13737 => x"34",
         13738 => x"05",
         13739 => x"99",
         13740 => x"61",
         13741 => x"80",
         13742 => x"34",
         13743 => x"05",
         13744 => x"2a",
         13745 => x"9d",
         13746 => x"90",
         13747 => x"61",
         13748 => x"7e",
         13749 => x"b9",
         13750 => x"b9",
         13751 => x"9f",
         13752 => x"83",
         13753 => x"38",
         13754 => x"05",
         13755 => x"a8",
         13756 => x"61",
         13757 => x"80",
         13758 => x"05",
         13759 => x"ff",
         13760 => x"74",
         13761 => x"34",
         13762 => x"4b",
         13763 => x"05",
         13764 => x"61",
         13765 => x"a9",
         13766 => x"34",
         13767 => x"05",
         13768 => x"59",
         13769 => x"70",
         13770 => x"33",
         13771 => x"05",
         13772 => x"15",
         13773 => x"38",
         13774 => x"05",
         13775 => x"69",
         13776 => x"ff",
         13777 => x"aa",
         13778 => x"54",
         13779 => x"52",
         13780 => x"c6",
         13781 => x"57",
         13782 => x"08",
         13783 => x"60",
         13784 => x"83",
         13785 => x"38",
         13786 => x"55",
         13787 => x"81",
         13788 => x"ff",
         13789 => x"f4",
         13790 => x"41",
         13791 => x"2e",
         13792 => x"87",
         13793 => x"57",
         13794 => x"83",
         13795 => x"76",
         13796 => x"88",
         13797 => x"55",
         13798 => x"81",
         13799 => x"76",
         13800 => x"78",
         13801 => x"05",
         13802 => x"98",
         13803 => x"64",
         13804 => x"65",
         13805 => x"26",
         13806 => x"59",
         13807 => x"53",
         13808 => x"51",
         13809 => x"3f",
         13810 => x"08",
         13811 => x"84",
         13812 => x"55",
         13813 => x"81",
         13814 => x"ff",
         13815 => x"f4",
         13816 => x"77",
         13817 => x"5b",
         13818 => x"7f",
         13819 => x"7f",
         13820 => x"89",
         13821 => x"62",
         13822 => x"38",
         13823 => x"55",
         13824 => x"83",
         13825 => x"74",
         13826 => x"60",
         13827 => x"fe",
         13828 => x"84",
         13829 => x"85",
         13830 => x"1b",
         13831 => x"57",
         13832 => x"38",
         13833 => x"83",
         13834 => x"86",
         13835 => x"ff",
         13836 => x"38",
         13837 => x"82",
         13838 => x"81",
         13839 => x"c1",
         13840 => x"2a",
         13841 => x"7d",
         13842 => x"84",
         13843 => x"59",
         13844 => x"81",
         13845 => x"ff",
         13846 => x"f4",
         13847 => x"69",
         13848 => x"6b",
         13849 => x"be",
         13850 => x"67",
         13851 => x"81",
         13852 => x"67",
         13853 => x"78",
         13854 => x"34",
         13855 => x"05",
         13856 => x"80",
         13857 => x"62",
         13858 => x"f8",
         13859 => x"67",
         13860 => x"84",
         13861 => x"82",
         13862 => x"57",
         13863 => x"05",
         13864 => x"c8",
         13865 => x"05",
         13866 => x"83",
         13867 => x"67",
         13868 => x"05",
         13869 => x"83",
         13870 => x"84",
         13871 => x"61",
         13872 => x"34",
         13873 => x"ca",
         13874 => x"88",
         13875 => x"61",
         13876 => x"34",
         13877 => x"58",
         13878 => x"cc",
         13879 => x"98",
         13880 => x"61",
         13881 => x"34",
         13882 => x"53",
         13883 => x"51",
         13884 => x"3f",
         13885 => x"b9",
         13886 => x"c9",
         13887 => x"80",
         13888 => x"fe",
         13889 => x"81",
         13890 => x"c8",
         13891 => x"38",
         13892 => x"08",
         13893 => x"0c",
         13894 => x"84",
         13895 => x"04",
         13896 => x"e4",
         13897 => x"64",
         13898 => x"f6",
         13899 => x"ae",
         13900 => x"2a",
         13901 => x"83",
         13902 => x"56",
         13903 => x"2e",
         13904 => x"77",
         13905 => x"83",
         13906 => x"77",
         13907 => x"70",
         13908 => x"58",
         13909 => x"86",
         13910 => x"27",
         13911 => x"52",
         13912 => x"f6",
         13913 => x"b9",
         13914 => x"10",
         13915 => x"70",
         13916 => x"5c",
         13917 => x"0b",
         13918 => x"08",
         13919 => x"05",
         13920 => x"ff",
         13921 => x"27",
         13922 => x"8e",
         13923 => x"39",
         13924 => x"08",
         13925 => x"26",
         13926 => x"7a",
         13927 => x"77",
         13928 => x"7a",
         13929 => x"8e",
         13930 => x"39",
         13931 => x"44",
         13932 => x"f8",
         13933 => x"43",
         13934 => x"75",
         13935 => x"34",
         13936 => x"49",
         13937 => x"05",
         13938 => x"2a",
         13939 => x"a2",
         13940 => x"98",
         13941 => x"61",
         13942 => x"f9",
         13943 => x"61",
         13944 => x"34",
         13945 => x"c4",
         13946 => x"61",
         13947 => x"34",
         13948 => x"80",
         13949 => x"7c",
         13950 => x"34",
         13951 => x"5c",
         13952 => x"05",
         13953 => x"2a",
         13954 => x"a6",
         13955 => x"98",
         13956 => x"61",
         13957 => x"82",
         13958 => x"34",
         13959 => x"05",
         13960 => x"ae",
         13961 => x"61",
         13962 => x"81",
         13963 => x"34",
         13964 => x"05",
         13965 => x"b2",
         13966 => x"61",
         13967 => x"ff",
         13968 => x"c0",
         13969 => x"61",
         13970 => x"34",
         13971 => x"c7",
         13972 => x"a4",
         13973 => x"76",
         13974 => x"58",
         13975 => x"81",
         13976 => x"ff",
         13977 => x"80",
         13978 => x"38",
         13979 => x"05",
         13980 => x"70",
         13981 => x"34",
         13982 => x"74",
         13983 => x"b8",
         13984 => x"80",
         13985 => x"79",
         13986 => x"d9",
         13987 => x"84",
         13988 => x"f4",
         13989 => x"90",
         13990 => x"42",
         13991 => x"b2",
         13992 => x"54",
         13993 => x"08",
         13994 => x"79",
         13995 => x"b4",
         13996 => x"39",
         13997 => x"b9",
         13998 => x"3d",
         13999 => x"d4",
         14000 => x"61",
         14001 => x"ff",
         14002 => x"05",
         14003 => x"6a",
         14004 => x"4c",
         14005 => x"34",
         14006 => x"05",
         14007 => x"85",
         14008 => x"61",
         14009 => x"ff",
         14010 => x"34",
         14011 => x"05",
         14012 => x"89",
         14013 => x"61",
         14014 => x"8f",
         14015 => x"57",
         14016 => x"76",
         14017 => x"53",
         14018 => x"51",
         14019 => x"3f",
         14020 => x"56",
         14021 => x"70",
         14022 => x"34",
         14023 => x"76",
         14024 => x"5c",
         14025 => x"70",
         14026 => x"34",
         14027 => x"d2",
         14028 => x"05",
         14029 => x"e1",
         14030 => x"05",
         14031 => x"c1",
         14032 => x"f2",
         14033 => x"05",
         14034 => x"61",
         14035 => x"34",
         14036 => x"83",
         14037 => x"80",
         14038 => x"e7",
         14039 => x"ff",
         14040 => x"61",
         14041 => x"34",
         14042 => x"59",
         14043 => x"e9",
         14044 => x"90",
         14045 => x"61",
         14046 => x"34",
         14047 => x"40",
         14048 => x"eb",
         14049 => x"61",
         14050 => x"34",
         14051 => x"ed",
         14052 => x"61",
         14053 => x"34",
         14054 => x"ef",
         14055 => x"d5",
         14056 => x"aa",
         14057 => x"54",
         14058 => x"60",
         14059 => x"fe",
         14060 => x"81",
         14061 => x"53",
         14062 => x"51",
         14063 => x"3f",
         14064 => x"55",
         14065 => x"f4",
         14066 => x"61",
         14067 => x"7b",
         14068 => x"5a",
         14069 => x"78",
         14070 => x"8d",
         14071 => x"3d",
         14072 => x"81",
         14073 => x"79",
         14074 => x"b4",
         14075 => x"2e",
         14076 => x"9e",
         14077 => x"33",
         14078 => x"2e",
         14079 => x"76",
         14080 => x"58",
         14081 => x"57",
         14082 => x"86",
         14083 => x"24",
         14084 => x"76",
         14085 => x"76",
         14086 => x"55",
         14087 => x"c8",
         14088 => x"0d",
         14089 => x"0d",
         14090 => x"05",
         14091 => x"59",
         14092 => x"2e",
         14093 => x"84",
         14094 => x"80",
         14095 => x"38",
         14096 => x"77",
         14097 => x"56",
         14098 => x"34",
         14099 => x"74",
         14100 => x"38",
         14101 => x"0c",
         14102 => x"18",
         14103 => x"0d",
         14104 => x"fc",
         14105 => x"53",
         14106 => x"76",
         14107 => x"9e",
         14108 => x"7a",
         14109 => x"70",
         14110 => x"2a",
         14111 => x"1b",
         14112 => x"88",
         14113 => x"56",
         14114 => x"8d",
         14115 => x"ff",
         14116 => x"a3",
         14117 => x"0d",
         14118 => x"05",
         14119 => x"58",
         14120 => x"77",
         14121 => x"76",
         14122 => x"58",
         14123 => x"55",
         14124 => x"a1",
         14125 => x"0c",
         14126 => x"80",
         14127 => x"56",
         14128 => x"80",
         14129 => x"77",
         14130 => x"56",
         14131 => x"34",
         14132 => x"74",
         14133 => x"38",
         14134 => x"0c",
         14135 => x"18",
         14136 => x"80",
         14137 => x"38",
         14138 => x"ac",
         14139 => x"54",
         14140 => x"76",
         14141 => x"9d",
         14142 => x"b9",
         14143 => x"38",
         14144 => x"ba",
         14145 => x"84",
         14146 => x"9f",
         14147 => x"9f",
         14148 => x"11",
         14149 => x"c0",
         14150 => x"08",
         14151 => x"a2",
         14152 => x"32",
         14153 => x"72",
         14154 => x"70",
         14155 => x"56",
         14156 => x"39",
         14157 => x"51",
         14158 => x"ff",
         14159 => x"84",
         14160 => x"9f",
         14161 => x"fd",
         14162 => x"02",
         14163 => x"05",
         14164 => x"80",
         14165 => x"ff",
         14166 => x"72",
         14167 => x"06",
         14168 => x"b9",
         14169 => x"3d",
         14170 => x"ff",
         14171 => x"54",
         14172 => x"2e",
         14173 => x"e9",
         14174 => x"2e",
         14175 => x"e7",
         14176 => x"72",
         14177 => x"38",
         14178 => x"83",
         14179 => x"53",
         14180 => x"ff",
         14181 => x"71",
         14182 => x"8c",
         14183 => x"51",
         14184 => x"81",
         14185 => x"81",
         14186 => x"b9",
         14187 => x"85",
         14188 => x"fe",
         14189 => x"92",
         14190 => x"84",
         14191 => x"22",
         14192 => x"53",
         14193 => x"26",
         14194 => x"53",
         14195 => x"c8",
         14196 => x"0d",
         14197 => x"b5",
         14198 => x"06",
         14199 => x"81",
         14200 => x"38",
         14201 => x"e5",
         14202 => x"22",
         14203 => x"0c",
         14204 => x"0d",
         14205 => x"0d",
         14206 => x"83",
         14207 => x"80",
         14208 => x"83",
         14209 => x"83",
         14210 => x"56",
         14211 => x"26",
         14212 => x"74",
         14213 => x"56",
         14214 => x"30",
         14215 => x"73",
         14216 => x"54",
         14217 => x"70",
         14218 => x"70",
         14219 => x"22",
         14220 => x"2a",
         14221 => x"ff",
         14222 => x"52",
         14223 => x"24",
         14224 => x"cf",
         14225 => x"15",
         14226 => x"05",
         14227 => x"73",
         14228 => x"25",
         14229 => x"07",
         14230 => x"70",
         14231 => x"38",
         14232 => x"84",
         14233 => x"87",
         14234 => x"83",
         14235 => x"ff",
         14236 => x"88",
         14237 => x"71",
         14238 => x"c9",
         14239 => x"73",
         14240 => x"a0",
         14241 => x"ff",
         14242 => x"51",
         14243 => x"39",
         14244 => x"70",
         14245 => x"06",
         14246 => x"39",
         14247 => x"83",
         14248 => x"57",
         14249 => x"e6",
         14250 => x"ff",
         14251 => x"51",
         14252 => x"16",
         14253 => x"ff",
         14254 => x"d0",
         14255 => x"70",
         14256 => x"06",
         14257 => x"39",
         14258 => x"83",
         14259 => x"57",
         14260 => x"39",
         14261 => x"81",
         14262 => x"31",
         14263 => x"ff",
         14264 => x"55",
         14265 => x"75",
         14266 => x"75",
         14267 => x"52",
         14268 => x"39",
         14269 => x"ff",
         14270 => x"00",
         14271 => x"ff",
         14272 => x"ff",
         14273 => x"00",
         14274 => x"00",
         14275 => x"00",
         14276 => x"00",
         14277 => x"00",
         14278 => x"00",
         14279 => x"00",
         14280 => x"00",
         14281 => x"00",
         14282 => x"00",
         14283 => x"00",
         14284 => x"00",
         14285 => x"00",
         14286 => x"00",
         14287 => x"00",
         14288 => x"00",
         14289 => x"00",
         14290 => x"00",
         14291 => x"00",
         14292 => x"00",
         14293 => x"00",
         14294 => x"00",
         14295 => x"00",
         14296 => x"00",
         14297 => x"00",
         14298 => x"00",
         14299 => x"00",
         14300 => x"00",
         14301 => x"00",
         14302 => x"00",
         14303 => x"00",
         14304 => x"00",
         14305 => x"00",
         14306 => x"00",
         14307 => x"00",
         14308 => x"00",
         14309 => x"00",
         14310 => x"00",
         14311 => x"00",
         14312 => x"00",
         14313 => x"00",
         14314 => x"00",
         14315 => x"00",
         14316 => x"00",
         14317 => x"00",
         14318 => x"00",
         14319 => x"00",
         14320 => x"00",
         14321 => x"00",
         14322 => x"00",
         14323 => x"00",
         14324 => x"00",
         14325 => x"00",
         14326 => x"00",
         14327 => x"00",
         14328 => x"00",
         14329 => x"00",
         14330 => x"00",
         14331 => x"00",
         14332 => x"00",
         14333 => x"00",
         14334 => x"00",
         14335 => x"00",
         14336 => x"00",
         14337 => x"00",
         14338 => x"00",
         14339 => x"00",
         14340 => x"00",
         14341 => x"00",
         14342 => x"00",
         14343 => x"00",
         14344 => x"00",
         14345 => x"00",
         14346 => x"00",
         14347 => x"00",
         14348 => x"00",
         14349 => x"00",
         14350 => x"00",
         14351 => x"00",
         14352 => x"00",
         14353 => x"00",
         14354 => x"00",
         14355 => x"00",
         14356 => x"00",
         14357 => x"00",
         14358 => x"00",
         14359 => x"00",
         14360 => x"00",
         14361 => x"00",
         14362 => x"00",
         14363 => x"00",
         14364 => x"00",
         14365 => x"00",
         14366 => x"00",
         14367 => x"00",
         14368 => x"00",
         14369 => x"00",
         14370 => x"00",
         14371 => x"00",
         14372 => x"00",
         14373 => x"00",
         14374 => x"00",
         14375 => x"00",
         14376 => x"00",
         14377 => x"00",
         14378 => x"00",
         14379 => x"00",
         14380 => x"00",
         14381 => x"00",
         14382 => x"00",
         14383 => x"00",
         14384 => x"00",
         14385 => x"00",
         14386 => x"00",
         14387 => x"00",
         14388 => x"00",
         14389 => x"00",
         14390 => x"00",
         14391 => x"00",
         14392 => x"00",
         14393 => x"00",
         14394 => x"00",
         14395 => x"00",
         14396 => x"00",
         14397 => x"00",
         14398 => x"00",
         14399 => x"00",
         14400 => x"00",
         14401 => x"00",
         14402 => x"00",
         14403 => x"00",
         14404 => x"00",
         14405 => x"00",
         14406 => x"00",
         14407 => x"00",
         14408 => x"00",
         14409 => x"00",
         14410 => x"00",
         14411 => x"00",
         14412 => x"00",
         14413 => x"00",
         14414 => x"00",
         14415 => x"00",
         14416 => x"00",
         14417 => x"00",
         14418 => x"00",
         14419 => x"00",
         14420 => x"00",
         14421 => x"00",
         14422 => x"00",
         14423 => x"00",
         14424 => x"00",
         14425 => x"00",
         14426 => x"00",
         14427 => x"00",
         14428 => x"00",
         14429 => x"00",
         14430 => x"00",
         14431 => x"00",
         14432 => x"00",
         14433 => x"00",
         14434 => x"00",
         14435 => x"00",
         14436 => x"00",
         14437 => x"00",
         14438 => x"00",
         14439 => x"00",
         14440 => x"00",
         14441 => x"00",
         14442 => x"00",
         14443 => x"00",
         14444 => x"00",
         14445 => x"00",
         14446 => x"00",
         14447 => x"00",
         14448 => x"00",
         14449 => x"00",
         14450 => x"00",
         14451 => x"00",
         14452 => x"00",
         14453 => x"00",
         14454 => x"00",
         14455 => x"00",
         14456 => x"00",
         14457 => x"00",
         14458 => x"00",
         14459 => x"00",
         14460 => x"00",
         14461 => x"00",
         14462 => x"00",
         14463 => x"00",
         14464 => x"00",
         14465 => x"00",
         14466 => x"00",
         14467 => x"00",
         14468 => x"00",
         14469 => x"00",
         14470 => x"00",
         14471 => x"00",
         14472 => x"00",
         14473 => x"00",
         14474 => x"00",
         14475 => x"00",
         14476 => x"00",
         14477 => x"00",
         14478 => x"00",
         14479 => x"00",
         14480 => x"00",
         14481 => x"00",
         14482 => x"00",
         14483 => x"00",
         14484 => x"00",
         14485 => x"00",
         14486 => x"00",
         14487 => x"00",
         14488 => x"00",
         14489 => x"00",
         14490 => x"00",
         14491 => x"00",
         14492 => x"00",
         14493 => x"00",
         14494 => x"00",
         14495 => x"00",
         14496 => x"00",
         14497 => x"00",
         14498 => x"00",
         14499 => x"00",
         14500 => x"00",
         14501 => x"00",
         14502 => x"00",
         14503 => x"00",
         14504 => x"00",
         14505 => x"00",
         14506 => x"00",
         14507 => x"00",
         14508 => x"00",
         14509 => x"00",
         14510 => x"00",
         14511 => x"00",
         14512 => x"00",
         14513 => x"00",
         14514 => x"00",
         14515 => x"00",
         14516 => x"00",
         14517 => x"00",
         14518 => x"00",
         14519 => x"00",
         14520 => x"00",
         14521 => x"00",
         14522 => x"00",
         14523 => x"00",
         14524 => x"00",
         14525 => x"00",
         14526 => x"00",
         14527 => x"00",
         14528 => x"00",
         14529 => x"00",
         14530 => x"00",
         14531 => x"00",
         14532 => x"00",
         14533 => x"00",
         14534 => x"00",
         14535 => x"00",
         14536 => x"00",
         14537 => x"00",
         14538 => x"00",
         14539 => x"00",
         14540 => x"00",
         14541 => x"00",
         14542 => x"00",
         14543 => x"00",
         14544 => x"00",
         14545 => x"00",
         14546 => x"00",
         14547 => x"00",
         14548 => x"00",
         14549 => x"00",
         14550 => x"00",
         14551 => x"00",
         14552 => x"00",
         14553 => x"00",
         14554 => x"00",
         14555 => x"00",
         14556 => x"00",
         14557 => x"00",
         14558 => x"00",
         14559 => x"00",
         14560 => x"00",
         14561 => x"00",
         14562 => x"00",
         14563 => x"00",
         14564 => x"00",
         14565 => x"00",
         14566 => x"00",
         14567 => x"00",
         14568 => x"00",
         14569 => x"00",
         14570 => x"00",
         14571 => x"00",
         14572 => x"00",
         14573 => x"00",
         14574 => x"00",
         14575 => x"00",
         14576 => x"00",
         14577 => x"00",
         14578 => x"00",
         14579 => x"00",
         14580 => x"00",
         14581 => x"00",
         14582 => x"00",
         14583 => x"00",
         14584 => x"00",
         14585 => x"00",
         14586 => x"00",
         14587 => x"00",
         14588 => x"00",
         14589 => x"00",
         14590 => x"00",
         14591 => x"00",
         14592 => x"00",
         14593 => x"00",
         14594 => x"00",
         14595 => x"00",
         14596 => x"00",
         14597 => x"00",
         14598 => x"00",
         14599 => x"00",
         14600 => x"00",
         14601 => x"00",
         14602 => x"00",
         14603 => x"00",
         14604 => x"00",
         14605 => x"00",
         14606 => x"00",
         14607 => x"00",
         14608 => x"00",
         14609 => x"00",
         14610 => x"00",
         14611 => x"00",
         14612 => x"00",
         14613 => x"00",
         14614 => x"00",
         14615 => x"00",
         14616 => x"00",
         14617 => x"00",
         14618 => x"00",
         14619 => x"00",
         14620 => x"00",
         14621 => x"00",
         14622 => x"00",
         14623 => x"00",
         14624 => x"00",
         14625 => x"00",
         14626 => x"00",
         14627 => x"00",
         14628 => x"00",
         14629 => x"00",
         14630 => x"00",
         14631 => x"00",
         14632 => x"00",
         14633 => x"00",
         14634 => x"00",
         14635 => x"00",
         14636 => x"00",
         14637 => x"00",
         14638 => x"00",
         14639 => x"00",
         14640 => x"00",
         14641 => x"00",
         14642 => x"00",
         14643 => x"00",
         14644 => x"00",
         14645 => x"00",
         14646 => x"00",
         14647 => x"00",
         14648 => x"00",
         14649 => x"00",
         14650 => x"00",
         14651 => x"00",
         14652 => x"00",
         14653 => x"00",
         14654 => x"00",
         14655 => x"00",
         14656 => x"00",
         14657 => x"00",
         14658 => x"00",
         14659 => x"00",
         14660 => x"00",
         14661 => x"00",
         14662 => x"00",
         14663 => x"00",
         14664 => x"00",
         14665 => x"00",
         14666 => x"00",
         14667 => x"00",
         14668 => x"00",
         14669 => x"00",
         14670 => x"00",
         14671 => x"00",
         14672 => x"00",
         14673 => x"00",
         14674 => x"00",
         14675 => x"00",
         14676 => x"00",
         14677 => x"00",
         14678 => x"00",
         14679 => x"00",
         14680 => x"00",
         14681 => x"00",
         14682 => x"00",
         14683 => x"00",
         14684 => x"00",
         14685 => x"00",
         14686 => x"00",
         14687 => x"00",
         14688 => x"00",
         14689 => x"00",
         14690 => x"00",
         14691 => x"00",
         14692 => x"00",
         14693 => x"00",
         14694 => x"00",
         14695 => x"00",
         14696 => x"00",
         14697 => x"00",
         14698 => x"00",
         14699 => x"00",
         14700 => x"00",
         14701 => x"00",
         14702 => x"00",
         14703 => x"00",
         14704 => x"00",
         14705 => x"00",
         14706 => x"00",
         14707 => x"00",
         14708 => x"00",
         14709 => x"00",
         14710 => x"00",
         14711 => x"00",
         14712 => x"00",
         14713 => x"00",
         14714 => x"00",
         14715 => x"00",
         14716 => x"00",
         14717 => x"00",
         14718 => x"00",
         14719 => x"00",
         14720 => x"00",
         14721 => x"00",
         14722 => x"00",
         14723 => x"00",
         14724 => x"00",
         14725 => x"00",
         14726 => x"00",
         14727 => x"00",
         14728 => x"00",
         14729 => x"00",
         14730 => x"00",
         14731 => x"00",
         14732 => x"00",
         14733 => x"00",
         14734 => x"00",
         14735 => x"00",
         14736 => x"00",
         14737 => x"00",
         14738 => x"00",
         14739 => x"00",
         14740 => x"00",
         14741 => x"00",
         14742 => x"00",
         14743 => x"00",
         14744 => x"00",
         14745 => x"00",
         14746 => x"69",
         14747 => x"00",
         14748 => x"69",
         14749 => x"6c",
         14750 => x"69",
         14751 => x"00",
         14752 => x"6c",
         14753 => x"00",
         14754 => x"65",
         14755 => x"00",
         14756 => x"63",
         14757 => x"72",
         14758 => x"63",
         14759 => x"00",
         14760 => x"64",
         14761 => x"00",
         14762 => x"64",
         14763 => x"00",
         14764 => x"65",
         14765 => x"65",
         14766 => x"65",
         14767 => x"69",
         14768 => x"69",
         14769 => x"66",
         14770 => x"66",
         14771 => x"61",
         14772 => x"00",
         14773 => x"6d",
         14774 => x"65",
         14775 => x"72",
         14776 => x"65",
         14777 => x"00",
         14778 => x"6e",
         14779 => x"00",
         14780 => x"65",
         14781 => x"00",
         14782 => x"6c",
         14783 => x"38",
         14784 => x"62",
         14785 => x"63",
         14786 => x"62",
         14787 => x"63",
         14788 => x"69",
         14789 => x"00",
         14790 => x"64",
         14791 => x"6e",
         14792 => x"77",
         14793 => x"72",
         14794 => x"2e",
         14795 => x"61",
         14796 => x"65",
         14797 => x"73",
         14798 => x"63",
         14799 => x"65",
         14800 => x"00",
         14801 => x"6f",
         14802 => x"61",
         14803 => x"6f",
         14804 => x"20",
         14805 => x"65",
         14806 => x"00",
         14807 => x"6e",
         14808 => x"66",
         14809 => x"65",
         14810 => x"6d",
         14811 => x"72",
         14812 => x"00",
         14813 => x"69",
         14814 => x"69",
         14815 => x"6f",
         14816 => x"64",
         14817 => x"69",
         14818 => x"75",
         14819 => x"6f",
         14820 => x"61",
         14821 => x"6e",
         14822 => x"6e",
         14823 => x"6c",
         14824 => x"00",
         14825 => x"6f",
         14826 => x"74",
         14827 => x"6f",
         14828 => x"64",
         14829 => x"6f",
         14830 => x"6d",
         14831 => x"69",
         14832 => x"20",
         14833 => x"65",
         14834 => x"74",
         14835 => x"66",
         14836 => x"64",
         14837 => x"20",
         14838 => x"6b",
         14839 => x"69",
         14840 => x"6e",
         14841 => x"65",
         14842 => x"6c",
         14843 => x"00",
         14844 => x"72",
         14845 => x"20",
         14846 => x"62",
         14847 => x"69",
         14848 => x"6e",
         14849 => x"69",
         14850 => x"00",
         14851 => x"44",
         14852 => x"20",
         14853 => x"74",
         14854 => x"72",
         14855 => x"63",
         14856 => x"2e",
         14857 => x"69",
         14858 => x"68",
         14859 => x"6c",
         14860 => x"6e",
         14861 => x"69",
         14862 => x"00",
         14863 => x"69",
         14864 => x"61",
         14865 => x"61",
         14866 => x"65",
         14867 => x"74",
         14868 => x"00",
         14869 => x"63",
         14870 => x"73",
         14871 => x"6e",
         14872 => x"2e",
         14873 => x"6e",
         14874 => x"69",
         14875 => x"69",
         14876 => x"61",
         14877 => x"00",
         14878 => x"6f",
         14879 => x"74",
         14880 => x"6f",
         14881 => x"2e",
         14882 => x"6f",
         14883 => x"6c",
         14884 => x"6f",
         14885 => x"2e",
         14886 => x"69",
         14887 => x"6e",
         14888 => x"72",
         14889 => x"79",
         14890 => x"6e",
         14891 => x"6e",
         14892 => x"65",
         14893 => x"72",
         14894 => x"69",
         14895 => x"45",
         14896 => x"72",
         14897 => x"75",
         14898 => x"73",
         14899 => x"00",
         14900 => x"25",
         14901 => x"62",
         14902 => x"73",
         14903 => x"20",
         14904 => x"25",
         14905 => x"62",
         14906 => x"73",
         14907 => x"63",
         14908 => x"00",
         14909 => x"65",
         14910 => x"00",
         14911 => x"30",
         14912 => x"00",
         14913 => x"20",
         14914 => x"30",
         14915 => x"00",
         14916 => x"7c",
         14917 => x"00",
         14918 => x"20",
         14919 => x"30",
         14920 => x"00",
         14921 => x"20",
         14922 => x"20",
         14923 => x"00",
         14924 => x"4f",
         14925 => x"2a",
         14926 => x"20",
         14927 => x"37",
         14928 => x"2f",
         14929 => x"31",
         14930 => x"31",
         14931 => x"00",
         14932 => x"5a",
         14933 => x"20",
         14934 => x"20",
         14935 => x"78",
         14936 => x"73",
         14937 => x"20",
         14938 => x"0a",
         14939 => x"53",
         14940 => x"20",
         14941 => x"61",
         14942 => x"41",
         14943 => x"65",
         14944 => x"20",
         14945 => x"20",
         14946 => x"20",
         14947 => x"3d",
         14948 => x"38",
         14949 => x"00",
         14950 => x"20",
         14951 => x"70",
         14952 => x"64",
         14953 => x"73",
         14954 => x"20",
         14955 => x"20",
         14956 => x"20",
         14957 => x"3d",
         14958 => x"38",
         14959 => x"00",
         14960 => x"50",
         14961 => x"6e",
         14962 => x"72",
         14963 => x"20",
         14964 => x"64",
         14965 => x"00",
         14966 => x"41",
         14967 => x"20",
         14968 => x"69",
         14969 => x"72",
         14970 => x"74",
         14971 => x"41",
         14972 => x"20",
         14973 => x"69",
         14974 => x"72",
         14975 => x"74",
         14976 => x"41",
         14977 => x"20",
         14978 => x"69",
         14979 => x"72",
         14980 => x"74",
         14981 => x"41",
         14982 => x"20",
         14983 => x"69",
         14984 => x"72",
         14985 => x"74",
         14986 => x"4f",
         14987 => x"20",
         14988 => x"69",
         14989 => x"72",
         14990 => x"74",
         14991 => x"4f",
         14992 => x"20",
         14993 => x"69",
         14994 => x"72",
         14995 => x"74",
         14996 => x"53",
         14997 => x"6e",
         14998 => x"72",
         14999 => x"00",
         15000 => x"69",
         15001 => x"20",
         15002 => x"65",
         15003 => x"70",
         15004 => x"65",
         15005 => x"6e",
         15006 => x"70",
         15007 => x"6d",
         15008 => x"2e",
         15009 => x"6e",
         15010 => x"69",
         15011 => x"74",
         15012 => x"72",
         15013 => x"00",
         15014 => x"75",
         15015 => x"78",
         15016 => x"62",
         15017 => x"00",
         15018 => x"4f",
         15019 => x"70",
         15020 => x"73",
         15021 => x"61",
         15022 => x"64",
         15023 => x"20",
         15024 => x"74",
         15025 => x"69",
         15026 => x"73",
         15027 => x"61",
         15028 => x"30",
         15029 => x"6c",
         15030 => x"65",
         15031 => x"69",
         15032 => x"61",
         15033 => x"6c",
         15034 => x"00",
         15035 => x"20",
         15036 => x"64",
         15037 => x"73",
         15038 => x"3a",
         15039 => x"61",
         15040 => x"6f",
         15041 => x"6e",
         15042 => x"00",
         15043 => x"50",
         15044 => x"69",
         15045 => x"64",
         15046 => x"73",
         15047 => x"2e",
         15048 => x"00",
         15049 => x"6f",
         15050 => x"72",
         15051 => x"6f",
         15052 => x"67",
         15053 => x"00",
         15054 => x"65",
         15055 => x"72",
         15056 => x"67",
         15057 => x"70",
         15058 => x"61",
         15059 => x"6e",
         15060 => x"00",
         15061 => x"61",
         15062 => x"6e",
         15063 => x"6f",
         15064 => x"40",
         15065 => x"38",
         15066 => x"2e",
         15067 => x"00",
         15068 => x"61",
         15069 => x"72",
         15070 => x"72",
         15071 => x"20",
         15072 => x"65",
         15073 => x"64",
         15074 => x"00",
         15075 => x"78",
         15076 => x"74",
         15077 => x"20",
         15078 => x"65",
         15079 => x"25",
         15080 => x"78",
         15081 => x"2e",
         15082 => x"30",
         15083 => x"20",
         15084 => x"6c",
         15085 => x"00",
         15086 => x"30",
         15087 => x"20",
         15088 => x"58",
         15089 => x"6f",
         15090 => x"72",
         15091 => x"2e",
         15092 => x"00",
         15093 => x"30",
         15094 => x"28",
         15095 => x"78",
         15096 => x"25",
         15097 => x"78",
         15098 => x"38",
         15099 => x"00",
         15100 => x"6f",
         15101 => x"6e",
         15102 => x"2e",
         15103 => x"30",
         15104 => x"20",
         15105 => x"58",
         15106 => x"6c",
         15107 => x"69",
         15108 => x"2e",
         15109 => x"00",
         15110 => x"75",
         15111 => x"4d",
         15112 => x"72",
         15113 => x"43",
         15114 => x"6c",
         15115 => x"2e",
         15116 => x"64",
         15117 => x"73",
         15118 => x"00",
         15119 => x"65",
         15120 => x"79",
         15121 => x"68",
         15122 => x"74",
         15123 => x"20",
         15124 => x"6e",
         15125 => x"70",
         15126 => x"65",
         15127 => x"63",
         15128 => x"61",
         15129 => x"00",
         15130 => x"3f",
         15131 => x"64",
         15132 => x"2f",
         15133 => x"25",
         15134 => x"64",
         15135 => x"2e",
         15136 => x"64",
         15137 => x"6f",
         15138 => x"6f",
         15139 => x"67",
         15140 => x"74",
         15141 => x"00",
         15142 => x"0a",
         15143 => x"69",
         15144 => x"20",
         15145 => x"6c",
         15146 => x"6e",
         15147 => x"3a",
         15148 => x"64",
         15149 => x"73",
         15150 => x"3a",
         15151 => x"20",
         15152 => x"50",
         15153 => x"65",
         15154 => x"20",
         15155 => x"74",
         15156 => x"41",
         15157 => x"65",
         15158 => x"3d",
         15159 => x"38",
         15160 => x"00",
         15161 => x"20",
         15162 => x"50",
         15163 => x"65",
         15164 => x"79",
         15165 => x"61",
         15166 => x"41",
         15167 => x"65",
         15168 => x"3d",
         15169 => x"38",
         15170 => x"00",
         15171 => x"20",
         15172 => x"74",
         15173 => x"20",
         15174 => x"72",
         15175 => x"64",
         15176 => x"73",
         15177 => x"20",
         15178 => x"3d",
         15179 => x"38",
         15180 => x"00",
         15181 => x"69",
         15182 => x"00",
         15183 => x"20",
         15184 => x"50",
         15185 => x"64",
         15186 => x"20",
         15187 => x"20",
         15188 => x"20",
         15189 => x"20",
         15190 => x"3d",
         15191 => x"34",
         15192 => x"00",
         15193 => x"20",
         15194 => x"79",
         15195 => x"6d",
         15196 => x"6f",
         15197 => x"46",
         15198 => x"20",
         15199 => x"20",
         15200 => x"3d",
         15201 => x"2e",
         15202 => x"64",
         15203 => x"0a",
         15204 => x"20",
         15205 => x"69",
         15206 => x"6f",
         15207 => x"53",
         15208 => x"4d",
         15209 => x"6f",
         15210 => x"46",
         15211 => x"3d",
         15212 => x"2e",
         15213 => x"64",
         15214 => x"0a",
         15215 => x"20",
         15216 => x"44",
         15217 => x"20",
         15218 => x"63",
         15219 => x"72",
         15220 => x"20",
         15221 => x"20",
         15222 => x"3d",
         15223 => x"2e",
         15224 => x"64",
         15225 => x"0a",
         15226 => x"20",
         15227 => x"50",
         15228 => x"20",
         15229 => x"53",
         15230 => x"20",
         15231 => x"4f",
         15232 => x"00",
         15233 => x"20",
         15234 => x"42",
         15235 => x"43",
         15236 => x"20",
         15237 => x"49",
         15238 => x"4f",
         15239 => x"42",
         15240 => x"00",
         15241 => x"20",
         15242 => x"4e",
         15243 => x"43",
         15244 => x"20",
         15245 => x"61",
         15246 => x"6c",
         15247 => x"30",
         15248 => x"2e",
         15249 => x"20",
         15250 => x"49",
         15251 => x"31",
         15252 => x"20",
         15253 => x"6d",
         15254 => x"20",
         15255 => x"30",
         15256 => x"2e",
         15257 => x"20",
         15258 => x"44",
         15259 => x"52",
         15260 => x"20",
         15261 => x"76",
         15262 => x"73",
         15263 => x"30",
         15264 => x"2e",
         15265 => x"20",
         15266 => x"41",
         15267 => x"20",
         15268 => x"20",
         15269 => x"38",
         15270 => x"30",
         15271 => x"2e",
         15272 => x"20",
         15273 => x"52",
         15274 => x"20",
         15275 => x"20",
         15276 => x"38",
         15277 => x"30",
         15278 => x"2e",
         15279 => x"20",
         15280 => x"4e",
         15281 => x"42",
         15282 => x"20",
         15283 => x"38",
         15284 => x"30",
         15285 => x"2e",
         15286 => x"20",
         15287 => x"44",
         15288 => x"20",
         15289 => x"20",
         15290 => x"38",
         15291 => x"30",
         15292 => x"2e",
         15293 => x"20",
         15294 => x"42",
         15295 => x"52",
         15296 => x"20",
         15297 => x"38",
         15298 => x"30",
         15299 => x"2e",
         15300 => x"28",
         15301 => x"6d",
         15302 => x"43",
         15303 => x"6e",
         15304 => x"29",
         15305 => x"6e",
         15306 => x"77",
         15307 => x"56",
         15308 => x"00",
         15309 => x"6d",
         15310 => x"00",
         15311 => x"65",
         15312 => x"6d",
         15313 => x"6c",
         15314 => x"00",
         15315 => x"56",
         15316 => x"00",
         15317 => x"00",
         15318 => x"00",
         15319 => x"00",
         15320 => x"00",
         15321 => x"00",
         15322 => x"00",
         15323 => x"00",
         15324 => x"00",
         15325 => x"00",
         15326 => x"00",
         15327 => x"00",
         15328 => x"00",
         15329 => x"00",
         15330 => x"00",
         15331 => x"00",
         15332 => x"00",
         15333 => x"00",
         15334 => x"00",
         15335 => x"00",
         15336 => x"00",
         15337 => x"00",
         15338 => x"00",
         15339 => x"00",
         15340 => x"00",
         15341 => x"00",
         15342 => x"00",
         15343 => x"00",
         15344 => x"00",
         15345 => x"00",
         15346 => x"00",
         15347 => x"00",
         15348 => x"00",
         15349 => x"00",
         15350 => x"00",
         15351 => x"00",
         15352 => x"00",
         15353 => x"00",
         15354 => x"00",
         15355 => x"00",
         15356 => x"00",
         15357 => x"00",
         15358 => x"00",
         15359 => x"00",
         15360 => x"00",
         15361 => x"00",
         15362 => x"00",
         15363 => x"00",
         15364 => x"00",
         15365 => x"00",
         15366 => x"00",
         15367 => x"00",
         15368 => x"00",
         15369 => x"00",
         15370 => x"00",
         15371 => x"00",
         15372 => x"00",
         15373 => x"00",
         15374 => x"00",
         15375 => x"00",
         15376 => x"00",
         15377 => x"00",
         15378 => x"00",
         15379 => x"00",
         15380 => x"00",
         15381 => x"00",
         15382 => x"5b",
         15383 => x"5b",
         15384 => x"5b",
         15385 => x"5b",
         15386 => x"5b",
         15387 => x"5b",
         15388 => x"5b",
         15389 => x"30",
         15390 => x"5b",
         15391 => x"5b",
         15392 => x"5b",
         15393 => x"00",
         15394 => x"00",
         15395 => x"00",
         15396 => x"00",
         15397 => x"00",
         15398 => x"00",
         15399 => x"00",
         15400 => x"00",
         15401 => x"00",
         15402 => x"00",
         15403 => x"00",
         15404 => x"61",
         15405 => x"74",
         15406 => x"65",
         15407 => x"72",
         15408 => x"65",
         15409 => x"73",
         15410 => x"79",
         15411 => x"6c",
         15412 => x"64",
         15413 => x"62",
         15414 => x"67",
         15415 => x"69",
         15416 => x"72",
         15417 => x"69",
         15418 => x"00",
         15419 => x"00",
         15420 => x"30",
         15421 => x"20",
         15422 => x"0a",
         15423 => x"61",
         15424 => x"64",
         15425 => x"20",
         15426 => x"65",
         15427 => x"68",
         15428 => x"69",
         15429 => x"72",
         15430 => x"69",
         15431 => x"74",
         15432 => x"4f",
         15433 => x"00",
         15434 => x"25",
         15435 => x"00",
         15436 => x"5b",
         15437 => x"00",
         15438 => x"5b",
         15439 => x"5b",
         15440 => x"5b",
         15441 => x"5b",
         15442 => x"5b",
         15443 => x"00",
         15444 => x"5b",
         15445 => x"00",
         15446 => x"5b",
         15447 => x"00",
         15448 => x"5b",
         15449 => x"00",
         15450 => x"5b",
         15451 => x"00",
         15452 => x"5b",
         15453 => x"00",
         15454 => x"5b",
         15455 => x"00",
         15456 => x"5b",
         15457 => x"00",
         15458 => x"5b",
         15459 => x"00",
         15460 => x"5b",
         15461 => x"00",
         15462 => x"5b",
         15463 => x"00",
         15464 => x"5b",
         15465 => x"00",
         15466 => x"5b",
         15467 => x"5b",
         15468 => x"00",
         15469 => x"5b",
         15470 => x"00",
         15471 => x"3a",
         15472 => x"25",
         15473 => x"64",
         15474 => x"2c",
         15475 => x"25",
         15476 => x"30",
         15477 => x"00",
         15478 => x"3a",
         15479 => x"25",
         15480 => x"64",
         15481 => x"3a",
         15482 => x"25",
         15483 => x"64",
         15484 => x"64",
         15485 => x"3a",
         15486 => x"00",
         15487 => x"30",
         15488 => x"00",
         15489 => x"63",
         15490 => x"3b",
         15491 => x"00",
         15492 => x"65",
         15493 => x"74",
         15494 => x"72",
         15495 => x"3a",
         15496 => x"70",
         15497 => x"32",
         15498 => x"30",
         15499 => x"00",
         15500 => x"77",
         15501 => x"32",
         15502 => x"30",
         15503 => x"00",
         15504 => x"64",
         15505 => x"32",
         15506 => x"00",
         15507 => x"6f",
         15508 => x"73",
         15509 => x"65",
         15510 => x"65",
         15511 => x"00",
         15512 => x"44",
         15513 => x"2a",
         15514 => x"3f",
         15515 => x"00",
         15516 => x"2c",
         15517 => x"5d",
         15518 => x"41",
         15519 => x"41",
         15520 => x"00",
         15521 => x"fe",
         15522 => x"44",
         15523 => x"2e",
         15524 => x"4f",
         15525 => x"4d",
         15526 => x"20",
         15527 => x"54",
         15528 => x"20",
         15529 => x"4f",
         15530 => x"4d",
         15531 => x"20",
         15532 => x"54",
         15533 => x"20",
         15534 => x"00",
         15535 => x"00",
         15536 => x"00",
         15537 => x"00",
         15538 => x"03",
         15539 => x"0e",
         15540 => x"16",
         15541 => x"00",
         15542 => x"9a",
         15543 => x"41",
         15544 => x"45",
         15545 => x"49",
         15546 => x"92",
         15547 => x"4f",
         15548 => x"99",
         15549 => x"9d",
         15550 => x"49",
         15551 => x"a5",
         15552 => x"a9",
         15553 => x"ad",
         15554 => x"b1",
         15555 => x"b5",
         15556 => x"b9",
         15557 => x"bd",
         15558 => x"c1",
         15559 => x"c5",
         15560 => x"c9",
         15561 => x"cd",
         15562 => x"d1",
         15563 => x"d5",
         15564 => x"d9",
         15565 => x"dd",
         15566 => x"e1",
         15567 => x"e5",
         15568 => x"e9",
         15569 => x"ed",
         15570 => x"f1",
         15571 => x"f5",
         15572 => x"f9",
         15573 => x"fd",
         15574 => x"2e",
         15575 => x"5b",
         15576 => x"22",
         15577 => x"3e",
         15578 => x"00",
         15579 => x"01",
         15580 => x"10",
         15581 => x"00",
         15582 => x"00",
         15583 => x"01",
         15584 => x"04",
         15585 => x"10",
         15586 => x"00",
         15587 => x"c7",
         15588 => x"e9",
         15589 => x"e4",
         15590 => x"e5",
         15591 => x"ea",
         15592 => x"e8",
         15593 => x"ee",
         15594 => x"c4",
         15595 => x"c9",
         15596 => x"c6",
         15597 => x"f6",
         15598 => x"fb",
         15599 => x"ff",
         15600 => x"dc",
         15601 => x"a3",
         15602 => x"a7",
         15603 => x"e1",
         15604 => x"f3",
         15605 => x"f1",
         15606 => x"aa",
         15607 => x"bf",
         15608 => x"ac",
         15609 => x"bc",
         15610 => x"ab",
         15611 => x"91",
         15612 => x"93",
         15613 => x"24",
         15614 => x"62",
         15615 => x"55",
         15616 => x"51",
         15617 => x"5d",
         15618 => x"5b",
         15619 => x"14",
         15620 => x"2c",
         15621 => x"00",
         15622 => x"5e",
         15623 => x"5a",
         15624 => x"69",
         15625 => x"60",
         15626 => x"6c",
         15627 => x"68",
         15628 => x"65",
         15629 => x"58",
         15630 => x"53",
         15631 => x"6a",
         15632 => x"0c",
         15633 => x"84",
         15634 => x"90",
         15635 => x"b1",
         15636 => x"93",
         15637 => x"a3",
         15638 => x"b5",
         15639 => x"a6",
         15640 => x"a9",
         15641 => x"1e",
         15642 => x"b5",
         15643 => x"61",
         15644 => x"65",
         15645 => x"20",
         15646 => x"f7",
         15647 => x"b0",
         15648 => x"b7",
         15649 => x"7f",
         15650 => x"a0",
         15651 => x"61",
         15652 => x"e0",
         15653 => x"f8",
         15654 => x"ff",
         15655 => x"78",
         15656 => x"30",
         15657 => x"06",
         15658 => x"10",
         15659 => x"2e",
         15660 => x"06",
         15661 => x"4d",
         15662 => x"81",
         15663 => x"82",
         15664 => x"84",
         15665 => x"87",
         15666 => x"89",
         15667 => x"8b",
         15668 => x"8d",
         15669 => x"8f",
         15670 => x"91",
         15671 => x"93",
         15672 => x"f6",
         15673 => x"97",
         15674 => x"98",
         15675 => x"9b",
         15676 => x"9d",
         15677 => x"9f",
         15678 => x"a0",
         15679 => x"a2",
         15680 => x"a4",
         15681 => x"a7",
         15682 => x"a9",
         15683 => x"ab",
         15684 => x"ac",
         15685 => x"af",
         15686 => x"b1",
         15687 => x"b3",
         15688 => x"b5",
         15689 => x"b7",
         15690 => x"b8",
         15691 => x"bb",
         15692 => x"bc",
         15693 => x"f7",
         15694 => x"c1",
         15695 => x"c3",
         15696 => x"c5",
         15697 => x"c7",
         15698 => x"c7",
         15699 => x"cb",
         15700 => x"cd",
         15701 => x"dd",
         15702 => x"8e",
         15703 => x"12",
         15704 => x"03",
         15705 => x"f4",
         15706 => x"f8",
         15707 => x"22",
         15708 => x"3a",
         15709 => x"65",
         15710 => x"3b",
         15711 => x"66",
         15712 => x"40",
         15713 => x"41",
         15714 => x"0a",
         15715 => x"40",
         15716 => x"86",
         15717 => x"89",
         15718 => x"58",
         15719 => x"5a",
         15720 => x"5c",
         15721 => x"5e",
         15722 => x"93",
         15723 => x"62",
         15724 => x"64",
         15725 => x"66",
         15726 => x"97",
         15727 => x"6a",
         15728 => x"6c",
         15729 => x"6e",
         15730 => x"70",
         15731 => x"9d",
         15732 => x"74",
         15733 => x"76",
         15734 => x"78",
         15735 => x"7a",
         15736 => x"7c",
         15737 => x"7e",
         15738 => x"a6",
         15739 => x"82",
         15740 => x"84",
         15741 => x"86",
         15742 => x"ae",
         15743 => x"b1",
         15744 => x"45",
         15745 => x"8e",
         15746 => x"90",
         15747 => x"b7",
         15748 => x"03",
         15749 => x"fe",
         15750 => x"ac",
         15751 => x"86",
         15752 => x"89",
         15753 => x"b1",
         15754 => x"c2",
         15755 => x"a3",
         15756 => x"c4",
         15757 => x"cc",
         15758 => x"8c",
         15759 => x"8f",
         15760 => x"18",
         15761 => x"0a",
         15762 => x"f3",
         15763 => x"f5",
         15764 => x"f7",
         15765 => x"f9",
         15766 => x"fa",
         15767 => x"20",
         15768 => x"10",
         15769 => x"22",
         15770 => x"36",
         15771 => x"0e",
         15772 => x"01",
         15773 => x"d0",
         15774 => x"61",
         15775 => x"00",
         15776 => x"7d",
         15777 => x"63",
         15778 => x"96",
         15779 => x"5a",
         15780 => x"08",
         15781 => x"06",
         15782 => x"08",
         15783 => x"08",
         15784 => x"06",
         15785 => x"07",
         15786 => x"52",
         15787 => x"54",
         15788 => x"56",
         15789 => x"60",
         15790 => x"70",
         15791 => x"ba",
         15792 => x"c8",
         15793 => x"ca",
         15794 => x"da",
         15795 => x"f8",
         15796 => x"ea",
         15797 => x"fa",
         15798 => x"80",
         15799 => x"90",
         15800 => x"a0",
         15801 => x"b0",
         15802 => x"b8",
         15803 => x"b2",
         15804 => x"cc",
         15805 => x"c3",
         15806 => x"02",
         15807 => x"02",
         15808 => x"01",
         15809 => x"f3",
         15810 => x"fc",
         15811 => x"01",
         15812 => x"70",
         15813 => x"84",
         15814 => x"83",
         15815 => x"1a",
         15816 => x"2f",
         15817 => x"02",
         15818 => x"06",
         15819 => x"02",
         15820 => x"64",
         15821 => x"26",
         15822 => x"1a",
         15823 => x"00",
         15824 => x"00",
         15825 => x"02",
         15826 => x"00",
         15827 => x"00",
         15828 => x"00",
         15829 => x"04",
         15830 => x"00",
         15831 => x"00",
         15832 => x"00",
         15833 => x"14",
         15834 => x"00",
         15835 => x"00",
         15836 => x"00",
         15837 => x"2b",
         15838 => x"00",
         15839 => x"00",
         15840 => x"00",
         15841 => x"30",
         15842 => x"00",
         15843 => x"00",
         15844 => x"00",
         15845 => x"3c",
         15846 => x"00",
         15847 => x"00",
         15848 => x"00",
         15849 => x"3d",
         15850 => x"00",
         15851 => x"00",
         15852 => x"00",
         15853 => x"3f",
         15854 => x"00",
         15855 => x"00",
         15856 => x"00",
         15857 => x"40",
         15858 => x"00",
         15859 => x"00",
         15860 => x"00",
         15861 => x"41",
         15862 => x"00",
         15863 => x"00",
         15864 => x"00",
         15865 => x"42",
         15866 => x"00",
         15867 => x"00",
         15868 => x"00",
         15869 => x"43",
         15870 => x"00",
         15871 => x"00",
         15872 => x"00",
         15873 => x"50",
         15874 => x"00",
         15875 => x"00",
         15876 => x"00",
         15877 => x"51",
         15878 => x"00",
         15879 => x"00",
         15880 => x"00",
         15881 => x"54",
         15882 => x"00",
         15883 => x"00",
         15884 => x"00",
         15885 => x"55",
         15886 => x"00",
         15887 => x"00",
         15888 => x"00",
         15889 => x"79",
         15890 => x"00",
         15891 => x"00",
         15892 => x"00",
         15893 => x"78",
         15894 => x"00",
         15895 => x"00",
         15896 => x"00",
         15897 => x"82",
         15898 => x"00",
         15899 => x"00",
         15900 => x"00",
         15901 => x"83",
         15902 => x"00",
         15903 => x"00",
         15904 => x"00",
         15905 => x"85",
         15906 => x"00",
         15907 => x"00",
         15908 => x"00",
         15909 => x"87",
         15910 => x"00",
         15911 => x"00",
         15912 => x"00",
         15913 => x"88",
         15914 => x"00",
         15915 => x"00",
         15916 => x"00",
         15917 => x"89",
         15918 => x"00",
         15919 => x"00",
         15920 => x"00",
         15921 => x"8c",
         15922 => x"00",
         15923 => x"00",
         15924 => x"00",
         15925 => x"8d",
         15926 => x"00",
         15927 => x"00",
         15928 => x"00",
         15929 => x"8e",
         15930 => x"00",
         15931 => x"00",
         15932 => x"00",
         15933 => x"8f",
         15934 => x"00",
         15935 => x"00",
         15936 => x"00",
         15937 => x"00",
         15938 => x"00",
         15939 => x"00",
         15940 => x"00",
         15941 => x"01",
         15942 => x"00",
         15943 => x"01",
         15944 => x"81",
         15945 => x"00",
         15946 => x"7f",
         15947 => x"00",
         15948 => x"00",
         15949 => x"00",
         15950 => x"00",
         15951 => x"f5",
         15952 => x"f5",
         15953 => x"f5",
         15954 => x"00",
         15955 => x"01",
         15956 => x"01",
         15957 => x"01",
         15958 => x"00",
         15959 => x"00",
         15960 => x"00",
         15961 => x"00",
         15962 => x"00",
         15963 => x"00",
         15964 => x"00",
         15965 => x"00",
         15966 => x"00",
         15967 => x"00",
         15968 => x"00",
         15969 => x"00",
         15970 => x"00",
         15971 => x"00",
         15972 => x"00",
         15973 => x"00",
         15974 => x"00",
         15975 => x"00",
         15976 => x"00",
         15977 => x"00",
         15978 => x"00",
         15979 => x"00",
         15980 => x"00",
         15981 => x"00",
         15982 => x"00",
         15983 => x"00",
         15984 => x"00",
         15985 => x"00",
         15986 => x"00",
         15987 => x"00",
         15988 => x"00",
         15989 => x"01",
         15990 => x"fc",
         15991 => x"3b",
         15992 => x"7a",
         15993 => x"f0",
         15994 => x"72",
         15995 => x"76",
         15996 => x"6a",
         15997 => x"6e",
         15998 => x"62",
         15999 => x"66",
         16000 => x"32",
         16001 => x"36",
         16002 => x"f3",
         16003 => x"39",
         16004 => x"7f",
         16005 => x"f2",
         16006 => x"f0",
         16007 => x"f0",
         16008 => x"81",
         16009 => x"f0",
         16010 => x"fc",
         16011 => x"3a",
         16012 => x"5a",
         16013 => x"f0",
         16014 => x"52",
         16015 => x"56",
         16016 => x"4a",
         16017 => x"4e",
         16018 => x"42",
         16019 => x"46",
         16020 => x"32",
         16021 => x"36",
         16022 => x"f3",
         16023 => x"39",
         16024 => x"7f",
         16025 => x"f2",
         16026 => x"f0",
         16027 => x"f0",
         16028 => x"81",
         16029 => x"f0",
         16030 => x"fc",
         16031 => x"2b",
         16032 => x"5a",
         16033 => x"f0",
         16034 => x"52",
         16035 => x"56",
         16036 => x"4a",
         16037 => x"4e",
         16038 => x"42",
         16039 => x"46",
         16040 => x"22",
         16041 => x"26",
         16042 => x"7e",
         16043 => x"29",
         16044 => x"e2",
         16045 => x"f8",
         16046 => x"f0",
         16047 => x"f0",
         16048 => x"86",
         16049 => x"f0",
         16050 => x"fe",
         16051 => x"f0",
         16052 => x"1a",
         16053 => x"f0",
         16054 => x"12",
         16055 => x"16",
         16056 => x"0a",
         16057 => x"0e",
         16058 => x"02",
         16059 => x"06",
         16060 => x"f0",
         16061 => x"f0",
         16062 => x"1e",
         16063 => x"1f",
         16064 => x"f0",
         16065 => x"f0",
         16066 => x"f0",
         16067 => x"f0",
         16068 => x"81",
         16069 => x"f0",
         16070 => x"f0",
         16071 => x"b5",
         16072 => x"77",
         16073 => x"f0",
         16074 => x"70",
         16075 => x"a6",
         16076 => x"5d",
         16077 => x"33",
         16078 => x"6e",
         16079 => x"43",
         16080 => x"36",
         16081 => x"1e",
         16082 => x"9f",
         16083 => x"a3",
         16084 => x"c5",
         16085 => x"c4",
         16086 => x"f0",
         16087 => x"f0",
         16088 => x"81",
         16089 => x"f0",
         16090 => x"00",
         16091 => x"00",
         16092 => x"00",
         16093 => x"00",
         16094 => x"00",
         16095 => x"00",
         16096 => x"00",
         16097 => x"00",
         16098 => x"00",
         16099 => x"00",
         16100 => x"00",
         16101 => x"00",
         16102 => x"00",
         16103 => x"00",
         16104 => x"00",
         16105 => x"00",
         16106 => x"00",
         16107 => x"00",
         16108 => x"00",
         16109 => x"00",
         16110 => x"00",
         16111 => x"00",
         16112 => x"00",
         16113 => x"00",
         16114 => x"00",
         16115 => x"01",
         16116 => x"00",
         16117 => x"00",
         16118 => x"00",
         16119 => x"00",
         16120 => x"00",
         16121 => x"00",
         16122 => x"00",
         16123 => x"00",
         16124 => x"00",
         16125 => x"00",
         16126 => x"00",
         16127 => x"00",
         16128 => x"00",
         16129 => x"00",
         16130 => x"00",
         16131 => x"00",
         16132 => x"00",
         16133 => x"00",
         16134 => x"00",
         16135 => x"00",
         16136 => x"00",
         16137 => x"00",
         16138 => x"00",
         16139 => x"00",
         16140 => x"00",
         16141 => x"00",
         16142 => x"00",
         16143 => x"00",
         16144 => x"00",
         16145 => x"00",
         16146 => x"00",
         16147 => x"00",
         16148 => x"00",
         16149 => x"00",
         16150 => x"00",
         16151 => x"00",
         16152 => x"00",
         16153 => x"00",
         16154 => x"00",
         16155 => x"00",
         16156 => x"00",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"00",
         16166 => x"00",
         16167 => x"00",
         16168 => x"00",
         16169 => x"00",
         16170 => x"00",
         16171 => x"00",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"00",
         18159 => x"00",
         18160 => x"00",
         18161 => x"e0",
         18162 => x"cf",
         18163 => x"f9",
         18164 => x"fd",
         18165 => x"c1",
         18166 => x"c5",
         18167 => x"e4",
         18168 => x"ee",
         18169 => x"61",
         18170 => x"65",
         18171 => x"69",
         18172 => x"2a",
         18173 => x"21",
         18174 => x"25",
         18175 => x"29",
         18176 => x"2b",
         18177 => x"01",
         18178 => x"05",
         18179 => x"09",
         18180 => x"0d",
         18181 => x"11",
         18182 => x"15",
         18183 => x"19",
         18184 => x"54",
         18185 => x"81",
         18186 => x"85",
         18187 => x"89",
         18188 => x"8d",
         18189 => x"91",
         18190 => x"95",
         18191 => x"99",
         18192 => x"40",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"00",
         18199 => x"00",
         18200 => x"00",
         18201 => x"00",
         18202 => x"00",
         18203 => x"00",
         18204 => x"00",
         18205 => x"00",
         18206 => x"00",
         18207 => x"00",
         18208 => x"00",
         18209 => x"00",
         18210 => x"00",
         18211 => x"00",
         18212 => x"00",
         18213 => x"00",
         18214 => x"00",
         18215 => x"00",
         18216 => x"00",
         18217 => x"00",
         18218 => x"00",
         18219 => x"00",
         18220 => x"00",
         18221 => x"00",
         18222 => x"00",
         18223 => x"02",
         18224 => x"04",
         18225 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"cd",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"f4",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"cc",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"ab",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"96",
           269 => x"0b",
           270 => x"0b",
           271 => x"b6",
           272 => x"0b",
           273 => x"0b",
           274 => x"d6",
           275 => x"0b",
           276 => x"0b",
           277 => x"f6",
           278 => x"0b",
           279 => x"0b",
           280 => x"96",
           281 => x"0b",
           282 => x"0b",
           283 => x"b6",
           284 => x"0b",
           285 => x"0b",
           286 => x"d7",
           287 => x"0b",
           288 => x"0b",
           289 => x"f9",
           290 => x"0b",
           291 => x"0b",
           292 => x"9b",
           293 => x"0b",
           294 => x"0b",
           295 => x"bd",
           296 => x"0b",
           297 => x"0b",
           298 => x"df",
           299 => x"0b",
           300 => x"0b",
           301 => x"81",
           302 => x"0b",
           303 => x"0b",
           304 => x"a3",
           305 => x"0b",
           306 => x"0b",
           307 => x"c5",
           308 => x"0b",
           309 => x"0b",
           310 => x"e7",
           311 => x"0b",
           312 => x"0b",
           313 => x"89",
           314 => x"0b",
           315 => x"0b",
           316 => x"ab",
           317 => x"0b",
           318 => x"0b",
           319 => x"cd",
           320 => x"0b",
           321 => x"0b",
           322 => x"ef",
           323 => x"0b",
           324 => x"0b",
           325 => x"91",
           326 => x"0b",
           327 => x"0b",
           328 => x"b3",
           329 => x"0b",
           330 => x"0b",
           331 => x"d5",
           332 => x"0b",
           333 => x"0b",
           334 => x"f7",
           335 => x"0b",
           336 => x"0b",
           337 => x"99",
           338 => x"0b",
           339 => x"0b",
           340 => x"bb",
           341 => x"0b",
           342 => x"0b",
           343 => x"dc",
           344 => x"0b",
           345 => x"0b",
           346 => x"fe",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"90",
           390 => x"d4",
           391 => x"2d",
           392 => x"08",
           393 => x"90",
           394 => x"d4",
           395 => x"2d",
           396 => x"08",
           397 => x"90",
           398 => x"d4",
           399 => x"2d",
           400 => x"08",
           401 => x"90",
           402 => x"d4",
           403 => x"2d",
           404 => x"08",
           405 => x"90",
           406 => x"d4",
           407 => x"2d",
           408 => x"08",
           409 => x"90",
           410 => x"d4",
           411 => x"2d",
           412 => x"08",
           413 => x"90",
           414 => x"d4",
           415 => x"2d",
           416 => x"08",
           417 => x"90",
           418 => x"d4",
           419 => x"2d",
           420 => x"08",
           421 => x"90",
           422 => x"d4",
           423 => x"2d",
           424 => x"08",
           425 => x"90",
           426 => x"d4",
           427 => x"2d",
           428 => x"08",
           429 => x"90",
           430 => x"d4",
           431 => x"2d",
           432 => x"08",
           433 => x"90",
           434 => x"d4",
           435 => x"ec",
           436 => x"d4",
           437 => x"80",
           438 => x"b9",
           439 => x"d5",
           440 => x"b9",
           441 => x"c0",
           442 => x"84",
           443 => x"80",
           444 => x"84",
           445 => x"80",
           446 => x"04",
           447 => x"0c",
           448 => x"2d",
           449 => x"08",
           450 => x"90",
           451 => x"d4",
           452 => x"ae",
           453 => x"d4",
           454 => x"80",
           455 => x"b9",
           456 => x"e3",
           457 => x"b9",
           458 => x"c0",
           459 => x"84",
           460 => x"82",
           461 => x"84",
           462 => x"80",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"90",
           468 => x"d4",
           469 => x"9d",
           470 => x"d4",
           471 => x"80",
           472 => x"b9",
           473 => x"fa",
           474 => x"b9",
           475 => x"c0",
           476 => x"84",
           477 => x"82",
           478 => x"84",
           479 => x"80",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"90",
           485 => x"d4",
           486 => x"8b",
           487 => x"d4",
           488 => x"80",
           489 => x"b9",
           490 => x"f3",
           491 => x"b9",
           492 => x"c0",
           493 => x"84",
           494 => x"83",
           495 => x"84",
           496 => x"80",
           497 => x"04",
           498 => x"0c",
           499 => x"2d",
           500 => x"08",
           501 => x"90",
           502 => x"d4",
           503 => x"86",
           504 => x"d4",
           505 => x"80",
           506 => x"b9",
           507 => x"f5",
           508 => x"b9",
           509 => x"c0",
           510 => x"84",
           511 => x"83",
           512 => x"84",
           513 => x"80",
           514 => x"04",
           515 => x"0c",
           516 => x"2d",
           517 => x"08",
           518 => x"90",
           519 => x"d4",
           520 => x"d0",
           521 => x"d4",
           522 => x"80",
           523 => x"b9",
           524 => x"e3",
           525 => x"b9",
           526 => x"c0",
           527 => x"84",
           528 => x"82",
           529 => x"84",
           530 => x"80",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"90",
           536 => x"d4",
           537 => x"9a",
           538 => x"d4",
           539 => x"80",
           540 => x"b9",
           541 => x"99",
           542 => x"b9",
           543 => x"c0",
           544 => x"84",
           545 => x"83",
           546 => x"84",
           547 => x"80",
           548 => x"04",
           549 => x"0c",
           550 => x"2d",
           551 => x"08",
           552 => x"90",
           553 => x"d4",
           554 => x"92",
           555 => x"d4",
           556 => x"80",
           557 => x"b9",
           558 => x"b9",
           559 => x"b9",
           560 => x"c0",
           561 => x"84",
           562 => x"83",
           563 => x"84",
           564 => x"80",
           565 => x"04",
           566 => x"0c",
           567 => x"2d",
           568 => x"08",
           569 => x"90",
           570 => x"d4",
           571 => x"e2",
           572 => x"d4",
           573 => x"80",
           574 => x"b9",
           575 => x"f5",
           576 => x"b9",
           577 => x"c0",
           578 => x"84",
           579 => x"80",
           580 => x"84",
           581 => x"80",
           582 => x"04",
           583 => x"0c",
           584 => x"2d",
           585 => x"08",
           586 => x"90",
           587 => x"d4",
           588 => x"a5",
           589 => x"d4",
           590 => x"80",
           591 => x"b9",
           592 => x"9a",
           593 => x"d4",
           594 => x"80",
           595 => x"b9",
           596 => x"db",
           597 => x"b9",
           598 => x"c0",
           599 => x"84",
           600 => x"81",
           601 => x"84",
           602 => x"80",
           603 => x"04",
           604 => x"0c",
           605 => x"2d",
           606 => x"08",
           607 => x"90",
           608 => x"d4",
           609 => x"91",
           610 => x"d4",
           611 => x"80",
           612 => x"04",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"53",
           621 => x"00",
           622 => x"06",
           623 => x"09",
           624 => x"05",
           625 => x"2b",
           626 => x"06",
           627 => x"04",
           628 => x"72",
           629 => x"05",
           630 => x"05",
           631 => x"72",
           632 => x"53",
           633 => x"51",
           634 => x"04",
           635 => x"70",
           636 => x"27",
           637 => x"71",
           638 => x"53",
           639 => x"0b",
           640 => x"8c",
           641 => x"ce",
           642 => x"fc",
           643 => x"3d",
           644 => x"05",
           645 => x"53",
           646 => x"d5",
           647 => x"81",
           648 => x"3d",
           649 => x"3d",
           650 => x"7c",
           651 => x"81",
           652 => x"80",
           653 => x"56",
           654 => x"80",
           655 => x"2e",
           656 => x"80",
           657 => x"14",
           658 => x"32",
           659 => x"72",
           660 => x"51",
           661 => x"54",
           662 => x"b7",
           663 => x"2e",
           664 => x"51",
           665 => x"84",
           666 => x"53",
           667 => x"08",
           668 => x"38",
           669 => x"08",
           670 => x"05",
           671 => x"14",
           672 => x"70",
           673 => x"07",
           674 => x"54",
           675 => x"80",
           676 => x"80",
           677 => x"52",
           678 => x"c8",
           679 => x"0d",
           680 => x"84",
           681 => x"88",
           682 => x"f5",
           683 => x"54",
           684 => x"05",
           685 => x"73",
           686 => x"58",
           687 => x"05",
           688 => x"8d",
           689 => x"51",
           690 => x"19",
           691 => x"34",
           692 => x"04",
           693 => x"86",
           694 => x"53",
           695 => x"51",
           696 => x"3d",
           697 => x"3d",
           698 => x"65",
           699 => x"80",
           700 => x"0c",
           701 => x"70",
           702 => x"32",
           703 => x"55",
           704 => x"72",
           705 => x"81",
           706 => x"38",
           707 => x"76",
           708 => x"c5",
           709 => x"7b",
           710 => x"5c",
           711 => x"81",
           712 => x"17",
           713 => x"26",
           714 => x"76",
           715 => x"30",
           716 => x"51",
           717 => x"ae",
           718 => x"2e",
           719 => x"83",
           720 => x"32",
           721 => x"54",
           722 => x"9e",
           723 => x"80",
           724 => x"33",
           725 => x"bd",
           726 => x"08",
           727 => x"b9",
           728 => x"3d",
           729 => x"83",
           730 => x"10",
           731 => x"10",
           732 => x"2b",
           733 => x"19",
           734 => x"0a",
           735 => x"05",
           736 => x"52",
           737 => x"5f",
           738 => x"81",
           739 => x"81",
           740 => x"ff",
           741 => x"7c",
           742 => x"76",
           743 => x"ff",
           744 => x"a5",
           745 => x"06",
           746 => x"73",
           747 => x"5b",
           748 => x"58",
           749 => x"dd",
           750 => x"39",
           751 => x"51",
           752 => x"7b",
           753 => x"fe",
           754 => x"8d",
           755 => x"2a",
           756 => x"54",
           757 => x"38",
           758 => x"06",
           759 => x"95",
           760 => x"53",
           761 => x"26",
           762 => x"10",
           763 => x"84",
           764 => x"08",
           765 => x"18",
           766 => x"d8",
           767 => x"38",
           768 => x"51",
           769 => x"80",
           770 => x"5b",
           771 => x"38",
           772 => x"80",
           773 => x"f6",
           774 => x"7f",
           775 => x"71",
           776 => x"ff",
           777 => x"58",
           778 => x"b9",
           779 => x"52",
           780 => x"9a",
           781 => x"c8",
           782 => x"06",
           783 => x"08",
           784 => x"56",
           785 => x"26",
           786 => x"b9",
           787 => x"05",
           788 => x"70",
           789 => x"34",
           790 => x"51",
           791 => x"84",
           792 => x"56",
           793 => x"08",
           794 => x"84",
           795 => x"98",
           796 => x"06",
           797 => x"80",
           798 => x"77",
           799 => x"29",
           800 => x"05",
           801 => x"59",
           802 => x"2a",
           803 => x"55",
           804 => x"2e",
           805 => x"84",
           806 => x"f8",
           807 => x"53",
           808 => x"8b",
           809 => x"80",
           810 => x"80",
           811 => x"72",
           812 => x"7a",
           813 => x"81",
           814 => x"72",
           815 => x"38",
           816 => x"70",
           817 => x"54",
           818 => x"24",
           819 => x"7a",
           820 => x"06",
           821 => x"71",
           822 => x"56",
           823 => x"06",
           824 => x"2e",
           825 => x"77",
           826 => x"2b",
           827 => x"7c",
           828 => x"56",
           829 => x"80",
           830 => x"38",
           831 => x"81",
           832 => x"85",
           833 => x"84",
           834 => x"54",
           835 => x"38",
           836 => x"81",
           837 => x"86",
           838 => x"81",
           839 => x"85",
           840 => x"88",
           841 => x"5f",
           842 => x"b2",
           843 => x"84",
           844 => x"fc",
           845 => x"70",
           846 => x"40",
           847 => x"25",
           848 => x"52",
           849 => x"a9",
           850 => x"84",
           851 => x"fc",
           852 => x"70",
           853 => x"40",
           854 => x"24",
           855 => x"81",
           856 => x"80",
           857 => x"78",
           858 => x"0a",
           859 => x"0a",
           860 => x"2c",
           861 => x"80",
           862 => x"38",
           863 => x"51",
           864 => x"78",
           865 => x"0a",
           866 => x"0a",
           867 => x"2c",
           868 => x"74",
           869 => x"38",
           870 => x"70",
           871 => x"55",
           872 => x"81",
           873 => x"80",
           874 => x"d8",
           875 => x"f3",
           876 => x"38",
           877 => x"2e",
           878 => x"7d",
           879 => x"2e",
           880 => x"52",
           881 => x"33",
           882 => x"a5",
           883 => x"b9",
           884 => x"81",
           885 => x"74",
           886 => x"7a",
           887 => x"a7",
           888 => x"84",
           889 => x"fc",
           890 => x"70",
           891 => x"40",
           892 => x"25",
           893 => x"7c",
           894 => x"86",
           895 => x"39",
           896 => x"5b",
           897 => x"7c",
           898 => x"76",
           899 => x"fa",
           900 => x"80",
           901 => x"80",
           902 => x"60",
           903 => x"71",
           904 => x"ff",
           905 => x"59",
           906 => x"fb",
           907 => x"60",
           908 => x"fe",
           909 => x"83",
           910 => x"98",
           911 => x"7c",
           912 => x"29",
           913 => x"05",
           914 => x"5e",
           915 => x"57",
           916 => x"87",
           917 => x"06",
           918 => x"fe",
           919 => x"78",
           920 => x"29",
           921 => x"05",
           922 => x"5a",
           923 => x"7f",
           924 => x"38",
           925 => x"51",
           926 => x"e2",
           927 => x"70",
           928 => x"06",
           929 => x"83",
           930 => x"fe",
           931 => x"52",
           932 => x"05",
           933 => x"85",
           934 => x"39",
           935 => x"83",
           936 => x"5b",
           937 => x"ff",
           938 => x"ab",
           939 => x"75",
           940 => x"57",
           941 => x"b9",
           942 => x"75",
           943 => x"81",
           944 => x"78",
           945 => x"29",
           946 => x"05",
           947 => x"5a",
           948 => x"e3",
           949 => x"70",
           950 => x"56",
           951 => x"c6",
           952 => x"39",
           953 => x"05",
           954 => x"53",
           955 => x"80",
           956 => x"df",
           957 => x"ff",
           958 => x"84",
           959 => x"fa",
           960 => x"84",
           961 => x"58",
           962 => x"89",
           963 => x"39",
           964 => x"5b",
           965 => x"58",
           966 => x"f9",
           967 => x"39",
           968 => x"05",
           969 => x"81",
           970 => x"41",
           971 => x"8a",
           972 => x"87",
           973 => x"b9",
           974 => x"ff",
           975 => x"71",
           976 => x"54",
           977 => x"2c",
           978 => x"39",
           979 => x"07",
           980 => x"5b",
           981 => x"38",
           982 => x"7f",
           983 => x"71",
           984 => x"06",
           985 => x"54",
           986 => x"38",
           987 => x"bb",
           988 => x"c8",
           989 => x"ff",
           990 => x"31",
           991 => x"5a",
           992 => x"81",
           993 => x"33",
           994 => x"f7",
           995 => x"c9",
           996 => x"84",
           997 => x"fc",
           998 => x"70",
           999 => x"54",
          1000 => x"25",
          1001 => x"7c",
          1002 => x"83",
          1003 => x"39",
          1004 => x"51",
          1005 => x"79",
          1006 => x"81",
          1007 => x"38",
          1008 => x"51",
          1009 => x"7a",
          1010 => x"06",
          1011 => x"2e",
          1012 => x"fa",
          1013 => x"98",
          1014 => x"31",
          1015 => x"90",
          1016 => x"80",
          1017 => x"51",
          1018 => x"90",
          1019 => x"39",
          1020 => x"51",
          1021 => x"7e",
          1022 => x"73",
          1023 => x"a2",
          1024 => x"39",
          1025 => x"98",
          1026 => x"e5",
          1027 => x"06",
          1028 => x"2e",
          1029 => x"fb",
          1030 => x"74",
          1031 => x"70",
          1032 => x"53",
          1033 => x"7c",
          1034 => x"82",
          1035 => x"39",
          1036 => x"51",
          1037 => x"ff",
          1038 => x"52",
          1039 => x"8b",
          1040 => x"c8",
          1041 => x"ff",
          1042 => x"31",
          1043 => x"5a",
          1044 => x"7a",
          1045 => x"30",
          1046 => x"bf",
          1047 => x"5b",
          1048 => x"fe",
          1049 => x"d5",
          1050 => x"75",
          1051 => x"f3",
          1052 => x"3d",
          1053 => x"3d",
          1054 => x"80",
          1055 => x"ac",
          1056 => x"33",
          1057 => x"81",
          1058 => x"06",
          1059 => x"55",
          1060 => x"72",
          1061 => x"81",
          1062 => x"38",
          1063 => x"05",
          1064 => x"72",
          1065 => x"38",
          1066 => x"08",
          1067 => x"90",
          1068 => x"72",
          1069 => x"c8",
          1070 => x"83",
          1071 => x"74",
          1072 => x"56",
          1073 => x"80",
          1074 => x"84",
          1075 => x"54",
          1076 => x"d5",
          1077 => x"84",
          1078 => x"52",
          1079 => x"14",
          1080 => x"2d",
          1081 => x"08",
          1082 => x"38",
          1083 => x"56",
          1084 => x"c8",
          1085 => x"0d",
          1086 => x"0d",
          1087 => x"54",
          1088 => x"16",
          1089 => x"2a",
          1090 => x"81",
          1091 => x"57",
          1092 => x"72",
          1093 => x"81",
          1094 => x"73",
          1095 => x"55",
          1096 => x"77",
          1097 => x"06",
          1098 => x"56",
          1099 => x"c8",
          1100 => x"0d",
          1101 => x"81",
          1102 => x"53",
          1103 => x"ea",
          1104 => x"72",
          1105 => x"08",
          1106 => x"84",
          1107 => x"80",
          1108 => x"ff",
          1109 => x"05",
          1110 => x"57",
          1111 => x"ca",
          1112 => x"0d",
          1113 => x"08",
          1114 => x"85",
          1115 => x"0d",
          1116 => x"0d",
          1117 => x"11",
          1118 => x"2a",
          1119 => x"06",
          1120 => x"57",
          1121 => x"ae",
          1122 => x"2a",
          1123 => x"73",
          1124 => x"38",
          1125 => x"53",
          1126 => x"08",
          1127 => x"74",
          1128 => x"76",
          1129 => x"81",
          1130 => x"8c",
          1131 => x"81",
          1132 => x"0c",
          1133 => x"84",
          1134 => x"88",
          1135 => x"74",
          1136 => x"ff",
          1137 => x"15",
          1138 => x"2d",
          1139 => x"b9",
          1140 => x"38",
          1141 => x"81",
          1142 => x"0c",
          1143 => x"39",
          1144 => x"77",
          1145 => x"70",
          1146 => x"70",
          1147 => x"06",
          1148 => x"56",
          1149 => x"b3",
          1150 => x"2a",
          1151 => x"71",
          1152 => x"82",
          1153 => x"52",
          1154 => x"80",
          1155 => x"08",
          1156 => x"53",
          1157 => x"80",
          1158 => x"13",
          1159 => x"16",
          1160 => x"8c",
          1161 => x"81",
          1162 => x"73",
          1163 => x"0c",
          1164 => x"04",
          1165 => x"06",
          1166 => x"17",
          1167 => x"08",
          1168 => x"17",
          1169 => x"33",
          1170 => x"0c",
          1171 => x"04",
          1172 => x"16",
          1173 => x"2d",
          1174 => x"08",
          1175 => x"c8",
          1176 => x"ff",
          1177 => x"16",
          1178 => x"07",
          1179 => x"b9",
          1180 => x"2e",
          1181 => x"a0",
          1182 => x"85",
          1183 => x"54",
          1184 => x"c8",
          1185 => x"0d",
          1186 => x"07",
          1187 => x"17",
          1188 => x"ec",
          1189 => x"0d",
          1190 => x"54",
          1191 => x"70",
          1192 => x"33",
          1193 => x"38",
          1194 => x"72",
          1195 => x"54",
          1196 => x"72",
          1197 => x"54",
          1198 => x"38",
          1199 => x"c8",
          1200 => x"0d",
          1201 => x"0d",
          1202 => x"7a",
          1203 => x"54",
          1204 => x"9d",
          1205 => x"27",
          1206 => x"80",
          1207 => x"71",
          1208 => x"53",
          1209 => x"81",
          1210 => x"ff",
          1211 => x"ef",
          1212 => x"b9",
          1213 => x"3d",
          1214 => x"12",
          1215 => x"27",
          1216 => x"14",
          1217 => x"ff",
          1218 => x"53",
          1219 => x"73",
          1220 => x"51",
          1221 => x"d9",
          1222 => x"ff",
          1223 => x"71",
          1224 => x"ff",
          1225 => x"df",
          1226 => x"fe",
          1227 => x"70",
          1228 => x"70",
          1229 => x"33",
          1230 => x"38",
          1231 => x"74",
          1232 => x"c8",
          1233 => x"3d",
          1234 => x"3d",
          1235 => x"71",
          1236 => x"72",
          1237 => x"54",
          1238 => x"72",
          1239 => x"54",
          1240 => x"38",
          1241 => x"c8",
          1242 => x"0d",
          1243 => x"0d",
          1244 => x"79",
          1245 => x"54",
          1246 => x"93",
          1247 => x"81",
          1248 => x"73",
          1249 => x"55",
          1250 => x"51",
          1251 => x"73",
          1252 => x"0c",
          1253 => x"04",
          1254 => x"76",
          1255 => x"56",
          1256 => x"2e",
          1257 => x"33",
          1258 => x"05",
          1259 => x"52",
          1260 => x"09",
          1261 => x"38",
          1262 => x"71",
          1263 => x"38",
          1264 => x"72",
          1265 => x"51",
          1266 => x"c8",
          1267 => x"0d",
          1268 => x"2e",
          1269 => x"33",
          1270 => x"72",
          1271 => x"38",
          1272 => x"52",
          1273 => x"80",
          1274 => x"72",
          1275 => x"b9",
          1276 => x"3d",
          1277 => x"84",
          1278 => x"86",
          1279 => x"fb",
          1280 => x"79",
          1281 => x"56",
          1282 => x"84",
          1283 => x"84",
          1284 => x"81",
          1285 => x"81",
          1286 => x"84",
          1287 => x"54",
          1288 => x"08",
          1289 => x"38",
          1290 => x"08",
          1291 => x"74",
          1292 => x"75",
          1293 => x"c8",
          1294 => x"b1",
          1295 => x"c8",
          1296 => x"84",
          1297 => x"87",
          1298 => x"fd",
          1299 => x"77",
          1300 => x"55",
          1301 => x"80",
          1302 => x"72",
          1303 => x"54",
          1304 => x"80",
          1305 => x"ff",
          1306 => x"ff",
          1307 => x"06",
          1308 => x"13",
          1309 => x"52",
          1310 => x"b9",
          1311 => x"3d",
          1312 => x"3d",
          1313 => x"79",
          1314 => x"54",
          1315 => x"2e",
          1316 => x"72",
          1317 => x"54",
          1318 => x"51",
          1319 => x"73",
          1320 => x"0c",
          1321 => x"04",
          1322 => x"78",
          1323 => x"a0",
          1324 => x"2e",
          1325 => x"51",
          1326 => x"84",
          1327 => x"52",
          1328 => x"73",
          1329 => x"38",
          1330 => x"e3",
          1331 => x"b9",
          1332 => x"53",
          1333 => x"9f",
          1334 => x"38",
          1335 => x"9f",
          1336 => x"38",
          1337 => x"71",
          1338 => x"31",
          1339 => x"57",
          1340 => x"80",
          1341 => x"2e",
          1342 => x"10",
          1343 => x"07",
          1344 => x"07",
          1345 => x"ff",
          1346 => x"70",
          1347 => x"72",
          1348 => x"31",
          1349 => x"56",
          1350 => x"58",
          1351 => x"da",
          1352 => x"76",
          1353 => x"84",
          1354 => x"88",
          1355 => x"fc",
          1356 => x"70",
          1357 => x"06",
          1358 => x"72",
          1359 => x"70",
          1360 => x"71",
          1361 => x"2a",
          1362 => x"80",
          1363 => x"70",
          1364 => x"2b",
          1365 => x"74",
          1366 => x"81",
          1367 => x"30",
          1368 => x"82",
          1369 => x"31",
          1370 => x"55",
          1371 => x"05",
          1372 => x"70",
          1373 => x"25",
          1374 => x"31",
          1375 => x"70",
          1376 => x"32",
          1377 => x"70",
          1378 => x"31",
          1379 => x"05",
          1380 => x"0c",
          1381 => x"55",
          1382 => x"5a",
          1383 => x"55",
          1384 => x"56",
          1385 => x"56",
          1386 => x"3d",
          1387 => x"3d",
          1388 => x"70",
          1389 => x"54",
          1390 => x"3f",
          1391 => x"08",
          1392 => x"71",
          1393 => x"c8",
          1394 => x"3d",
          1395 => x"3d",
          1396 => x"58",
          1397 => x"76",
          1398 => x"38",
          1399 => x"cf",
          1400 => x"c8",
          1401 => x"13",
          1402 => x"2e",
          1403 => x"51",
          1404 => x"72",
          1405 => x"08",
          1406 => x"53",
          1407 => x"80",
          1408 => x"53",
          1409 => x"be",
          1410 => x"74",
          1411 => x"72",
          1412 => x"2b",
          1413 => x"55",
          1414 => x"76",
          1415 => x"72",
          1416 => x"2a",
          1417 => x"77",
          1418 => x"31",
          1419 => x"2c",
          1420 => x"7b",
          1421 => x"71",
          1422 => x"5c",
          1423 => x"55",
          1424 => x"74",
          1425 => x"84",
          1426 => x"88",
          1427 => x"fa",
          1428 => x"9f",
          1429 => x"2c",
          1430 => x"7b",
          1431 => x"2c",
          1432 => x"73",
          1433 => x"31",
          1434 => x"31",
          1435 => x"59",
          1436 => x"b4",
          1437 => x"c8",
          1438 => x"75",
          1439 => x"c8",
          1440 => x"0d",
          1441 => x"0d",
          1442 => x"57",
          1443 => x"0c",
          1444 => x"33",
          1445 => x"73",
          1446 => x"81",
          1447 => x"81",
          1448 => x"0c",
          1449 => x"55",
          1450 => x"f3",
          1451 => x"2e",
          1452 => x"73",
          1453 => x"83",
          1454 => x"58",
          1455 => x"89",
          1456 => x"38",
          1457 => x"56",
          1458 => x"80",
          1459 => x"e0",
          1460 => x"38",
          1461 => x"81",
          1462 => x"53",
          1463 => x"81",
          1464 => x"53",
          1465 => x"8f",
          1466 => x"70",
          1467 => x"54",
          1468 => x"27",
          1469 => x"72",
          1470 => x"83",
          1471 => x"29",
          1472 => x"70",
          1473 => x"33",
          1474 => x"73",
          1475 => x"be",
          1476 => x"2e",
          1477 => x"30",
          1478 => x"0c",
          1479 => x"84",
          1480 => x"8b",
          1481 => x"81",
          1482 => x"79",
          1483 => x"56",
          1484 => x"b0",
          1485 => x"06",
          1486 => x"81",
          1487 => x"0c",
          1488 => x"55",
          1489 => x"2e",
          1490 => x"58",
          1491 => x"2e",
          1492 => x"56",
          1493 => x"c6",
          1494 => x"53",
          1495 => x"58",
          1496 => x"fe",
          1497 => x"84",
          1498 => x"8b",
          1499 => x"82",
          1500 => x"70",
          1501 => x"33",
          1502 => x"56",
          1503 => x"80",
          1504 => x"c8",
          1505 => x"0d",
          1506 => x"0d",
          1507 => x"57",
          1508 => x"0c",
          1509 => x"33",
          1510 => x"73",
          1511 => x"81",
          1512 => x"81",
          1513 => x"0c",
          1514 => x"55",
          1515 => x"f3",
          1516 => x"2e",
          1517 => x"73",
          1518 => x"83",
          1519 => x"58",
          1520 => x"89",
          1521 => x"38",
          1522 => x"56",
          1523 => x"80",
          1524 => x"e0",
          1525 => x"38",
          1526 => x"81",
          1527 => x"53",
          1528 => x"81",
          1529 => x"53",
          1530 => x"8f",
          1531 => x"70",
          1532 => x"54",
          1533 => x"27",
          1534 => x"72",
          1535 => x"83",
          1536 => x"29",
          1537 => x"70",
          1538 => x"33",
          1539 => x"73",
          1540 => x"be",
          1541 => x"2e",
          1542 => x"30",
          1543 => x"0c",
          1544 => x"84",
          1545 => x"8b",
          1546 => x"81",
          1547 => x"79",
          1548 => x"56",
          1549 => x"b0",
          1550 => x"06",
          1551 => x"81",
          1552 => x"0c",
          1553 => x"55",
          1554 => x"2e",
          1555 => x"58",
          1556 => x"2e",
          1557 => x"56",
          1558 => x"c6",
          1559 => x"53",
          1560 => x"58",
          1561 => x"fe",
          1562 => x"84",
          1563 => x"8b",
          1564 => x"82",
          1565 => x"70",
          1566 => x"33",
          1567 => x"56",
          1568 => x"80",
          1569 => x"c8",
          1570 => x"0d",
          1571 => x"e2",
          1572 => x"c8",
          1573 => x"06",
          1574 => x"0c",
          1575 => x"0d",
          1576 => x"93",
          1577 => x"71",
          1578 => x"be",
          1579 => x"71",
          1580 => x"ce",
          1581 => x"be",
          1582 => x"0d",
          1583 => x"ac",
          1584 => x"3f",
          1585 => x"04",
          1586 => x"51",
          1587 => x"83",
          1588 => x"83",
          1589 => x"ef",
          1590 => x"3d",
          1591 => x"ce",
          1592 => x"92",
          1593 => x"0d",
          1594 => x"84",
          1595 => x"3f",
          1596 => x"04",
          1597 => x"51",
          1598 => x"83",
          1599 => x"83",
          1600 => x"ee",
          1601 => x"3d",
          1602 => x"cf",
          1603 => x"e6",
          1604 => x"0d",
          1605 => x"f0",
          1606 => x"3f",
          1607 => x"04",
          1608 => x"51",
          1609 => x"83",
          1610 => x"83",
          1611 => x"ee",
          1612 => x"3d",
          1613 => x"d0",
          1614 => x"ba",
          1615 => x"0d",
          1616 => x"d4",
          1617 => x"3f",
          1618 => x"04",
          1619 => x"51",
          1620 => x"83",
          1621 => x"83",
          1622 => x"ee",
          1623 => x"3d",
          1624 => x"d1",
          1625 => x"8e",
          1626 => x"0d",
          1627 => x"98",
          1628 => x"3f",
          1629 => x"04",
          1630 => x"51",
          1631 => x"83",
          1632 => x"83",
          1633 => x"ed",
          1634 => x"3d",
          1635 => x"d1",
          1636 => x"e2",
          1637 => x"0d",
          1638 => x"0d",
          1639 => x"05",
          1640 => x"33",
          1641 => x"68",
          1642 => x"7b",
          1643 => x"51",
          1644 => x"78",
          1645 => x"ff",
          1646 => x"81",
          1647 => x"07",
          1648 => x"06",
          1649 => x"57",
          1650 => x"38",
          1651 => x"52",
          1652 => x"52",
          1653 => x"d9",
          1654 => x"c8",
          1655 => x"b9",
          1656 => x"2e",
          1657 => x"77",
          1658 => x"97",
          1659 => x"70",
          1660 => x"25",
          1661 => x"9f",
          1662 => x"53",
          1663 => x"77",
          1664 => x"38",
          1665 => x"88",
          1666 => x"87",
          1667 => x"e0",
          1668 => x"78",
          1669 => x"51",
          1670 => x"84",
          1671 => x"54",
          1672 => x"53",
          1673 => x"d1",
          1674 => x"df",
          1675 => x"b9",
          1676 => x"3d",
          1677 => x"b9",
          1678 => x"c0",
          1679 => x"84",
          1680 => x"59",
          1681 => x"05",
          1682 => x"53",
          1683 => x"51",
          1684 => x"3f",
          1685 => x"08",
          1686 => x"c8",
          1687 => x"38",
          1688 => x"80",
          1689 => x"38",
          1690 => x"17",
          1691 => x"39",
          1692 => x"74",
          1693 => x"3f",
          1694 => x"08",
          1695 => x"f4",
          1696 => x"b9",
          1697 => x"83",
          1698 => x"78",
          1699 => x"d0",
          1700 => x"3f",
          1701 => x"f8",
          1702 => x"02",
          1703 => x"05",
          1704 => x"ff",
          1705 => x"7b",
          1706 => x"fd",
          1707 => x"b9",
          1708 => x"38",
          1709 => x"91",
          1710 => x"2e",
          1711 => x"84",
          1712 => x"8a",
          1713 => x"78",
          1714 => x"a8",
          1715 => x"60",
          1716 => x"c8",
          1717 => x"7e",
          1718 => x"84",
          1719 => x"84",
          1720 => x"8a",
          1721 => x"f3",
          1722 => x"61",
          1723 => x"05",
          1724 => x"33",
          1725 => x"68",
          1726 => x"5c",
          1727 => x"78",
          1728 => x"82",
          1729 => x"83",
          1730 => x"dd",
          1731 => x"d2",
          1732 => x"f7",
          1733 => x"73",
          1734 => x"38",
          1735 => x"81",
          1736 => x"a0",
          1737 => x"38",
          1738 => x"72",
          1739 => x"a7",
          1740 => x"52",
          1741 => x"51",
          1742 => x"81",
          1743 => x"ac",
          1744 => x"a0",
          1745 => x"3f",
          1746 => x"dc",
          1747 => x"90",
          1748 => x"3f",
          1749 => x"79",
          1750 => x"38",
          1751 => x"33",
          1752 => x"55",
          1753 => x"83",
          1754 => x"80",
          1755 => x"27",
          1756 => x"53",
          1757 => x"70",
          1758 => x"56",
          1759 => x"2e",
          1760 => x"fe",
          1761 => x"ee",
          1762 => x"ac",
          1763 => x"51",
          1764 => x"81",
          1765 => x"76",
          1766 => x"83",
          1767 => x"e9",
          1768 => x"18",
          1769 => x"58",
          1770 => x"c3",
          1771 => x"c8",
          1772 => x"70",
          1773 => x"54",
          1774 => x"81",
          1775 => x"9b",
          1776 => x"38",
          1777 => x"76",
          1778 => x"b9",
          1779 => x"84",
          1780 => x"8f",
          1781 => x"83",
          1782 => x"dc",
          1783 => x"14",
          1784 => x"08",
          1785 => x"51",
          1786 => x"78",
          1787 => x"b8",
          1788 => x"39",
          1789 => x"51",
          1790 => x"82",
          1791 => x"ac",
          1792 => x"a0",
          1793 => x"3f",
          1794 => x"fe",
          1795 => x"18",
          1796 => x"27",
          1797 => x"22",
          1798 => x"9c",
          1799 => x"3f",
          1800 => x"d5",
          1801 => x"54",
          1802 => x"c5",
          1803 => x"26",
          1804 => x"99",
          1805 => x"a4",
          1806 => x"3f",
          1807 => x"d5",
          1808 => x"54",
          1809 => x"a9",
          1810 => x"27",
          1811 => x"73",
          1812 => x"7a",
          1813 => x"72",
          1814 => x"d1",
          1815 => x"ab",
          1816 => x"84",
          1817 => x"53",
          1818 => x"ea",
          1819 => x"74",
          1820 => x"fd",
          1821 => x"d5",
          1822 => x"73",
          1823 => x"3f",
          1824 => x"fe",
          1825 => x"ce",
          1826 => x"b9",
          1827 => x"ff",
          1828 => x"59",
          1829 => x"fc",
          1830 => x"59",
          1831 => x"2e",
          1832 => x"fc",
          1833 => x"59",
          1834 => x"80",
          1835 => x"3f",
          1836 => x"08",
          1837 => x"98",
          1838 => x"32",
          1839 => x"9b",
          1840 => x"70",
          1841 => x"75",
          1842 => x"55",
          1843 => x"58",
          1844 => x"25",
          1845 => x"80",
          1846 => x"3f",
          1847 => x"08",
          1848 => x"98",
          1849 => x"32",
          1850 => x"9b",
          1851 => x"70",
          1852 => x"75",
          1853 => x"55",
          1854 => x"58",
          1855 => x"24",
          1856 => x"fd",
          1857 => x"0b",
          1858 => x"0c",
          1859 => x"04",
          1860 => x"87",
          1861 => x"08",
          1862 => x"3f",
          1863 => x"88",
          1864 => x"c0",
          1865 => x"3f",
          1866 => x"fc",
          1867 => x"2a",
          1868 => x"51",
          1869 => x"b7",
          1870 => x"2a",
          1871 => x"51",
          1872 => x"89",
          1873 => x"2a",
          1874 => x"51",
          1875 => x"db",
          1876 => x"2a",
          1877 => x"51",
          1878 => x"ad",
          1879 => x"2a",
          1880 => x"51",
          1881 => x"ff",
          1882 => x"2a",
          1883 => x"51",
          1884 => x"d2",
          1885 => x"2a",
          1886 => x"51",
          1887 => x"38",
          1888 => x"81",
          1889 => x"88",
          1890 => x"3f",
          1891 => x"04",
          1892 => x"94",
          1893 => x"d8",
          1894 => x"3f",
          1895 => x"88",
          1896 => x"3f",
          1897 => x"04",
          1898 => x"fc",
          1899 => x"ec",
          1900 => x"3f",
          1901 => x"f0",
          1902 => x"2a",
          1903 => x"72",
          1904 => x"38",
          1905 => x"51",
          1906 => x"83",
          1907 => x"9b",
          1908 => x"51",
          1909 => x"72",
          1910 => x"81",
          1911 => x"71",
          1912 => x"9c",
          1913 => x"81",
          1914 => x"3f",
          1915 => x"51",
          1916 => x"80",
          1917 => x"3f",
          1918 => x"70",
          1919 => x"52",
          1920 => x"fe",
          1921 => x"be",
          1922 => x"9b",
          1923 => x"d4",
          1924 => x"ac",
          1925 => x"9b",
          1926 => x"85",
          1927 => x"06",
          1928 => x"80",
          1929 => x"38",
          1930 => x"81",
          1931 => x"3f",
          1932 => x"51",
          1933 => x"80",
          1934 => x"3f",
          1935 => x"70",
          1936 => x"52",
          1937 => x"fe",
          1938 => x"bd",
          1939 => x"9a",
          1940 => x"d4",
          1941 => x"e8",
          1942 => x"9a",
          1943 => x"83",
          1944 => x"06",
          1945 => x"80",
          1946 => x"38",
          1947 => x"81",
          1948 => x"3f",
          1949 => x"51",
          1950 => x"80",
          1951 => x"3f",
          1952 => x"70",
          1953 => x"52",
          1954 => x"fd",
          1955 => x"bd",
          1956 => x"0d",
          1957 => x"41",
          1958 => x"d0",
          1959 => x"81",
          1960 => x"81",
          1961 => x"84",
          1962 => x"81",
          1963 => x"3d",
          1964 => x"61",
          1965 => x"38",
          1966 => x"51",
          1967 => x"98",
          1968 => x"d5",
          1969 => x"c3",
          1970 => x"80",
          1971 => x"52",
          1972 => x"ae",
          1973 => x"83",
          1974 => x"70",
          1975 => x"5b",
          1976 => x"2e",
          1977 => x"79",
          1978 => x"88",
          1979 => x"ff",
          1980 => x"82",
          1981 => x"38",
          1982 => x"5a",
          1983 => x"83",
          1984 => x"33",
          1985 => x"2e",
          1986 => x"8c",
          1987 => x"70",
          1988 => x"7b",
          1989 => x"38",
          1990 => x"9b",
          1991 => x"7b",
          1992 => x"ee",
          1993 => x"08",
          1994 => x"ff",
          1995 => x"c8",
          1996 => x"c8",
          1997 => x"53",
          1998 => x"5d",
          1999 => x"84",
          2000 => x"8b",
          2001 => x"33",
          2002 => x"2e",
          2003 => x"81",
          2004 => x"ff",
          2005 => x"9b",
          2006 => x"38",
          2007 => x"5c",
          2008 => x"fe",
          2009 => x"f8",
          2010 => x"e9",
          2011 => x"b9",
          2012 => x"84",
          2013 => x"80",
          2014 => x"38",
          2015 => x"08",
          2016 => x"ff",
          2017 => x"91",
          2018 => x"b9",
          2019 => x"62",
          2020 => x"7a",
          2021 => x"84",
          2022 => x"c8",
          2023 => x"8b",
          2024 => x"c8",
          2025 => x"80",
          2026 => x"0b",
          2027 => x"5b",
          2028 => x"8d",
          2029 => x"82",
          2030 => x"38",
          2031 => x"82",
          2032 => x"54",
          2033 => x"d5",
          2034 => x"51",
          2035 => x"83",
          2036 => x"84",
          2037 => x"7d",
          2038 => x"80",
          2039 => x"0a",
          2040 => x"0a",
          2041 => x"f5",
          2042 => x"b9",
          2043 => x"b9",
          2044 => x"70",
          2045 => x"07",
          2046 => x"5b",
          2047 => x"5a",
          2048 => x"83",
          2049 => x"78",
          2050 => x"78",
          2051 => x"38",
          2052 => x"81",
          2053 => x"5a",
          2054 => x"38",
          2055 => x"61",
          2056 => x"5d",
          2057 => x"38",
          2058 => x"81",
          2059 => x"51",
          2060 => x"3f",
          2061 => x"51",
          2062 => x"7e",
          2063 => x"53",
          2064 => x"51",
          2065 => x"0b",
          2066 => x"bc",
          2067 => x"ff",
          2068 => x"79",
          2069 => x"81",
          2070 => x"98",
          2071 => x"d8",
          2072 => x"cd",
          2073 => x"c8",
          2074 => x"38",
          2075 => x"0b",
          2076 => x"34",
          2077 => x"53",
          2078 => x"7e",
          2079 => x"c8",
          2080 => x"c8",
          2081 => x"a0",
          2082 => x"c8",
          2083 => x"e6",
          2084 => x"83",
          2085 => x"70",
          2086 => x"5f",
          2087 => x"2e",
          2088 => x"fc",
          2089 => x"39",
          2090 => x"51",
          2091 => x"3f",
          2092 => x"0b",
          2093 => x"34",
          2094 => x"53",
          2095 => x"7e",
          2096 => x"3f",
          2097 => x"5a",
          2098 => x"38",
          2099 => x"1a",
          2100 => x"1b",
          2101 => x"81",
          2102 => x"80",
          2103 => x"10",
          2104 => x"05",
          2105 => x"04",
          2106 => x"d5",
          2107 => x"51",
          2108 => x"60",
          2109 => x"84",
          2110 => x"82",
          2111 => x"84",
          2112 => x"61",
          2113 => x"06",
          2114 => x"81",
          2115 => x"45",
          2116 => x"ae",
          2117 => x"fc",
          2118 => x"3f",
          2119 => x"92",
          2120 => x"90",
          2121 => x"8c",
          2122 => x"83",
          2123 => x"80",
          2124 => x"94",
          2125 => x"d2",
          2126 => x"93",
          2127 => x"ab",
          2128 => x"39",
          2129 => x"fa",
          2130 => x"52",
          2131 => x"a4",
          2132 => x"39",
          2133 => x"3f",
          2134 => x"83",
          2135 => x"de",
          2136 => x"59",
          2137 => x"d6",
          2138 => x"8a",
          2139 => x"3f",
          2140 => x"b8",
          2141 => x"11",
          2142 => x"05",
          2143 => x"3f",
          2144 => x"08",
          2145 => x"ba",
          2146 => x"83",
          2147 => x"d0",
          2148 => x"5a",
          2149 => x"b9",
          2150 => x"2e",
          2151 => x"84",
          2152 => x"52",
          2153 => x"51",
          2154 => x"fa",
          2155 => x"3d",
          2156 => x"53",
          2157 => x"51",
          2158 => x"84",
          2159 => x"80",
          2160 => x"38",
          2161 => x"d7",
          2162 => x"bf",
          2163 => x"78",
          2164 => x"fe",
          2165 => x"ff",
          2166 => x"e9",
          2167 => x"b9",
          2168 => x"2e",
          2169 => x"b8",
          2170 => x"11",
          2171 => x"05",
          2172 => x"3f",
          2173 => x"08",
          2174 => x"64",
          2175 => x"53",
          2176 => x"d7",
          2177 => x"83",
          2178 => x"a8",
          2179 => x"f8",
          2180 => x"d0",
          2181 => x"48",
          2182 => x"78",
          2183 => x"a2",
          2184 => x"26",
          2185 => x"64",
          2186 => x"46",
          2187 => x"b8",
          2188 => x"11",
          2189 => x"05",
          2190 => x"3f",
          2191 => x"08",
          2192 => x"fe",
          2193 => x"fe",
          2194 => x"ff",
          2195 => x"e8",
          2196 => x"b9",
          2197 => x"b0",
          2198 => x"78",
          2199 => x"52",
          2200 => x"51",
          2201 => x"84",
          2202 => x"53",
          2203 => x"7e",
          2204 => x"3f",
          2205 => x"33",
          2206 => x"2e",
          2207 => x"78",
          2208 => x"ca",
          2209 => x"05",
          2210 => x"cf",
          2211 => x"ff",
          2212 => x"ff",
          2213 => x"e9",
          2214 => x"b9",
          2215 => x"2e",
          2216 => x"b8",
          2217 => x"11",
          2218 => x"05",
          2219 => x"3f",
          2220 => x"08",
          2221 => x"8a",
          2222 => x"fe",
          2223 => x"ff",
          2224 => x"e9",
          2225 => x"b9",
          2226 => x"2e",
          2227 => x"83",
          2228 => x"ce",
          2229 => x"67",
          2230 => x"7c",
          2231 => x"38",
          2232 => x"7a",
          2233 => x"5a",
          2234 => x"95",
          2235 => x"79",
          2236 => x"53",
          2237 => x"d7",
          2238 => x"8f",
          2239 => x"5b",
          2240 => x"81",
          2241 => x"d2",
          2242 => x"ff",
          2243 => x"ff",
          2244 => x"e8",
          2245 => x"b9",
          2246 => x"2e",
          2247 => x"b8",
          2248 => x"11",
          2249 => x"05",
          2250 => x"3f",
          2251 => x"08",
          2252 => x"8e",
          2253 => x"fe",
          2254 => x"ff",
          2255 => x"e8",
          2256 => x"b9",
          2257 => x"2e",
          2258 => x"83",
          2259 => x"cd",
          2260 => x"5a",
          2261 => x"82",
          2262 => x"5c",
          2263 => x"05",
          2264 => x"34",
          2265 => x"46",
          2266 => x"3d",
          2267 => x"53",
          2268 => x"51",
          2269 => x"84",
          2270 => x"80",
          2271 => x"38",
          2272 => x"fc",
          2273 => x"80",
          2274 => x"fd",
          2275 => x"c8",
          2276 => x"68",
          2277 => x"52",
          2278 => x"51",
          2279 => x"84",
          2280 => x"53",
          2281 => x"7e",
          2282 => x"3f",
          2283 => x"33",
          2284 => x"2e",
          2285 => x"78",
          2286 => x"97",
          2287 => x"05",
          2288 => x"68",
          2289 => x"db",
          2290 => x"34",
          2291 => x"49",
          2292 => x"fc",
          2293 => x"80",
          2294 => x"ad",
          2295 => x"c8",
          2296 => x"f5",
          2297 => x"59",
          2298 => x"05",
          2299 => x"68",
          2300 => x"b8",
          2301 => x"11",
          2302 => x"05",
          2303 => x"3f",
          2304 => x"08",
          2305 => x"f5",
          2306 => x"3d",
          2307 => x"53",
          2308 => x"51",
          2309 => x"84",
          2310 => x"80",
          2311 => x"38",
          2312 => x"fc",
          2313 => x"80",
          2314 => x"dd",
          2315 => x"c8",
          2316 => x"f5",
          2317 => x"3d",
          2318 => x"53",
          2319 => x"51",
          2320 => x"84",
          2321 => x"86",
          2322 => x"c8",
          2323 => x"d8",
          2324 => x"b7",
          2325 => x"5b",
          2326 => x"27",
          2327 => x"5b",
          2328 => x"84",
          2329 => x"79",
          2330 => x"38",
          2331 => x"f1",
          2332 => x"39",
          2333 => x"80",
          2334 => x"b1",
          2335 => x"c8",
          2336 => x"ff",
          2337 => x"59",
          2338 => x"81",
          2339 => x"c8",
          2340 => x"51",
          2341 => x"84",
          2342 => x"80",
          2343 => x"38",
          2344 => x"08",
          2345 => x"3f",
          2346 => x"b8",
          2347 => x"11",
          2348 => x"05",
          2349 => x"3f",
          2350 => x"08",
          2351 => x"f2",
          2352 => x"79",
          2353 => x"c0",
          2354 => x"84",
          2355 => x"3d",
          2356 => x"53",
          2357 => x"51",
          2358 => x"84",
          2359 => x"91",
          2360 => x"cc",
          2361 => x"80",
          2362 => x"38",
          2363 => x"08",
          2364 => x"fe",
          2365 => x"ff",
          2366 => x"e5",
          2367 => x"b9",
          2368 => x"2e",
          2369 => x"66",
          2370 => x"88",
          2371 => x"81",
          2372 => x"32",
          2373 => x"72",
          2374 => x"7e",
          2375 => x"5d",
          2376 => x"88",
          2377 => x"2e",
          2378 => x"46",
          2379 => x"51",
          2380 => x"80",
          2381 => x"65",
          2382 => x"68",
          2383 => x"3f",
          2384 => x"51",
          2385 => x"f2",
          2386 => x"64",
          2387 => x"64",
          2388 => x"b8",
          2389 => x"11",
          2390 => x"05",
          2391 => x"3f",
          2392 => x"08",
          2393 => x"da",
          2394 => x"71",
          2395 => x"84",
          2396 => x"3d",
          2397 => x"53",
          2398 => x"51",
          2399 => x"84",
          2400 => x"c6",
          2401 => x"39",
          2402 => x"80",
          2403 => x"7e",
          2404 => x"40",
          2405 => x"b8",
          2406 => x"11",
          2407 => x"05",
          2408 => x"3f",
          2409 => x"08",
          2410 => x"96",
          2411 => x"02",
          2412 => x"22",
          2413 => x"05",
          2414 => x"45",
          2415 => x"f0",
          2416 => x"80",
          2417 => x"bd",
          2418 => x"c8",
          2419 => x"38",
          2420 => x"b8",
          2421 => x"11",
          2422 => x"05",
          2423 => x"3f",
          2424 => x"08",
          2425 => x"dc",
          2426 => x"02",
          2427 => x"33",
          2428 => x"81",
          2429 => x"9b",
          2430 => x"fe",
          2431 => x"ff",
          2432 => x"e1",
          2433 => x"b9",
          2434 => x"2e",
          2435 => x"64",
          2436 => x"5d",
          2437 => x"70",
          2438 => x"e1",
          2439 => x"2e",
          2440 => x"f3",
          2441 => x"55",
          2442 => x"54",
          2443 => x"d8",
          2444 => x"51",
          2445 => x"f3",
          2446 => x"52",
          2447 => x"8a",
          2448 => x"39",
          2449 => x"51",
          2450 => x"f0",
          2451 => x"3d",
          2452 => x"53",
          2453 => x"51",
          2454 => x"84",
          2455 => x"80",
          2456 => x"64",
          2457 => x"ce",
          2458 => x"70",
          2459 => x"23",
          2460 => x"e7",
          2461 => x"cd",
          2462 => x"80",
          2463 => x"38",
          2464 => x"08",
          2465 => x"39",
          2466 => x"33",
          2467 => x"2e",
          2468 => x"f2",
          2469 => x"fc",
          2470 => x"d8",
          2471 => x"d6",
          2472 => x"f7",
          2473 => x"d8",
          2474 => x"ca",
          2475 => x"f6",
          2476 => x"f2",
          2477 => x"78",
          2478 => x"38",
          2479 => x"08",
          2480 => x"39",
          2481 => x"51",
          2482 => x"f9",
          2483 => x"f2",
          2484 => x"78",
          2485 => x"38",
          2486 => x"08",
          2487 => x"39",
          2488 => x"33",
          2489 => x"2e",
          2490 => x"f2",
          2491 => x"fb",
          2492 => x"f2",
          2493 => x"7d",
          2494 => x"38",
          2495 => x"08",
          2496 => x"39",
          2497 => x"33",
          2498 => x"2e",
          2499 => x"f2",
          2500 => x"fb",
          2501 => x"f2",
          2502 => x"7c",
          2503 => x"38",
          2504 => x"08",
          2505 => x"39",
          2506 => x"08",
          2507 => x"49",
          2508 => x"83",
          2509 => x"88",
          2510 => x"b5",
          2511 => x"0d",
          2512 => x"b9",
          2513 => x"c0",
          2514 => x"08",
          2515 => x"84",
          2516 => x"51",
          2517 => x"84",
          2518 => x"90",
          2519 => x"57",
          2520 => x"80",
          2521 => x"da",
          2522 => x"84",
          2523 => x"07",
          2524 => x"c0",
          2525 => x"08",
          2526 => x"84",
          2527 => x"51",
          2528 => x"84",
          2529 => x"90",
          2530 => x"57",
          2531 => x"80",
          2532 => x"da",
          2533 => x"84",
          2534 => x"07",
          2535 => x"80",
          2536 => x"c0",
          2537 => x"8c",
          2538 => x"87",
          2539 => x"0c",
          2540 => x"5c",
          2541 => x"5d",
          2542 => x"05",
          2543 => x"80",
          2544 => x"a8",
          2545 => x"70",
          2546 => x"70",
          2547 => x"d5",
          2548 => x"b7",
          2549 => x"9e",
          2550 => x"3f",
          2551 => x"95",
          2552 => x"d2",
          2553 => x"d2",
          2554 => x"9f",
          2555 => x"b8",
          2556 => x"55",
          2557 => x"83",
          2558 => x"83",
          2559 => x"81",
          2560 => x"83",
          2561 => x"c4",
          2562 => x"b2",
          2563 => x"ec",
          2564 => x"3f",
          2565 => x"d2",
          2566 => x"ef",
          2567 => x"0a",
          2568 => x"98",
          2569 => x"3f",
          2570 => x"80",
          2571 => x"0d",
          2572 => x"56",
          2573 => x"52",
          2574 => x"2e",
          2575 => x"74",
          2576 => x"ff",
          2577 => x"70",
          2578 => x"81",
          2579 => x"81",
          2580 => x"70",
          2581 => x"53",
          2582 => x"a0",
          2583 => x"71",
          2584 => x"54",
          2585 => x"81",
          2586 => x"52",
          2587 => x"80",
          2588 => x"72",
          2589 => x"ff",
          2590 => x"54",
          2591 => x"83",
          2592 => x"70",
          2593 => x"38",
          2594 => x"86",
          2595 => x"52",
          2596 => x"73",
          2597 => x"52",
          2598 => x"2e",
          2599 => x"83",
          2600 => x"70",
          2601 => x"30",
          2602 => x"76",
          2603 => x"53",
          2604 => x"88",
          2605 => x"70",
          2606 => x"34",
          2607 => x"74",
          2608 => x"b9",
          2609 => x"3d",
          2610 => x"80",
          2611 => x"73",
          2612 => x"be",
          2613 => x"52",
          2614 => x"70",
          2615 => x"53",
          2616 => x"a2",
          2617 => x"81",
          2618 => x"81",
          2619 => x"75",
          2620 => x"81",
          2621 => x"06",
          2622 => x"dc",
          2623 => x"0d",
          2624 => x"08",
          2625 => x"0b",
          2626 => x"0c",
          2627 => x"04",
          2628 => x"05",
          2629 => x"da",
          2630 => x"b9",
          2631 => x"2e",
          2632 => x"84",
          2633 => x"86",
          2634 => x"fc",
          2635 => x"82",
          2636 => x"05",
          2637 => x"52",
          2638 => x"81",
          2639 => x"13",
          2640 => x"54",
          2641 => x"9e",
          2642 => x"38",
          2643 => x"51",
          2644 => x"97",
          2645 => x"38",
          2646 => x"54",
          2647 => x"bb",
          2648 => x"38",
          2649 => x"55",
          2650 => x"bb",
          2651 => x"38",
          2652 => x"55",
          2653 => x"87",
          2654 => x"d9",
          2655 => x"22",
          2656 => x"73",
          2657 => x"80",
          2658 => x"0b",
          2659 => x"9c",
          2660 => x"87",
          2661 => x"0c",
          2662 => x"87",
          2663 => x"0c",
          2664 => x"87",
          2665 => x"0c",
          2666 => x"87",
          2667 => x"0c",
          2668 => x"87",
          2669 => x"0c",
          2670 => x"87",
          2671 => x"0c",
          2672 => x"98",
          2673 => x"87",
          2674 => x"0c",
          2675 => x"c0",
          2676 => x"80",
          2677 => x"b9",
          2678 => x"3d",
          2679 => x"3d",
          2680 => x"87",
          2681 => x"5d",
          2682 => x"87",
          2683 => x"08",
          2684 => x"23",
          2685 => x"b8",
          2686 => x"82",
          2687 => x"c0",
          2688 => x"5a",
          2689 => x"34",
          2690 => x"b0",
          2691 => x"84",
          2692 => x"c0",
          2693 => x"5a",
          2694 => x"34",
          2695 => x"a8",
          2696 => x"86",
          2697 => x"c0",
          2698 => x"5c",
          2699 => x"23",
          2700 => x"a0",
          2701 => x"8a",
          2702 => x"7d",
          2703 => x"ff",
          2704 => x"7b",
          2705 => x"06",
          2706 => x"33",
          2707 => x"33",
          2708 => x"33",
          2709 => x"33",
          2710 => x"33",
          2711 => x"ff",
          2712 => x"83",
          2713 => x"ff",
          2714 => x"8f",
          2715 => x"fe",
          2716 => x"93",
          2717 => x"72",
          2718 => x"38",
          2719 => x"e8",
          2720 => x"b9",
          2721 => x"2b",
          2722 => x"51",
          2723 => x"2e",
          2724 => x"86",
          2725 => x"2e",
          2726 => x"84",
          2727 => x"84",
          2728 => x"72",
          2729 => x"ff",
          2730 => x"c8",
          2731 => x"70",
          2732 => x"52",
          2733 => x"09",
          2734 => x"38",
          2735 => x"e7",
          2736 => x"b9",
          2737 => x"2b",
          2738 => x"51",
          2739 => x"2e",
          2740 => x"39",
          2741 => x"80",
          2742 => x"71",
          2743 => x"81",
          2744 => x"c3",
          2745 => x"c8",
          2746 => x"70",
          2747 => x"52",
          2748 => x"eb",
          2749 => x"07",
          2750 => x"52",
          2751 => x"db",
          2752 => x"b9",
          2753 => x"3d",
          2754 => x"3d",
          2755 => x"05",
          2756 => x"80",
          2757 => x"ff",
          2758 => x"55",
          2759 => x"80",
          2760 => x"c0",
          2761 => x"70",
          2762 => x"81",
          2763 => x"52",
          2764 => x"8c",
          2765 => x"2a",
          2766 => x"51",
          2767 => x"38",
          2768 => x"81",
          2769 => x"80",
          2770 => x"71",
          2771 => x"06",
          2772 => x"38",
          2773 => x"06",
          2774 => x"94",
          2775 => x"80",
          2776 => x"87",
          2777 => x"52",
          2778 => x"74",
          2779 => x"0c",
          2780 => x"04",
          2781 => x"70",
          2782 => x"51",
          2783 => x"72",
          2784 => x"06",
          2785 => x"2e",
          2786 => x"93",
          2787 => x"52",
          2788 => x"c0",
          2789 => x"94",
          2790 => x"96",
          2791 => x"06",
          2792 => x"70",
          2793 => x"39",
          2794 => x"02",
          2795 => x"70",
          2796 => x"2a",
          2797 => x"70",
          2798 => x"34",
          2799 => x"04",
          2800 => x"78",
          2801 => x"33",
          2802 => x"57",
          2803 => x"80",
          2804 => x"15",
          2805 => x"33",
          2806 => x"06",
          2807 => x"71",
          2808 => x"ff",
          2809 => x"94",
          2810 => x"96",
          2811 => x"06",
          2812 => x"70",
          2813 => x"38",
          2814 => x"70",
          2815 => x"51",
          2816 => x"72",
          2817 => x"06",
          2818 => x"2e",
          2819 => x"93",
          2820 => x"52",
          2821 => x"75",
          2822 => x"51",
          2823 => x"80",
          2824 => x"2e",
          2825 => x"c0",
          2826 => x"73",
          2827 => x"17",
          2828 => x"57",
          2829 => x"38",
          2830 => x"c8",
          2831 => x"0d",
          2832 => x"2a",
          2833 => x"51",
          2834 => x"38",
          2835 => x"81",
          2836 => x"80",
          2837 => x"71",
          2838 => x"06",
          2839 => x"2e",
          2840 => x"87",
          2841 => x"08",
          2842 => x"70",
          2843 => x"54",
          2844 => x"38",
          2845 => x"3d",
          2846 => x"9e",
          2847 => x"9c",
          2848 => x"52",
          2849 => x"2e",
          2850 => x"87",
          2851 => x"08",
          2852 => x"0c",
          2853 => x"a8",
          2854 => x"88",
          2855 => x"9e",
          2856 => x"f2",
          2857 => x"c0",
          2858 => x"83",
          2859 => x"87",
          2860 => x"08",
          2861 => x"0c",
          2862 => x"a0",
          2863 => x"98",
          2864 => x"9e",
          2865 => x"f2",
          2866 => x"c0",
          2867 => x"83",
          2868 => x"87",
          2869 => x"08",
          2870 => x"0c",
          2871 => x"b8",
          2872 => x"a8",
          2873 => x"9e",
          2874 => x"f2",
          2875 => x"c0",
          2876 => x"83",
          2877 => x"87",
          2878 => x"08",
          2879 => x"0c",
          2880 => x"80",
          2881 => x"83",
          2882 => x"87",
          2883 => x"08",
          2884 => x"0c",
          2885 => x"88",
          2886 => x"c0",
          2887 => x"9e",
          2888 => x"f2",
          2889 => x"0b",
          2890 => x"34",
          2891 => x"c0",
          2892 => x"70",
          2893 => x"06",
          2894 => x"70",
          2895 => x"71",
          2896 => x"34",
          2897 => x"c0",
          2898 => x"70",
          2899 => x"06",
          2900 => x"70",
          2901 => x"38",
          2902 => x"83",
          2903 => x"80",
          2904 => x"9e",
          2905 => x"90",
          2906 => x"51",
          2907 => x"80",
          2908 => x"81",
          2909 => x"f2",
          2910 => x"0b",
          2911 => x"90",
          2912 => x"80",
          2913 => x"52",
          2914 => x"2e",
          2915 => x"52",
          2916 => x"cc",
          2917 => x"87",
          2918 => x"08",
          2919 => x"80",
          2920 => x"52",
          2921 => x"83",
          2922 => x"71",
          2923 => x"34",
          2924 => x"c0",
          2925 => x"70",
          2926 => x"06",
          2927 => x"70",
          2928 => x"38",
          2929 => x"83",
          2930 => x"80",
          2931 => x"9e",
          2932 => x"84",
          2933 => x"51",
          2934 => x"80",
          2935 => x"81",
          2936 => x"f2",
          2937 => x"0b",
          2938 => x"90",
          2939 => x"80",
          2940 => x"52",
          2941 => x"2e",
          2942 => x"52",
          2943 => x"d0",
          2944 => x"87",
          2945 => x"08",
          2946 => x"80",
          2947 => x"52",
          2948 => x"83",
          2949 => x"71",
          2950 => x"34",
          2951 => x"c0",
          2952 => x"70",
          2953 => x"06",
          2954 => x"70",
          2955 => x"38",
          2956 => x"83",
          2957 => x"80",
          2958 => x"9e",
          2959 => x"a0",
          2960 => x"52",
          2961 => x"2e",
          2962 => x"52",
          2963 => x"d3",
          2964 => x"9e",
          2965 => x"80",
          2966 => x"2a",
          2967 => x"83",
          2968 => x"80",
          2969 => x"9e",
          2970 => x"84",
          2971 => x"52",
          2972 => x"2e",
          2973 => x"52",
          2974 => x"d5",
          2975 => x"9e",
          2976 => x"f0",
          2977 => x"2a",
          2978 => x"83",
          2979 => x"80",
          2980 => x"9e",
          2981 => x"88",
          2982 => x"52",
          2983 => x"83",
          2984 => x"71",
          2985 => x"34",
          2986 => x"90",
          2987 => x"51",
          2988 => x"d8",
          2989 => x"0d",
          2990 => x"fd",
          2991 => x"3d",
          2992 => x"84",
          2993 => x"c3",
          2994 => x"c8",
          2995 => x"86",
          2996 => x"d9",
          2997 => x"9e",
          2998 => x"ca",
          2999 => x"85",
          3000 => x"f2",
          3001 => x"73",
          3002 => x"83",
          3003 => x"56",
          3004 => x"38",
          3005 => x"33",
          3006 => x"f4",
          3007 => x"ce",
          3008 => x"84",
          3009 => x"f2",
          3010 => x"75",
          3011 => x"83",
          3012 => x"54",
          3013 => x"38",
          3014 => x"33",
          3015 => x"e2",
          3016 => x"c9",
          3017 => x"83",
          3018 => x"f2",
          3019 => x"73",
          3020 => x"83",
          3021 => x"55",
          3022 => x"38",
          3023 => x"33",
          3024 => x"e9",
          3025 => x"d2",
          3026 => x"81",
          3027 => x"d9",
          3028 => x"a2",
          3029 => x"ac",
          3030 => x"d9",
          3031 => x"b5",
          3032 => x"f2",
          3033 => x"83",
          3034 => x"ff",
          3035 => x"83",
          3036 => x"52",
          3037 => x"51",
          3038 => x"3f",
          3039 => x"51",
          3040 => x"83",
          3041 => x"52",
          3042 => x"51",
          3043 => x"3f",
          3044 => x"08",
          3045 => x"c0",
          3046 => x"ca",
          3047 => x"b9",
          3048 => x"84",
          3049 => x"71",
          3050 => x"84",
          3051 => x"52",
          3052 => x"51",
          3053 => x"3f",
          3054 => x"33",
          3055 => x"38",
          3056 => x"33",
          3057 => x"38",
          3058 => x"04",
          3059 => x"08",
          3060 => x"c0",
          3061 => x"c9",
          3062 => x"b9",
          3063 => x"84",
          3064 => x"71",
          3065 => x"84",
          3066 => x"52",
          3067 => x"51",
          3068 => x"3f",
          3069 => x"04",
          3070 => x"08",
          3071 => x"c0",
          3072 => x"c9",
          3073 => x"b9",
          3074 => x"84",
          3075 => x"71",
          3076 => x"84",
          3077 => x"52",
          3078 => x"51",
          3079 => x"3f",
          3080 => x"33",
          3081 => x"2e",
          3082 => x"ff",
          3083 => x"db",
          3084 => x"c2",
          3085 => x"b0",
          3086 => x"3f",
          3087 => x"08",
          3088 => x"bc",
          3089 => x"c3",
          3090 => x"b0",
          3091 => x"d9",
          3092 => x"b3",
          3093 => x"f2",
          3094 => x"83",
          3095 => x"ff",
          3096 => x"83",
          3097 => x"c0",
          3098 => x"f2",
          3099 => x"83",
          3100 => x"ff",
          3101 => x"83",
          3102 => x"56",
          3103 => x"52",
          3104 => x"a4",
          3105 => x"c8",
          3106 => x"c0",
          3107 => x"31",
          3108 => x"b9",
          3109 => x"83",
          3110 => x"ff",
          3111 => x"83",
          3112 => x"55",
          3113 => x"fe",
          3114 => x"cc",
          3115 => x"f0",
          3116 => x"c2",
          3117 => x"d2",
          3118 => x"80",
          3119 => x"38",
          3120 => x"83",
          3121 => x"ff",
          3122 => x"83",
          3123 => x"56",
          3124 => x"fc",
          3125 => x"39",
          3126 => x"51",
          3127 => x"3f",
          3128 => x"33",
          3129 => x"2e",
          3130 => x"d7",
          3131 => x"90",
          3132 => x"82",
          3133 => x"cb",
          3134 => x"80",
          3135 => x"38",
          3136 => x"f2",
          3137 => x"83",
          3138 => x"ff",
          3139 => x"83",
          3140 => x"56",
          3141 => x"fc",
          3142 => x"39",
          3143 => x"33",
          3144 => x"c4",
          3145 => x"e3",
          3146 => x"d5",
          3147 => x"80",
          3148 => x"38",
          3149 => x"f2",
          3150 => x"83",
          3151 => x"ff",
          3152 => x"83",
          3153 => x"54",
          3154 => x"fb",
          3155 => x"39",
          3156 => x"08",
          3157 => x"08",
          3158 => x"83",
          3159 => x"ff",
          3160 => x"83",
          3161 => x"56",
          3162 => x"fb",
          3163 => x"39",
          3164 => x"08",
          3165 => x"08",
          3166 => x"83",
          3167 => x"ff",
          3168 => x"83",
          3169 => x"54",
          3170 => x"fa",
          3171 => x"39",
          3172 => x"08",
          3173 => x"08",
          3174 => x"83",
          3175 => x"ff",
          3176 => x"83",
          3177 => x"55",
          3178 => x"fa",
          3179 => x"39",
          3180 => x"08",
          3181 => x"08",
          3182 => x"83",
          3183 => x"ff",
          3184 => x"83",
          3185 => x"56",
          3186 => x"fa",
          3187 => x"39",
          3188 => x"08",
          3189 => x"08",
          3190 => x"83",
          3191 => x"ff",
          3192 => x"83",
          3193 => x"54",
          3194 => x"f9",
          3195 => x"39",
          3196 => x"51",
          3197 => x"3f",
          3198 => x"51",
          3199 => x"3f",
          3200 => x"33",
          3201 => x"2e",
          3202 => x"c4",
          3203 => x"0d",
          3204 => x"33",
          3205 => x"26",
          3206 => x"10",
          3207 => x"fc",
          3208 => x"08",
          3209 => x"a4",
          3210 => x"df",
          3211 => x"0d",
          3212 => x"ac",
          3213 => x"d3",
          3214 => x"0d",
          3215 => x"b4",
          3216 => x"c7",
          3217 => x"0d",
          3218 => x"bc",
          3219 => x"bb",
          3220 => x"0d",
          3221 => x"c4",
          3222 => x"af",
          3223 => x"0d",
          3224 => x"cc",
          3225 => x"a3",
          3226 => x"0d",
          3227 => x"80",
          3228 => x"0b",
          3229 => x"84",
          3230 => x"f2",
          3231 => x"c0",
          3232 => x"04",
          3233 => x"aa",
          3234 => x"3d",
          3235 => x"81",
          3236 => x"80",
          3237 => x"b4",
          3238 => x"88",
          3239 => x"b9",
          3240 => x"ed",
          3241 => x"57",
          3242 => x"f3",
          3243 => x"55",
          3244 => x"76",
          3245 => x"90",
          3246 => x"c8",
          3247 => x"a4",
          3248 => x"c0",
          3249 => x"b9",
          3250 => x"17",
          3251 => x"0b",
          3252 => x"08",
          3253 => x"84",
          3254 => x"ff",
          3255 => x"55",
          3256 => x"34",
          3257 => x"30",
          3258 => x"9f",
          3259 => x"55",
          3260 => x"85",
          3261 => x"b0",
          3262 => x"b4",
          3263 => x"08",
          3264 => x"87",
          3265 => x"b9",
          3266 => x"38",
          3267 => x"9a",
          3268 => x"b9",
          3269 => x"3d",
          3270 => x"e1",
          3271 => x"ad",
          3272 => x"76",
          3273 => x"06",
          3274 => x"52",
          3275 => x"9a",
          3276 => x"ff",
          3277 => x"ab",
          3278 => x"84",
          3279 => x"76",
          3280 => x"83",
          3281 => x"ff",
          3282 => x"80",
          3283 => x"c8",
          3284 => x"0d",
          3285 => x"0d",
          3286 => x"ad",
          3287 => x"72",
          3288 => x"57",
          3289 => x"73",
          3290 => x"91",
          3291 => x"8d",
          3292 => x"75",
          3293 => x"83",
          3294 => x"70",
          3295 => x"ff",
          3296 => x"84",
          3297 => x"53",
          3298 => x"08",
          3299 => x"3f",
          3300 => x"08",
          3301 => x"14",
          3302 => x"81",
          3303 => x"38",
          3304 => x"99",
          3305 => x"70",
          3306 => x"57",
          3307 => x"27",
          3308 => x"54",
          3309 => x"c8",
          3310 => x"0d",
          3311 => x"5a",
          3312 => x"84",
          3313 => x"80",
          3314 => x"bd",
          3315 => x"c8",
          3316 => x"d1",
          3317 => x"53",
          3318 => x"51",
          3319 => x"84",
          3320 => x"81",
          3321 => x"73",
          3322 => x"38",
          3323 => x"81",
          3324 => x"54",
          3325 => x"fe",
          3326 => x"b6",
          3327 => x"77",
          3328 => x"76",
          3329 => x"38",
          3330 => x"5b",
          3331 => x"55",
          3332 => x"09",
          3333 => x"d5",
          3334 => x"26",
          3335 => x"0b",
          3336 => x"56",
          3337 => x"73",
          3338 => x"08",
          3339 => x"b4",
          3340 => x"82",
          3341 => x"84",
          3342 => x"80",
          3343 => x"f3",
          3344 => x"80",
          3345 => x"51",
          3346 => x"3f",
          3347 => x"08",
          3348 => x"38",
          3349 => x"bd",
          3350 => x"b9",
          3351 => x"80",
          3352 => x"c8",
          3353 => x"38",
          3354 => x"08",
          3355 => x"19",
          3356 => x"77",
          3357 => x"75",
          3358 => x"83",
          3359 => x"56",
          3360 => x"3f",
          3361 => x"09",
          3362 => x"b2",
          3363 => x"84",
          3364 => x"aa",
          3365 => x"ce",
          3366 => x"3d",
          3367 => x"08",
          3368 => x"5a",
          3369 => x"0b",
          3370 => x"83",
          3371 => x"83",
          3372 => x"56",
          3373 => x"38",
          3374 => x"b0",
          3375 => x"74",
          3376 => x"cb",
          3377 => x"2e",
          3378 => x"81",
          3379 => x"5a",
          3380 => x"a0",
          3381 => x"2e",
          3382 => x"93",
          3383 => x"5f",
          3384 => x"eb",
          3385 => x"b9",
          3386 => x"2b",
          3387 => x"5b",
          3388 => x"2e",
          3389 => x"81",
          3390 => x"d1",
          3391 => x"98",
          3392 => x"2c",
          3393 => x"33",
          3394 => x"70",
          3395 => x"98",
          3396 => x"10",
          3397 => x"d0",
          3398 => x"15",
          3399 => x"53",
          3400 => x"52",
          3401 => x"59",
          3402 => x"79",
          3403 => x"38",
          3404 => x"81",
          3405 => x"81",
          3406 => x"81",
          3407 => x"70",
          3408 => x"55",
          3409 => x"81",
          3410 => x"10",
          3411 => x"2b",
          3412 => x"0b",
          3413 => x"16",
          3414 => x"77",
          3415 => x"38",
          3416 => x"15",
          3417 => x"33",
          3418 => x"75",
          3419 => x"38",
          3420 => x"c2",
          3421 => x"d1",
          3422 => x"57",
          3423 => x"81",
          3424 => x"1b",
          3425 => x"70",
          3426 => x"d1",
          3427 => x"98",
          3428 => x"2c",
          3429 => x"05",
          3430 => x"83",
          3431 => x"33",
          3432 => x"5d",
          3433 => x"57",
          3434 => x"81",
          3435 => x"84",
          3436 => x"fe",
          3437 => x"57",
          3438 => x"38",
          3439 => x"0a",
          3440 => x"0a",
          3441 => x"2c",
          3442 => x"06",
          3443 => x"76",
          3444 => x"c0",
          3445 => x"16",
          3446 => x"51",
          3447 => x"83",
          3448 => x"33",
          3449 => x"61",
          3450 => x"83",
          3451 => x"08",
          3452 => x"42",
          3453 => x"2e",
          3454 => x"76",
          3455 => x"bc",
          3456 => x"39",
          3457 => x"80",
          3458 => x"38",
          3459 => x"81",
          3460 => x"39",
          3461 => x"fe",
          3462 => x"84",
          3463 => x"76",
          3464 => x"34",
          3465 => x"76",
          3466 => x"55",
          3467 => x"fd",
          3468 => x"10",
          3469 => x"94",
          3470 => x"08",
          3471 => x"d8",
          3472 => x"0c",
          3473 => x"d1",
          3474 => x"0b",
          3475 => x"34",
          3476 => x"d1",
          3477 => x"75",
          3478 => x"85",
          3479 => x"ac",
          3480 => x"51",
          3481 => x"3f",
          3482 => x"33",
          3483 => x"76",
          3484 => x"34",
          3485 => x"84",
          3486 => x"70",
          3487 => x"84",
          3488 => x"5b",
          3489 => x"79",
          3490 => x"38",
          3491 => x"08",
          3492 => x"58",
          3493 => x"8c",
          3494 => x"70",
          3495 => x"ff",
          3496 => x"fc",
          3497 => x"93",
          3498 => x"38",
          3499 => x"83",
          3500 => x"70",
          3501 => x"75",
          3502 => x"75",
          3503 => x"34",
          3504 => x"84",
          3505 => x"84",
          3506 => x"56",
          3507 => x"2e",
          3508 => x"d5",
          3509 => x"88",
          3510 => x"95",
          3511 => x"ac",
          3512 => x"51",
          3513 => x"3f",
          3514 => x"08",
          3515 => x"ff",
          3516 => x"84",
          3517 => x"ff",
          3518 => x"84",
          3519 => x"7a",
          3520 => x"55",
          3521 => x"7b",
          3522 => x"ff",
          3523 => x"d1",
          3524 => x"cd",
          3525 => x"38",
          3526 => x"08",
          3527 => x"9e",
          3528 => x"10",
          3529 => x"05",
          3530 => x"57",
          3531 => x"f9",
          3532 => x"56",
          3533 => x"fb",
          3534 => x"51",
          3535 => x"3f",
          3536 => x"08",
          3537 => x"34",
          3538 => x"08",
          3539 => x"81",
          3540 => x"52",
          3541 => x"b8",
          3542 => x"d1",
          3543 => x"d1",
          3544 => x"56",
          3545 => x"ff",
          3546 => x"d5",
          3547 => x"88",
          3548 => x"fd",
          3549 => x"ac",
          3550 => x"51",
          3551 => x"3f",
          3552 => x"08",
          3553 => x"ff",
          3554 => x"84",
          3555 => x"ff",
          3556 => x"84",
          3557 => x"74",
          3558 => x"55",
          3559 => x"d1",
          3560 => x"81",
          3561 => x"d1",
          3562 => x"57",
          3563 => x"27",
          3564 => x"84",
          3565 => x"52",
          3566 => x"76",
          3567 => x"34",
          3568 => x"33",
          3569 => x"b3",
          3570 => x"d1",
          3571 => x"81",
          3572 => x"d1",
          3573 => x"57",
          3574 => x"27",
          3575 => x"84",
          3576 => x"52",
          3577 => x"76",
          3578 => x"34",
          3579 => x"33",
          3580 => x"b2",
          3581 => x"d1",
          3582 => x"81",
          3583 => x"d1",
          3584 => x"57",
          3585 => x"26",
          3586 => x"f9",
          3587 => x"d1",
          3588 => x"d1",
          3589 => x"56",
          3590 => x"f9",
          3591 => x"15",
          3592 => x"d1",
          3593 => x"98",
          3594 => x"2c",
          3595 => x"06",
          3596 => x"60",
          3597 => x"ef",
          3598 => x"ac",
          3599 => x"51",
          3600 => x"3f",
          3601 => x"33",
          3602 => x"70",
          3603 => x"d1",
          3604 => x"57",
          3605 => x"77",
          3606 => x"38",
          3607 => x"08",
          3608 => x"ff",
          3609 => x"74",
          3610 => x"29",
          3611 => x"05",
          3612 => x"84",
          3613 => x"5d",
          3614 => x"7b",
          3615 => x"38",
          3616 => x"08",
          3617 => x"ff",
          3618 => x"74",
          3619 => x"29",
          3620 => x"05",
          3621 => x"84",
          3622 => x"5d",
          3623 => x"75",
          3624 => x"38",
          3625 => x"7b",
          3626 => x"18",
          3627 => x"84",
          3628 => x"52",
          3629 => x"ff",
          3630 => x"75",
          3631 => x"29",
          3632 => x"05",
          3633 => x"84",
          3634 => x"5b",
          3635 => x"79",
          3636 => x"38",
          3637 => x"81",
          3638 => x"34",
          3639 => x"08",
          3640 => x"51",
          3641 => x"3f",
          3642 => x"0a",
          3643 => x"0a",
          3644 => x"2c",
          3645 => x"33",
          3646 => x"78",
          3647 => x"a7",
          3648 => x"39",
          3649 => x"33",
          3650 => x"2e",
          3651 => x"84",
          3652 => x"52",
          3653 => x"b0",
          3654 => x"d1",
          3655 => x"05",
          3656 => x"d1",
          3657 => x"81",
          3658 => x"dd",
          3659 => x"88",
          3660 => x"5f",
          3661 => x"84",
          3662 => x"52",
          3663 => x"b0",
          3664 => x"d1",
          3665 => x"51",
          3666 => x"84",
          3667 => x"81",
          3668 => x"77",
          3669 => x"84",
          3670 => x"57",
          3671 => x"80",
          3672 => x"f3",
          3673 => x"10",
          3674 => x"e0",
          3675 => x"57",
          3676 => x"8b",
          3677 => x"82",
          3678 => x"06",
          3679 => x"05",
          3680 => x"53",
          3681 => x"e7",
          3682 => x"b9",
          3683 => x"0c",
          3684 => x"33",
          3685 => x"83",
          3686 => x"70",
          3687 => x"41",
          3688 => x"38",
          3689 => x"08",
          3690 => x"2e",
          3691 => x"f3",
          3692 => x"77",
          3693 => x"bc",
          3694 => x"84",
          3695 => x"80",
          3696 => x"88",
          3697 => x"b9",
          3698 => x"3d",
          3699 => x"d1",
          3700 => x"74",
          3701 => x"38",
          3702 => x"08",
          3703 => x"ff",
          3704 => x"84",
          3705 => x"52",
          3706 => x"af",
          3707 => x"d5",
          3708 => x"88",
          3709 => x"f9",
          3710 => x"8c",
          3711 => x"56",
          3712 => x"8c",
          3713 => x"ff",
          3714 => x"cc",
          3715 => x"f0",
          3716 => x"f7",
          3717 => x"84",
          3718 => x"80",
          3719 => x"88",
          3720 => x"39",
          3721 => x"80",
          3722 => x"34",
          3723 => x"33",
          3724 => x"2e",
          3725 => x"d5",
          3726 => x"88",
          3727 => x"b1",
          3728 => x"ac",
          3729 => x"51",
          3730 => x"3f",
          3731 => x"08",
          3732 => x"ff",
          3733 => x"84",
          3734 => x"ff",
          3735 => x"84",
          3736 => x"7c",
          3737 => x"55",
          3738 => x"83",
          3739 => x"ff",
          3740 => x"80",
          3741 => x"8c",
          3742 => x"84",
          3743 => x"7b",
          3744 => x"0c",
          3745 => x"04",
          3746 => x"33",
          3747 => x"06",
          3748 => x"80",
          3749 => x"38",
          3750 => x"33",
          3751 => x"78",
          3752 => x"34",
          3753 => x"77",
          3754 => x"34",
          3755 => x"08",
          3756 => x"ff",
          3757 => x"84",
          3758 => x"70",
          3759 => x"98",
          3760 => x"88",
          3761 => x"5b",
          3762 => x"24",
          3763 => x"84",
          3764 => x"52",
          3765 => x"ad",
          3766 => x"d1",
          3767 => x"98",
          3768 => x"2c",
          3769 => x"33",
          3770 => x"56",
          3771 => x"f3",
          3772 => x"d5",
          3773 => x"88",
          3774 => x"f5",
          3775 => x"80",
          3776 => x"80",
          3777 => x"98",
          3778 => x"88",
          3779 => x"55",
          3780 => x"f3",
          3781 => x"d5",
          3782 => x"88",
          3783 => x"d1",
          3784 => x"80",
          3785 => x"80",
          3786 => x"98",
          3787 => x"88",
          3788 => x"55",
          3789 => x"ff",
          3790 => x"a5",
          3791 => x"57",
          3792 => x"77",
          3793 => x"ac",
          3794 => x"33",
          3795 => x"a1",
          3796 => x"80",
          3797 => x"80",
          3798 => x"98",
          3799 => x"88",
          3800 => x"5b",
          3801 => x"fe",
          3802 => x"16",
          3803 => x"33",
          3804 => x"d5",
          3805 => x"76",
          3806 => x"ab",
          3807 => x"81",
          3808 => x"81",
          3809 => x"70",
          3810 => x"d1",
          3811 => x"57",
          3812 => x"24",
          3813 => x"fe",
          3814 => x"d1",
          3815 => x"81",
          3816 => x"58",
          3817 => x"f2",
          3818 => x"d1",
          3819 => x"76",
          3820 => x"38",
          3821 => x"70",
          3822 => x"41",
          3823 => x"a1",
          3824 => x"5b",
          3825 => x"1c",
          3826 => x"80",
          3827 => x"ff",
          3828 => x"98",
          3829 => x"8c",
          3830 => x"58",
          3831 => x"e1",
          3832 => x"55",
          3833 => x"8c",
          3834 => x"ff",
          3835 => x"5a",
          3836 => x"7a",
          3837 => x"88",
          3838 => x"60",
          3839 => x"81",
          3840 => x"84",
          3841 => x"75",
          3842 => x"8c",
          3843 => x"80",
          3844 => x"ff",
          3845 => x"98",
          3846 => x"ff",
          3847 => x"5c",
          3848 => x"24",
          3849 => x"77",
          3850 => x"98",
          3851 => x"ff",
          3852 => x"59",
          3853 => x"f1",
          3854 => x"d5",
          3855 => x"88",
          3856 => x"ad",
          3857 => x"80",
          3858 => x"80",
          3859 => x"98",
          3860 => x"88",
          3861 => x"41",
          3862 => x"f1",
          3863 => x"d5",
          3864 => x"88",
          3865 => x"89",
          3866 => x"80",
          3867 => x"80",
          3868 => x"98",
          3869 => x"88",
          3870 => x"41",
          3871 => x"ff",
          3872 => x"dd",
          3873 => x"e0",
          3874 => x"80",
          3875 => x"38",
          3876 => x"ad",
          3877 => x"b9",
          3878 => x"d1",
          3879 => x"b9",
          3880 => x"ff",
          3881 => x"53",
          3882 => x"51",
          3883 => x"3f",
          3884 => x"33",
          3885 => x"33",
          3886 => x"80",
          3887 => x"38",
          3888 => x"08",
          3889 => x"ff",
          3890 => x"84",
          3891 => x"52",
          3892 => x"a9",
          3893 => x"d5",
          3894 => x"88",
          3895 => x"91",
          3896 => x"8c",
          3897 => x"5b",
          3898 => x"8c",
          3899 => x"ff",
          3900 => x"39",
          3901 => x"e1",
          3902 => x"b9",
          3903 => x"f3",
          3904 => x"b9",
          3905 => x"a5",
          3906 => x"f3",
          3907 => x"ef",
          3908 => x"c3",
          3909 => x"ac",
          3910 => x"16",
          3911 => x"58",
          3912 => x"3f",
          3913 => x"0a",
          3914 => x"0a",
          3915 => x"2c",
          3916 => x"33",
          3917 => x"76",
          3918 => x"38",
          3919 => x"33",
          3920 => x"70",
          3921 => x"81",
          3922 => x"58",
          3923 => x"7a",
          3924 => x"38",
          3925 => x"83",
          3926 => x"80",
          3927 => x"38",
          3928 => x"57",
          3929 => x"08",
          3930 => x"38",
          3931 => x"18",
          3932 => x"80",
          3933 => x"80",
          3934 => x"b8",
          3935 => x"b4",
          3936 => x"80",
          3937 => x"38",
          3938 => x"e7",
          3939 => x"f3",
          3940 => x"80",
          3941 => x"80",
          3942 => x"b4",
          3943 => x"b4",
          3944 => x"ee",
          3945 => x"51",
          3946 => x"3f",
          3947 => x"ff",
          3948 => x"58",
          3949 => x"25",
          3950 => x"ff",
          3951 => x"51",
          3952 => x"3f",
          3953 => x"08",
          3954 => x"34",
          3955 => x"08",
          3956 => x"81",
          3957 => x"52",
          3958 => x"ab",
          3959 => x"0b",
          3960 => x"33",
          3961 => x"33",
          3962 => x"74",
          3963 => x"97",
          3964 => x"ac",
          3965 => x"51",
          3966 => x"3f",
          3967 => x"08",
          3968 => x"ff",
          3969 => x"84",
          3970 => x"52",
          3971 => x"a6",
          3972 => x"d1",
          3973 => x"05",
          3974 => x"d1",
          3975 => x"81",
          3976 => x"c7",
          3977 => x"34",
          3978 => x"d1",
          3979 => x"0b",
          3980 => x"34",
          3981 => x"c8",
          3982 => x"0d",
          3983 => x"ff",
          3984 => x"84",
          3985 => x"84",
          3986 => x"84",
          3987 => x"81",
          3988 => x"05",
          3989 => x"7b",
          3990 => x"91",
          3991 => x"70",
          3992 => x"84",
          3993 => x"84",
          3994 => x"58",
          3995 => x"74",
          3996 => x"93",
          3997 => x"ac",
          3998 => x"51",
          3999 => x"3f",
          4000 => x"08",
          4001 => x"ff",
          4002 => x"84",
          4003 => x"52",
          4004 => x"a5",
          4005 => x"d1",
          4006 => x"05",
          4007 => x"d1",
          4008 => x"81",
          4009 => x"c7",
          4010 => x"ff",
          4011 => x"84",
          4012 => x"84",
          4013 => x"84",
          4014 => x"81",
          4015 => x"05",
          4016 => x"7b",
          4017 => x"a5",
          4018 => x"70",
          4019 => x"84",
          4020 => x"84",
          4021 => x"58",
          4022 => x"74",
          4023 => x"a7",
          4024 => x"ac",
          4025 => x"51",
          4026 => x"3f",
          4027 => x"08",
          4028 => x"ff",
          4029 => x"84",
          4030 => x"52",
          4031 => x"a4",
          4032 => x"d1",
          4033 => x"05",
          4034 => x"d1",
          4035 => x"81",
          4036 => x"c7",
          4037 => x"80",
          4038 => x"83",
          4039 => x"70",
          4040 => x"fc",
          4041 => x"e0",
          4042 => x"70",
          4043 => x"56",
          4044 => x"3f",
          4045 => x"08",
          4046 => x"f3",
          4047 => x"10",
          4048 => x"e0",
          4049 => x"57",
          4050 => x"80",
          4051 => x"38",
          4052 => x"52",
          4053 => x"a8",
          4054 => x"f3",
          4055 => x"05",
          4056 => x"06",
          4057 => x"79",
          4058 => x"38",
          4059 => x"b8",
          4060 => x"39",
          4061 => x"f8",
          4062 => x"53",
          4063 => x"51",
          4064 => x"3f",
          4065 => x"08",
          4066 => x"82",
          4067 => x"83",
          4068 => x"51",
          4069 => x"3f",
          4070 => x"d1",
          4071 => x"0b",
          4072 => x"34",
          4073 => x"c8",
          4074 => x"0d",
          4075 => x"77",
          4076 => x"c8",
          4077 => x"c9",
          4078 => x"b9",
          4079 => x"a5",
          4080 => x"c8",
          4081 => x"5c",
          4082 => x"b4",
          4083 => x"f8",
          4084 => x"82",
          4085 => x"84",
          4086 => x"5a",
          4087 => x"08",
          4088 => x"81",
          4089 => x"38",
          4090 => x"08",
          4091 => x"bb",
          4092 => x"c8",
          4093 => x"0b",
          4094 => x"08",
          4095 => x"38",
          4096 => x"08",
          4097 => x"1b",
          4098 => x"77",
          4099 => x"ff",
          4100 => x"b8",
          4101 => x"10",
          4102 => x"05",
          4103 => x"40",
          4104 => x"80",
          4105 => x"82",
          4106 => x"06",
          4107 => x"05",
          4108 => x"53",
          4109 => x"da",
          4110 => x"b9",
          4111 => x"0c",
          4112 => x"33",
          4113 => x"83",
          4114 => x"70",
          4115 => x"41",
          4116 => x"81",
          4117 => x"ff",
          4118 => x"93",
          4119 => x"38",
          4120 => x"ff",
          4121 => x"06",
          4122 => x"77",
          4123 => x"f9",
          4124 => x"53",
          4125 => x"51",
          4126 => x"3f",
          4127 => x"33",
          4128 => x"81",
          4129 => x"57",
          4130 => x"80",
          4131 => x"0b",
          4132 => x"34",
          4133 => x"74",
          4134 => x"f8",
          4135 => x"b8",
          4136 => x"2b",
          4137 => x"83",
          4138 => x"81",
          4139 => x"52",
          4140 => x"d9",
          4141 => x"b9",
          4142 => x"0c",
          4143 => x"33",
          4144 => x"83",
          4145 => x"70",
          4146 => x"41",
          4147 => x"ff",
          4148 => x"9e",
          4149 => x"f3",
          4150 => x"f7",
          4151 => x"f3",
          4152 => x"c0",
          4153 => x"b0",
          4154 => x"8a",
          4155 => x"eb",
          4156 => x"39",
          4157 => x"02",
          4158 => x"33",
          4159 => x"80",
          4160 => x"5b",
          4161 => x"26",
          4162 => x"72",
          4163 => x"8b",
          4164 => x"25",
          4165 => x"72",
          4166 => x"a8",
          4167 => x"a0",
          4168 => x"a7",
          4169 => x"5e",
          4170 => x"9f",
          4171 => x"76",
          4172 => x"75",
          4173 => x"34",
          4174 => x"f9",
          4175 => x"f8",
          4176 => x"f8",
          4177 => x"98",
          4178 => x"2b",
          4179 => x"2b",
          4180 => x"7a",
          4181 => x"56",
          4182 => x"27",
          4183 => x"74",
          4184 => x"56",
          4185 => x"70",
          4186 => x"0c",
          4187 => x"ee",
          4188 => x"27",
          4189 => x"f8",
          4190 => x"98",
          4191 => x"78",
          4192 => x"55",
          4193 => x"e0",
          4194 => x"74",
          4195 => x"56",
          4196 => x"53",
          4197 => x"90",
          4198 => x"86",
          4199 => x"0b",
          4200 => x"33",
          4201 => x"11",
          4202 => x"33",
          4203 => x"11",
          4204 => x"41",
          4205 => x"86",
          4206 => x"0b",
          4207 => x"33",
          4208 => x"06",
          4209 => x"33",
          4210 => x"06",
          4211 => x"22",
          4212 => x"ff",
          4213 => x"29",
          4214 => x"58",
          4215 => x"5d",
          4216 => x"87",
          4217 => x"31",
          4218 => x"79",
          4219 => x"7e",
          4220 => x"7c",
          4221 => x"7a",
          4222 => x"06",
          4223 => x"06",
          4224 => x"14",
          4225 => x"57",
          4226 => x"74",
          4227 => x"83",
          4228 => x"74",
          4229 => x"70",
          4230 => x"59",
          4231 => x"06",
          4232 => x"2e",
          4233 => x"78",
          4234 => x"72",
          4235 => x"c1",
          4236 => x"70",
          4237 => x"34",
          4238 => x"33",
          4239 => x"05",
          4240 => x"39",
          4241 => x"80",
          4242 => x"b0",
          4243 => x"b7",
          4244 => x"81",
          4245 => x"b7",
          4246 => x"81",
          4247 => x"f8",
          4248 => x"74",
          4249 => x"5d",
          4250 => x"5e",
          4251 => x"27",
          4252 => x"73",
          4253 => x"73",
          4254 => x"71",
          4255 => x"5a",
          4256 => x"80",
          4257 => x"38",
          4258 => x"f8",
          4259 => x"0b",
          4260 => x"34",
          4261 => x"33",
          4262 => x"71",
          4263 => x"71",
          4264 => x"71",
          4265 => x"56",
          4266 => x"76",
          4267 => x"ae",
          4268 => x"39",
          4269 => x"38",
          4270 => x"33",
          4271 => x"06",
          4272 => x"11",
          4273 => x"33",
          4274 => x"11",
          4275 => x"80",
          4276 => x"5b",
          4277 => x"86",
          4278 => x"70",
          4279 => x"bc",
          4280 => x"ff",
          4281 => x"bb",
          4282 => x"ff",
          4283 => x"f6",
          4284 => x"ff",
          4285 => x"75",
          4286 => x"5e",
          4287 => x"58",
          4288 => x"57",
          4289 => x"8b",
          4290 => x"31",
          4291 => x"29",
          4292 => x"7d",
          4293 => x"74",
          4294 => x"71",
          4295 => x"83",
          4296 => x"62",
          4297 => x"70",
          4298 => x"5f",
          4299 => x"55",
          4300 => x"85",
          4301 => x"29",
          4302 => x"31",
          4303 => x"06",
          4304 => x"fd",
          4305 => x"83",
          4306 => x"fd",
          4307 => x"f2",
          4308 => x"31",
          4309 => x"fe",
          4310 => x"3d",
          4311 => x"80",
          4312 => x"8a",
          4313 => x"73",
          4314 => x"34",
          4315 => x"87",
          4316 => x"55",
          4317 => x"34",
          4318 => x"34",
          4319 => x"98",
          4320 => x"34",
          4321 => x"87",
          4322 => x"54",
          4323 => x"80",
          4324 => x"80",
          4325 => x"52",
          4326 => x"d8",
          4327 => x"87",
          4328 => x"54",
          4329 => x"56",
          4330 => x"f8",
          4331 => x"84",
          4332 => x"72",
          4333 => x"08",
          4334 => x"06",
          4335 => x"51",
          4336 => x"34",
          4337 => x"cc",
          4338 => x"06",
          4339 => x"53",
          4340 => x"81",
          4341 => x"08",
          4342 => x"88",
          4343 => x"75",
          4344 => x"0b",
          4345 => x"34",
          4346 => x"b9",
          4347 => x"3d",
          4348 => x"b7",
          4349 => x"b9",
          4350 => x"f7",
          4351 => x"af",
          4352 => x"84",
          4353 => x"33",
          4354 => x"33",
          4355 => x"81",
          4356 => x"26",
          4357 => x"84",
          4358 => x"83",
          4359 => x"83",
          4360 => x"72",
          4361 => x"86",
          4362 => x"11",
          4363 => x"22",
          4364 => x"59",
          4365 => x"05",
          4366 => x"ff",
          4367 => x"ce",
          4368 => x"58",
          4369 => x"2e",
          4370 => x"83",
          4371 => x"76",
          4372 => x"83",
          4373 => x"83",
          4374 => x"76",
          4375 => x"ff",
          4376 => x"ff",
          4377 => x"55",
          4378 => x"82",
          4379 => x"19",
          4380 => x"f8",
          4381 => x"f8",
          4382 => x"83",
          4383 => x"84",
          4384 => x"5c",
          4385 => x"74",
          4386 => x"38",
          4387 => x"33",
          4388 => x"54",
          4389 => x"72",
          4390 => x"ac",
          4391 => x"9a",
          4392 => x"55",
          4393 => x"33",
          4394 => x"34",
          4395 => x"05",
          4396 => x"70",
          4397 => x"34",
          4398 => x"84",
          4399 => x"27",
          4400 => x"9f",
          4401 => x"38",
          4402 => x"33",
          4403 => x"15",
          4404 => x"0b",
          4405 => x"34",
          4406 => x"81",
          4407 => x"81",
          4408 => x"9f",
          4409 => x"38",
          4410 => x"33",
          4411 => x"75",
          4412 => x"23",
          4413 => x"81",
          4414 => x"83",
          4415 => x"54",
          4416 => x"26",
          4417 => x"72",
          4418 => x"05",
          4419 => x"33",
          4420 => x"58",
          4421 => x"55",
          4422 => x"80",
          4423 => x"b0",
          4424 => x"ff",
          4425 => x"ff",
          4426 => x"29",
          4427 => x"54",
          4428 => x"27",
          4429 => x"98",
          4430 => x"e0",
          4431 => x"53",
          4432 => x"13",
          4433 => x"81",
          4434 => x"73",
          4435 => x"55",
          4436 => x"81",
          4437 => x"81",
          4438 => x"bc",
          4439 => x"bb",
          4440 => x"29",
          4441 => x"5a",
          4442 => x"26",
          4443 => x"53",
          4444 => x"c8",
          4445 => x"0d",
          4446 => x"f8",
          4447 => x"f8",
          4448 => x"83",
          4449 => x"84",
          4450 => x"5c",
          4451 => x"7a",
          4452 => x"38",
          4453 => x"fe",
          4454 => x"81",
          4455 => x"05",
          4456 => x"33",
          4457 => x"75",
          4458 => x"06",
          4459 => x"73",
          4460 => x"05",
          4461 => x"33",
          4462 => x"78",
          4463 => x"56",
          4464 => x"73",
          4465 => x"ae",
          4466 => x"f4",
          4467 => x"9a",
          4468 => x"31",
          4469 => x"a0",
          4470 => x"16",
          4471 => x"70",
          4472 => x"34",
          4473 => x"72",
          4474 => x"8a",
          4475 => x"e0",
          4476 => x"75",
          4477 => x"05",
          4478 => x"13",
          4479 => x"38",
          4480 => x"80",
          4481 => x"bc",
          4482 => x"fe",
          4483 => x"f8",
          4484 => x"59",
          4485 => x"19",
          4486 => x"84",
          4487 => x"59",
          4488 => x"fc",
          4489 => x"02",
          4490 => x"05",
          4491 => x"70",
          4492 => x"38",
          4493 => x"83",
          4494 => x"51",
          4495 => x"84",
          4496 => x"51",
          4497 => x"86",
          4498 => x"f8",
          4499 => x"0b",
          4500 => x"0c",
          4501 => x"04",
          4502 => x"f8",
          4503 => x"f8",
          4504 => x"81",
          4505 => x"52",
          4506 => x"e2",
          4507 => x"51",
          4508 => x"f8",
          4509 => x"84",
          4510 => x"86",
          4511 => x"83",
          4512 => x"70",
          4513 => x"09",
          4514 => x"72",
          4515 => x"53",
          4516 => x"f8",
          4517 => x"39",
          4518 => x"33",
          4519 => x"b7",
          4520 => x"11",
          4521 => x"70",
          4522 => x"38",
          4523 => x"83",
          4524 => x"80",
          4525 => x"c8",
          4526 => x"0d",
          4527 => x"f9",
          4528 => x"31",
          4529 => x"9f",
          4530 => x"54",
          4531 => x"70",
          4532 => x"34",
          4533 => x"b9",
          4534 => x"3d",
          4535 => x"f8",
          4536 => x"05",
          4537 => x"33",
          4538 => x"55",
          4539 => x"25",
          4540 => x"53",
          4541 => x"f9",
          4542 => x"84",
          4543 => x"86",
          4544 => x"80",
          4545 => x"f9",
          4546 => x"f8",
          4547 => x"bb",
          4548 => x"56",
          4549 => x"25",
          4550 => x"81",
          4551 => x"83",
          4552 => x"fe",
          4553 => x"3d",
          4554 => x"05",
          4555 => x"b1",
          4556 => x"70",
          4557 => x"c4",
          4558 => x"70",
          4559 => x"f8",
          4560 => x"80",
          4561 => x"84",
          4562 => x"06",
          4563 => x"2a",
          4564 => x"53",
          4565 => x"f0",
          4566 => x"06",
          4567 => x"f2",
          4568 => x"f4",
          4569 => x"84",
          4570 => x"83",
          4571 => x"83",
          4572 => x"81",
          4573 => x"07",
          4574 => x"f8",
          4575 => x"0b",
          4576 => x"0c",
          4577 => x"04",
          4578 => x"33",
          4579 => x"51",
          4580 => x"f4",
          4581 => x"83",
          4582 => x"81",
          4583 => x"07",
          4584 => x"f8",
          4585 => x"39",
          4586 => x"83",
          4587 => x"80",
          4588 => x"c8",
          4589 => x"0d",
          4590 => x"f4",
          4591 => x"06",
          4592 => x"70",
          4593 => x"34",
          4594 => x"83",
          4595 => x"87",
          4596 => x"83",
          4597 => x"ff",
          4598 => x"f8",
          4599 => x"fd",
          4600 => x"51",
          4601 => x"f4",
          4602 => x"39",
          4603 => x"33",
          4604 => x"83",
          4605 => x"83",
          4606 => x"ff",
          4607 => x"f8",
          4608 => x"f9",
          4609 => x"51",
          4610 => x"f4",
          4611 => x"39",
          4612 => x"33",
          4613 => x"51",
          4614 => x"f4",
          4615 => x"39",
          4616 => x"33",
          4617 => x"80",
          4618 => x"70",
          4619 => x"34",
          4620 => x"83",
          4621 => x"81",
          4622 => x"07",
          4623 => x"f8",
          4624 => x"ba",
          4625 => x"f4",
          4626 => x"06",
          4627 => x"51",
          4628 => x"f4",
          4629 => x"39",
          4630 => x"33",
          4631 => x"80",
          4632 => x"70",
          4633 => x"34",
          4634 => x"83",
          4635 => x"81",
          4636 => x"07",
          4637 => x"f8",
          4638 => x"82",
          4639 => x"f4",
          4640 => x"06",
          4641 => x"f8",
          4642 => x"f2",
          4643 => x"f4",
          4644 => x"06",
          4645 => x"70",
          4646 => x"34",
          4647 => x"f3",
          4648 => x"bf",
          4649 => x"84",
          4650 => x"05",
          4651 => x"f8",
          4652 => x"f7",
          4653 => x"f9",
          4654 => x"be",
          4655 => x"5f",
          4656 => x"78",
          4657 => x"a1",
          4658 => x"24",
          4659 => x"81",
          4660 => x"38",
          4661 => x"be",
          4662 => x"84",
          4663 => x"7a",
          4664 => x"34",
          4665 => x"f6",
          4666 => x"f8",
          4667 => x"3d",
          4668 => x"83",
          4669 => x"06",
          4670 => x"0b",
          4671 => x"34",
          4672 => x"b7",
          4673 => x"0b",
          4674 => x"34",
          4675 => x"f8",
          4676 => x"0b",
          4677 => x"23",
          4678 => x"b7",
          4679 => x"84",
          4680 => x"56",
          4681 => x"33",
          4682 => x"7c",
          4683 => x"83",
          4684 => x"ff",
          4685 => x"7d",
          4686 => x"34",
          4687 => x"b7",
          4688 => x"83",
          4689 => x"7b",
          4690 => x"23",
          4691 => x"f9",
          4692 => x"0d",
          4693 => x"84",
          4694 => x"81",
          4695 => x"c0",
          4696 => x"83",
          4697 => x"a8",
          4698 => x"f9",
          4699 => x"83",
          4700 => x"84",
          4701 => x"58",
          4702 => x"33",
          4703 => x"c9",
          4704 => x"55",
          4705 => x"53",
          4706 => x"e3",
          4707 => x"80",
          4708 => x"0b",
          4709 => x"33",
          4710 => x"79",
          4711 => x"79",
          4712 => x"9c",
          4713 => x"53",
          4714 => x"f0",
          4715 => x"db",
          4716 => x"70",
          4717 => x"84",
          4718 => x"52",
          4719 => x"7a",
          4720 => x"83",
          4721 => x"ff",
          4722 => x"7d",
          4723 => x"34",
          4724 => x"b7",
          4725 => x"83",
          4726 => x"7b",
          4727 => x"23",
          4728 => x"f9",
          4729 => x"0d",
          4730 => x"84",
          4731 => x"81",
          4732 => x"c0",
          4733 => x"83",
          4734 => x"a8",
          4735 => x"f9",
          4736 => x"83",
          4737 => x"83",
          4738 => x"ff",
          4739 => x"84",
          4740 => x"52",
          4741 => x"51",
          4742 => x"3f",
          4743 => x"f7",
          4744 => x"92",
          4745 => x"84",
          4746 => x"27",
          4747 => x"83",
          4748 => x"33",
          4749 => x"fc",
          4750 => x"cf",
          4751 => x"70",
          4752 => x"5a",
          4753 => x"f9",
          4754 => x"02",
          4755 => x"05",
          4756 => x"bc",
          4757 => x"f9",
          4758 => x"f8",
          4759 => x"29",
          4760 => x"a0",
          4761 => x"f8",
          4762 => x"51",
          4763 => x"7c",
          4764 => x"83",
          4765 => x"83",
          4766 => x"52",
          4767 => x"57",
          4768 => x"2e",
          4769 => x"75",
          4770 => x"f9",
          4771 => x"24",
          4772 => x"75",
          4773 => x"85",
          4774 => x"2e",
          4775 => x"84",
          4776 => x"83",
          4777 => x"83",
          4778 => x"72",
          4779 => x"55",
          4780 => x"b7",
          4781 => x"86",
          4782 => x"14",
          4783 => x"bc",
          4784 => x"f9",
          4785 => x"f6",
          4786 => x"29",
          4787 => x"56",
          4788 => x"f8",
          4789 => x"83",
          4790 => x"73",
          4791 => x"58",
          4792 => x"f4",
          4793 => x"b0",
          4794 => x"84",
          4795 => x"70",
          4796 => x"83",
          4797 => x"83",
          4798 => x"72",
          4799 => x"57",
          4800 => x"57",
          4801 => x"33",
          4802 => x"14",
          4803 => x"70",
          4804 => x"59",
          4805 => x"26",
          4806 => x"84",
          4807 => x"58",
          4808 => x"38",
          4809 => x"72",
          4810 => x"34",
          4811 => x"33",
          4812 => x"2e",
          4813 => x"b7",
          4814 => x"76",
          4815 => x"fb",
          4816 => x"84",
          4817 => x"89",
          4818 => x"75",
          4819 => x"38",
          4820 => x"80",
          4821 => x"8a",
          4822 => x"06",
          4823 => x"81",
          4824 => x"f1",
          4825 => x"0b",
          4826 => x"34",
          4827 => x"83",
          4828 => x"33",
          4829 => x"c4",
          4830 => x"34",
          4831 => x"09",
          4832 => x"89",
          4833 => x"76",
          4834 => x"fd",
          4835 => x"13",
          4836 => x"06",
          4837 => x"83",
          4838 => x"38",
          4839 => x"51",
          4840 => x"81",
          4841 => x"ff",
          4842 => x"83",
          4843 => x"38",
          4844 => x"74",
          4845 => x"34",
          4846 => x"75",
          4847 => x"f9",
          4848 => x"0b",
          4849 => x"0c",
          4850 => x"04",
          4851 => x"2e",
          4852 => x"fd",
          4853 => x"f8",
          4854 => x"81",
          4855 => x"ff",
          4856 => x"83",
          4857 => x"72",
          4858 => x"34",
          4859 => x"51",
          4860 => x"83",
          4861 => x"70",
          4862 => x"55",
          4863 => x"73",
          4864 => x"73",
          4865 => x"f8",
          4866 => x"a0",
          4867 => x"83",
          4868 => x"81",
          4869 => x"ef",
          4870 => x"90",
          4871 => x"75",
          4872 => x"3f",
          4873 => x"e6",
          4874 => x"80",
          4875 => x"84",
          4876 => x"57",
          4877 => x"2e",
          4878 => x"75",
          4879 => x"82",
          4880 => x"2e",
          4881 => x"78",
          4882 => x"d1",
          4883 => x"2e",
          4884 => x"78",
          4885 => x"8f",
          4886 => x"bc",
          4887 => x"f8",
          4888 => x"f9",
          4889 => x"29",
          4890 => x"5c",
          4891 => x"19",
          4892 => x"a0",
          4893 => x"84",
          4894 => x"83",
          4895 => x"83",
          4896 => x"72",
          4897 => x"5a",
          4898 => x"78",
          4899 => x"18",
          4900 => x"f8",
          4901 => x"29",
          4902 => x"5a",
          4903 => x"33",
          4904 => x"b0",
          4905 => x"84",
          4906 => x"70",
          4907 => x"83",
          4908 => x"83",
          4909 => x"72",
          4910 => x"42",
          4911 => x"59",
          4912 => x"33",
          4913 => x"1f",
          4914 => x"70",
          4915 => x"42",
          4916 => x"26",
          4917 => x"84",
          4918 => x"5a",
          4919 => x"38",
          4920 => x"75",
          4921 => x"34",
          4922 => x"b9",
          4923 => x"3d",
          4924 => x"b7",
          4925 => x"38",
          4926 => x"81",
          4927 => x"b8",
          4928 => x"38",
          4929 => x"2e",
          4930 => x"80",
          4931 => x"c4",
          4932 => x"bc",
          4933 => x"f8",
          4934 => x"f9",
          4935 => x"29",
          4936 => x"40",
          4937 => x"19",
          4938 => x"a0",
          4939 => x"84",
          4940 => x"83",
          4941 => x"83",
          4942 => x"72",
          4943 => x"41",
          4944 => x"78",
          4945 => x"1f",
          4946 => x"f8",
          4947 => x"29",
          4948 => x"83",
          4949 => x"86",
          4950 => x"1b",
          4951 => x"bc",
          4952 => x"ff",
          4953 => x"f6",
          4954 => x"f9",
          4955 => x"29",
          4956 => x"43",
          4957 => x"f8",
          4958 => x"84",
          4959 => x"34",
          4960 => x"77",
          4961 => x"41",
          4962 => x"fe",
          4963 => x"83",
          4964 => x"80",
          4965 => x"c8",
          4966 => x"0d",
          4967 => x"2e",
          4968 => x"78",
          4969 => x"81",
          4970 => x"2e",
          4971 => x"fd",
          4972 => x"0b",
          4973 => x"34",
          4974 => x"b9",
          4975 => x"3d",
          4976 => x"9b",
          4977 => x"38",
          4978 => x"75",
          4979 => x"d0",
          4980 => x"c8",
          4981 => x"59",
          4982 => x"b8",
          4983 => x"84",
          4984 => x"34",
          4985 => x"06",
          4986 => x"84",
          4987 => x"34",
          4988 => x"b9",
          4989 => x"3d",
          4990 => x"9b",
          4991 => x"38",
          4992 => x"b8",
          4993 => x"b7",
          4994 => x"f8",
          4995 => x"f8",
          4996 => x"72",
          4997 => x"40",
          4998 => x"c4",
          4999 => x"a7",
          5000 => x"34",
          5001 => x"33",
          5002 => x"33",
          5003 => x"22",
          5004 => x"12",
          5005 => x"56",
          5006 => x"fa",
          5007 => x"f8",
          5008 => x"71",
          5009 => x"57",
          5010 => x"33",
          5011 => x"80",
          5012 => x"b7",
          5013 => x"81",
          5014 => x"f8",
          5015 => x"f8",
          5016 => x"72",
          5017 => x"42",
          5018 => x"83",
          5019 => x"60",
          5020 => x"05",
          5021 => x"58",
          5022 => x"81",
          5023 => x"ea",
          5024 => x"0b",
          5025 => x"34",
          5026 => x"84",
          5027 => x"83",
          5028 => x"70",
          5029 => x"83",
          5030 => x"73",
          5031 => x"86",
          5032 => x"05",
          5033 => x"22",
          5034 => x"72",
          5035 => x"70",
          5036 => x"06",
          5037 => x"33",
          5038 => x"5a",
          5039 => x"2e",
          5040 => x"78",
          5041 => x"ff",
          5042 => x"76",
          5043 => x"76",
          5044 => x"f8",
          5045 => x"90",
          5046 => x"84",
          5047 => x"80",
          5048 => x"c9",
          5049 => x"84",
          5050 => x"80",
          5051 => x"cb",
          5052 => x"84",
          5053 => x"80",
          5054 => x"c8",
          5055 => x"0d",
          5056 => x"f8",
          5057 => x"b0",
          5058 => x"f9",
          5059 => x"b1",
          5060 => x"f7",
          5061 => x"b2",
          5062 => x"84",
          5063 => x"80",
          5064 => x"c8",
          5065 => x"0d",
          5066 => x"ff",
          5067 => x"06",
          5068 => x"83",
          5069 => x"84",
          5070 => x"70",
          5071 => x"83",
          5072 => x"70",
          5073 => x"72",
          5074 => x"86",
          5075 => x"05",
          5076 => x"22",
          5077 => x"7b",
          5078 => x"83",
          5079 => x"83",
          5080 => x"44",
          5081 => x"42",
          5082 => x"81",
          5083 => x"38",
          5084 => x"06",
          5085 => x"56",
          5086 => x"75",
          5087 => x"f8",
          5088 => x"81",
          5089 => x"81",
          5090 => x"81",
          5091 => x"72",
          5092 => x"40",
          5093 => x"e4",
          5094 => x"a0",
          5095 => x"84",
          5096 => x"83",
          5097 => x"83",
          5098 => x"72",
          5099 => x"5a",
          5100 => x"a0",
          5101 => x"fa",
          5102 => x"f8",
          5103 => x"71",
          5104 => x"5a",
          5105 => x"f4",
          5106 => x"b0",
          5107 => x"84",
          5108 => x"70",
          5109 => x"83",
          5110 => x"83",
          5111 => x"72",
          5112 => x"43",
          5113 => x"59",
          5114 => x"33",
          5115 => x"9a",
          5116 => x"1a",
          5117 => x"06",
          5118 => x"7b",
          5119 => x"38",
          5120 => x"33",
          5121 => x"d0",
          5122 => x"58",
          5123 => x"f9",
          5124 => x"f9",
          5125 => x"ff",
          5126 => x"05",
          5127 => x"39",
          5128 => x"95",
          5129 => x"bd",
          5130 => x"38",
          5131 => x"95",
          5132 => x"b8",
          5133 => x"7e",
          5134 => x"ff",
          5135 => x"75",
          5136 => x"c8",
          5137 => x"10",
          5138 => x"05",
          5139 => x"04",
          5140 => x"f8",
          5141 => x"52",
          5142 => x"9f",
          5143 => x"84",
          5144 => x"9c",
          5145 => x"83",
          5146 => x"84",
          5147 => x"70",
          5148 => x"83",
          5149 => x"70",
          5150 => x"72",
          5151 => x"86",
          5152 => x"05",
          5153 => x"22",
          5154 => x"7b",
          5155 => x"83",
          5156 => x"83",
          5157 => x"46",
          5158 => x"59",
          5159 => x"81",
          5160 => x"38",
          5161 => x"81",
          5162 => x"81",
          5163 => x"81",
          5164 => x"72",
          5165 => x"58",
          5166 => x"e4",
          5167 => x"a0",
          5168 => x"84",
          5169 => x"83",
          5170 => x"83",
          5171 => x"72",
          5172 => x"5e",
          5173 => x"a0",
          5174 => x"fa",
          5175 => x"f8",
          5176 => x"71",
          5177 => x"5e",
          5178 => x"33",
          5179 => x"80",
          5180 => x"b7",
          5181 => x"81",
          5182 => x"f8",
          5183 => x"f8",
          5184 => x"72",
          5185 => x"44",
          5186 => x"83",
          5187 => x"84",
          5188 => x"34",
          5189 => x"70",
          5190 => x"5b",
          5191 => x"26",
          5192 => x"84",
          5193 => x"58",
          5194 => x"38",
          5195 => x"75",
          5196 => x"34",
          5197 => x"81",
          5198 => x"59",
          5199 => x"f7",
          5200 => x"f8",
          5201 => x"b7",
          5202 => x"f8",
          5203 => x"81",
          5204 => x"81",
          5205 => x"81",
          5206 => x"72",
          5207 => x"5b",
          5208 => x"5b",
          5209 => x"33",
          5210 => x"80",
          5211 => x"b7",
          5212 => x"f8",
          5213 => x"f8",
          5214 => x"71",
          5215 => x"41",
          5216 => x"0b",
          5217 => x"1c",
          5218 => x"f8",
          5219 => x"29",
          5220 => x"83",
          5221 => x"86",
          5222 => x"1a",
          5223 => x"bc",
          5224 => x"ff",
          5225 => x"f6",
          5226 => x"f9",
          5227 => x"29",
          5228 => x"5a",
          5229 => x"f8",
          5230 => x"98",
          5231 => x"60",
          5232 => x"81",
          5233 => x"58",
          5234 => x"fe",
          5235 => x"83",
          5236 => x"fe",
          5237 => x"0b",
          5238 => x"0c",
          5239 => x"b9",
          5240 => x"3d",
          5241 => x"f8",
          5242 => x"59",
          5243 => x"19",
          5244 => x"83",
          5245 => x"70",
          5246 => x"58",
          5247 => x"f9",
          5248 => x"0b",
          5249 => x"34",
          5250 => x"b9",
          5251 => x"3d",
          5252 => x"f8",
          5253 => x"5b",
          5254 => x"1b",
          5255 => x"83",
          5256 => x"84",
          5257 => x"83",
          5258 => x"5b",
          5259 => x"5c",
          5260 => x"84",
          5261 => x"9c",
          5262 => x"53",
          5263 => x"ff",
          5264 => x"84",
          5265 => x"80",
          5266 => x"38",
          5267 => x"33",
          5268 => x"5a",
          5269 => x"c9",
          5270 => x"83",
          5271 => x"02",
          5272 => x"22",
          5273 => x"9c",
          5274 => x"cf",
          5275 => x"fa",
          5276 => x"84",
          5277 => x"33",
          5278 => x"f8",
          5279 => x"b7",
          5280 => x"f8",
          5281 => x"5b",
          5282 => x"39",
          5283 => x"33",
          5284 => x"33",
          5285 => x"33",
          5286 => x"05",
          5287 => x"84",
          5288 => x"33",
          5289 => x"a0",
          5290 => x"84",
          5291 => x"83",
          5292 => x"83",
          5293 => x"72",
          5294 => x"5a",
          5295 => x"78",
          5296 => x"18",
          5297 => x"f8",
          5298 => x"29",
          5299 => x"83",
          5300 => x"60",
          5301 => x"80",
          5302 => x"b7",
          5303 => x"81",
          5304 => x"f8",
          5305 => x"f8",
          5306 => x"72",
          5307 => x"5f",
          5308 => x"83",
          5309 => x"84",
          5310 => x"34",
          5311 => x"81",
          5312 => x"58",
          5313 => x"90",
          5314 => x"b7",
          5315 => x"77",
          5316 => x"ff",
          5317 => x"83",
          5318 => x"80",
          5319 => x"c4",
          5320 => x"bf",
          5321 => x"80",
          5322 => x"38",
          5323 => x"33",
          5324 => x"b4",
          5325 => x"81",
          5326 => x"3f",
          5327 => x"b9",
          5328 => x"3d",
          5329 => x"b9",
          5330 => x"f8",
          5331 => x"b9",
          5332 => x"f8",
          5333 => x"b9",
          5334 => x"76",
          5335 => x"23",
          5336 => x"83",
          5337 => x"84",
          5338 => x"83",
          5339 => x"84",
          5340 => x"83",
          5341 => x"84",
          5342 => x"ff",
          5343 => x"b8",
          5344 => x"7a",
          5345 => x"93",
          5346 => x"9c",
          5347 => x"86",
          5348 => x"06",
          5349 => x"83",
          5350 => x"81",
          5351 => x"f8",
          5352 => x"05",
          5353 => x"83",
          5354 => x"94",
          5355 => x"57",
          5356 => x"3f",
          5357 => x"fe",
          5358 => x"b9",
          5359 => x"ff",
          5360 => x"cc",
          5361 => x"05",
          5362 => x"24",
          5363 => x"76",
          5364 => x"ac",
          5365 => x"bd",
          5366 => x"39",
          5367 => x"b8",
          5368 => x"58",
          5369 => x"06",
          5370 => x"27",
          5371 => x"77",
          5372 => x"9c",
          5373 => x"33",
          5374 => x"b1",
          5375 => x"38",
          5376 => x"83",
          5377 => x"5f",
          5378 => x"84",
          5379 => x"5e",
          5380 => x"8f",
          5381 => x"f8",
          5382 => x"b9",
          5383 => x"71",
          5384 => x"70",
          5385 => x"06",
          5386 => x"5e",
          5387 => x"f8",
          5388 => x"e7",
          5389 => x"c9",
          5390 => x"80",
          5391 => x"38",
          5392 => x"33",
          5393 => x"81",
          5394 => x"b7",
          5395 => x"57",
          5396 => x"27",
          5397 => x"75",
          5398 => x"34",
          5399 => x"80",
          5400 => x"f9",
          5401 => x"f8",
          5402 => x"ff",
          5403 => x"7b",
          5404 => x"a7",
          5405 => x"56",
          5406 => x"f8",
          5407 => x"39",
          5408 => x"f8",
          5409 => x"f8",
          5410 => x"b7",
          5411 => x"05",
          5412 => x"76",
          5413 => x"38",
          5414 => x"75",
          5415 => x"34",
          5416 => x"84",
          5417 => x"40",
          5418 => x"8d",
          5419 => x"f8",
          5420 => x"b9",
          5421 => x"71",
          5422 => x"70",
          5423 => x"06",
          5424 => x"42",
          5425 => x"f8",
          5426 => x"cf",
          5427 => x"c9",
          5428 => x"80",
          5429 => x"38",
          5430 => x"22",
          5431 => x"2e",
          5432 => x"fc",
          5433 => x"b7",
          5434 => x"f8",
          5435 => x"f8",
          5436 => x"71",
          5437 => x"a7",
          5438 => x"83",
          5439 => x"43",
          5440 => x"71",
          5441 => x"70",
          5442 => x"06",
          5443 => x"08",
          5444 => x"80",
          5445 => x"5d",
          5446 => x"82",
          5447 => x"bf",
          5448 => x"83",
          5449 => x"fb",
          5450 => x"b8",
          5451 => x"79",
          5452 => x"e7",
          5453 => x"9c",
          5454 => x"99",
          5455 => x"06",
          5456 => x"81",
          5457 => x"cd",
          5458 => x"39",
          5459 => x"33",
          5460 => x"2e",
          5461 => x"84",
          5462 => x"83",
          5463 => x"5d",
          5464 => x"b7",
          5465 => x"11",
          5466 => x"75",
          5467 => x"38",
          5468 => x"83",
          5469 => x"fb",
          5470 => x"b8",
          5471 => x"76",
          5472 => x"c8",
          5473 => x"9d",
          5474 => x"f8",
          5475 => x"05",
          5476 => x"33",
          5477 => x"41",
          5478 => x"25",
          5479 => x"57",
          5480 => x"f8",
          5481 => x"39",
          5482 => x"51",
          5483 => x"3f",
          5484 => x"b8",
          5485 => x"57",
          5486 => x"8b",
          5487 => x"10",
          5488 => x"05",
          5489 => x"5a",
          5490 => x"51",
          5491 => x"3f",
          5492 => x"81",
          5493 => x"b8",
          5494 => x"58",
          5495 => x"82",
          5496 => x"c9",
          5497 => x"7d",
          5498 => x"38",
          5499 => x"22",
          5500 => x"26",
          5501 => x"57",
          5502 => x"81",
          5503 => x"d5",
          5504 => x"97",
          5505 => x"c9",
          5506 => x"77",
          5507 => x"38",
          5508 => x"33",
          5509 => x"81",
          5510 => x"b9",
          5511 => x"05",
          5512 => x"06",
          5513 => x"33",
          5514 => x"06",
          5515 => x"43",
          5516 => x"5c",
          5517 => x"27",
          5518 => x"5a",
          5519 => x"f6",
          5520 => x"ff",
          5521 => x"58",
          5522 => x"27",
          5523 => x"57",
          5524 => x"f8",
          5525 => x"bc",
          5526 => x"57",
          5527 => x"27",
          5528 => x"7a",
          5529 => x"f8",
          5530 => x"af",
          5531 => x"c9",
          5532 => x"80",
          5533 => x"38",
          5534 => x"33",
          5535 => x"33",
          5536 => x"7f",
          5537 => x"38",
          5538 => x"33",
          5539 => x"33",
          5540 => x"06",
          5541 => x"33",
          5542 => x"11",
          5543 => x"80",
          5544 => x"f6",
          5545 => x"71",
          5546 => x"70",
          5547 => x"06",
          5548 => x"33",
          5549 => x"59",
          5550 => x"81",
          5551 => x"38",
          5552 => x"ff",
          5553 => x"31",
          5554 => x"7c",
          5555 => x"38",
          5556 => x"33",
          5557 => x"27",
          5558 => x"ff",
          5559 => x"83",
          5560 => x"7c",
          5561 => x"70",
          5562 => x"57",
          5563 => x"8e",
          5564 => x"b7",
          5565 => x"76",
          5566 => x"ee",
          5567 => x"56",
          5568 => x"f8",
          5569 => x"ff",
          5570 => x"f6",
          5571 => x"80",
          5572 => x"26",
          5573 => x"77",
          5574 => x"7e",
          5575 => x"71",
          5576 => x"5e",
          5577 => x"86",
          5578 => x"5b",
          5579 => x"80",
          5580 => x"06",
          5581 => x"06",
          5582 => x"1d",
          5583 => x"5c",
          5584 => x"f7",
          5585 => x"98",
          5586 => x"e0",
          5587 => x"5f",
          5588 => x"1f",
          5589 => x"81",
          5590 => x"76",
          5591 => x"58",
          5592 => x"81",
          5593 => x"81",
          5594 => x"bc",
          5595 => x"bb",
          5596 => x"29",
          5597 => x"5e",
          5598 => x"27",
          5599 => x"e0",
          5600 => x"5f",
          5601 => x"1f",
          5602 => x"81",
          5603 => x"76",
          5604 => x"58",
          5605 => x"81",
          5606 => x"81",
          5607 => x"bc",
          5608 => x"bb",
          5609 => x"29",
          5610 => x"5e",
          5611 => x"26",
          5612 => x"f6",
          5613 => x"b8",
          5614 => x"75",
          5615 => x"e0",
          5616 => x"84",
          5617 => x"51",
          5618 => x"f6",
          5619 => x"0b",
          5620 => x"33",
          5621 => x"b8",
          5622 => x"59",
          5623 => x"78",
          5624 => x"84",
          5625 => x"56",
          5626 => x"09",
          5627 => x"be",
          5628 => x"f9",
          5629 => x"81",
          5630 => x"f8",
          5631 => x"43",
          5632 => x"ff",
          5633 => x"38",
          5634 => x"33",
          5635 => x"26",
          5636 => x"7e",
          5637 => x"56",
          5638 => x"f5",
          5639 => x"76",
          5640 => x"27",
          5641 => x"f5",
          5642 => x"10",
          5643 => x"90",
          5644 => x"86",
          5645 => x"11",
          5646 => x"5a",
          5647 => x"80",
          5648 => x"06",
          5649 => x"75",
          5650 => x"79",
          5651 => x"76",
          5652 => x"83",
          5653 => x"70",
          5654 => x"90",
          5655 => x"88",
          5656 => x"07",
          5657 => x"52",
          5658 => x"7a",
          5659 => x"80",
          5660 => x"05",
          5661 => x"76",
          5662 => x"58",
          5663 => x"26",
          5664 => x"b7",
          5665 => x"b7",
          5666 => x"5f",
          5667 => x"06",
          5668 => x"06",
          5669 => x"22",
          5670 => x"64",
          5671 => x"59",
          5672 => x"26",
          5673 => x"78",
          5674 => x"7b",
          5675 => x"57",
          5676 => x"1d",
          5677 => x"76",
          5678 => x"38",
          5679 => x"33",
          5680 => x"18",
          5681 => x"0b",
          5682 => x"34",
          5683 => x"81",
          5684 => x"81",
          5685 => x"76",
          5686 => x"38",
          5687 => x"e0",
          5688 => x"78",
          5689 => x"5a",
          5690 => x"57",
          5691 => x"d6",
          5692 => x"39",
          5693 => x"81",
          5694 => x"58",
          5695 => x"83",
          5696 => x"70",
          5697 => x"71",
          5698 => x"f0",
          5699 => x"2a",
          5700 => x"57",
          5701 => x"2e",
          5702 => x"be",
          5703 => x"0b",
          5704 => x"34",
          5705 => x"81",
          5706 => x"56",
          5707 => x"83",
          5708 => x"33",
          5709 => x"c4",
          5710 => x"34",
          5711 => x"33",
          5712 => x"33",
          5713 => x"22",
          5714 => x"33",
          5715 => x"5d",
          5716 => x"83",
          5717 => x"87",
          5718 => x"83",
          5719 => x"81",
          5720 => x"ff",
          5721 => x"f4",
          5722 => x"f8",
          5723 => x"fd",
          5724 => x"56",
          5725 => x"f4",
          5726 => x"83",
          5727 => x"81",
          5728 => x"07",
          5729 => x"f8",
          5730 => x"39",
          5731 => x"33",
          5732 => x"81",
          5733 => x"83",
          5734 => x"c3",
          5735 => x"f4",
          5736 => x"06",
          5737 => x"75",
          5738 => x"34",
          5739 => x"80",
          5740 => x"f8",
          5741 => x"18",
          5742 => x"06",
          5743 => x"a4",
          5744 => x"f4",
          5745 => x"06",
          5746 => x"f8",
          5747 => x"8f",
          5748 => x"f4",
          5749 => x"06",
          5750 => x"75",
          5751 => x"34",
          5752 => x"83",
          5753 => x"81",
          5754 => x"e0",
          5755 => x"83",
          5756 => x"fe",
          5757 => x"f8",
          5758 => x"cf",
          5759 => x"07",
          5760 => x"f8",
          5761 => x"d7",
          5762 => x"f4",
          5763 => x"06",
          5764 => x"75",
          5765 => x"34",
          5766 => x"83",
          5767 => x"81",
          5768 => x"07",
          5769 => x"f8",
          5770 => x"b3",
          5771 => x"f4",
          5772 => x"06",
          5773 => x"75",
          5774 => x"34",
          5775 => x"83",
          5776 => x"81",
          5777 => x"07",
          5778 => x"f8",
          5779 => x"8f",
          5780 => x"f4",
          5781 => x"06",
          5782 => x"f8",
          5783 => x"ff",
          5784 => x"f4",
          5785 => x"07",
          5786 => x"f8",
          5787 => x"ef",
          5788 => x"f4",
          5789 => x"07",
          5790 => x"f8",
          5791 => x"df",
          5792 => x"f4",
          5793 => x"06",
          5794 => x"56",
          5795 => x"f4",
          5796 => x"39",
          5797 => x"33",
          5798 => x"b0",
          5799 => x"83",
          5800 => x"fd",
          5801 => x"0b",
          5802 => x"34",
          5803 => x"51",
          5804 => x"ec",
          5805 => x"b9",
          5806 => x"f8",
          5807 => x"b9",
          5808 => x"f8",
          5809 => x"b9",
          5810 => x"78",
          5811 => x"23",
          5812 => x"b8",
          5813 => x"c7",
          5814 => x"84",
          5815 => x"80",
          5816 => x"c8",
          5817 => x"0d",
          5818 => x"f8",
          5819 => x"f8",
          5820 => x"81",
          5821 => x"ff",
          5822 => x"cf",
          5823 => x"cc",
          5824 => x"dc",
          5825 => x"05",
          5826 => x"fd",
          5827 => x"c8",
          5828 => x"84",
          5829 => x"84",
          5830 => x"80",
          5831 => x"c8",
          5832 => x"84",
          5833 => x"9c",
          5834 => x"77",
          5835 => x"34",
          5836 => x"84",
          5837 => x"81",
          5838 => x"7a",
          5839 => x"34",
          5840 => x"fe",
          5841 => x"80",
          5842 => x"84",
          5843 => x"23",
          5844 => x"b8",
          5845 => x"39",
          5846 => x"f8",
          5847 => x"52",
          5848 => x"97",
          5849 => x"f9",
          5850 => x"ff",
          5851 => x"05",
          5852 => x"39",
          5853 => x"f8",
          5854 => x"52",
          5855 => x"fb",
          5856 => x"39",
          5857 => x"eb",
          5858 => x"8f",
          5859 => x"f9",
          5860 => x"70",
          5861 => x"2c",
          5862 => x"5f",
          5863 => x"39",
          5864 => x"51",
          5865 => x"b7",
          5866 => x"75",
          5867 => x"eb",
          5868 => x"f8",
          5869 => x"e3",
          5870 => x"f8",
          5871 => x"70",
          5872 => x"2c",
          5873 => x"40",
          5874 => x"39",
          5875 => x"33",
          5876 => x"b7",
          5877 => x"11",
          5878 => x"75",
          5879 => x"c0",
          5880 => x"f3",
          5881 => x"b7",
          5882 => x"81",
          5883 => x"5c",
          5884 => x"ee",
          5885 => x"f8",
          5886 => x"b7",
          5887 => x"81",
          5888 => x"f8",
          5889 => x"74",
          5890 => x"a7",
          5891 => x"83",
          5892 => x"5f",
          5893 => x"29",
          5894 => x"ff",
          5895 => x"f7",
          5896 => x"5b",
          5897 => x"5d",
          5898 => x"81",
          5899 => x"83",
          5900 => x"ff",
          5901 => x"80",
          5902 => x"89",
          5903 => x"bb",
          5904 => x"76",
          5905 => x"38",
          5906 => x"75",
          5907 => x"23",
          5908 => x"06",
          5909 => x"57",
          5910 => x"83",
          5911 => x"b7",
          5912 => x"76",
          5913 => x"ec",
          5914 => x"56",
          5915 => x"f8",
          5916 => x"ff",
          5917 => x"f6",
          5918 => x"80",
          5919 => x"26",
          5920 => x"77",
          5921 => x"7e",
          5922 => x"71",
          5923 => x"5e",
          5924 => x"86",
          5925 => x"5b",
          5926 => x"80",
          5927 => x"06",
          5928 => x"06",
          5929 => x"1d",
          5930 => x"5d",
          5931 => x"ec",
          5932 => x"98",
          5933 => x"e0",
          5934 => x"5e",
          5935 => x"1e",
          5936 => x"81",
          5937 => x"76",
          5938 => x"58",
          5939 => x"81",
          5940 => x"81",
          5941 => x"bc",
          5942 => x"bb",
          5943 => x"29",
          5944 => x"5d",
          5945 => x"27",
          5946 => x"e0",
          5947 => x"5e",
          5948 => x"1e",
          5949 => x"81",
          5950 => x"76",
          5951 => x"58",
          5952 => x"81",
          5953 => x"81",
          5954 => x"bc",
          5955 => x"bb",
          5956 => x"29",
          5957 => x"5d",
          5958 => x"26",
          5959 => x"eb",
          5960 => x"f8",
          5961 => x"5c",
          5962 => x"1c",
          5963 => x"83",
          5964 => x"84",
          5965 => x"83",
          5966 => x"84",
          5967 => x"5f",
          5968 => x"fd",
          5969 => x"eb",
          5970 => x"b7",
          5971 => x"81",
          5972 => x"11",
          5973 => x"76",
          5974 => x"38",
          5975 => x"83",
          5976 => x"77",
          5977 => x"ff",
          5978 => x"80",
          5979 => x"38",
          5980 => x"83",
          5981 => x"84",
          5982 => x"70",
          5983 => x"ff",
          5984 => x"56",
          5985 => x"eb",
          5986 => x"56",
          5987 => x"f9",
          5988 => x"39",
          5989 => x"33",
          5990 => x"b7",
          5991 => x"11",
          5992 => x"75",
          5993 => x"ca",
          5994 => x"ef",
          5995 => x"81",
          5996 => x"06",
          5997 => x"83",
          5998 => x"70",
          5999 => x"83",
          6000 => x"7a",
          6001 => x"57",
          6002 => x"09",
          6003 => x"b8",
          6004 => x"39",
          6005 => x"75",
          6006 => x"34",
          6007 => x"ff",
          6008 => x"83",
          6009 => x"fc",
          6010 => x"7b",
          6011 => x"83",
          6012 => x"f2",
          6013 => x"7d",
          6014 => x"7a",
          6015 => x"38",
          6016 => x"81",
          6017 => x"83",
          6018 => x"77",
          6019 => x"59",
          6020 => x"26",
          6021 => x"80",
          6022 => x"05",
          6023 => x"f8",
          6024 => x"70",
          6025 => x"34",
          6026 => x"d4",
          6027 => x"39",
          6028 => x"56",
          6029 => x"f6",
          6030 => x"39",
          6031 => x"f8",
          6032 => x"ad",
          6033 => x"f8",
          6034 => x"84",
          6035 => x"83",
          6036 => x"f1",
          6037 => x"0b",
          6038 => x"34",
          6039 => x"83",
          6040 => x"33",
          6041 => x"c4",
          6042 => x"34",
          6043 => x"f7",
          6044 => x"a7",
          6045 => x"0d",
          6046 => x"33",
          6047 => x"33",
          6048 => x"80",
          6049 => x"73",
          6050 => x"3f",
          6051 => x"b9",
          6052 => x"3d",
          6053 => x"52",
          6054 => x"ab",
          6055 => x"84",
          6056 => x"85",
          6057 => x"f3",
          6058 => x"bf",
          6059 => x"ff",
          6060 => x"cc",
          6061 => x"ff",
          6062 => x"ac",
          6063 => x"55",
          6064 => x"80",
          6065 => x"38",
          6066 => x"75",
          6067 => x"34",
          6068 => x"84",
          6069 => x"8f",
          6070 => x"83",
          6071 => x"54",
          6072 => x"80",
          6073 => x"73",
          6074 => x"30",
          6075 => x"09",
          6076 => x"56",
          6077 => x"72",
          6078 => x"0c",
          6079 => x"54",
          6080 => x"09",
          6081 => x"38",
          6082 => x"83",
          6083 => x"70",
          6084 => x"07",
          6085 => x"79",
          6086 => x"c4",
          6087 => x"bc",
          6088 => x"f9",
          6089 => x"f8",
          6090 => x"29",
          6091 => x"a0",
          6092 => x"f8",
          6093 => x"59",
          6094 => x"29",
          6095 => x"ff",
          6096 => x"f7",
          6097 => x"59",
          6098 => x"81",
          6099 => x"38",
          6100 => x"73",
          6101 => x"80",
          6102 => x"87",
          6103 => x"0c",
          6104 => x"88",
          6105 => x"80",
          6106 => x"87",
          6107 => x"08",
          6108 => x"f4",
          6109 => x"81",
          6110 => x"ff",
          6111 => x"81",
          6112 => x"cf",
          6113 => x"83",
          6114 => x"33",
          6115 => x"06",
          6116 => x"16",
          6117 => x"55",
          6118 => x"85",
          6119 => x"81",
          6120 => x"b4",
          6121 => x"f6",
          6122 => x"75",
          6123 => x"5a",
          6124 => x"2e",
          6125 => x"75",
          6126 => x"15",
          6127 => x"e8",
          6128 => x"f6",
          6129 => x"81",
          6130 => x"ff",
          6131 => x"89",
          6132 => x"b3",
          6133 => x"f0",
          6134 => x"2b",
          6135 => x"58",
          6136 => x"83",
          6137 => x"73",
          6138 => x"70",
          6139 => x"32",
          6140 => x"51",
          6141 => x"80",
          6142 => x"38",
          6143 => x"f7",
          6144 => x"09",
          6145 => x"72",
          6146 => x"e4",
          6147 => x"83",
          6148 => x"80",
          6149 => x"a1",
          6150 => x"a8",
          6151 => x"a2",
          6152 => x"f7",
          6153 => x"f7",
          6154 => x"5d",
          6155 => x"5e",
          6156 => x"fc",
          6157 => x"74",
          6158 => x"8d",
          6159 => x"90",
          6160 => x"73",
          6161 => x"82",
          6162 => x"86",
          6163 => x"72",
          6164 => x"8b",
          6165 => x"90",
          6166 => x"73",
          6167 => x"74",
          6168 => x"54",
          6169 => x"2e",
          6170 => x"f7",
          6171 => x"53",
          6172 => x"81",
          6173 => x"81",
          6174 => x"72",
          6175 => x"84",
          6176 => x"f7",
          6177 => x"54",
          6178 => x"84",
          6179 => x"f7",
          6180 => x"e8",
          6181 => x"98",
          6182 => x"54",
          6183 => x"83",
          6184 => x"0b",
          6185 => x"9c",
          6186 => x"9c",
          6187 => x"16",
          6188 => x"06",
          6189 => x"76",
          6190 => x"38",
          6191 => x"a3",
          6192 => x"f7",
          6193 => x"9e",
          6194 => x"9c",
          6195 => x"38",
          6196 => x"83",
          6197 => x"5a",
          6198 => x"83",
          6199 => x"54",
          6200 => x"91",
          6201 => x"14",
          6202 => x"9c",
          6203 => x"7d",
          6204 => x"dc",
          6205 => x"83",
          6206 => x"54",
          6207 => x"2e",
          6208 => x"54",
          6209 => x"ce",
          6210 => x"98",
          6211 => x"f7",
          6212 => x"81",
          6213 => x"77",
          6214 => x"38",
          6215 => x"17",
          6216 => x"b7",
          6217 => x"76",
          6218 => x"54",
          6219 => x"83",
          6220 => x"53",
          6221 => x"82",
          6222 => x"81",
          6223 => x"38",
          6224 => x"34",
          6225 => x"fc",
          6226 => x"58",
          6227 => x"80",
          6228 => x"83",
          6229 => x"2e",
          6230 => x"77",
          6231 => x"06",
          6232 => x"7d",
          6233 => x"ed",
          6234 => x"2e",
          6235 => x"79",
          6236 => x"59",
          6237 => x"75",
          6238 => x"54",
          6239 => x"a1",
          6240 => x"2e",
          6241 => x"17",
          6242 => x"06",
          6243 => x"fe",
          6244 => x"27",
          6245 => x"57",
          6246 => x"54",
          6247 => x"e1",
          6248 => x"10",
          6249 => x"05",
          6250 => x"2b",
          6251 => x"f3",
          6252 => x"33",
          6253 => x"78",
          6254 => x"9c",
          6255 => x"9c",
          6256 => x"ea",
          6257 => x"7d",
          6258 => x"a8",
          6259 => x"ff",
          6260 => x"a0",
          6261 => x"ff",
          6262 => x"ff",
          6263 => x"38",
          6264 => x"b7",
          6265 => x"54",
          6266 => x"83",
          6267 => x"82",
          6268 => x"70",
          6269 => x"07",
          6270 => x"7d",
          6271 => x"83",
          6272 => x"06",
          6273 => x"78",
          6274 => x"c6",
          6275 => x"72",
          6276 => x"83",
          6277 => x"70",
          6278 => x"78",
          6279 => x"ba",
          6280 => x"70",
          6281 => x"54",
          6282 => x"27",
          6283 => x"b7",
          6284 => x"72",
          6285 => x"9a",
          6286 => x"c0",
          6287 => x"f9",
          6288 => x"81",
          6289 => x"82",
          6290 => x"3f",
          6291 => x"c8",
          6292 => x"0d",
          6293 => x"34",
          6294 => x"f9",
          6295 => x"81",
          6296 => x"38",
          6297 => x"14",
          6298 => x"5b",
          6299 => x"90",
          6300 => x"c9",
          6301 => x"83",
          6302 => x"34",
          6303 => x"f6",
          6304 => x"ff",
          6305 => x"86",
          6306 => x"b1",
          6307 => x"ff",
          6308 => x"81",
          6309 => x"96",
          6310 => x"90",
          6311 => x"81",
          6312 => x"8a",
          6313 => x"ff",
          6314 => x"81",
          6315 => x"06",
          6316 => x"83",
          6317 => x"81",
          6318 => x"c0",
          6319 => x"54",
          6320 => x"27",
          6321 => x"87",
          6322 => x"08",
          6323 => x"0c",
          6324 => x"06",
          6325 => x"39",
          6326 => x"f6",
          6327 => x"f9",
          6328 => x"83",
          6329 => x"73",
          6330 => x"53",
          6331 => x"38",
          6332 => x"a2",
          6333 => x"83",
          6334 => x"83",
          6335 => x"83",
          6336 => x"70",
          6337 => x"33",
          6338 => x"33",
          6339 => x"5e",
          6340 => x"fa",
          6341 => x"82",
          6342 => x"06",
          6343 => x"7a",
          6344 => x"2e",
          6345 => x"79",
          6346 => x"81",
          6347 => x"38",
          6348 => x"ef",
          6349 => x"f0",
          6350 => x"39",
          6351 => x"b7",
          6352 => x"54",
          6353 => x"81",
          6354 => x"b7",
          6355 => x"59",
          6356 => x"80",
          6357 => x"be",
          6358 => x"76",
          6359 => x"54",
          6360 => x"be",
          6361 => x"f7",
          6362 => x"53",
          6363 => x"08",
          6364 => x"83",
          6365 => x"83",
          6366 => x"f6",
          6367 => x"b7",
          6368 => x"81",
          6369 => x"11",
          6370 => x"80",
          6371 => x"38",
          6372 => x"83",
          6373 => x"73",
          6374 => x"ff",
          6375 => x"80",
          6376 => x"38",
          6377 => x"83",
          6378 => x"84",
          6379 => x"70",
          6380 => x"56",
          6381 => x"80",
          6382 => x"38",
          6383 => x"83",
          6384 => x"ff",
          6385 => x"39",
          6386 => x"51",
          6387 => x"3f",
          6388 => x"aa",
          6389 => x"fc",
          6390 => x"14",
          6391 => x"f7",
          6392 => x"de",
          6393 => x"0b",
          6394 => x"34",
          6395 => x"33",
          6396 => x"39",
          6397 => x"81",
          6398 => x"3f",
          6399 => x"04",
          6400 => x"80",
          6401 => x"d4",
          6402 => x"02",
          6403 => x"82",
          6404 => x"f3",
          6405 => x"80",
          6406 => x"85",
          6407 => x"d4",
          6408 => x"fe",
          6409 => x"34",
          6410 => x"90",
          6411 => x"87",
          6412 => x"08",
          6413 => x"08",
          6414 => x"90",
          6415 => x"c0",
          6416 => x"52",
          6417 => x"9c",
          6418 => x"72",
          6419 => x"81",
          6420 => x"c0",
          6421 => x"56",
          6422 => x"27",
          6423 => x"81",
          6424 => x"38",
          6425 => x"a4",
          6426 => x"55",
          6427 => x"80",
          6428 => x"55",
          6429 => x"80",
          6430 => x"c0",
          6431 => x"80",
          6432 => x"53",
          6433 => x"9c",
          6434 => x"c0",
          6435 => x"55",
          6436 => x"f6",
          6437 => x"33",
          6438 => x"9c",
          6439 => x"70",
          6440 => x"38",
          6441 => x"2e",
          6442 => x"c0",
          6443 => x"55",
          6444 => x"83",
          6445 => x"71",
          6446 => x"70",
          6447 => x"57",
          6448 => x"2e",
          6449 => x"81",
          6450 => x"71",
          6451 => x"74",
          6452 => x"38",
          6453 => x"c8",
          6454 => x"0d",
          6455 => x"84",
          6456 => x"88",
          6457 => x"fa",
          6458 => x"02",
          6459 => x"05",
          6460 => x"80",
          6461 => x"d4",
          6462 => x"2b",
          6463 => x"80",
          6464 => x"98",
          6465 => x"55",
          6466 => x"83",
          6467 => x"90",
          6468 => x"84",
          6469 => x"90",
          6470 => x"85",
          6471 => x"86",
          6472 => x"f3",
          6473 => x"74",
          6474 => x"83",
          6475 => x"51",
          6476 => x"34",
          6477 => x"f3",
          6478 => x"56",
          6479 => x"15",
          6480 => x"87",
          6481 => x"34",
          6482 => x"9c",
          6483 => x"d4",
          6484 => x"ce",
          6485 => x"87",
          6486 => x"08",
          6487 => x"98",
          6488 => x"70",
          6489 => x"38",
          6490 => x"87",
          6491 => x"08",
          6492 => x"73",
          6493 => x"71",
          6494 => x"db",
          6495 => x"98",
          6496 => x"ff",
          6497 => x"27",
          6498 => x"71",
          6499 => x"2e",
          6500 => x"87",
          6501 => x"08",
          6502 => x"05",
          6503 => x"98",
          6504 => x"87",
          6505 => x"08",
          6506 => x"2e",
          6507 => x"14",
          6508 => x"98",
          6509 => x"52",
          6510 => x"87",
          6511 => x"ff",
          6512 => x"87",
          6513 => x"08",
          6514 => x"26",
          6515 => x"52",
          6516 => x"16",
          6517 => x"06",
          6518 => x"80",
          6519 => x"38",
          6520 => x"06",
          6521 => x"d4",
          6522 => x"70",
          6523 => x"56",
          6524 => x"80",
          6525 => x"84",
          6526 => x"52",
          6527 => x"27",
          6528 => x"70",
          6529 => x"33",
          6530 => x"05",
          6531 => x"71",
          6532 => x"76",
          6533 => x"0c",
          6534 => x"04",
          6535 => x"b9",
          6536 => x"3d",
          6537 => x"51",
          6538 => x"3d",
          6539 => x"84",
          6540 => x"33",
          6541 => x"0b",
          6542 => x"08",
          6543 => x"87",
          6544 => x"06",
          6545 => x"2a",
          6546 => x"55",
          6547 => x"15",
          6548 => x"2a",
          6549 => x"15",
          6550 => x"2a",
          6551 => x"15",
          6552 => x"15",
          6553 => x"f3",
          6554 => x"c6",
          6555 => x"13",
          6556 => x"51",
          6557 => x"97",
          6558 => x"81",
          6559 => x"72",
          6560 => x"54",
          6561 => x"26",
          6562 => x"f3",
          6563 => x"74",
          6564 => x"83",
          6565 => x"55",
          6566 => x"34",
          6567 => x"f3",
          6568 => x"56",
          6569 => x"15",
          6570 => x"87",
          6571 => x"34",
          6572 => x"9c",
          6573 => x"d4",
          6574 => x"ce",
          6575 => x"87",
          6576 => x"08",
          6577 => x"98",
          6578 => x"70",
          6579 => x"38",
          6580 => x"87",
          6581 => x"08",
          6582 => x"73",
          6583 => x"71",
          6584 => x"db",
          6585 => x"98",
          6586 => x"ff",
          6587 => x"27",
          6588 => x"71",
          6589 => x"2e",
          6590 => x"87",
          6591 => x"08",
          6592 => x"05",
          6593 => x"98",
          6594 => x"87",
          6595 => x"08",
          6596 => x"2e",
          6597 => x"14",
          6598 => x"98",
          6599 => x"52",
          6600 => x"87",
          6601 => x"ff",
          6602 => x"87",
          6603 => x"08",
          6604 => x"26",
          6605 => x"52",
          6606 => x"16",
          6607 => x"06",
          6608 => x"80",
          6609 => x"74",
          6610 => x"52",
          6611 => x"38",
          6612 => x"81",
          6613 => x"73",
          6614 => x"38",
          6615 => x"84",
          6616 => x"88",
          6617 => x"ff",
          6618 => x"fb",
          6619 => x"f3",
          6620 => x"80",
          6621 => x"85",
          6622 => x"d4",
          6623 => x"fe",
          6624 => x"34",
          6625 => x"90",
          6626 => x"87",
          6627 => x"08",
          6628 => x"08",
          6629 => x"90",
          6630 => x"c0",
          6631 => x"52",
          6632 => x"9c",
          6633 => x"72",
          6634 => x"81",
          6635 => x"c0",
          6636 => x"52",
          6637 => x"27",
          6638 => x"81",
          6639 => x"38",
          6640 => x"a4",
          6641 => x"53",
          6642 => x"80",
          6643 => x"53",
          6644 => x"80",
          6645 => x"c0",
          6646 => x"80",
          6647 => x"53",
          6648 => x"9c",
          6649 => x"c0",
          6650 => x"51",
          6651 => x"f6",
          6652 => x"33",
          6653 => x"9c",
          6654 => x"73",
          6655 => x"38",
          6656 => x"2e",
          6657 => x"c0",
          6658 => x"51",
          6659 => x"83",
          6660 => x"71",
          6661 => x"70",
          6662 => x"57",
          6663 => x"2e",
          6664 => x"81",
          6665 => x"73",
          6666 => x"ff",
          6667 => x"0d",
          6668 => x"51",
          6669 => x"3f",
          6670 => x"04",
          6671 => x"84",
          6672 => x"7a",
          6673 => x"2a",
          6674 => x"ff",
          6675 => x"2b",
          6676 => x"33",
          6677 => x"71",
          6678 => x"83",
          6679 => x"11",
          6680 => x"12",
          6681 => x"2b",
          6682 => x"07",
          6683 => x"53",
          6684 => x"59",
          6685 => x"53",
          6686 => x"81",
          6687 => x"16",
          6688 => x"83",
          6689 => x"8b",
          6690 => x"2b",
          6691 => x"70",
          6692 => x"33",
          6693 => x"71",
          6694 => x"57",
          6695 => x"59",
          6696 => x"71",
          6697 => x"38",
          6698 => x"85",
          6699 => x"8b",
          6700 => x"2b",
          6701 => x"76",
          6702 => x"54",
          6703 => x"86",
          6704 => x"81",
          6705 => x"73",
          6706 => x"84",
          6707 => x"70",
          6708 => x"33",
          6709 => x"71",
          6710 => x"70",
          6711 => x"55",
          6712 => x"77",
          6713 => x"71",
          6714 => x"84",
          6715 => x"16",
          6716 => x"86",
          6717 => x"0b",
          6718 => x"84",
          6719 => x"53",
          6720 => x"34",
          6721 => x"34",
          6722 => x"08",
          6723 => x"81",
          6724 => x"88",
          6725 => x"80",
          6726 => x"88",
          6727 => x"52",
          6728 => x"34",
          6729 => x"34",
          6730 => x"04",
          6731 => x"87",
          6732 => x"8b",
          6733 => x"2b",
          6734 => x"84",
          6735 => x"17",
          6736 => x"2b",
          6737 => x"2a",
          6738 => x"51",
          6739 => x"71",
          6740 => x"72",
          6741 => x"84",
          6742 => x"70",
          6743 => x"33",
          6744 => x"71",
          6745 => x"83",
          6746 => x"5a",
          6747 => x"05",
          6748 => x"87",
          6749 => x"88",
          6750 => x"88",
          6751 => x"59",
          6752 => x"13",
          6753 => x"13",
          6754 => x"b8",
          6755 => x"33",
          6756 => x"71",
          6757 => x"81",
          6758 => x"70",
          6759 => x"5a",
          6760 => x"72",
          6761 => x"13",
          6762 => x"b8",
          6763 => x"70",
          6764 => x"33",
          6765 => x"71",
          6766 => x"74",
          6767 => x"81",
          6768 => x"88",
          6769 => x"83",
          6770 => x"f8",
          6771 => x"7b",
          6772 => x"52",
          6773 => x"5a",
          6774 => x"77",
          6775 => x"73",
          6776 => x"84",
          6777 => x"70",
          6778 => x"81",
          6779 => x"8b",
          6780 => x"2b",
          6781 => x"70",
          6782 => x"33",
          6783 => x"07",
          6784 => x"06",
          6785 => x"5f",
          6786 => x"5a",
          6787 => x"77",
          6788 => x"81",
          6789 => x"b9",
          6790 => x"17",
          6791 => x"83",
          6792 => x"8b",
          6793 => x"2b",
          6794 => x"70",
          6795 => x"33",
          6796 => x"71",
          6797 => x"58",
          6798 => x"5a",
          6799 => x"70",
          6800 => x"e4",
          6801 => x"81",
          6802 => x"88",
          6803 => x"80",
          6804 => x"88",
          6805 => x"54",
          6806 => x"77",
          6807 => x"84",
          6808 => x"70",
          6809 => x"81",
          6810 => x"8b",
          6811 => x"2b",
          6812 => x"82",
          6813 => x"15",
          6814 => x"2b",
          6815 => x"2a",
          6816 => x"52",
          6817 => x"53",
          6818 => x"34",
          6819 => x"34",
          6820 => x"04",
          6821 => x"79",
          6822 => x"08",
          6823 => x"80",
          6824 => x"77",
          6825 => x"38",
          6826 => x"90",
          6827 => x"0d",
          6828 => x"f4",
          6829 => x"b8",
          6830 => x"0b",
          6831 => x"23",
          6832 => x"53",
          6833 => x"ff",
          6834 => x"d3",
          6835 => x"b9",
          6836 => x"76",
          6837 => x"0b",
          6838 => x"84",
          6839 => x"54",
          6840 => x"34",
          6841 => x"15",
          6842 => x"b8",
          6843 => x"86",
          6844 => x"0b",
          6845 => x"84",
          6846 => x"84",
          6847 => x"ff",
          6848 => x"80",
          6849 => x"ff",
          6850 => x"88",
          6851 => x"55",
          6852 => x"17",
          6853 => x"17",
          6854 => x"b4",
          6855 => x"10",
          6856 => x"b8",
          6857 => x"05",
          6858 => x"82",
          6859 => x"0b",
          6860 => x"fe",
          6861 => x"3d",
          6862 => x"80",
          6863 => x"84",
          6864 => x"38",
          6865 => x"2a",
          6866 => x"83",
          6867 => x"51",
          6868 => x"ff",
          6869 => x"b9",
          6870 => x"11",
          6871 => x"33",
          6872 => x"07",
          6873 => x"5a",
          6874 => x"ff",
          6875 => x"80",
          6876 => x"38",
          6877 => x"10",
          6878 => x"81",
          6879 => x"88",
          6880 => x"81",
          6881 => x"79",
          6882 => x"ff",
          6883 => x"7a",
          6884 => x"5c",
          6885 => x"72",
          6886 => x"38",
          6887 => x"85",
          6888 => x"55",
          6889 => x"33",
          6890 => x"71",
          6891 => x"57",
          6892 => x"38",
          6893 => x"ff",
          6894 => x"77",
          6895 => x"80",
          6896 => x"78",
          6897 => x"81",
          6898 => x"88",
          6899 => x"81",
          6900 => x"56",
          6901 => x"59",
          6902 => x"2e",
          6903 => x"59",
          6904 => x"73",
          6905 => x"38",
          6906 => x"80",
          6907 => x"38",
          6908 => x"82",
          6909 => x"16",
          6910 => x"78",
          6911 => x"80",
          6912 => x"88",
          6913 => x"56",
          6914 => x"74",
          6915 => x"15",
          6916 => x"b8",
          6917 => x"88",
          6918 => x"71",
          6919 => x"75",
          6920 => x"84",
          6921 => x"70",
          6922 => x"81",
          6923 => x"88",
          6924 => x"83",
          6925 => x"f8",
          6926 => x"7e",
          6927 => x"06",
          6928 => x"5c",
          6929 => x"59",
          6930 => x"82",
          6931 => x"81",
          6932 => x"72",
          6933 => x"84",
          6934 => x"18",
          6935 => x"34",
          6936 => x"34",
          6937 => x"08",
          6938 => x"11",
          6939 => x"33",
          6940 => x"71",
          6941 => x"74",
          6942 => x"5c",
          6943 => x"84",
          6944 => x"85",
          6945 => x"b9",
          6946 => x"16",
          6947 => x"86",
          6948 => x"12",
          6949 => x"2b",
          6950 => x"2a",
          6951 => x"59",
          6952 => x"34",
          6953 => x"34",
          6954 => x"08",
          6955 => x"11",
          6956 => x"33",
          6957 => x"71",
          6958 => x"74",
          6959 => x"5c",
          6960 => x"86",
          6961 => x"87",
          6962 => x"b9",
          6963 => x"16",
          6964 => x"84",
          6965 => x"12",
          6966 => x"2b",
          6967 => x"2a",
          6968 => x"59",
          6969 => x"34",
          6970 => x"34",
          6971 => x"08",
          6972 => x"51",
          6973 => x"c8",
          6974 => x"0d",
          6975 => x"33",
          6976 => x"71",
          6977 => x"83",
          6978 => x"05",
          6979 => x"85",
          6980 => x"88",
          6981 => x"88",
          6982 => x"59",
          6983 => x"74",
          6984 => x"76",
          6985 => x"84",
          6986 => x"70",
          6987 => x"33",
          6988 => x"71",
          6989 => x"83",
          6990 => x"05",
          6991 => x"87",
          6992 => x"88",
          6993 => x"88",
          6994 => x"5f",
          6995 => x"57",
          6996 => x"1a",
          6997 => x"1a",
          6998 => x"b8",
          6999 => x"33",
          7000 => x"71",
          7001 => x"81",
          7002 => x"70",
          7003 => x"57",
          7004 => x"77",
          7005 => x"18",
          7006 => x"b8",
          7007 => x"05",
          7008 => x"39",
          7009 => x"79",
          7010 => x"08",
          7011 => x"80",
          7012 => x"77",
          7013 => x"38",
          7014 => x"c8",
          7015 => x"0d",
          7016 => x"fb",
          7017 => x"b9",
          7018 => x"b9",
          7019 => x"3d",
          7020 => x"ff",
          7021 => x"b9",
          7022 => x"80",
          7023 => x"b4",
          7024 => x"80",
          7025 => x"84",
          7026 => x"fe",
          7027 => x"84",
          7028 => x"55",
          7029 => x"81",
          7030 => x"34",
          7031 => x"08",
          7032 => x"15",
          7033 => x"85",
          7034 => x"b9",
          7035 => x"76",
          7036 => x"81",
          7037 => x"34",
          7038 => x"08",
          7039 => x"22",
          7040 => x"80",
          7041 => x"83",
          7042 => x"70",
          7043 => x"51",
          7044 => x"88",
          7045 => x"89",
          7046 => x"b9",
          7047 => x"10",
          7048 => x"b9",
          7049 => x"f8",
          7050 => x"76",
          7051 => x"81",
          7052 => x"34",
          7053 => x"80",
          7054 => x"38",
          7055 => x"ed",
          7056 => x"67",
          7057 => x"70",
          7058 => x"08",
          7059 => x"76",
          7060 => x"aa",
          7061 => x"2e",
          7062 => x"7f",
          7063 => x"d7",
          7064 => x"84",
          7065 => x"38",
          7066 => x"83",
          7067 => x"70",
          7068 => x"06",
          7069 => x"83",
          7070 => x"7f",
          7071 => x"2a",
          7072 => x"ff",
          7073 => x"2b",
          7074 => x"33",
          7075 => x"71",
          7076 => x"70",
          7077 => x"83",
          7078 => x"70",
          7079 => x"fc",
          7080 => x"2b",
          7081 => x"33",
          7082 => x"71",
          7083 => x"70",
          7084 => x"90",
          7085 => x"45",
          7086 => x"54",
          7087 => x"48",
          7088 => x"5f",
          7089 => x"24",
          7090 => x"82",
          7091 => x"16",
          7092 => x"2b",
          7093 => x"10",
          7094 => x"33",
          7095 => x"71",
          7096 => x"90",
          7097 => x"5c",
          7098 => x"56",
          7099 => x"85",
          7100 => x"62",
          7101 => x"38",
          7102 => x"77",
          7103 => x"a2",
          7104 => x"2e",
          7105 => x"60",
          7106 => x"62",
          7107 => x"38",
          7108 => x"61",
          7109 => x"f7",
          7110 => x"70",
          7111 => x"33",
          7112 => x"71",
          7113 => x"7a",
          7114 => x"81",
          7115 => x"98",
          7116 => x"2b",
          7117 => x"59",
          7118 => x"5b",
          7119 => x"24",
          7120 => x"76",
          7121 => x"33",
          7122 => x"71",
          7123 => x"83",
          7124 => x"11",
          7125 => x"87",
          7126 => x"8b",
          7127 => x"2b",
          7128 => x"84",
          7129 => x"15",
          7130 => x"2b",
          7131 => x"2a",
          7132 => x"52",
          7133 => x"53",
          7134 => x"77",
          7135 => x"79",
          7136 => x"84",
          7137 => x"70",
          7138 => x"33",
          7139 => x"71",
          7140 => x"83",
          7141 => x"05",
          7142 => x"87",
          7143 => x"88",
          7144 => x"88",
          7145 => x"5e",
          7146 => x"41",
          7147 => x"16",
          7148 => x"16",
          7149 => x"b8",
          7150 => x"33",
          7151 => x"71",
          7152 => x"81",
          7153 => x"70",
          7154 => x"5c",
          7155 => x"79",
          7156 => x"1a",
          7157 => x"b8",
          7158 => x"82",
          7159 => x"12",
          7160 => x"2b",
          7161 => x"07",
          7162 => x"33",
          7163 => x"71",
          7164 => x"70",
          7165 => x"5c",
          7166 => x"5a",
          7167 => x"79",
          7168 => x"1a",
          7169 => x"b8",
          7170 => x"70",
          7171 => x"33",
          7172 => x"71",
          7173 => x"74",
          7174 => x"33",
          7175 => x"71",
          7176 => x"70",
          7177 => x"5c",
          7178 => x"5a",
          7179 => x"82",
          7180 => x"83",
          7181 => x"b9",
          7182 => x"1f",
          7183 => x"83",
          7184 => x"88",
          7185 => x"57",
          7186 => x"83",
          7187 => x"5a",
          7188 => x"84",
          7189 => x"c4",
          7190 => x"b9",
          7191 => x"84",
          7192 => x"05",
          7193 => x"ff",
          7194 => x"44",
          7195 => x"26",
          7196 => x"7e",
          7197 => x"b9",
          7198 => x"3d",
          7199 => x"ff",
          7200 => x"b9",
          7201 => x"80",
          7202 => x"b4",
          7203 => x"80",
          7204 => x"84",
          7205 => x"fe",
          7206 => x"84",
          7207 => x"5e",
          7208 => x"81",
          7209 => x"34",
          7210 => x"08",
          7211 => x"1e",
          7212 => x"85",
          7213 => x"b9",
          7214 => x"60",
          7215 => x"81",
          7216 => x"34",
          7217 => x"08",
          7218 => x"22",
          7219 => x"80",
          7220 => x"83",
          7221 => x"70",
          7222 => x"5a",
          7223 => x"88",
          7224 => x"89",
          7225 => x"b9",
          7226 => x"10",
          7227 => x"b9",
          7228 => x"f8",
          7229 => x"60",
          7230 => x"81",
          7231 => x"34",
          7232 => x"08",
          7233 => x"d3",
          7234 => x"2e",
          7235 => x"7e",
          7236 => x"2e",
          7237 => x"7f",
          7238 => x"3f",
          7239 => x"08",
          7240 => x"0c",
          7241 => x"04",
          7242 => x"b9",
          7243 => x"83",
          7244 => x"5e",
          7245 => x"70",
          7246 => x"33",
          7247 => x"07",
          7248 => x"06",
          7249 => x"48",
          7250 => x"40",
          7251 => x"60",
          7252 => x"61",
          7253 => x"08",
          7254 => x"2a",
          7255 => x"82",
          7256 => x"83",
          7257 => x"b9",
          7258 => x"1f",
          7259 => x"12",
          7260 => x"2b",
          7261 => x"2b",
          7262 => x"06",
          7263 => x"83",
          7264 => x"70",
          7265 => x"5c",
          7266 => x"5b",
          7267 => x"82",
          7268 => x"81",
          7269 => x"60",
          7270 => x"34",
          7271 => x"08",
          7272 => x"7b",
          7273 => x"1c",
          7274 => x"b9",
          7275 => x"84",
          7276 => x"88",
          7277 => x"fd",
          7278 => x"75",
          7279 => x"ff",
          7280 => x"54",
          7281 => x"77",
          7282 => x"06",
          7283 => x"83",
          7284 => x"82",
          7285 => x"18",
          7286 => x"2b",
          7287 => x"10",
          7288 => x"33",
          7289 => x"71",
          7290 => x"90",
          7291 => x"5e",
          7292 => x"58",
          7293 => x"80",
          7294 => x"38",
          7295 => x"61",
          7296 => x"83",
          7297 => x"24",
          7298 => x"77",
          7299 => x"06",
          7300 => x"27",
          7301 => x"fe",
          7302 => x"ff",
          7303 => x"b9",
          7304 => x"80",
          7305 => x"b4",
          7306 => x"80",
          7307 => x"84",
          7308 => x"fe",
          7309 => x"84",
          7310 => x"5a",
          7311 => x"81",
          7312 => x"34",
          7313 => x"08",
          7314 => x"1a",
          7315 => x"85",
          7316 => x"b9",
          7317 => x"7e",
          7318 => x"81",
          7319 => x"34",
          7320 => x"08",
          7321 => x"22",
          7322 => x"80",
          7323 => x"83",
          7324 => x"70",
          7325 => x"56",
          7326 => x"64",
          7327 => x"73",
          7328 => x"34",
          7329 => x"22",
          7330 => x"10",
          7331 => x"08",
          7332 => x"42",
          7333 => x"82",
          7334 => x"61",
          7335 => x"fc",
          7336 => x"7a",
          7337 => x"38",
          7338 => x"ff",
          7339 => x"7b",
          7340 => x"38",
          7341 => x"76",
          7342 => x"bd",
          7343 => x"ea",
          7344 => x"54",
          7345 => x"c8",
          7346 => x"0d",
          7347 => x"82",
          7348 => x"12",
          7349 => x"2b",
          7350 => x"07",
          7351 => x"11",
          7352 => x"33",
          7353 => x"71",
          7354 => x"7e",
          7355 => x"33",
          7356 => x"71",
          7357 => x"70",
          7358 => x"44",
          7359 => x"46",
          7360 => x"45",
          7361 => x"84",
          7362 => x"64",
          7363 => x"84",
          7364 => x"70",
          7365 => x"33",
          7366 => x"71",
          7367 => x"83",
          7368 => x"05",
          7369 => x"87",
          7370 => x"88",
          7371 => x"88",
          7372 => x"42",
          7373 => x"5d",
          7374 => x"86",
          7375 => x"64",
          7376 => x"84",
          7377 => x"16",
          7378 => x"12",
          7379 => x"2b",
          7380 => x"ff",
          7381 => x"2a",
          7382 => x"5d",
          7383 => x"79",
          7384 => x"84",
          7385 => x"70",
          7386 => x"33",
          7387 => x"71",
          7388 => x"83",
          7389 => x"05",
          7390 => x"15",
          7391 => x"2b",
          7392 => x"2a",
          7393 => x"40",
          7394 => x"54",
          7395 => x"75",
          7396 => x"84",
          7397 => x"70",
          7398 => x"81",
          7399 => x"8b",
          7400 => x"2b",
          7401 => x"82",
          7402 => x"15",
          7403 => x"2b",
          7404 => x"2a",
          7405 => x"5b",
          7406 => x"55",
          7407 => x"34",
          7408 => x"34",
          7409 => x"08",
          7410 => x"11",
          7411 => x"33",
          7412 => x"07",
          7413 => x"56",
          7414 => x"42",
          7415 => x"7e",
          7416 => x"51",
          7417 => x"3f",
          7418 => x"08",
          7419 => x"78",
          7420 => x"06",
          7421 => x"99",
          7422 => x"f4",
          7423 => x"b8",
          7424 => x"0b",
          7425 => x"23",
          7426 => x"53",
          7427 => x"ff",
          7428 => x"c0",
          7429 => x"b9",
          7430 => x"7f",
          7431 => x"0b",
          7432 => x"84",
          7433 => x"55",
          7434 => x"34",
          7435 => x"16",
          7436 => x"b8",
          7437 => x"86",
          7438 => x"0b",
          7439 => x"84",
          7440 => x"84",
          7441 => x"ff",
          7442 => x"80",
          7443 => x"ff",
          7444 => x"88",
          7445 => x"44",
          7446 => x"1f",
          7447 => x"1f",
          7448 => x"b4",
          7449 => x"10",
          7450 => x"b8",
          7451 => x"05",
          7452 => x"82",
          7453 => x"0b",
          7454 => x"7e",
          7455 => x"3f",
          7456 => x"c0",
          7457 => x"33",
          7458 => x"71",
          7459 => x"83",
          7460 => x"05",
          7461 => x"85",
          7462 => x"88",
          7463 => x"88",
          7464 => x"5e",
          7465 => x"76",
          7466 => x"34",
          7467 => x"05",
          7468 => x"b8",
          7469 => x"84",
          7470 => x"12",
          7471 => x"2b",
          7472 => x"07",
          7473 => x"14",
          7474 => x"33",
          7475 => x"07",
          7476 => x"41",
          7477 => x"59",
          7478 => x"79",
          7479 => x"34",
          7480 => x"05",
          7481 => x"b8",
          7482 => x"33",
          7483 => x"71",
          7484 => x"81",
          7485 => x"70",
          7486 => x"42",
          7487 => x"78",
          7488 => x"19",
          7489 => x"b8",
          7490 => x"70",
          7491 => x"33",
          7492 => x"71",
          7493 => x"74",
          7494 => x"81",
          7495 => x"88",
          7496 => x"83",
          7497 => x"f8",
          7498 => x"63",
          7499 => x"5d",
          7500 => x"40",
          7501 => x"7f",
          7502 => x"7b",
          7503 => x"84",
          7504 => x"70",
          7505 => x"81",
          7506 => x"8b",
          7507 => x"2b",
          7508 => x"70",
          7509 => x"33",
          7510 => x"07",
          7511 => x"06",
          7512 => x"48",
          7513 => x"46",
          7514 => x"60",
          7515 => x"60",
          7516 => x"61",
          7517 => x"06",
          7518 => x"39",
          7519 => x"87",
          7520 => x"8b",
          7521 => x"2b",
          7522 => x"84",
          7523 => x"19",
          7524 => x"2b",
          7525 => x"2a",
          7526 => x"52",
          7527 => x"84",
          7528 => x"85",
          7529 => x"b9",
          7530 => x"19",
          7531 => x"85",
          7532 => x"8b",
          7533 => x"2b",
          7534 => x"86",
          7535 => x"15",
          7536 => x"2b",
          7537 => x"2a",
          7538 => x"52",
          7539 => x"56",
          7540 => x"05",
          7541 => x"87",
          7542 => x"b9",
          7543 => x"70",
          7544 => x"33",
          7545 => x"07",
          7546 => x"06",
          7547 => x"5b",
          7548 => x"77",
          7549 => x"81",
          7550 => x"b9",
          7551 => x"1f",
          7552 => x"12",
          7553 => x"2b",
          7554 => x"07",
          7555 => x"33",
          7556 => x"71",
          7557 => x"70",
          7558 => x"ff",
          7559 => x"05",
          7560 => x"56",
          7561 => x"58",
          7562 => x"55",
          7563 => x"34",
          7564 => x"34",
          7565 => x"08",
          7566 => x"33",
          7567 => x"71",
          7568 => x"83",
          7569 => x"05",
          7570 => x"12",
          7571 => x"2b",
          7572 => x"ff",
          7573 => x"2a",
          7574 => x"58",
          7575 => x"55",
          7576 => x"76",
          7577 => x"84",
          7578 => x"70",
          7579 => x"33",
          7580 => x"71",
          7581 => x"83",
          7582 => x"11",
          7583 => x"87",
          7584 => x"8b",
          7585 => x"2b",
          7586 => x"84",
          7587 => x"15",
          7588 => x"2b",
          7589 => x"2a",
          7590 => x"52",
          7591 => x"53",
          7592 => x"57",
          7593 => x"34",
          7594 => x"34",
          7595 => x"08",
          7596 => x"11",
          7597 => x"33",
          7598 => x"71",
          7599 => x"74",
          7600 => x"33",
          7601 => x"71",
          7602 => x"70",
          7603 => x"42",
          7604 => x"57",
          7605 => x"86",
          7606 => x"87",
          7607 => x"b9",
          7608 => x"70",
          7609 => x"33",
          7610 => x"07",
          7611 => x"06",
          7612 => x"5a",
          7613 => x"76",
          7614 => x"81",
          7615 => x"b9",
          7616 => x"1f",
          7617 => x"83",
          7618 => x"8b",
          7619 => x"2b",
          7620 => x"73",
          7621 => x"33",
          7622 => x"07",
          7623 => x"41",
          7624 => x"5f",
          7625 => x"79",
          7626 => x"81",
          7627 => x"b9",
          7628 => x"1f",
          7629 => x"12",
          7630 => x"2b",
          7631 => x"07",
          7632 => x"14",
          7633 => x"33",
          7634 => x"07",
          7635 => x"41",
          7636 => x"5f",
          7637 => x"79",
          7638 => x"75",
          7639 => x"84",
          7640 => x"70",
          7641 => x"33",
          7642 => x"71",
          7643 => x"66",
          7644 => x"70",
          7645 => x"52",
          7646 => x"05",
          7647 => x"fe",
          7648 => x"84",
          7649 => x"1e",
          7650 => x"65",
          7651 => x"83",
          7652 => x"5d",
          7653 => x"d5",
          7654 => x"33",
          7655 => x"71",
          7656 => x"83",
          7657 => x"05",
          7658 => x"85",
          7659 => x"88",
          7660 => x"88",
          7661 => x"5d",
          7662 => x"7a",
          7663 => x"34",
          7664 => x"05",
          7665 => x"b8",
          7666 => x"84",
          7667 => x"12",
          7668 => x"2b",
          7669 => x"07",
          7670 => x"14",
          7671 => x"33",
          7672 => x"07",
          7673 => x"5b",
          7674 => x"5c",
          7675 => x"73",
          7676 => x"34",
          7677 => x"05",
          7678 => x"b8",
          7679 => x"33",
          7680 => x"71",
          7681 => x"81",
          7682 => x"70",
          7683 => x"5f",
          7684 => x"75",
          7685 => x"16",
          7686 => x"b8",
          7687 => x"70",
          7688 => x"33",
          7689 => x"71",
          7690 => x"74",
          7691 => x"81",
          7692 => x"88",
          7693 => x"83",
          7694 => x"f8",
          7695 => x"63",
          7696 => x"44",
          7697 => x"5e",
          7698 => x"74",
          7699 => x"7b",
          7700 => x"84",
          7701 => x"70",
          7702 => x"81",
          7703 => x"8b",
          7704 => x"2b",
          7705 => x"70",
          7706 => x"33",
          7707 => x"07",
          7708 => x"06",
          7709 => x"47",
          7710 => x"46",
          7711 => x"7f",
          7712 => x"81",
          7713 => x"83",
          7714 => x"5b",
          7715 => x"7e",
          7716 => x"e5",
          7717 => x"b9",
          7718 => x"84",
          7719 => x"80",
          7720 => x"62",
          7721 => x"84",
          7722 => x"51",
          7723 => x"3f",
          7724 => x"88",
          7725 => x"61",
          7726 => x"b7",
          7727 => x"39",
          7728 => x"7a",
          7729 => x"b9",
          7730 => x"58",
          7731 => x"b7",
          7732 => x"77",
          7733 => x"84",
          7734 => x"89",
          7735 => x"77",
          7736 => x"3f",
          7737 => x"08",
          7738 => x"c8",
          7739 => x"e6",
          7740 => x"80",
          7741 => x"c8",
          7742 => x"b7",
          7743 => x"84",
          7744 => x"89",
          7745 => x"84",
          7746 => x"84",
          7747 => x"a0",
          7748 => x"b9",
          7749 => x"80",
          7750 => x"52",
          7751 => x"51",
          7752 => x"3f",
          7753 => x"08",
          7754 => x"34",
          7755 => x"16",
          7756 => x"b8",
          7757 => x"84",
          7758 => x"0b",
          7759 => x"84",
          7760 => x"56",
          7761 => x"34",
          7762 => x"17",
          7763 => x"b8",
          7764 => x"b4",
          7765 => x"fe",
          7766 => x"70",
          7767 => x"06",
          7768 => x"58",
          7769 => x"74",
          7770 => x"73",
          7771 => x"84",
          7772 => x"70",
          7773 => x"84",
          7774 => x"05",
          7775 => x"55",
          7776 => x"34",
          7777 => x"15",
          7778 => x"77",
          7779 => x"c6",
          7780 => x"39",
          7781 => x"02",
          7782 => x"51",
          7783 => x"72",
          7784 => x"84",
          7785 => x"33",
          7786 => x"b9",
          7787 => x"3d",
          7788 => x"3d",
          7789 => x"05",
          7790 => x"53",
          7791 => x"9d",
          7792 => x"d4",
          7793 => x"b9",
          7794 => x"ff",
          7795 => x"87",
          7796 => x"b9",
          7797 => x"84",
          7798 => x"33",
          7799 => x"b9",
          7800 => x"3d",
          7801 => x"3d",
          7802 => x"60",
          7803 => x"af",
          7804 => x"5c",
          7805 => x"54",
          7806 => x"87",
          7807 => x"c4",
          7808 => x"73",
          7809 => x"83",
          7810 => x"38",
          7811 => x"0b",
          7812 => x"8c",
          7813 => x"75",
          7814 => x"d5",
          7815 => x"b9",
          7816 => x"ff",
          7817 => x"80",
          7818 => x"87",
          7819 => x"08",
          7820 => x"38",
          7821 => x"d6",
          7822 => x"80",
          7823 => x"73",
          7824 => x"38",
          7825 => x"55",
          7826 => x"c8",
          7827 => x"0d",
          7828 => x"16",
          7829 => x"81",
          7830 => x"55",
          7831 => x"26",
          7832 => x"d5",
          7833 => x"0d",
          7834 => x"02",
          7835 => x"05",
          7836 => x"57",
          7837 => x"76",
          7838 => x"38",
          7839 => x"17",
          7840 => x"81",
          7841 => x"55",
          7842 => x"73",
          7843 => x"87",
          7844 => x"0c",
          7845 => x"52",
          7846 => x"8e",
          7847 => x"c8",
          7848 => x"06",
          7849 => x"2e",
          7850 => x"c0",
          7851 => x"54",
          7852 => x"79",
          7853 => x"38",
          7854 => x"80",
          7855 => x"80",
          7856 => x"81",
          7857 => x"74",
          7858 => x"0c",
          7859 => x"04",
          7860 => x"81",
          7861 => x"ff",
          7862 => x"56",
          7863 => x"ff",
          7864 => x"39",
          7865 => x"78",
          7866 => x"9b",
          7867 => x"88",
          7868 => x"33",
          7869 => x"81",
          7870 => x"26",
          7871 => x"b9",
          7872 => x"53",
          7873 => x"54",
          7874 => x"9b",
          7875 => x"87",
          7876 => x"0c",
          7877 => x"73",
          7878 => x"72",
          7879 => x"38",
          7880 => x"9a",
          7881 => x"72",
          7882 => x"0c",
          7883 => x"04",
          7884 => x"75",
          7885 => x"b9",
          7886 => x"3d",
          7887 => x"80",
          7888 => x"0b",
          7889 => x"0c",
          7890 => x"04",
          7891 => x"87",
          7892 => x"11",
          7893 => x"cd",
          7894 => x"70",
          7895 => x"06",
          7896 => x"80",
          7897 => x"87",
          7898 => x"08",
          7899 => x"38",
          7900 => x"8c",
          7901 => x"ca",
          7902 => x"0c",
          7903 => x"8c",
          7904 => x"08",
          7905 => x"73",
          7906 => x"9b",
          7907 => x"82",
          7908 => x"ee",
          7909 => x"39",
          7910 => x"7c",
          7911 => x"83",
          7912 => x"5b",
          7913 => x"77",
          7914 => x"06",
          7915 => x"33",
          7916 => x"2e",
          7917 => x"80",
          7918 => x"81",
          7919 => x"fe",
          7920 => x"b9",
          7921 => x"2e",
          7922 => x"59",
          7923 => x"c8",
          7924 => x"0d",
          7925 => x"b4",
          7926 => x"b8",
          7927 => x"81",
          7928 => x"5a",
          7929 => x"81",
          7930 => x"c8",
          7931 => x"09",
          7932 => x"38",
          7933 => x"08",
          7934 => x"b4",
          7935 => x"a8",
          7936 => x"a0",
          7937 => x"b9",
          7938 => x"58",
          7939 => x"76",
          7940 => x"38",
          7941 => x"55",
          7942 => x"09",
          7943 => x"8e",
          7944 => x"75",
          7945 => x"52",
          7946 => x"51",
          7947 => x"76",
          7948 => x"59",
          7949 => x"09",
          7950 => x"fb",
          7951 => x"33",
          7952 => x"2e",
          7953 => x"fe",
          7954 => x"18",
          7955 => x"7a",
          7956 => x"75",
          7957 => x"57",
          7958 => x"57",
          7959 => x"80",
          7960 => x"b6",
          7961 => x"aa",
          7962 => x"19",
          7963 => x"7a",
          7964 => x"0b",
          7965 => x"80",
          7966 => x"19",
          7967 => x"0b",
          7968 => x"80",
          7969 => x"9c",
          7970 => x"f2",
          7971 => x"19",
          7972 => x"0b",
          7973 => x"34",
          7974 => x"84",
          7975 => x"94",
          7976 => x"74",
          7977 => x"34",
          7978 => x"5b",
          7979 => x"19",
          7980 => x"2a",
          7981 => x"a2",
          7982 => x"98",
          7983 => x"84",
          7984 => x"90",
          7985 => x"7a",
          7986 => x"34",
          7987 => x"55",
          7988 => x"19",
          7989 => x"2a",
          7990 => x"a6",
          7991 => x"98",
          7992 => x"84",
          7993 => x"a4",
          7994 => x"05",
          7995 => x"0c",
          7996 => x"7a",
          7997 => x"81",
          7998 => x"fa",
          7999 => x"84",
          8000 => x"53",
          8001 => x"18",
          8002 => x"d8",
          8003 => x"c8",
          8004 => x"fd",
          8005 => x"b2",
          8006 => x"0d",
          8007 => x"08",
          8008 => x"81",
          8009 => x"38",
          8010 => x"76",
          8011 => x"81",
          8012 => x"b9",
          8013 => x"3d",
          8014 => x"77",
          8015 => x"74",
          8016 => x"cc",
          8017 => x"24",
          8018 => x"74",
          8019 => x"81",
          8020 => x"75",
          8021 => x"70",
          8022 => x"19",
          8023 => x"5a",
          8024 => x"17",
          8025 => x"b0",
          8026 => x"33",
          8027 => x"2e",
          8028 => x"83",
          8029 => x"54",
          8030 => x"17",
          8031 => x"33",
          8032 => x"3f",
          8033 => x"08",
          8034 => x"38",
          8035 => x"5b",
          8036 => x"0c",
          8037 => x"38",
          8038 => x"06",
          8039 => x"33",
          8040 => x"89",
          8041 => x"08",
          8042 => x"5d",
          8043 => x"08",
          8044 => x"38",
          8045 => x"18",
          8046 => x"56",
          8047 => x"2e",
          8048 => x"84",
          8049 => x"54",
          8050 => x"17",
          8051 => x"33",
          8052 => x"3f",
          8053 => x"08",
          8054 => x"38",
          8055 => x"5a",
          8056 => x"0c",
          8057 => x"38",
          8058 => x"06",
          8059 => x"33",
          8060 => x"7e",
          8061 => x"06",
          8062 => x"53",
          8063 => x"5d",
          8064 => x"38",
          8065 => x"06",
          8066 => x"0c",
          8067 => x"04",
          8068 => x"a8",
          8069 => x"59",
          8070 => x"79",
          8071 => x"80",
          8072 => x"33",
          8073 => x"5b",
          8074 => x"09",
          8075 => x"c2",
          8076 => x"78",
          8077 => x"52",
          8078 => x"51",
          8079 => x"84",
          8080 => x"80",
          8081 => x"ff",
          8082 => x"78",
          8083 => x"79",
          8084 => x"75",
          8085 => x"06",
          8086 => x"05",
          8087 => x"71",
          8088 => x"2b",
          8089 => x"c8",
          8090 => x"8f",
          8091 => x"74",
          8092 => x"81",
          8093 => x"38",
          8094 => x"a8",
          8095 => x"59",
          8096 => x"79",
          8097 => x"80",
          8098 => x"33",
          8099 => x"5b",
          8100 => x"09",
          8101 => x"81",
          8102 => x"78",
          8103 => x"52",
          8104 => x"51",
          8105 => x"84",
          8106 => x"80",
          8107 => x"ff",
          8108 => x"78",
          8109 => x"79",
          8110 => x"75",
          8111 => x"fc",
          8112 => x"b8",
          8113 => x"33",
          8114 => x"71",
          8115 => x"88",
          8116 => x"14",
          8117 => x"07",
          8118 => x"33",
          8119 => x"ff",
          8120 => x"07",
          8121 => x"0c",
          8122 => x"59",
          8123 => x"3d",
          8124 => x"54",
          8125 => x"53",
          8126 => x"53",
          8127 => x"52",
          8128 => x"3f",
          8129 => x"b9",
          8130 => x"2e",
          8131 => x"fe",
          8132 => x"b9",
          8133 => x"18",
          8134 => x"08",
          8135 => x"31",
          8136 => x"08",
          8137 => x"a0",
          8138 => x"fe",
          8139 => x"17",
          8140 => x"82",
          8141 => x"06",
          8142 => x"81",
          8143 => x"08",
          8144 => x"05",
          8145 => x"81",
          8146 => x"f6",
          8147 => x"5a",
          8148 => x"81",
          8149 => x"08",
          8150 => x"70",
          8151 => x"33",
          8152 => x"81",
          8153 => x"c8",
          8154 => x"09",
          8155 => x"81",
          8156 => x"c8",
          8157 => x"34",
          8158 => x"a8",
          8159 => x"5d",
          8160 => x"08",
          8161 => x"82",
          8162 => x"7d",
          8163 => x"cb",
          8164 => x"c8",
          8165 => x"de",
          8166 => x"b4",
          8167 => x"b8",
          8168 => x"81",
          8169 => x"5c",
          8170 => x"81",
          8171 => x"c8",
          8172 => x"09",
          8173 => x"ff",
          8174 => x"c8",
          8175 => x"34",
          8176 => x"a8",
          8177 => x"84",
          8178 => x"5b",
          8179 => x"18",
          8180 => x"c5",
          8181 => x"33",
          8182 => x"2e",
          8183 => x"fd",
          8184 => x"54",
          8185 => x"a0",
          8186 => x"53",
          8187 => x"17",
          8188 => x"f1",
          8189 => x"fd",
          8190 => x"54",
          8191 => x"53",
          8192 => x"53",
          8193 => x"52",
          8194 => x"3f",
          8195 => x"b9",
          8196 => x"2e",
          8197 => x"fb",
          8198 => x"b9",
          8199 => x"18",
          8200 => x"08",
          8201 => x"31",
          8202 => x"08",
          8203 => x"a0",
          8204 => x"fb",
          8205 => x"17",
          8206 => x"82",
          8207 => x"06",
          8208 => x"81",
          8209 => x"08",
          8210 => x"05",
          8211 => x"81",
          8212 => x"f4",
          8213 => x"5a",
          8214 => x"81",
          8215 => x"08",
          8216 => x"05",
          8217 => x"81",
          8218 => x"f3",
          8219 => x"86",
          8220 => x"7a",
          8221 => x"fa",
          8222 => x"3d",
          8223 => x"64",
          8224 => x"82",
          8225 => x"27",
          8226 => x"9c",
          8227 => x"95",
          8228 => x"55",
          8229 => x"96",
          8230 => x"24",
          8231 => x"74",
          8232 => x"8a",
          8233 => x"b9",
          8234 => x"3d",
          8235 => x"88",
          8236 => x"08",
          8237 => x"0b",
          8238 => x"58",
          8239 => x"2e",
          8240 => x"83",
          8241 => x"5b",
          8242 => x"2e",
          8243 => x"83",
          8244 => x"54",
          8245 => x"19",
          8246 => x"33",
          8247 => x"3f",
          8248 => x"08",
          8249 => x"38",
          8250 => x"5a",
          8251 => x"0c",
          8252 => x"ff",
          8253 => x"10",
          8254 => x"79",
          8255 => x"ff",
          8256 => x"5e",
          8257 => x"34",
          8258 => x"5a",
          8259 => x"34",
          8260 => x"1a",
          8261 => x"b9",
          8262 => x"3d",
          8263 => x"83",
          8264 => x"06",
          8265 => x"75",
          8266 => x"1a",
          8267 => x"80",
          8268 => x"08",
          8269 => x"78",
          8270 => x"38",
          8271 => x"7c",
          8272 => x"7c",
          8273 => x"06",
          8274 => x"81",
          8275 => x"b8",
          8276 => x"19",
          8277 => x"8e",
          8278 => x"c8",
          8279 => x"85",
          8280 => x"81",
          8281 => x"1a",
          8282 => x"79",
          8283 => x"75",
          8284 => x"fc",
          8285 => x"b8",
          8286 => x"33",
          8287 => x"8f",
          8288 => x"f0",
          8289 => x"41",
          8290 => x"7d",
          8291 => x"88",
          8292 => x"b9",
          8293 => x"90",
          8294 => x"ba",
          8295 => x"98",
          8296 => x"bb",
          8297 => x"0b",
          8298 => x"fe",
          8299 => x"81",
          8300 => x"89",
          8301 => x"08",
          8302 => x"08",
          8303 => x"76",
          8304 => x"38",
          8305 => x"1a",
          8306 => x"56",
          8307 => x"2e",
          8308 => x"82",
          8309 => x"54",
          8310 => x"19",
          8311 => x"33",
          8312 => x"3f",
          8313 => x"08",
          8314 => x"38",
          8315 => x"5c",
          8316 => x"0c",
          8317 => x"fd",
          8318 => x"83",
          8319 => x"b8",
          8320 => x"77",
          8321 => x"5f",
          8322 => x"7c",
          8323 => x"38",
          8324 => x"9f",
          8325 => x"33",
          8326 => x"07",
          8327 => x"77",
          8328 => x"83",
          8329 => x"89",
          8330 => x"08",
          8331 => x"0b",
          8332 => x"56",
          8333 => x"2e",
          8334 => x"81",
          8335 => x"b8",
          8336 => x"81",
          8337 => x"57",
          8338 => x"81",
          8339 => x"c8",
          8340 => x"09",
          8341 => x"c7",
          8342 => x"c8",
          8343 => x"34",
          8344 => x"70",
          8345 => x"31",
          8346 => x"84",
          8347 => x"5b",
          8348 => x"74",
          8349 => x"38",
          8350 => x"55",
          8351 => x"82",
          8352 => x"54",
          8353 => x"52",
          8354 => x"51",
          8355 => x"84",
          8356 => x"80",
          8357 => x"ff",
          8358 => x"75",
          8359 => x"77",
          8360 => x"7d",
          8361 => x"19",
          8362 => x"84",
          8363 => x"7c",
          8364 => x"88",
          8365 => x"81",
          8366 => x"8f",
          8367 => x"5c",
          8368 => x"81",
          8369 => x"34",
          8370 => x"81",
          8371 => x"b8",
          8372 => x"81",
          8373 => x"5d",
          8374 => x"81",
          8375 => x"c8",
          8376 => x"09",
          8377 => x"88",
          8378 => x"c8",
          8379 => x"34",
          8380 => x"70",
          8381 => x"31",
          8382 => x"84",
          8383 => x"5d",
          8384 => x"7e",
          8385 => x"ca",
          8386 => x"33",
          8387 => x"2e",
          8388 => x"fb",
          8389 => x"54",
          8390 => x"7c",
          8391 => x"33",
          8392 => x"3f",
          8393 => x"aa",
          8394 => x"76",
          8395 => x"70",
          8396 => x"33",
          8397 => x"ad",
          8398 => x"84",
          8399 => x"7d",
          8400 => x"06",
          8401 => x"84",
          8402 => x"83",
          8403 => x"19",
          8404 => x"1b",
          8405 => x"1b",
          8406 => x"c8",
          8407 => x"56",
          8408 => x"27",
          8409 => x"82",
          8410 => x"74",
          8411 => x"81",
          8412 => x"38",
          8413 => x"1f",
          8414 => x"81",
          8415 => x"ed",
          8416 => x"5c",
          8417 => x"81",
          8418 => x"b8",
          8419 => x"81",
          8420 => x"57",
          8421 => x"81",
          8422 => x"c8",
          8423 => x"09",
          8424 => x"c5",
          8425 => x"c8",
          8426 => x"34",
          8427 => x"70",
          8428 => x"31",
          8429 => x"84",
          8430 => x"5d",
          8431 => x"7e",
          8432 => x"87",
          8433 => x"33",
          8434 => x"2e",
          8435 => x"fa",
          8436 => x"54",
          8437 => x"76",
          8438 => x"33",
          8439 => x"3f",
          8440 => x"e7",
          8441 => x"79",
          8442 => x"52",
          8443 => x"51",
          8444 => x"7e",
          8445 => x"39",
          8446 => x"83",
          8447 => x"05",
          8448 => x"ff",
          8449 => x"58",
          8450 => x"34",
          8451 => x"5a",
          8452 => x"34",
          8453 => x"7e",
          8454 => x"39",
          8455 => x"2b",
          8456 => x"7a",
          8457 => x"83",
          8458 => x"98",
          8459 => x"06",
          8460 => x"06",
          8461 => x"5f",
          8462 => x"7d",
          8463 => x"2a",
          8464 => x"1d",
          8465 => x"2a",
          8466 => x"1d",
          8467 => x"2a",
          8468 => x"1d",
          8469 => x"39",
          8470 => x"7c",
          8471 => x"5b",
          8472 => x"81",
          8473 => x"19",
          8474 => x"80",
          8475 => x"38",
          8476 => x"08",
          8477 => x"38",
          8478 => x"70",
          8479 => x"80",
          8480 => x"38",
          8481 => x"81",
          8482 => x"56",
          8483 => x"9c",
          8484 => x"26",
          8485 => x"56",
          8486 => x"82",
          8487 => x"52",
          8488 => x"f5",
          8489 => x"c8",
          8490 => x"81",
          8491 => x"58",
          8492 => x"08",
          8493 => x"38",
          8494 => x"08",
          8495 => x"70",
          8496 => x"25",
          8497 => x"51",
          8498 => x"73",
          8499 => x"75",
          8500 => x"81",
          8501 => x"38",
          8502 => x"84",
          8503 => x"8c",
          8504 => x"81",
          8505 => x"39",
          8506 => x"08",
          8507 => x"7a",
          8508 => x"f0",
          8509 => x"55",
          8510 => x"c8",
          8511 => x"38",
          8512 => x"08",
          8513 => x"c8",
          8514 => x"ce",
          8515 => x"08",
          8516 => x"08",
          8517 => x"7a",
          8518 => x"39",
          8519 => x"9c",
          8520 => x"26",
          8521 => x"56",
          8522 => x"51",
          8523 => x"80",
          8524 => x"c8",
          8525 => x"81",
          8526 => x"b9",
          8527 => x"70",
          8528 => x"07",
          8529 => x"7b",
          8530 => x"c8",
          8531 => x"51",
          8532 => x"ff",
          8533 => x"b9",
          8534 => x"2e",
          8535 => x"19",
          8536 => x"74",
          8537 => x"38",
          8538 => x"08",
          8539 => x"38",
          8540 => x"57",
          8541 => x"75",
          8542 => x"8e",
          8543 => x"75",
          8544 => x"f5",
          8545 => x"b9",
          8546 => x"b9",
          8547 => x"70",
          8548 => x"08",
          8549 => x"56",
          8550 => x"80",
          8551 => x"80",
          8552 => x"90",
          8553 => x"19",
          8554 => x"94",
          8555 => x"58",
          8556 => x"86",
          8557 => x"94",
          8558 => x"19",
          8559 => x"5a",
          8560 => x"34",
          8561 => x"84",
          8562 => x"8c",
          8563 => x"80",
          8564 => x"c8",
          8565 => x"0d",
          8566 => x"c8",
          8567 => x"da",
          8568 => x"2e",
          8569 => x"75",
          8570 => x"78",
          8571 => x"3f",
          8572 => x"08",
          8573 => x"39",
          8574 => x"08",
          8575 => x"0c",
          8576 => x"04",
          8577 => x"81",
          8578 => x"38",
          8579 => x"b6",
          8580 => x"0d",
          8581 => x"08",
          8582 => x"73",
          8583 => x"26",
          8584 => x"73",
          8585 => x"72",
          8586 => x"73",
          8587 => x"88",
          8588 => x"74",
          8589 => x"76",
          8590 => x"82",
          8591 => x"38",
          8592 => x"53",
          8593 => x"18",
          8594 => x"72",
          8595 => x"38",
          8596 => x"98",
          8597 => x"94",
          8598 => x"18",
          8599 => x"56",
          8600 => x"94",
          8601 => x"2a",
          8602 => x"0c",
          8603 => x"06",
          8604 => x"9c",
          8605 => x"56",
          8606 => x"c8",
          8607 => x"0d",
          8608 => x"84",
          8609 => x"8a",
          8610 => x"ac",
          8611 => x"74",
          8612 => x"ac",
          8613 => x"22",
          8614 => x"57",
          8615 => x"27",
          8616 => x"17",
          8617 => x"15",
          8618 => x"56",
          8619 => x"73",
          8620 => x"8a",
          8621 => x"71",
          8622 => x"08",
          8623 => x"78",
          8624 => x"ff",
          8625 => x"52",
          8626 => x"cd",
          8627 => x"c8",
          8628 => x"b9",
          8629 => x"2e",
          8630 => x"0b",
          8631 => x"08",
          8632 => x"38",
          8633 => x"53",
          8634 => x"08",
          8635 => x"91",
          8636 => x"31",
          8637 => x"27",
          8638 => x"aa",
          8639 => x"84",
          8640 => x"8a",
          8641 => x"f3",
          8642 => x"70",
          8643 => x"08",
          8644 => x"5a",
          8645 => x"0a",
          8646 => x"38",
          8647 => x"18",
          8648 => x"08",
          8649 => x"74",
          8650 => x"38",
          8651 => x"06",
          8652 => x"38",
          8653 => x"18",
          8654 => x"75",
          8655 => x"85",
          8656 => x"22",
          8657 => x"76",
          8658 => x"38",
          8659 => x"0c",
          8660 => x"0c",
          8661 => x"05",
          8662 => x"80",
          8663 => x"b9",
          8664 => x"3d",
          8665 => x"98",
          8666 => x"19",
          8667 => x"7a",
          8668 => x"5c",
          8669 => x"75",
          8670 => x"eb",
          8671 => x"b9",
          8672 => x"82",
          8673 => x"84",
          8674 => x"27",
          8675 => x"56",
          8676 => x"08",
          8677 => x"38",
          8678 => x"84",
          8679 => x"26",
          8680 => x"60",
          8681 => x"98",
          8682 => x"08",
          8683 => x"f9",
          8684 => x"b9",
          8685 => x"87",
          8686 => x"c8",
          8687 => x"ff",
          8688 => x"56",
          8689 => x"08",
          8690 => x"91",
          8691 => x"84",
          8692 => x"ff",
          8693 => x"38",
          8694 => x"08",
          8695 => x"5f",
          8696 => x"ea",
          8697 => x"9c",
          8698 => x"05",
          8699 => x"5c",
          8700 => x"8d",
          8701 => x"22",
          8702 => x"b0",
          8703 => x"5d",
          8704 => x"1a",
          8705 => x"58",
          8706 => x"57",
          8707 => x"70",
          8708 => x"34",
          8709 => x"74",
          8710 => x"56",
          8711 => x"55",
          8712 => x"81",
          8713 => x"54",
          8714 => x"77",
          8715 => x"33",
          8716 => x"3f",
          8717 => x"08",
          8718 => x"81",
          8719 => x"39",
          8720 => x"0c",
          8721 => x"b9",
          8722 => x"3d",
          8723 => x"54",
          8724 => x"53",
          8725 => x"53",
          8726 => x"52",
          8727 => x"3f",
          8728 => x"08",
          8729 => x"84",
          8730 => x"83",
          8731 => x"19",
          8732 => x"08",
          8733 => x"a0",
          8734 => x"fe",
          8735 => x"19",
          8736 => x"82",
          8737 => x"06",
          8738 => x"81",
          8739 => x"08",
          8740 => x"05",
          8741 => x"81",
          8742 => x"e3",
          8743 => x"c5",
          8744 => x"22",
          8745 => x"ff",
          8746 => x"74",
          8747 => x"81",
          8748 => x"7c",
          8749 => x"fe",
          8750 => x"08",
          8751 => x"56",
          8752 => x"7d",
          8753 => x"38",
          8754 => x"76",
          8755 => x"1b",
          8756 => x"19",
          8757 => x"f8",
          8758 => x"84",
          8759 => x"8f",
          8760 => x"ee",
          8761 => x"66",
          8762 => x"7c",
          8763 => x"81",
          8764 => x"1e",
          8765 => x"5e",
          8766 => x"82",
          8767 => x"19",
          8768 => x"80",
          8769 => x"08",
          8770 => x"d1",
          8771 => x"33",
          8772 => x"74",
          8773 => x"81",
          8774 => x"38",
          8775 => x"53",
          8776 => x"81",
          8777 => x"e1",
          8778 => x"b9",
          8779 => x"2e",
          8780 => x"5a",
          8781 => x"b4",
          8782 => x"5b",
          8783 => x"38",
          8784 => x"70",
          8785 => x"76",
          8786 => x"81",
          8787 => x"33",
          8788 => x"81",
          8789 => x"41",
          8790 => x"34",
          8791 => x"32",
          8792 => x"ae",
          8793 => x"72",
          8794 => x"80",
          8795 => x"45",
          8796 => x"74",
          8797 => x"7a",
          8798 => x"56",
          8799 => x"81",
          8800 => x"60",
          8801 => x"38",
          8802 => x"80",
          8803 => x"fa",
          8804 => x"b9",
          8805 => x"84",
          8806 => x"81",
          8807 => x"1c",
          8808 => x"fe",
          8809 => x"84",
          8810 => x"94",
          8811 => x"81",
          8812 => x"08",
          8813 => x"81",
          8814 => x"e1",
          8815 => x"57",
          8816 => x"08",
          8817 => x"81",
          8818 => x"38",
          8819 => x"08",
          8820 => x"b4",
          8821 => x"1a",
          8822 => x"b9",
          8823 => x"5b",
          8824 => x"08",
          8825 => x"38",
          8826 => x"41",
          8827 => x"09",
          8828 => x"a8",
          8829 => x"b4",
          8830 => x"1a",
          8831 => x"7e",
          8832 => x"33",
          8833 => x"3f",
          8834 => x"90",
          8835 => x"2e",
          8836 => x"81",
          8837 => x"86",
          8838 => x"5b",
          8839 => x"93",
          8840 => x"33",
          8841 => x"06",
          8842 => x"08",
          8843 => x"0c",
          8844 => x"76",
          8845 => x"38",
          8846 => x"74",
          8847 => x"39",
          8848 => x"60",
          8849 => x"06",
          8850 => x"c1",
          8851 => x"80",
          8852 => x"0c",
          8853 => x"c8",
          8854 => x"0d",
          8855 => x"fd",
          8856 => x"18",
          8857 => x"77",
          8858 => x"06",
          8859 => x"19",
          8860 => x"33",
          8861 => x"71",
          8862 => x"58",
          8863 => x"ff",
          8864 => x"33",
          8865 => x"06",
          8866 => x"05",
          8867 => x"76",
          8868 => x"e5",
          8869 => x"78",
          8870 => x"33",
          8871 => x"88",
          8872 => x"44",
          8873 => x"2e",
          8874 => x"79",
          8875 => x"ff",
          8876 => x"10",
          8877 => x"5c",
          8878 => x"23",
          8879 => x"81",
          8880 => x"77",
          8881 => x"77",
          8882 => x"2a",
          8883 => x"57",
          8884 => x"90",
          8885 => x"fe",
          8886 => x"38",
          8887 => x"05",
          8888 => x"23",
          8889 => x"81",
          8890 => x"41",
          8891 => x"75",
          8892 => x"2e",
          8893 => x"ff",
          8894 => x"39",
          8895 => x"7c",
          8896 => x"74",
          8897 => x"81",
          8898 => x"78",
          8899 => x"5a",
          8900 => x"05",
          8901 => x"06",
          8902 => x"56",
          8903 => x"38",
          8904 => x"fd",
          8905 => x"0b",
          8906 => x"7a",
          8907 => x"0c",
          8908 => x"04",
          8909 => x"63",
          8910 => x"5c",
          8911 => x"51",
          8912 => x"84",
          8913 => x"5a",
          8914 => x"08",
          8915 => x"81",
          8916 => x"5d",
          8917 => x"1d",
          8918 => x"5e",
          8919 => x"56",
          8920 => x"1b",
          8921 => x"82",
          8922 => x"1b",
          8923 => x"55",
          8924 => x"09",
          8925 => x"df",
          8926 => x"75",
          8927 => x"52",
          8928 => x"51",
          8929 => x"84",
          8930 => x"80",
          8931 => x"ff",
          8932 => x"75",
          8933 => x"76",
          8934 => x"b2",
          8935 => x"08",
          8936 => x"59",
          8937 => x"84",
          8938 => x"19",
          8939 => x"70",
          8940 => x"57",
          8941 => x"1d",
          8942 => x"e5",
          8943 => x"38",
          8944 => x"81",
          8945 => x"8f",
          8946 => x"38",
          8947 => x"38",
          8948 => x"81",
          8949 => x"aa",
          8950 => x"56",
          8951 => x"74",
          8952 => x"81",
          8953 => x"78",
          8954 => x"5a",
          8955 => x"05",
          8956 => x"06",
          8957 => x"56",
          8958 => x"38",
          8959 => x"80",
          8960 => x"1c",
          8961 => x"57",
          8962 => x"8b",
          8963 => x"59",
          8964 => x"81",
          8965 => x"78",
          8966 => x"5a",
          8967 => x"31",
          8968 => x"58",
          8969 => x"80",
          8970 => x"38",
          8971 => x"e1",
          8972 => x"5d",
          8973 => x"1d",
          8974 => x"7b",
          8975 => x"3f",
          8976 => x"08",
          8977 => x"c8",
          8978 => x"fe",
          8979 => x"84",
          8980 => x"93",
          8981 => x"81",
          8982 => x"08",
          8983 => x"81",
          8984 => x"dc",
          8985 => x"57",
          8986 => x"08",
          8987 => x"81",
          8988 => x"38",
          8989 => x"08",
          8990 => x"b4",
          8991 => x"1c",
          8992 => x"b9",
          8993 => x"59",
          8994 => x"08",
          8995 => x"38",
          8996 => x"5a",
          8997 => x"09",
          8998 => x"dd",
          8999 => x"b4",
          9000 => x"1c",
          9001 => x"7d",
          9002 => x"33",
          9003 => x"3f",
          9004 => x"c5",
          9005 => x"fd",
          9006 => x"1c",
          9007 => x"2a",
          9008 => x"55",
          9009 => x"38",
          9010 => x"81",
          9011 => x"80",
          9012 => x"8d",
          9013 => x"81",
          9014 => x"90",
          9015 => x"ac",
          9016 => x"5e",
          9017 => x"2e",
          9018 => x"ff",
          9019 => x"80",
          9020 => x"f4",
          9021 => x"b9",
          9022 => x"84",
          9023 => x"80",
          9024 => x"38",
          9025 => x"75",
          9026 => x"c2",
          9027 => x"5d",
          9028 => x"1d",
          9029 => x"39",
          9030 => x"57",
          9031 => x"09",
          9032 => x"38",
          9033 => x"9b",
          9034 => x"1b",
          9035 => x"2b",
          9036 => x"40",
          9037 => x"38",
          9038 => x"bf",
          9039 => x"f3",
          9040 => x"81",
          9041 => x"83",
          9042 => x"33",
          9043 => x"11",
          9044 => x"71",
          9045 => x"52",
          9046 => x"80",
          9047 => x"38",
          9048 => x"26",
          9049 => x"76",
          9050 => x"8a",
          9051 => x"c8",
          9052 => x"61",
          9053 => x"53",
          9054 => x"5b",
          9055 => x"f6",
          9056 => x"b9",
          9057 => x"09",
          9058 => x"de",
          9059 => x"81",
          9060 => x"78",
          9061 => x"38",
          9062 => x"86",
          9063 => x"56",
          9064 => x"2e",
          9065 => x"80",
          9066 => x"79",
          9067 => x"70",
          9068 => x"7f",
          9069 => x"ff",
          9070 => x"ff",
          9071 => x"fe",
          9072 => x"0b",
          9073 => x"0c",
          9074 => x"04",
          9075 => x"ff",
          9076 => x"38",
          9077 => x"fe",
          9078 => x"3d",
          9079 => x"08",
          9080 => x"33",
          9081 => x"58",
          9082 => x"86",
          9083 => x"b5",
          9084 => x"1d",
          9085 => x"57",
          9086 => x"80",
          9087 => x"81",
          9088 => x"17",
          9089 => x"56",
          9090 => x"38",
          9091 => x"1f",
          9092 => x"60",
          9093 => x"55",
          9094 => x"05",
          9095 => x"70",
          9096 => x"34",
          9097 => x"74",
          9098 => x"80",
          9099 => x"70",
          9100 => x"56",
          9101 => x"82",
          9102 => x"c0",
          9103 => x"34",
          9104 => x"3d",
          9105 => x"1c",
          9106 => x"59",
          9107 => x"5a",
          9108 => x"70",
          9109 => x"33",
          9110 => x"05",
          9111 => x"15",
          9112 => x"38",
          9113 => x"80",
          9114 => x"79",
          9115 => x"74",
          9116 => x"38",
          9117 => x"5a",
          9118 => x"75",
          9119 => x"10",
          9120 => x"2a",
          9121 => x"ff",
          9122 => x"2a",
          9123 => x"58",
          9124 => x"80",
          9125 => x"76",
          9126 => x"32",
          9127 => x"58",
          9128 => x"d7",
          9129 => x"55",
          9130 => x"87",
          9131 => x"80",
          9132 => x"58",
          9133 => x"bf",
          9134 => x"75",
          9135 => x"87",
          9136 => x"76",
          9137 => x"ff",
          9138 => x"2a",
          9139 => x"76",
          9140 => x"1f",
          9141 => x"79",
          9142 => x"58",
          9143 => x"27",
          9144 => x"33",
          9145 => x"2e",
          9146 => x"16",
          9147 => x"27",
          9148 => x"75",
          9149 => x"56",
          9150 => x"2e",
          9151 => x"ea",
          9152 => x"56",
          9153 => x"87",
          9154 => x"98",
          9155 => x"ec",
          9156 => x"71",
          9157 => x"41",
          9158 => x"87",
          9159 => x"f4",
          9160 => x"f8",
          9161 => x"b9",
          9162 => x"38",
          9163 => x"80",
          9164 => x"fe",
          9165 => x"56",
          9166 => x"2e",
          9167 => x"84",
          9168 => x"56",
          9169 => x"08",
          9170 => x"81",
          9171 => x"38",
          9172 => x"05",
          9173 => x"34",
          9174 => x"84",
          9175 => x"05",
          9176 => x"75",
          9177 => x"06",
          9178 => x"7e",
          9179 => x"38",
          9180 => x"1d",
          9181 => x"b0",
          9182 => x"c8",
          9183 => x"80",
          9184 => x"ed",
          9185 => x"b9",
          9186 => x"84",
          9187 => x"81",
          9188 => x"b9",
          9189 => x"19",
          9190 => x"1e",
          9191 => x"57",
          9192 => x"76",
          9193 => x"38",
          9194 => x"40",
          9195 => x"09",
          9196 => x"a3",
          9197 => x"75",
          9198 => x"52",
          9199 => x"51",
          9200 => x"84",
          9201 => x"80",
          9202 => x"ff",
          9203 => x"75",
          9204 => x"76",
          9205 => x"38",
          9206 => x"70",
          9207 => x"74",
          9208 => x"81",
          9209 => x"30",
          9210 => x"78",
          9211 => x"74",
          9212 => x"c9",
          9213 => x"59",
          9214 => x"86",
          9215 => x"52",
          9216 => x"83",
          9217 => x"c8",
          9218 => x"b9",
          9219 => x"2e",
          9220 => x"87",
          9221 => x"2e",
          9222 => x"75",
          9223 => x"83",
          9224 => x"40",
          9225 => x"38",
          9226 => x"57",
          9227 => x"77",
          9228 => x"83",
          9229 => x"57",
          9230 => x"82",
          9231 => x"76",
          9232 => x"52",
          9233 => x"51",
          9234 => x"84",
          9235 => x"80",
          9236 => x"ff",
          9237 => x"76",
          9238 => x"75",
          9239 => x"c3",
          9240 => x"9c",
          9241 => x"55",
          9242 => x"81",
          9243 => x"ff",
          9244 => x"f4",
          9245 => x"9c",
          9246 => x"58",
          9247 => x"70",
          9248 => x"33",
          9249 => x"05",
          9250 => x"15",
          9251 => x"38",
          9252 => x"ab",
          9253 => x"06",
          9254 => x"8c",
          9255 => x"0b",
          9256 => x"77",
          9257 => x"b9",
          9258 => x"3d",
          9259 => x"75",
          9260 => x"25",
          9261 => x"40",
          9262 => x"b9",
          9263 => x"81",
          9264 => x"ec",
          9265 => x"b9",
          9266 => x"84",
          9267 => x"80",
          9268 => x"38",
          9269 => x"81",
          9270 => x"08",
          9271 => x"81",
          9272 => x"d3",
          9273 => x"b9",
          9274 => x"2e",
          9275 => x"83",
          9276 => x"b9",
          9277 => x"19",
          9278 => x"08",
          9279 => x"31",
          9280 => x"19",
          9281 => x"38",
          9282 => x"41",
          9283 => x"84",
          9284 => x"b9",
          9285 => x"fd",
          9286 => x"85",
          9287 => x"08",
          9288 => x"58",
          9289 => x"e9",
          9290 => x"c8",
          9291 => x"b9",
          9292 => x"ef",
          9293 => x"b9",
          9294 => x"58",
          9295 => x"81",
          9296 => x"80",
          9297 => x"70",
          9298 => x"33",
          9299 => x"70",
          9300 => x"ff",
          9301 => x"5d",
          9302 => x"74",
          9303 => x"b8",
          9304 => x"98",
          9305 => x"80",
          9306 => x"08",
          9307 => x"38",
          9308 => x"5b",
          9309 => x"09",
          9310 => x"c9",
          9311 => x"76",
          9312 => x"52",
          9313 => x"51",
          9314 => x"84",
          9315 => x"80",
          9316 => x"ff",
          9317 => x"76",
          9318 => x"75",
          9319 => x"83",
          9320 => x"08",
          9321 => x"61",
          9322 => x"5f",
          9323 => x"8d",
          9324 => x"0b",
          9325 => x"75",
          9326 => x"75",
          9327 => x"75",
          9328 => x"7c",
          9329 => x"05",
          9330 => x"58",
          9331 => x"ff",
          9332 => x"38",
          9333 => x"70",
          9334 => x"5b",
          9335 => x"e5",
          9336 => x"7b",
          9337 => x"75",
          9338 => x"57",
          9339 => x"2a",
          9340 => x"34",
          9341 => x"83",
          9342 => x"81",
          9343 => x"78",
          9344 => x"76",
          9345 => x"2e",
          9346 => x"78",
          9347 => x"22",
          9348 => x"80",
          9349 => x"38",
          9350 => x"81",
          9351 => x"34",
          9352 => x"51",
          9353 => x"84",
          9354 => x"58",
          9355 => x"08",
          9356 => x"7f",
          9357 => x"7f",
          9358 => x"fb",
          9359 => x"54",
          9360 => x"53",
          9361 => x"53",
          9362 => x"52",
          9363 => x"3f",
          9364 => x"b9",
          9365 => x"83",
          9366 => x"c8",
          9367 => x"34",
          9368 => x"a8",
          9369 => x"84",
          9370 => x"57",
          9371 => x"1d",
          9372 => x"c9",
          9373 => x"33",
          9374 => x"2e",
          9375 => x"fb",
          9376 => x"54",
          9377 => x"a0",
          9378 => x"53",
          9379 => x"1c",
          9380 => x"d1",
          9381 => x"fb",
          9382 => x"9c",
          9383 => x"33",
          9384 => x"74",
          9385 => x"09",
          9386 => x"ba",
          9387 => x"39",
          9388 => x"57",
          9389 => x"fa",
          9390 => x"d7",
          9391 => x"c0",
          9392 => x"d4",
          9393 => x"b4",
          9394 => x"61",
          9395 => x"33",
          9396 => x"3f",
          9397 => x"08",
          9398 => x"81",
          9399 => x"84",
          9400 => x"83",
          9401 => x"1c",
          9402 => x"08",
          9403 => x"a0",
          9404 => x"8a",
          9405 => x"33",
          9406 => x"2e",
          9407 => x"b9",
          9408 => x"fc",
          9409 => x"ff",
          9410 => x"7f",
          9411 => x"98",
          9412 => x"39",
          9413 => x"f7",
          9414 => x"70",
          9415 => x"80",
          9416 => x"38",
          9417 => x"81",
          9418 => x"08",
          9419 => x"05",
          9420 => x"81",
          9421 => x"ce",
          9422 => x"c1",
          9423 => x"b4",
          9424 => x"19",
          9425 => x"7c",
          9426 => x"33",
          9427 => x"3f",
          9428 => x"f3",
          9429 => x"61",
          9430 => x"5e",
          9431 => x"96",
          9432 => x"1c",
          9433 => x"82",
          9434 => x"1c",
          9435 => x"80",
          9436 => x"70",
          9437 => x"05",
          9438 => x"57",
          9439 => x"58",
          9440 => x"bc",
          9441 => x"74",
          9442 => x"81",
          9443 => x"56",
          9444 => x"38",
          9445 => x"14",
          9446 => x"ff",
          9447 => x"76",
          9448 => x"82",
          9449 => x"79",
          9450 => x"70",
          9451 => x"55",
          9452 => x"38",
          9453 => x"80",
          9454 => x"7a",
          9455 => x"5e",
          9456 => x"05",
          9457 => x"82",
          9458 => x"70",
          9459 => x"57",
          9460 => x"08",
          9461 => x"81",
          9462 => x"53",
          9463 => x"b2",
          9464 => x"2e",
          9465 => x"75",
          9466 => x"30",
          9467 => x"80",
          9468 => x"54",
          9469 => x"90",
          9470 => x"2e",
          9471 => x"77",
          9472 => x"59",
          9473 => x"58",
          9474 => x"81",
          9475 => x"81",
          9476 => x"76",
          9477 => x"38",
          9478 => x"05",
          9479 => x"81",
          9480 => x"1d",
          9481 => x"a5",
          9482 => x"f3",
          9483 => x"96",
          9484 => x"57",
          9485 => x"05",
          9486 => x"82",
          9487 => x"1c",
          9488 => x"33",
          9489 => x"89",
          9490 => x"1e",
          9491 => x"08",
          9492 => x"33",
          9493 => x"9c",
          9494 => x"11",
          9495 => x"82",
          9496 => x"90",
          9497 => x"2b",
          9498 => x"33",
          9499 => x"88",
          9500 => x"71",
          9501 => x"59",
          9502 => x"96",
          9503 => x"88",
          9504 => x"41",
          9505 => x"56",
          9506 => x"86",
          9507 => x"15",
          9508 => x"33",
          9509 => x"07",
          9510 => x"84",
          9511 => x"3d",
          9512 => x"e5",
          9513 => x"39",
          9514 => x"11",
          9515 => x"31",
          9516 => x"83",
          9517 => x"90",
          9518 => x"51",
          9519 => x"3f",
          9520 => x"08",
          9521 => x"06",
          9522 => x"75",
          9523 => x"81",
          9524 => x"b3",
          9525 => x"2a",
          9526 => x"34",
          9527 => x"34",
          9528 => x"58",
          9529 => x"1f",
          9530 => x"78",
          9531 => x"70",
          9532 => x"54",
          9533 => x"38",
          9534 => x"74",
          9535 => x"70",
          9536 => x"25",
          9537 => x"07",
          9538 => x"75",
          9539 => x"74",
          9540 => x"78",
          9541 => x"0b",
          9542 => x"56",
          9543 => x"72",
          9544 => x"33",
          9545 => x"77",
          9546 => x"88",
          9547 => x"1e",
          9548 => x"54",
          9549 => x"ff",
          9550 => x"54",
          9551 => x"a4",
          9552 => x"08",
          9553 => x"54",
          9554 => x"27",
          9555 => x"84",
          9556 => x"81",
          9557 => x"80",
          9558 => x"a0",
          9559 => x"ff",
          9560 => x"53",
          9561 => x"81",
          9562 => x"81",
          9563 => x"81",
          9564 => x"13",
          9565 => x"59",
          9566 => x"ff",
          9567 => x"b4",
          9568 => x"2a",
          9569 => x"80",
          9570 => x"80",
          9571 => x"73",
          9572 => x"5f",
          9573 => x"39",
          9574 => x"63",
          9575 => x"42",
          9576 => x"65",
          9577 => x"55",
          9578 => x"2e",
          9579 => x"53",
          9580 => x"2e",
          9581 => x"72",
          9582 => x"d9",
          9583 => x"08",
          9584 => x"73",
          9585 => x"94",
          9586 => x"55",
          9587 => x"82",
          9588 => x"42",
          9589 => x"58",
          9590 => x"70",
          9591 => x"52",
          9592 => x"73",
          9593 => x"72",
          9594 => x"ff",
          9595 => x"38",
          9596 => x"74",
          9597 => x"76",
          9598 => x"80",
          9599 => x"17",
          9600 => x"ff",
          9601 => x"af",
          9602 => x"9f",
          9603 => x"80",
          9604 => x"5b",
          9605 => x"82",
          9606 => x"80",
          9607 => x"89",
          9608 => x"ff",
          9609 => x"83",
          9610 => x"83",
          9611 => x"70",
          9612 => x"56",
          9613 => x"80",
          9614 => x"38",
          9615 => x"8f",
          9616 => x"70",
          9617 => x"ff",
          9618 => x"56",
          9619 => x"72",
          9620 => x"5b",
          9621 => x"38",
          9622 => x"26",
          9623 => x"76",
          9624 => x"74",
          9625 => x"17",
          9626 => x"81",
          9627 => x"56",
          9628 => x"80",
          9629 => x"38",
          9630 => x"81",
          9631 => x"32",
          9632 => x"80",
          9633 => x"51",
          9634 => x"72",
          9635 => x"38",
          9636 => x"46",
          9637 => x"33",
          9638 => x"af",
          9639 => x"72",
          9640 => x"70",
          9641 => x"25",
          9642 => x"54",
          9643 => x"38",
          9644 => x"0c",
          9645 => x"3d",
          9646 => x"42",
          9647 => x"26",
          9648 => x"b4",
          9649 => x"52",
          9650 => x"8d",
          9651 => x"b9",
          9652 => x"ff",
          9653 => x"73",
          9654 => x"86",
          9655 => x"b9",
          9656 => x"3d",
          9657 => x"e4",
          9658 => x"81",
          9659 => x"53",
          9660 => x"fe",
          9661 => x"39",
          9662 => x"ab",
          9663 => x"52",
          9664 => x"8d",
          9665 => x"c8",
          9666 => x"c8",
          9667 => x"0d",
          9668 => x"80",
          9669 => x"30",
          9670 => x"73",
          9671 => x"5a",
          9672 => x"2e",
          9673 => x"14",
          9674 => x"70",
          9675 => x"56",
          9676 => x"dd",
          9677 => x"dc",
          9678 => x"70",
          9679 => x"07",
          9680 => x"7d",
          9681 => x"61",
          9682 => x"27",
          9683 => x"76",
          9684 => x"f8",
          9685 => x"2e",
          9686 => x"76",
          9687 => x"80",
          9688 => x"76",
          9689 => x"fe",
          9690 => x"70",
          9691 => x"30",
          9692 => x"52",
          9693 => x"56",
          9694 => x"2e",
          9695 => x"89",
          9696 => x"57",
          9697 => x"76",
          9698 => x"56",
          9699 => x"76",
          9700 => x"c7",
          9701 => x"22",
          9702 => x"ff",
          9703 => x"5d",
          9704 => x"a0",
          9705 => x"38",
          9706 => x"ff",
          9707 => x"ae",
          9708 => x"38",
          9709 => x"aa",
          9710 => x"fe",
          9711 => x"5a",
          9712 => x"2e",
          9713 => x"10",
          9714 => x"54",
          9715 => x"76",
          9716 => x"38",
          9717 => x"22",
          9718 => x"ae",
          9719 => x"06",
          9720 => x"0b",
          9721 => x"53",
          9722 => x"81",
          9723 => x"ff",
          9724 => x"f4",
          9725 => x"5c",
          9726 => x"16",
          9727 => x"19",
          9728 => x"5d",
          9729 => x"80",
          9730 => x"a0",
          9731 => x"38",
          9732 => x"70",
          9733 => x"25",
          9734 => x"75",
          9735 => x"ce",
          9736 => x"bb",
          9737 => x"7c",
          9738 => x"38",
          9739 => x"77",
          9740 => x"70",
          9741 => x"25",
          9742 => x"51",
          9743 => x"72",
          9744 => x"e0",
          9745 => x"2e",
          9746 => x"75",
          9747 => x"38",
          9748 => x"5a",
          9749 => x"9e",
          9750 => x"88",
          9751 => x"82",
          9752 => x"06",
          9753 => x"5f",
          9754 => x"70",
          9755 => x"58",
          9756 => x"ff",
          9757 => x"1c",
          9758 => x"81",
          9759 => x"84",
          9760 => x"2e",
          9761 => x"7d",
          9762 => x"77",
          9763 => x"ed",
          9764 => x"06",
          9765 => x"2e",
          9766 => x"79",
          9767 => x"06",
          9768 => x"38",
          9769 => x"5d",
          9770 => x"85",
          9771 => x"07",
          9772 => x"2a",
          9773 => x"7d",
          9774 => x"38",
          9775 => x"5a",
          9776 => x"34",
          9777 => x"ec",
          9778 => x"c8",
          9779 => x"33",
          9780 => x"b9",
          9781 => x"2e",
          9782 => x"84",
          9783 => x"84",
          9784 => x"06",
          9785 => x"74",
          9786 => x"06",
          9787 => x"2e",
          9788 => x"74",
          9789 => x"06",
          9790 => x"98",
          9791 => x"65",
          9792 => x"42",
          9793 => x"58",
          9794 => x"ce",
          9795 => x"70",
          9796 => x"70",
          9797 => x"56",
          9798 => x"2e",
          9799 => x"80",
          9800 => x"38",
          9801 => x"5a",
          9802 => x"82",
          9803 => x"75",
          9804 => x"81",
          9805 => x"38",
          9806 => x"73",
          9807 => x"81",
          9808 => x"38",
          9809 => x"5b",
          9810 => x"80",
          9811 => x"56",
          9812 => x"76",
          9813 => x"38",
          9814 => x"75",
          9815 => x"57",
          9816 => x"53",
          9817 => x"e9",
          9818 => x"07",
          9819 => x"1d",
          9820 => x"e3",
          9821 => x"b9",
          9822 => x"1d",
          9823 => x"84",
          9824 => x"fe",
          9825 => x"82",
          9826 => x"58",
          9827 => x"38",
          9828 => x"70",
          9829 => x"06",
          9830 => x"80",
          9831 => x"38",
          9832 => x"83",
          9833 => x"05",
          9834 => x"33",
          9835 => x"33",
          9836 => x"07",
          9837 => x"57",
          9838 => x"83",
          9839 => x"38",
          9840 => x"0c",
          9841 => x"55",
          9842 => x"39",
          9843 => x"74",
          9844 => x"f0",
          9845 => x"59",
          9846 => x"38",
          9847 => x"79",
          9848 => x"17",
          9849 => x"81",
          9850 => x"2b",
          9851 => x"70",
          9852 => x"5e",
          9853 => x"09",
          9854 => x"95",
          9855 => x"07",
          9856 => x"39",
          9857 => x"1d",
          9858 => x"2e",
          9859 => x"fc",
          9860 => x"39",
          9861 => x"ab",
          9862 => x"0b",
          9863 => x"0c",
          9864 => x"04",
          9865 => x"26",
          9866 => x"ff",
          9867 => x"c9",
          9868 => x"59",
          9869 => x"81",
          9870 => x"83",
          9871 => x"18",
          9872 => x"fc",
          9873 => x"82",
          9874 => x"b5",
          9875 => x"81",
          9876 => x"84",
          9877 => x"83",
          9878 => x"70",
          9879 => x"06",
          9880 => x"80",
          9881 => x"74",
          9882 => x"83",
          9883 => x"33",
          9884 => x"81",
          9885 => x"b9",
          9886 => x"2e",
          9887 => x"83",
          9888 => x"83",
          9889 => x"70",
          9890 => x"56",
          9891 => x"80",
          9892 => x"38",
          9893 => x"8f",
          9894 => x"70",
          9895 => x"ff",
          9896 => x"59",
          9897 => x"72",
          9898 => x"59",
          9899 => x"38",
          9900 => x"54",
          9901 => x"8a",
          9902 => x"07",
          9903 => x"06",
          9904 => x"9f",
          9905 => x"99",
          9906 => x"7d",
          9907 => x"81",
          9908 => x"17",
          9909 => x"ff",
          9910 => x"5f",
          9911 => x"a0",
          9912 => x"79",
          9913 => x"5b",
          9914 => x"fa",
          9915 => x"53",
          9916 => x"83",
          9917 => x"70",
          9918 => x"5a",
          9919 => x"2e",
          9920 => x"80",
          9921 => x"07",
          9922 => x"05",
          9923 => x"74",
          9924 => x"1b",
          9925 => x"80",
          9926 => x"80",
          9927 => x"71",
          9928 => x"90",
          9929 => x"07",
          9930 => x"5a",
          9931 => x"39",
          9932 => x"05",
          9933 => x"54",
          9934 => x"34",
          9935 => x"11",
          9936 => x"5b",
          9937 => x"81",
          9938 => x"9c",
          9939 => x"07",
          9940 => x"58",
          9941 => x"e5",
          9942 => x"06",
          9943 => x"fd",
          9944 => x"82",
          9945 => x"5c",
          9946 => x"38",
          9947 => x"b9",
          9948 => x"3d",
          9949 => x"3d",
          9950 => x"02",
          9951 => x"e7",
          9952 => x"42",
          9953 => x"0c",
          9954 => x"70",
          9955 => x"79",
          9956 => x"d7",
          9957 => x"81",
          9958 => x"70",
          9959 => x"56",
          9960 => x"85",
          9961 => x"ed",
          9962 => x"2e",
          9963 => x"84",
          9964 => x"56",
          9965 => x"85",
          9966 => x"10",
          9967 => x"90",
          9968 => x"58",
          9969 => x"76",
          9970 => x"96",
          9971 => x"0c",
          9972 => x"06",
          9973 => x"59",
          9974 => x"9b",
          9975 => x"33",
          9976 => x"b0",
          9977 => x"c8",
          9978 => x"06",
          9979 => x"5e",
          9980 => x"2e",
          9981 => x"80",
          9982 => x"16",
          9983 => x"bc",
          9984 => x"18",
          9985 => x"81",
          9986 => x"ff",
          9987 => x"84",
          9988 => x"81",
          9989 => x"81",
          9990 => x"83",
          9991 => x"c2",
          9992 => x"2e",
          9993 => x"82",
          9994 => x"41",
          9995 => x"84",
          9996 => x"5b",
          9997 => x"34",
          9998 => x"18",
          9999 => x"5a",
         10000 => x"7a",
         10001 => x"70",
         10002 => x"33",
         10003 => x"bb",
         10004 => x"b9",
         10005 => x"2e",
         10006 => x"55",
         10007 => x"b4",
         10008 => x"56",
         10009 => x"84",
         10010 => x"84",
         10011 => x"71",
         10012 => x"56",
         10013 => x"74",
         10014 => x"2e",
         10015 => x"75",
         10016 => x"38",
         10017 => x"1d",
         10018 => x"85",
         10019 => x"58",
         10020 => x"83",
         10021 => x"58",
         10022 => x"83",
         10023 => x"c4",
         10024 => x"c3",
         10025 => x"88",
         10026 => x"59",
         10027 => x"2e",
         10028 => x"83",
         10029 => x"cf",
         10030 => x"ce",
         10031 => x"88",
         10032 => x"5a",
         10033 => x"80",
         10034 => x"11",
         10035 => x"33",
         10036 => x"71",
         10037 => x"81",
         10038 => x"72",
         10039 => x"75",
         10040 => x"56",
         10041 => x"5e",
         10042 => x"a0",
         10043 => x"c8",
         10044 => x"18",
         10045 => x"17",
         10046 => x"70",
         10047 => x"5f",
         10048 => x"58",
         10049 => x"82",
         10050 => x"81",
         10051 => x"71",
         10052 => x"19",
         10053 => x"5a",
         10054 => x"23",
         10055 => x"80",
         10056 => x"38",
         10057 => x"06",
         10058 => x"bb",
         10059 => x"17",
         10060 => x"18",
         10061 => x"2b",
         10062 => x"74",
         10063 => x"74",
         10064 => x"5e",
         10065 => x"7c",
         10066 => x"80",
         10067 => x"80",
         10068 => x"71",
         10069 => x"56",
         10070 => x"38",
         10071 => x"83",
         10072 => x"12",
         10073 => x"2b",
         10074 => x"07",
         10075 => x"70",
         10076 => x"2b",
         10077 => x"07",
         10078 => x"58",
         10079 => x"80",
         10080 => x"80",
         10081 => x"71",
         10082 => x"5d",
         10083 => x"7b",
         10084 => x"ce",
         10085 => x"7a",
         10086 => x"5a",
         10087 => x"81",
         10088 => x"52",
         10089 => x"51",
         10090 => x"3f",
         10091 => x"08",
         10092 => x"c8",
         10093 => x"81",
         10094 => x"b9",
         10095 => x"ff",
         10096 => x"26",
         10097 => x"5d",
         10098 => x"f5",
         10099 => x"82",
         10100 => x"f5",
         10101 => x"38",
         10102 => x"16",
         10103 => x"0c",
         10104 => x"0c",
         10105 => x"a8",
         10106 => x"1d",
         10107 => x"57",
         10108 => x"2e",
         10109 => x"88",
         10110 => x"8d",
         10111 => x"2e",
         10112 => x"7d",
         10113 => x"0c",
         10114 => x"7c",
         10115 => x"38",
         10116 => x"70",
         10117 => x"81",
         10118 => x"5a",
         10119 => x"89",
         10120 => x"58",
         10121 => x"08",
         10122 => x"ff",
         10123 => x"0c",
         10124 => x"18",
         10125 => x"0b",
         10126 => x"7c",
         10127 => x"96",
         10128 => x"34",
         10129 => x"22",
         10130 => x"7c",
         10131 => x"23",
         10132 => x"23",
         10133 => x"0b",
         10134 => x"80",
         10135 => x"0c",
         10136 => x"84",
         10137 => x"97",
         10138 => x"8b",
         10139 => x"c8",
         10140 => x"0d",
         10141 => x"d0",
         10142 => x"ff",
         10143 => x"58",
         10144 => x"91",
         10145 => x"78",
         10146 => x"d0",
         10147 => x"78",
         10148 => x"fe",
         10149 => x"08",
         10150 => x"5f",
         10151 => x"08",
         10152 => x"7a",
         10153 => x"5c",
         10154 => x"81",
         10155 => x"ff",
         10156 => x"58",
         10157 => x"26",
         10158 => x"16",
         10159 => x"06",
         10160 => x"9f",
         10161 => x"99",
         10162 => x"e0",
         10163 => x"ff",
         10164 => x"75",
         10165 => x"2a",
         10166 => x"77",
         10167 => x"06",
         10168 => x"ff",
         10169 => x"7a",
         10170 => x"70",
         10171 => x"2a",
         10172 => x"58",
         10173 => x"2e",
         10174 => x"81",
         10175 => x"5e",
         10176 => x"25",
         10177 => x"61",
         10178 => x"39",
         10179 => x"fe",
         10180 => x"82",
         10181 => x"5e",
         10182 => x"fe",
         10183 => x"58",
         10184 => x"7a",
         10185 => x"59",
         10186 => x"2e",
         10187 => x"83",
         10188 => x"75",
         10189 => x"70",
         10190 => x"25",
         10191 => x"5b",
         10192 => x"ad",
         10193 => x"e8",
         10194 => x"38",
         10195 => x"57",
         10196 => x"83",
         10197 => x"70",
         10198 => x"80",
         10199 => x"84",
         10200 => x"84",
         10201 => x"71",
         10202 => x"88",
         10203 => x"ff",
         10204 => x"72",
         10205 => x"83",
         10206 => x"71",
         10207 => x"5b",
         10208 => x"77",
         10209 => x"05",
         10210 => x"19",
         10211 => x"59",
         10212 => x"ff",
         10213 => x"b9",
         10214 => x"70",
         10215 => x"2a",
         10216 => x"9b",
         10217 => x"10",
         10218 => x"84",
         10219 => x"5d",
         10220 => x"42",
         10221 => x"83",
         10222 => x"2e",
         10223 => x"80",
         10224 => x"34",
         10225 => x"18",
         10226 => x"80",
         10227 => x"2e",
         10228 => x"54",
         10229 => x"17",
         10230 => x"33",
         10231 => x"86",
         10232 => x"c8",
         10233 => x"85",
         10234 => x"81",
         10235 => x"18",
         10236 => x"75",
         10237 => x"1f",
         10238 => x"71",
         10239 => x"5d",
         10240 => x"7b",
         10241 => x"2e",
         10242 => x"a8",
         10243 => x"b8",
         10244 => x"58",
         10245 => x"2e",
         10246 => x"75",
         10247 => x"70",
         10248 => x"25",
         10249 => x"42",
         10250 => x"38",
         10251 => x"2e",
         10252 => x"58",
         10253 => x"06",
         10254 => x"84",
         10255 => x"33",
         10256 => x"78",
         10257 => x"06",
         10258 => x"58",
         10259 => x"f8",
         10260 => x"80",
         10261 => x"38",
         10262 => x"1a",
         10263 => x"7a",
         10264 => x"38",
         10265 => x"83",
         10266 => x"18",
         10267 => x"40",
         10268 => x"70",
         10269 => x"33",
         10270 => x"05",
         10271 => x"71",
         10272 => x"5b",
         10273 => x"77",
         10274 => x"c5",
         10275 => x"2e",
         10276 => x"0b",
         10277 => x"83",
         10278 => x"5d",
         10279 => x"81",
         10280 => x"7e",
         10281 => x"40",
         10282 => x"31",
         10283 => x"58",
         10284 => x"80",
         10285 => x"38",
         10286 => x"e1",
         10287 => x"fe",
         10288 => x"58",
         10289 => x"38",
         10290 => x"c8",
         10291 => x"0d",
         10292 => x"75",
         10293 => x"dc",
         10294 => x"81",
         10295 => x"e4",
         10296 => x"58",
         10297 => x"8d",
         10298 => x"c8",
         10299 => x"0d",
         10300 => x"80",
         10301 => x"e4",
         10302 => x"58",
         10303 => x"05",
         10304 => x"70",
         10305 => x"33",
         10306 => x"ff",
         10307 => x"5f",
         10308 => x"2e",
         10309 => x"74",
         10310 => x"38",
         10311 => x"8a",
         10312 => x"fc",
         10313 => x"78",
         10314 => x"5a",
         10315 => x"81",
         10316 => x"71",
         10317 => x"1b",
         10318 => x"40",
         10319 => x"84",
         10320 => x"80",
         10321 => x"93",
         10322 => x"5a",
         10323 => x"83",
         10324 => x"fd",
         10325 => x"e9",
         10326 => x"e8",
         10327 => x"88",
         10328 => x"55",
         10329 => x"09",
         10330 => x"d5",
         10331 => x"58",
         10332 => x"17",
         10333 => x"b1",
         10334 => x"33",
         10335 => x"2e",
         10336 => x"82",
         10337 => x"54",
         10338 => x"17",
         10339 => x"33",
         10340 => x"d2",
         10341 => x"c8",
         10342 => x"85",
         10343 => x"81",
         10344 => x"18",
         10345 => x"99",
         10346 => x"18",
         10347 => x"17",
         10348 => x"18",
         10349 => x"2b",
         10350 => x"75",
         10351 => x"2e",
         10352 => x"f8",
         10353 => x"17",
         10354 => x"82",
         10355 => x"90",
         10356 => x"2b",
         10357 => x"33",
         10358 => x"88",
         10359 => x"71",
         10360 => x"59",
         10361 => x"59",
         10362 => x"85",
         10363 => x"09",
         10364 => x"cd",
         10365 => x"17",
         10366 => x"82",
         10367 => x"90",
         10368 => x"2b",
         10369 => x"33",
         10370 => x"88",
         10371 => x"71",
         10372 => x"40",
         10373 => x"5e",
         10374 => x"85",
         10375 => x"09",
         10376 => x"9d",
         10377 => x"17",
         10378 => x"82",
         10379 => x"90",
         10380 => x"2b",
         10381 => x"33",
         10382 => x"88",
         10383 => x"71",
         10384 => x"0c",
         10385 => x"1c",
         10386 => x"82",
         10387 => x"90",
         10388 => x"2b",
         10389 => x"33",
         10390 => x"88",
         10391 => x"71",
         10392 => x"05",
         10393 => x"49",
         10394 => x"40",
         10395 => x"5a",
         10396 => x"84",
         10397 => x"81",
         10398 => x"84",
         10399 => x"7c",
         10400 => x"84",
         10401 => x"8c",
         10402 => x"0b",
         10403 => x"f7",
         10404 => x"83",
         10405 => x"38",
         10406 => x"0c",
         10407 => x"39",
         10408 => x"17",
         10409 => x"17",
         10410 => x"18",
         10411 => x"ff",
         10412 => x"84",
         10413 => x"7a",
         10414 => x"06",
         10415 => x"84",
         10416 => x"83",
         10417 => x"17",
         10418 => x"08",
         10419 => x"a0",
         10420 => x"8b",
         10421 => x"33",
         10422 => x"2e",
         10423 => x"84",
         10424 => x"5a",
         10425 => x"74",
         10426 => x"2e",
         10427 => x"85",
         10428 => x"18",
         10429 => x"5c",
         10430 => x"ab",
         10431 => x"17",
         10432 => x"18",
         10433 => x"2b",
         10434 => x"8d",
         10435 => x"d2",
         10436 => x"22",
         10437 => x"ca",
         10438 => x"17",
         10439 => x"82",
         10440 => x"90",
         10441 => x"2b",
         10442 => x"33",
         10443 => x"88",
         10444 => x"71",
         10445 => x"0c",
         10446 => x"2b",
         10447 => x"40",
         10448 => x"d8",
         10449 => x"75",
         10450 => x"e8",
         10451 => x"f9",
         10452 => x"80",
         10453 => x"38",
         10454 => x"57",
         10455 => x"f7",
         10456 => x"5a",
         10457 => x"38",
         10458 => x"75",
         10459 => x"08",
         10460 => x"05",
         10461 => x"81",
         10462 => x"ff",
         10463 => x"fc",
         10464 => x"3d",
         10465 => x"d3",
         10466 => x"70",
         10467 => x"41",
         10468 => x"76",
         10469 => x"80",
         10470 => x"38",
         10471 => x"05",
         10472 => x"9f",
         10473 => x"74",
         10474 => x"e2",
         10475 => x"38",
         10476 => x"80",
         10477 => x"d1",
         10478 => x"80",
         10479 => x"c4",
         10480 => x"10",
         10481 => x"05",
         10482 => x"55",
         10483 => x"84",
         10484 => x"34",
         10485 => x"80",
         10486 => x"80",
         10487 => x"54",
         10488 => x"7c",
         10489 => x"2e",
         10490 => x"53",
         10491 => x"53",
         10492 => x"ef",
         10493 => x"b9",
         10494 => x"73",
         10495 => x"0c",
         10496 => x"04",
         10497 => x"b9",
         10498 => x"3d",
         10499 => x"33",
         10500 => x"81",
         10501 => x"56",
         10502 => x"26",
         10503 => x"16",
         10504 => x"06",
         10505 => x"58",
         10506 => x"80",
         10507 => x"7f",
         10508 => x"b8",
         10509 => x"7b",
         10510 => x"5a",
         10511 => x"05",
         10512 => x"70",
         10513 => x"33",
         10514 => x"59",
         10515 => x"99",
         10516 => x"e0",
         10517 => x"ff",
         10518 => x"ff",
         10519 => x"76",
         10520 => x"38",
         10521 => x"81",
         10522 => x"54",
         10523 => x"9f",
         10524 => x"74",
         10525 => x"81",
         10526 => x"76",
         10527 => x"77",
         10528 => x"30",
         10529 => x"9f",
         10530 => x"5c",
         10531 => x"80",
         10532 => x"81",
         10533 => x"5d",
         10534 => x"25",
         10535 => x"7f",
         10536 => x"39",
         10537 => x"f7",
         10538 => x"60",
         10539 => x"8b",
         10540 => x"0d",
         10541 => x"05",
         10542 => x"33",
         10543 => x"56",
         10544 => x"a6",
         10545 => x"06",
         10546 => x"3d",
         10547 => x"9e",
         10548 => x"52",
         10549 => x"3f",
         10550 => x"08",
         10551 => x"c8",
         10552 => x"8f",
         10553 => x"0c",
         10554 => x"84",
         10555 => x"9c",
         10556 => x"7e",
         10557 => x"90",
         10558 => x"5a",
         10559 => x"84",
         10560 => x"57",
         10561 => x"08",
         10562 => x"ba",
         10563 => x"06",
         10564 => x"2e",
         10565 => x"76",
         10566 => x"c1",
         10567 => x"2e",
         10568 => x"77",
         10569 => x"76",
         10570 => x"77",
         10571 => x"06",
         10572 => x"2e",
         10573 => x"66",
         10574 => x"9a",
         10575 => x"88",
         10576 => x"70",
         10577 => x"5e",
         10578 => x"83",
         10579 => x"38",
         10580 => x"17",
         10581 => x"8f",
         10582 => x"0b",
         10583 => x"80",
         10584 => x"17",
         10585 => x"a0",
         10586 => x"34",
         10587 => x"5e",
         10588 => x"17",
         10589 => x"9b",
         10590 => x"33",
         10591 => x"2e",
         10592 => x"66",
         10593 => x"9c",
         10594 => x"0b",
         10595 => x"80",
         10596 => x"34",
         10597 => x"1c",
         10598 => x"81",
         10599 => x"34",
         10600 => x"80",
         10601 => x"b4",
         10602 => x"7c",
         10603 => x"5f",
         10604 => x"27",
         10605 => x"17",
         10606 => x"83",
         10607 => x"57",
         10608 => x"fe",
         10609 => x"80",
         10610 => x"70",
         10611 => x"5b",
         10612 => x"fe",
         10613 => x"78",
         10614 => x"57",
         10615 => x"38",
         10616 => x"38",
         10617 => x"05",
         10618 => x"2a",
         10619 => x"56",
         10620 => x"38",
         10621 => x"81",
         10622 => x"80",
         10623 => x"75",
         10624 => x"79",
         10625 => x"77",
         10626 => x"06",
         10627 => x"2e",
         10628 => x"80",
         10629 => x"7e",
         10630 => x"a0",
         10631 => x"a4",
         10632 => x"9b",
         10633 => x"12",
         10634 => x"2b",
         10635 => x"40",
         10636 => x"5a",
         10637 => x"81",
         10638 => x"88",
         10639 => x"16",
         10640 => x"82",
         10641 => x"90",
         10642 => x"2b",
         10643 => x"33",
         10644 => x"88",
         10645 => x"71",
         10646 => x"8c",
         10647 => x"60",
         10648 => x"41",
         10649 => x"5e",
         10650 => x"84",
         10651 => x"90",
         10652 => x"0b",
         10653 => x"80",
         10654 => x"0c",
         10655 => x"81",
         10656 => x"80",
         10657 => x"38",
         10658 => x"84",
         10659 => x"94",
         10660 => x"1a",
         10661 => x"2b",
         10662 => x"58",
         10663 => x"78",
         10664 => x"56",
         10665 => x"27",
         10666 => x"81",
         10667 => x"5f",
         10668 => x"2e",
         10669 => x"77",
         10670 => x"ff",
         10671 => x"84",
         10672 => x"58",
         10673 => x"08",
         10674 => x"38",
         10675 => x"b9",
         10676 => x"2e",
         10677 => x"75",
         10678 => x"c0",
         10679 => x"c2",
         10680 => x"06",
         10681 => x"38",
         10682 => x"81",
         10683 => x"80",
         10684 => x"38",
         10685 => x"79",
         10686 => x"39",
         10687 => x"79",
         10688 => x"39",
         10689 => x"79",
         10690 => x"39",
         10691 => x"ca",
         10692 => x"c8",
         10693 => x"07",
         10694 => x"fb",
         10695 => x"8b",
         10696 => x"7b",
         10697 => x"fe",
         10698 => x"16",
         10699 => x"33",
         10700 => x"71",
         10701 => x"7d",
         10702 => x"5c",
         10703 => x"7c",
         10704 => x"27",
         10705 => x"74",
         10706 => x"ff",
         10707 => x"84",
         10708 => x"5d",
         10709 => x"08",
         10710 => x"a7",
         10711 => x"c8",
         10712 => x"fc",
         10713 => x"b9",
         10714 => x"2e",
         10715 => x"80",
         10716 => x"76",
         10717 => x"82",
         10718 => x"c8",
         10719 => x"38",
         10720 => x"fe",
         10721 => x"08",
         10722 => x"75",
         10723 => x"af",
         10724 => x"94",
         10725 => x"17",
         10726 => x"55",
         10727 => x"34",
         10728 => x"7d",
         10729 => x"38",
         10730 => x"80",
         10731 => x"34",
         10732 => x"17",
         10733 => x"39",
         10734 => x"94",
         10735 => x"98",
         10736 => x"2b",
         10737 => x"5e",
         10738 => x"0b",
         10739 => x"80",
         10740 => x"34",
         10741 => x"17",
         10742 => x"0b",
         10743 => x"66",
         10744 => x"8b",
         10745 => x"67",
         10746 => x"0b",
         10747 => x"80",
         10748 => x"34",
         10749 => x"7c",
         10750 => x"81",
         10751 => x"38",
         10752 => x"80",
         10753 => x"5e",
         10754 => x"b4",
         10755 => x"2e",
         10756 => x"16",
         10757 => x"7d",
         10758 => x"06",
         10759 => x"54",
         10760 => x"16",
         10761 => x"33",
         10762 => x"ba",
         10763 => x"c8",
         10764 => x"85",
         10765 => x"81",
         10766 => x"17",
         10767 => x"7a",
         10768 => x"18",
         10769 => x"80",
         10770 => x"38",
         10771 => x"f9",
         10772 => x"54",
         10773 => x"53",
         10774 => x"53",
         10775 => x"52",
         10776 => x"81",
         10777 => x"c8",
         10778 => x"09",
         10779 => x"aa",
         10780 => x"c8",
         10781 => x"34",
         10782 => x"a8",
         10783 => x"84",
         10784 => x"5c",
         10785 => x"17",
         10786 => x"92",
         10787 => x"33",
         10788 => x"2e",
         10789 => x"ff",
         10790 => x"54",
         10791 => x"a0",
         10792 => x"53",
         10793 => x"16",
         10794 => x"a3",
         10795 => x"5b",
         10796 => x"74",
         10797 => x"76",
         10798 => x"39",
         10799 => x"0c",
         10800 => x"38",
         10801 => x"06",
         10802 => x"2e",
         10803 => x"7e",
         10804 => x"12",
         10805 => x"5f",
         10806 => x"7d",
         10807 => x"38",
         10808 => x"78",
         10809 => x"1c",
         10810 => x"5c",
         10811 => x"f9",
         10812 => x"89",
         10813 => x"1a",
         10814 => x"f7",
         10815 => x"94",
         10816 => x"56",
         10817 => x"81",
         10818 => x"0c",
         10819 => x"84",
         10820 => x"57",
         10821 => x"f7",
         10822 => x"7f",
         10823 => x"9f",
         10824 => x"0d",
         10825 => x"66",
         10826 => x"5a",
         10827 => x"89",
         10828 => x"2e",
         10829 => x"08",
         10830 => x"2e",
         10831 => x"33",
         10832 => x"2e",
         10833 => x"16",
         10834 => x"22",
         10835 => x"78",
         10836 => x"38",
         10837 => x"41",
         10838 => x"82",
         10839 => x"1a",
         10840 => x"82",
         10841 => x"1a",
         10842 => x"57",
         10843 => x"80",
         10844 => x"38",
         10845 => x"8c",
         10846 => x"31",
         10847 => x"75",
         10848 => x"38",
         10849 => x"81",
         10850 => x"59",
         10851 => x"06",
         10852 => x"e3",
         10853 => x"22",
         10854 => x"89",
         10855 => x"7a",
         10856 => x"83",
         10857 => x"1a",
         10858 => x"75",
         10859 => x"38",
         10860 => x"83",
         10861 => x"98",
         10862 => x"59",
         10863 => x"fe",
         10864 => x"08",
         10865 => x"57",
         10866 => x"83",
         10867 => x"19",
         10868 => x"29",
         10869 => x"05",
         10870 => x"80",
         10871 => x"38",
         10872 => x"89",
         10873 => x"77",
         10874 => x"81",
         10875 => x"55",
         10876 => x"85",
         10877 => x"31",
         10878 => x"76",
         10879 => x"81",
         10880 => x"ff",
         10881 => x"84",
         10882 => x"83",
         10883 => x"83",
         10884 => x"59",
         10885 => x"a9",
         10886 => x"08",
         10887 => x"75",
         10888 => x"38",
         10889 => x"71",
         10890 => x"1b",
         10891 => x"75",
         10892 => x"57",
         10893 => x"81",
         10894 => x"ff",
         10895 => x"ef",
         10896 => x"2b",
         10897 => x"31",
         10898 => x"7f",
         10899 => x"94",
         10900 => x"70",
         10901 => x"0c",
         10902 => x"fe",
         10903 => x"56",
         10904 => x"c8",
         10905 => x"0d",
         10906 => x"b9",
         10907 => x"3d",
         10908 => x"5c",
         10909 => x"9c",
         10910 => x"75",
         10911 => x"84",
         10912 => x"59",
         10913 => x"27",
         10914 => x"58",
         10915 => x"19",
         10916 => x"b6",
         10917 => x"83",
         10918 => x"5d",
         10919 => x"7f",
         10920 => x"06",
         10921 => x"81",
         10922 => x"b8",
         10923 => x"19",
         10924 => x"9e",
         10925 => x"b9",
         10926 => x"2e",
         10927 => x"56",
         10928 => x"b4",
         10929 => x"81",
         10930 => x"94",
         10931 => x"ff",
         10932 => x"7f",
         10933 => x"05",
         10934 => x"80",
         10935 => x"38",
         10936 => x"05",
         10937 => x"70",
         10938 => x"34",
         10939 => x"75",
         10940 => x"d1",
         10941 => x"81",
         10942 => x"77",
         10943 => x"59",
         10944 => x"56",
         10945 => x"fe",
         10946 => x"54",
         10947 => x"53",
         10948 => x"53",
         10949 => x"52",
         10950 => x"c9",
         10951 => x"84",
         10952 => x"7f",
         10953 => x"06",
         10954 => x"84",
         10955 => x"83",
         10956 => x"19",
         10957 => x"08",
         10958 => x"c8",
         10959 => x"74",
         10960 => x"27",
         10961 => x"82",
         10962 => x"74",
         10963 => x"81",
         10964 => x"38",
         10965 => x"19",
         10966 => x"08",
         10967 => x"52",
         10968 => x"51",
         10969 => x"3f",
         10970 => x"bb",
         10971 => x"1b",
         10972 => x"08",
         10973 => x"39",
         10974 => x"52",
         10975 => x"a3",
         10976 => x"b9",
         10977 => x"fc",
         10978 => x"16",
         10979 => x"9c",
         10980 => x"b9",
         10981 => x"06",
         10982 => x"b8",
         10983 => x"08",
         10984 => x"b2",
         10985 => x"91",
         10986 => x"0b",
         10987 => x"0c",
         10988 => x"04",
         10989 => x"1b",
         10990 => x"84",
         10991 => x"92",
         10992 => x"f0",
         10993 => x"65",
         10994 => x"40",
         10995 => x"7e",
         10996 => x"79",
         10997 => x"38",
         10998 => x"75",
         10999 => x"38",
         11000 => x"74",
         11001 => x"38",
         11002 => x"84",
         11003 => x"59",
         11004 => x"85",
         11005 => x"55",
         11006 => x"55",
         11007 => x"38",
         11008 => x"55",
         11009 => x"38",
         11010 => x"70",
         11011 => x"06",
         11012 => x"56",
         11013 => x"82",
         11014 => x"1a",
         11015 => x"5d",
         11016 => x"27",
         11017 => x"09",
         11018 => x"2e",
         11019 => x"76",
         11020 => x"5f",
         11021 => x"38",
         11022 => x"22",
         11023 => x"89",
         11024 => x"56",
         11025 => x"76",
         11026 => x"88",
         11027 => x"74",
         11028 => x"b1",
         11029 => x"2e",
         11030 => x"74",
         11031 => x"8c",
         11032 => x"1b",
         11033 => x"08",
         11034 => x"88",
         11035 => x"56",
         11036 => x"9c",
         11037 => x"81",
         11038 => x"1a",
         11039 => x"9c",
         11040 => x"05",
         11041 => x"77",
         11042 => x"38",
         11043 => x"70",
         11044 => x"18",
         11045 => x"57",
         11046 => x"85",
         11047 => x"15",
         11048 => x"59",
         11049 => x"2e",
         11050 => x"77",
         11051 => x"7f",
         11052 => x"76",
         11053 => x"77",
         11054 => x"7c",
         11055 => x"33",
         11056 => x"a1",
         11057 => x"c8",
         11058 => x"38",
         11059 => x"08",
         11060 => x"57",
         11061 => x"a5",
         11062 => x"0b",
         11063 => x"72",
         11064 => x"58",
         11065 => x"81",
         11066 => x"77",
         11067 => x"59",
         11068 => x"56",
         11069 => x"60",
         11070 => x"1a",
         11071 => x"2b",
         11072 => x"31",
         11073 => x"7f",
         11074 => x"94",
         11075 => x"70",
         11076 => x"0c",
         11077 => x"5a",
         11078 => x"5b",
         11079 => x"83",
         11080 => x"75",
         11081 => x"7a",
         11082 => x"90",
         11083 => x"77",
         11084 => x"5b",
         11085 => x"34",
         11086 => x"84",
         11087 => x"92",
         11088 => x"74",
         11089 => x"0c",
         11090 => x"04",
         11091 => x"55",
         11092 => x"38",
         11093 => x"a2",
         11094 => x"1b",
         11095 => x"76",
         11096 => x"84",
         11097 => x"5a",
         11098 => x"27",
         11099 => x"59",
         11100 => x"16",
         11101 => x"b6",
         11102 => x"83",
         11103 => x"5e",
         11104 => x"7f",
         11105 => x"06",
         11106 => x"81",
         11107 => x"b8",
         11108 => x"16",
         11109 => x"98",
         11110 => x"b9",
         11111 => x"2e",
         11112 => x"57",
         11113 => x"b4",
         11114 => x"83",
         11115 => x"94",
         11116 => x"ff",
         11117 => x"58",
         11118 => x"59",
         11119 => x"80",
         11120 => x"76",
         11121 => x"58",
         11122 => x"81",
         11123 => x"ff",
         11124 => x"ef",
         11125 => x"81",
         11126 => x"34",
         11127 => x"81",
         11128 => x"08",
         11129 => x"70",
         11130 => x"33",
         11131 => x"98",
         11132 => x"5c",
         11133 => x"08",
         11134 => x"81",
         11135 => x"38",
         11136 => x"08",
         11137 => x"b4",
         11138 => x"17",
         11139 => x"b9",
         11140 => x"55",
         11141 => x"08",
         11142 => x"38",
         11143 => x"55",
         11144 => x"09",
         11145 => x"e3",
         11146 => x"b4",
         11147 => x"17",
         11148 => x"7f",
         11149 => x"33",
         11150 => x"a9",
         11151 => x"fe",
         11152 => x"1a",
         11153 => x"1a",
         11154 => x"93",
         11155 => x"33",
         11156 => x"b9",
         11157 => x"b4",
         11158 => x"1b",
         11159 => x"7b",
         11160 => x"0c",
         11161 => x"39",
         11162 => x"52",
         11163 => x"ab",
         11164 => x"b9",
         11165 => x"84",
         11166 => x"fb",
         11167 => x"1a",
         11168 => x"ab",
         11169 => x"79",
         11170 => x"cc",
         11171 => x"c8",
         11172 => x"b9",
         11173 => x"bd",
         11174 => x"81",
         11175 => x"08",
         11176 => x"70",
         11177 => x"33",
         11178 => x"97",
         11179 => x"b9",
         11180 => x"b8",
         11181 => x"c8",
         11182 => x"34",
         11183 => x"a8",
         11184 => x"58",
         11185 => x"08",
         11186 => x"38",
         11187 => x"5c",
         11188 => x"09",
         11189 => x"fc",
         11190 => x"b4",
         11191 => x"17",
         11192 => x"76",
         11193 => x"33",
         11194 => x"f9",
         11195 => x"fb",
         11196 => x"16",
         11197 => x"95",
         11198 => x"b9",
         11199 => x"06",
         11200 => x"f2",
         11201 => x"08",
         11202 => x"ec",
         11203 => x"b4",
         11204 => x"b8",
         11205 => x"81",
         11206 => x"57",
         11207 => x"3f",
         11208 => x"08",
         11209 => x"84",
         11210 => x"83",
         11211 => x"16",
         11212 => x"08",
         11213 => x"a0",
         11214 => x"fe",
         11215 => x"16",
         11216 => x"82",
         11217 => x"06",
         11218 => x"81",
         11219 => x"08",
         11220 => x"05",
         11221 => x"81",
         11222 => x"ff",
         11223 => x"60",
         11224 => x"0c",
         11225 => x"58",
         11226 => x"39",
         11227 => x"1b",
         11228 => x"84",
         11229 => x"92",
         11230 => x"82",
         11231 => x"34",
         11232 => x"b9",
         11233 => x"3d",
         11234 => x"3d",
         11235 => x"89",
         11236 => x"2e",
         11237 => x"08",
         11238 => x"2e",
         11239 => x"33",
         11240 => x"2e",
         11241 => x"16",
         11242 => x"22",
         11243 => x"77",
         11244 => x"38",
         11245 => x"5c",
         11246 => x"81",
         11247 => x"18",
         11248 => x"2a",
         11249 => x"57",
         11250 => x"81",
         11251 => x"a0",
         11252 => x"57",
         11253 => x"79",
         11254 => x"83",
         11255 => x"7a",
         11256 => x"81",
         11257 => x"b8",
         11258 => x"17",
         11259 => x"93",
         11260 => x"b9",
         11261 => x"2e",
         11262 => x"59",
         11263 => x"b4",
         11264 => x"81",
         11265 => x"18",
         11266 => x"33",
         11267 => x"57",
         11268 => x"34",
         11269 => x"19",
         11270 => x"ff",
         11271 => x"5a",
         11272 => x"18",
         11273 => x"2a",
         11274 => x"18",
         11275 => x"76",
         11276 => x"5c",
         11277 => x"83",
         11278 => x"38",
         11279 => x"55",
         11280 => x"74",
         11281 => x"7a",
         11282 => x"74",
         11283 => x"75",
         11284 => x"74",
         11285 => x"78",
         11286 => x"80",
         11287 => x"0b",
         11288 => x"a1",
         11289 => x"34",
         11290 => x"99",
         11291 => x"0b",
         11292 => x"80",
         11293 => x"34",
         11294 => x"0b",
         11295 => x"7b",
         11296 => x"94",
         11297 => x"c8",
         11298 => x"33",
         11299 => x"5b",
         11300 => x"19",
         11301 => x"b9",
         11302 => x"3d",
         11303 => x"54",
         11304 => x"53",
         11305 => x"53",
         11306 => x"52",
         11307 => x"b5",
         11308 => x"84",
         11309 => x"fe",
         11310 => x"b9",
         11311 => x"18",
         11312 => x"08",
         11313 => x"31",
         11314 => x"08",
         11315 => x"a0",
         11316 => x"fe",
         11317 => x"17",
         11318 => x"82",
         11319 => x"06",
         11320 => x"81",
         11321 => x"08",
         11322 => x"05",
         11323 => x"81",
         11324 => x"ff",
         11325 => x"79",
         11326 => x"39",
         11327 => x"55",
         11328 => x"34",
         11329 => x"56",
         11330 => x"34",
         11331 => x"55",
         11332 => x"74",
         11333 => x"7a",
         11334 => x"74",
         11335 => x"75",
         11336 => x"74",
         11337 => x"78",
         11338 => x"80",
         11339 => x"0b",
         11340 => x"a1",
         11341 => x"34",
         11342 => x"99",
         11343 => x"0b",
         11344 => x"80",
         11345 => x"34",
         11346 => x"0b",
         11347 => x"7b",
         11348 => x"c4",
         11349 => x"c8",
         11350 => x"33",
         11351 => x"5b",
         11352 => x"19",
         11353 => x"39",
         11354 => x"51",
         11355 => x"3f",
         11356 => x"08",
         11357 => x"74",
         11358 => x"74",
         11359 => x"5a",
         11360 => x"f9",
         11361 => x"70",
         11362 => x"fe",
         11363 => x"c8",
         11364 => x"b9",
         11365 => x"38",
         11366 => x"80",
         11367 => x"74",
         11368 => x"80",
         11369 => x"72",
         11370 => x"80",
         11371 => x"86",
         11372 => x"16",
         11373 => x"71",
         11374 => x"38",
         11375 => x"58",
         11376 => x"84",
         11377 => x"0c",
         11378 => x"c8",
         11379 => x"0d",
         11380 => x"33",
         11381 => x"bc",
         11382 => x"c8",
         11383 => x"53",
         11384 => x"73",
         11385 => x"56",
         11386 => x"3d",
         11387 => x"70",
         11388 => x"75",
         11389 => x"38",
         11390 => x"05",
         11391 => x"9f",
         11392 => x"71",
         11393 => x"38",
         11394 => x"71",
         11395 => x"38",
         11396 => x"33",
         11397 => x"24",
         11398 => x"84",
         11399 => x"80",
         11400 => x"c8",
         11401 => x"0d",
         11402 => x"84",
         11403 => x"8c",
         11404 => x"78",
         11405 => x"70",
         11406 => x"53",
         11407 => x"89",
         11408 => x"82",
         11409 => x"ff",
         11410 => x"59",
         11411 => x"2e",
         11412 => x"80",
         11413 => x"b8",
         11414 => x"08",
         11415 => x"76",
         11416 => x"58",
         11417 => x"81",
         11418 => x"ff",
         11419 => x"54",
         11420 => x"26",
         11421 => x"12",
         11422 => x"06",
         11423 => x"9f",
         11424 => x"99",
         11425 => x"e0",
         11426 => x"ff",
         11427 => x"71",
         11428 => x"2a",
         11429 => x"73",
         11430 => x"06",
         11431 => x"ff",
         11432 => x"76",
         11433 => x"70",
         11434 => x"2a",
         11435 => x"52",
         11436 => x"2e",
         11437 => x"18",
         11438 => x"58",
         11439 => x"ff",
         11440 => x"51",
         11441 => x"77",
         11442 => x"38",
         11443 => x"51",
         11444 => x"ea",
         11445 => x"53",
         11446 => x"05",
         11447 => x"51",
         11448 => x"84",
         11449 => x"55",
         11450 => x"08",
         11451 => x"38",
         11452 => x"c8",
         11453 => x"0d",
         11454 => x"68",
         11455 => x"d0",
         11456 => x"94",
         11457 => x"c8",
         11458 => x"b9",
         11459 => x"c6",
         11460 => x"d7",
         11461 => x"98",
         11462 => x"80",
         11463 => x"e2",
         11464 => x"05",
         11465 => x"2a",
         11466 => x"59",
         11467 => x"b2",
         11468 => x"9b",
         11469 => x"12",
         11470 => x"2b",
         11471 => x"5e",
         11472 => x"58",
         11473 => x"a4",
         11474 => x"19",
         11475 => x"b9",
         11476 => x"3d",
         11477 => x"b9",
         11478 => x"2e",
         11479 => x"ff",
         11480 => x"0b",
         11481 => x"0c",
         11482 => x"04",
         11483 => x"94",
         11484 => x"98",
         11485 => x"2b",
         11486 => x"98",
         11487 => x"54",
         11488 => x"7e",
         11489 => x"58",
         11490 => x"c8",
         11491 => x"0d",
         11492 => x"3d",
         11493 => x"3d",
         11494 => x"3d",
         11495 => x"80",
         11496 => x"53",
         11497 => x"fd",
         11498 => x"80",
         11499 => x"cf",
         11500 => x"b9",
         11501 => x"84",
         11502 => x"83",
         11503 => x"80",
         11504 => x"7f",
         11505 => x"08",
         11506 => x"0c",
         11507 => x"3d",
         11508 => x"79",
         11509 => x"cc",
         11510 => x"3d",
         11511 => x"5b",
         11512 => x"51",
         11513 => x"3f",
         11514 => x"08",
         11515 => x"c8",
         11516 => x"38",
         11517 => x"3d",
         11518 => x"b4",
         11519 => x"2e",
         11520 => x"b9",
         11521 => x"17",
         11522 => x"7d",
         11523 => x"81",
         11524 => x"b8",
         11525 => x"16",
         11526 => x"8b",
         11527 => x"b9",
         11528 => x"2e",
         11529 => x"57",
         11530 => x"b4",
         11531 => x"82",
         11532 => x"df",
         11533 => x"11",
         11534 => x"33",
         11535 => x"07",
         11536 => x"5d",
         11537 => x"56",
         11538 => x"82",
         11539 => x"80",
         11540 => x"80",
         11541 => x"ff",
         11542 => x"84",
         11543 => x"59",
         11544 => x"08",
         11545 => x"80",
         11546 => x"ff",
         11547 => x"84",
         11548 => x"59",
         11549 => x"08",
         11550 => x"df",
         11551 => x"11",
         11552 => x"33",
         11553 => x"07",
         11554 => x"42",
         11555 => x"56",
         11556 => x"81",
         11557 => x"7a",
         11558 => x"84",
         11559 => x"52",
         11560 => x"a4",
         11561 => x"b9",
         11562 => x"84",
         11563 => x"80",
         11564 => x"38",
         11565 => x"83",
         11566 => x"81",
         11567 => x"e4",
         11568 => x"05",
         11569 => x"ff",
         11570 => x"78",
         11571 => x"33",
         11572 => x"80",
         11573 => x"82",
         11574 => x"17",
         11575 => x"33",
         11576 => x"7c",
         11577 => x"17",
         11578 => x"26",
         11579 => x"76",
         11580 => x"38",
         11581 => x"05",
         11582 => x"80",
         11583 => x"11",
         11584 => x"19",
         11585 => x"58",
         11586 => x"34",
         11587 => x"ff",
         11588 => x"3d",
         11589 => x"58",
         11590 => x"80",
         11591 => x"5a",
         11592 => x"38",
         11593 => x"82",
         11594 => x"0b",
         11595 => x"33",
         11596 => x"83",
         11597 => x"70",
         11598 => x"43",
         11599 => x"5a",
         11600 => x"8d",
         11601 => x"70",
         11602 => x"57",
         11603 => x"f5",
         11604 => x"5b",
         11605 => x"ab",
         11606 => x"76",
         11607 => x"38",
         11608 => x"7e",
         11609 => x"81",
         11610 => x"81",
         11611 => x"77",
         11612 => x"ba",
         11613 => x"05",
         11614 => x"ff",
         11615 => x"06",
         11616 => x"91",
         11617 => x"34",
         11618 => x"c8",
         11619 => x"3d",
         11620 => x"16",
         11621 => x"33",
         11622 => x"71",
         11623 => x"79",
         11624 => x"5e",
         11625 => x"95",
         11626 => x"17",
         11627 => x"2b",
         11628 => x"07",
         11629 => x"dd",
         11630 => x"5d",
         11631 => x"51",
         11632 => x"3f",
         11633 => x"08",
         11634 => x"c8",
         11635 => x"fd",
         11636 => x"b1",
         11637 => x"b4",
         11638 => x"b8",
         11639 => x"81",
         11640 => x"5e",
         11641 => x"3f",
         11642 => x"b9",
         11643 => x"be",
         11644 => x"c8",
         11645 => x"34",
         11646 => x"a8",
         11647 => x"84",
         11648 => x"5a",
         11649 => x"17",
         11650 => x"83",
         11651 => x"33",
         11652 => x"2e",
         11653 => x"fb",
         11654 => x"54",
         11655 => x"a0",
         11656 => x"53",
         11657 => x"16",
         11658 => x"88",
         11659 => x"59",
         11660 => x"ff",
         11661 => x"3d",
         11662 => x"58",
         11663 => x"80",
         11664 => x"a4",
         11665 => x"10",
         11666 => x"05",
         11667 => x"33",
         11668 => x"5e",
         11669 => x"2e",
         11670 => x"fd",
         11671 => x"f1",
         11672 => x"3d",
         11673 => x"19",
         11674 => x"33",
         11675 => x"05",
         11676 => x"60",
         11677 => x"38",
         11678 => x"08",
         11679 => x"59",
         11680 => x"7c",
         11681 => x"5e",
         11682 => x"26",
         11683 => x"f5",
         11684 => x"80",
         11685 => x"84",
         11686 => x"80",
         11687 => x"04",
         11688 => x"7b",
         11689 => x"89",
         11690 => x"2e",
         11691 => x"08",
         11692 => x"2e",
         11693 => x"33",
         11694 => x"2e",
         11695 => x"14",
         11696 => x"22",
         11697 => x"78",
         11698 => x"38",
         11699 => x"5a",
         11700 => x"81",
         11701 => x"15",
         11702 => x"81",
         11703 => x"15",
         11704 => x"76",
         11705 => x"38",
         11706 => x"54",
         11707 => x"78",
         11708 => x"38",
         11709 => x"22",
         11710 => x"52",
         11711 => x"78",
         11712 => x"38",
         11713 => x"17",
         11714 => x"9c",
         11715 => x"c8",
         11716 => x"77",
         11717 => x"55",
         11718 => x"8c",
         11719 => x"c8",
         11720 => x"81",
         11721 => x"30",
         11722 => x"94",
         11723 => x"71",
         11724 => x"08",
         11725 => x"73",
         11726 => x"98",
         11727 => x"27",
         11728 => x"76",
         11729 => x"16",
         11730 => x"17",
         11731 => x"33",
         11732 => x"81",
         11733 => x"57",
         11734 => x"81",
         11735 => x"52",
         11736 => x"99",
         11737 => x"b9",
         11738 => x"84",
         11739 => x"80",
         11740 => x"38",
         11741 => x"98",
         11742 => x"27",
         11743 => x"79",
         11744 => x"14",
         11745 => x"aa",
         11746 => x"16",
         11747 => x"39",
         11748 => x"16",
         11749 => x"72",
         11750 => x"0c",
         11751 => x"04",
         11752 => x"70",
         11753 => x"06",
         11754 => x"fe",
         11755 => x"94",
         11756 => x"57",
         11757 => x"78",
         11758 => x"06",
         11759 => x"77",
         11760 => x"94",
         11761 => x"75",
         11762 => x"38",
         11763 => x"0c",
         11764 => x"80",
         11765 => x"76",
         11766 => x"73",
         11767 => x"59",
         11768 => x"8c",
         11769 => x"08",
         11770 => x"38",
         11771 => x"0c",
         11772 => x"b9",
         11773 => x"3d",
         11774 => x"0b",
         11775 => x"88",
         11776 => x"73",
         11777 => x"fe",
         11778 => x"16",
         11779 => x"2e",
         11780 => x"fe",
         11781 => x"b9",
         11782 => x"94",
         11783 => x"94",
         11784 => x"83",
         11785 => x"75",
         11786 => x"38",
         11787 => x"9c",
         11788 => x"05",
         11789 => x"73",
         11790 => x"f6",
         11791 => x"22",
         11792 => x"b0",
         11793 => x"78",
         11794 => x"5a",
         11795 => x"80",
         11796 => x"38",
         11797 => x"56",
         11798 => x"73",
         11799 => x"ff",
         11800 => x"84",
         11801 => x"54",
         11802 => x"81",
         11803 => x"ff",
         11804 => x"84",
         11805 => x"81",
         11806 => x"fc",
         11807 => x"75",
         11808 => x"fc",
         11809 => x"52",
         11810 => x"97",
         11811 => x"b9",
         11812 => x"84",
         11813 => x"81",
         11814 => x"84",
         11815 => x"ff",
         11816 => x"38",
         11817 => x"08",
         11818 => x"73",
         11819 => x"fe",
         11820 => x"0b",
         11821 => x"82",
         11822 => x"c8",
         11823 => x"0d",
         11824 => x"0d",
         11825 => x"54",
         11826 => x"a2",
         11827 => x"8c",
         11828 => x"52",
         11829 => x"05",
         11830 => x"3f",
         11831 => x"08",
         11832 => x"c8",
         11833 => x"8f",
         11834 => x"0c",
         11835 => x"84",
         11836 => x"8c",
         11837 => x"7a",
         11838 => x"52",
         11839 => x"b9",
         11840 => x"b9",
         11841 => x"84",
         11842 => x"80",
         11843 => x"16",
         11844 => x"2b",
         11845 => x"78",
         11846 => x"86",
         11847 => x"84",
         11848 => x"5b",
         11849 => x"2e",
         11850 => x"9c",
         11851 => x"11",
         11852 => x"33",
         11853 => x"07",
         11854 => x"5d",
         11855 => x"57",
         11856 => x"b3",
         11857 => x"17",
         11858 => x"86",
         11859 => x"17",
         11860 => x"75",
         11861 => x"b9",
         11862 => x"c8",
         11863 => x"84",
         11864 => x"74",
         11865 => x"84",
         11866 => x"0c",
         11867 => x"85",
         11868 => x"0c",
         11869 => x"95",
         11870 => x"18",
         11871 => x"2b",
         11872 => x"07",
         11873 => x"19",
         11874 => x"ff",
         11875 => x"3d",
         11876 => x"89",
         11877 => x"2e",
         11878 => x"08",
         11879 => x"2e",
         11880 => x"33",
         11881 => x"2e",
         11882 => x"13",
         11883 => x"22",
         11884 => x"76",
         11885 => x"80",
         11886 => x"73",
         11887 => x"75",
         11888 => x"b9",
         11889 => x"3d",
         11890 => x"13",
         11891 => x"ff",
         11892 => x"b9",
         11893 => x"06",
         11894 => x"38",
         11895 => x"53",
         11896 => x"f8",
         11897 => x"7c",
         11898 => x"56",
         11899 => x"9f",
         11900 => x"54",
         11901 => x"97",
         11902 => x"53",
         11903 => x"8f",
         11904 => x"22",
         11905 => x"59",
         11906 => x"2e",
         11907 => x"80",
         11908 => x"75",
         11909 => x"c7",
         11910 => x"2e",
         11911 => x"75",
         11912 => x"ff",
         11913 => x"84",
         11914 => x"53",
         11915 => x"08",
         11916 => x"38",
         11917 => x"08",
         11918 => x"52",
         11919 => x"b2",
         11920 => x"52",
         11921 => x"99",
         11922 => x"b9",
         11923 => x"32",
         11924 => x"72",
         11925 => x"84",
         11926 => x"06",
         11927 => x"72",
         11928 => x"0c",
         11929 => x"04",
         11930 => x"75",
         11931 => x"b1",
         11932 => x"52",
         11933 => x"99",
         11934 => x"b9",
         11935 => x"32",
         11936 => x"72",
         11937 => x"84",
         11938 => x"06",
         11939 => x"cf",
         11940 => x"74",
         11941 => x"f9",
         11942 => x"c8",
         11943 => x"c8",
         11944 => x"0d",
         11945 => x"33",
         11946 => x"e8",
         11947 => x"c8",
         11948 => x"53",
         11949 => x"38",
         11950 => x"54",
         11951 => x"39",
         11952 => x"66",
         11953 => x"89",
         11954 => x"97",
         11955 => x"c1",
         11956 => x"b9",
         11957 => x"84",
         11958 => x"80",
         11959 => x"74",
         11960 => x"0c",
         11961 => x"04",
         11962 => x"51",
         11963 => x"3f",
         11964 => x"08",
         11965 => x"c8",
         11966 => x"02",
         11967 => x"33",
         11968 => x"55",
         11969 => x"24",
         11970 => x"80",
         11971 => x"76",
         11972 => x"ff",
         11973 => x"74",
         11974 => x"0c",
         11975 => x"04",
         11976 => x"b9",
         11977 => x"3d",
         11978 => x"3d",
         11979 => x"56",
         11980 => x"95",
         11981 => x"52",
         11982 => x"c0",
         11983 => x"b9",
         11984 => x"84",
         11985 => x"9a",
         11986 => x"0c",
         11987 => x"11",
         11988 => x"94",
         11989 => x"57",
         11990 => x"75",
         11991 => x"75",
         11992 => x"84",
         11993 => x"95",
         11994 => x"84",
         11995 => x"77",
         11996 => x"78",
         11997 => x"93",
         11998 => x"18",
         11999 => x"c8",
         12000 => x"59",
         12001 => x"38",
         12002 => x"71",
         12003 => x"b4",
         12004 => x"2e",
         12005 => x"83",
         12006 => x"5f",
         12007 => x"8d",
         12008 => x"75",
         12009 => x"52",
         12010 => x"51",
         12011 => x"3f",
         12012 => x"08",
         12013 => x"38",
         12014 => x"5e",
         12015 => x"0c",
         12016 => x"57",
         12017 => x"38",
         12018 => x"7d",
         12019 => x"8d",
         12020 => x"b8",
         12021 => x"33",
         12022 => x"71",
         12023 => x"88",
         12024 => x"14",
         12025 => x"07",
         12026 => x"33",
         12027 => x"ff",
         12028 => x"07",
         12029 => x"80",
         12030 => x"60",
         12031 => x"ff",
         12032 => x"05",
         12033 => x"53",
         12034 => x"58",
         12035 => x"78",
         12036 => x"7a",
         12037 => x"94",
         12038 => x"17",
         12039 => x"58",
         12040 => x"34",
         12041 => x"c8",
         12042 => x"0d",
         12043 => x"b4",
         12044 => x"b8",
         12045 => x"81",
         12046 => x"5d",
         12047 => x"3f",
         12048 => x"b9",
         12049 => x"f8",
         12050 => x"c8",
         12051 => x"34",
         12052 => x"a8",
         12053 => x"84",
         12054 => x"5f",
         12055 => x"18",
         12056 => x"bd",
         12057 => x"33",
         12058 => x"2e",
         12059 => x"fe",
         12060 => x"54",
         12061 => x"a0",
         12062 => x"53",
         12063 => x"17",
         12064 => x"fb",
         12065 => x"5e",
         12066 => x"82",
         12067 => x"3d",
         12068 => x"52",
         12069 => x"81",
         12070 => x"b9",
         12071 => x"2e",
         12072 => x"84",
         12073 => x"81",
         12074 => x"38",
         12075 => x"08",
         12076 => x"b9",
         12077 => x"80",
         12078 => x"81",
         12079 => x"58",
         12080 => x"17",
         12081 => x"ca",
         12082 => x"0c",
         12083 => x"0c",
         12084 => x"81",
         12085 => x"84",
         12086 => x"c8",
         12087 => x"b8",
         12088 => x"33",
         12089 => x"88",
         12090 => x"30",
         12091 => x"1f",
         12092 => x"ff",
         12093 => x"5f",
         12094 => x"5f",
         12095 => x"fd",
         12096 => x"8f",
         12097 => x"fd",
         12098 => x"60",
         12099 => x"7f",
         12100 => x"18",
         12101 => x"33",
         12102 => x"77",
         12103 => x"fe",
         12104 => x"60",
         12105 => x"39",
         12106 => x"7b",
         12107 => x"76",
         12108 => x"38",
         12109 => x"74",
         12110 => x"38",
         12111 => x"73",
         12112 => x"38",
         12113 => x"84",
         12114 => x"59",
         12115 => x"81",
         12116 => x"54",
         12117 => x"80",
         12118 => x"17",
         12119 => x"80",
         12120 => x"17",
         12121 => x"2a",
         12122 => x"58",
         12123 => x"80",
         12124 => x"38",
         12125 => x"54",
         12126 => x"08",
         12127 => x"73",
         12128 => x"88",
         12129 => x"08",
         12130 => x"74",
         12131 => x"9c",
         12132 => x"26",
         12133 => x"56",
         12134 => x"18",
         12135 => x"08",
         12136 => x"77",
         12137 => x"59",
         12138 => x"34",
         12139 => x"85",
         12140 => x"18",
         12141 => x"74",
         12142 => x"0c",
         12143 => x"04",
         12144 => x"78",
         12145 => x"38",
         12146 => x"51",
         12147 => x"3f",
         12148 => x"08",
         12149 => x"c8",
         12150 => x"80",
         12151 => x"b9",
         12152 => x"2e",
         12153 => x"84",
         12154 => x"ff",
         12155 => x"38",
         12156 => x"52",
         12157 => x"85",
         12158 => x"b9",
         12159 => x"c8",
         12160 => x"08",
         12161 => x"18",
         12162 => x"58",
         12163 => x"ff",
         12164 => x"15",
         12165 => x"84",
         12166 => x"07",
         12167 => x"17",
         12168 => x"77",
         12169 => x"a0",
         12170 => x"81",
         12171 => x"fe",
         12172 => x"84",
         12173 => x"81",
         12174 => x"fe",
         12175 => x"77",
         12176 => x"fe",
         12177 => x"0b",
         12178 => x"59",
         12179 => x"80",
         12180 => x"0c",
         12181 => x"98",
         12182 => x"76",
         12183 => x"b9",
         12184 => x"c8",
         12185 => x"81",
         12186 => x"b9",
         12187 => x"2e",
         12188 => x"75",
         12189 => x"79",
         12190 => x"c8",
         12191 => x"08",
         12192 => x"38",
         12193 => x"08",
         12194 => x"78",
         12195 => x"54",
         12196 => x"b9",
         12197 => x"81",
         12198 => x"b9",
         12199 => x"17",
         12200 => x"96",
         12201 => x"2e",
         12202 => x"53",
         12203 => x"51",
         12204 => x"3f",
         12205 => x"08",
         12206 => x"c8",
         12207 => x"38",
         12208 => x"51",
         12209 => x"3f",
         12210 => x"08",
         12211 => x"c8",
         12212 => x"80",
         12213 => x"b9",
         12214 => x"2e",
         12215 => x"84",
         12216 => x"ff",
         12217 => x"38",
         12218 => x"52",
         12219 => x"83",
         12220 => x"b9",
         12221 => x"e6",
         12222 => x"08",
         12223 => x"18",
         12224 => x"58",
         12225 => x"90",
         12226 => x"94",
         12227 => x"16",
         12228 => x"54",
         12229 => x"34",
         12230 => x"79",
         12231 => x"38",
         12232 => x"56",
         12233 => x"58",
         12234 => x"81",
         12235 => x"39",
         12236 => x"18",
         12237 => x"fc",
         12238 => x"56",
         12239 => x"0b",
         12240 => x"59",
         12241 => x"39",
         12242 => x"08",
         12243 => x"59",
         12244 => x"39",
         12245 => x"18",
         12246 => x"fd",
         12247 => x"b9",
         12248 => x"c0",
         12249 => x"ff",
         12250 => x"3d",
         12251 => x"a7",
         12252 => x"05",
         12253 => x"51",
         12254 => x"3f",
         12255 => x"08",
         12256 => x"c8",
         12257 => x"8a",
         12258 => x"b9",
         12259 => x"3d",
         12260 => x"4b",
         12261 => x"52",
         12262 => x"52",
         12263 => x"f8",
         12264 => x"c8",
         12265 => x"b9",
         12266 => x"38",
         12267 => x"05",
         12268 => x"2a",
         12269 => x"57",
         12270 => x"cd",
         12271 => x"2b",
         12272 => x"24",
         12273 => x"80",
         12274 => x"70",
         12275 => x"57",
         12276 => x"ff",
         12277 => x"a3",
         12278 => x"11",
         12279 => x"33",
         12280 => x"07",
         12281 => x"5e",
         12282 => x"7c",
         12283 => x"d5",
         12284 => x"2a",
         12285 => x"76",
         12286 => x"ed",
         12287 => x"98",
         12288 => x"2e",
         12289 => x"77",
         12290 => x"84",
         12291 => x"52",
         12292 => x"52",
         12293 => x"f9",
         12294 => x"c8",
         12295 => x"b9",
         12296 => x"e5",
         12297 => x"c8",
         12298 => x"51",
         12299 => x"3f",
         12300 => x"08",
         12301 => x"c8",
         12302 => x"87",
         12303 => x"c8",
         12304 => x"0d",
         12305 => x"33",
         12306 => x"71",
         12307 => x"90",
         12308 => x"07",
         12309 => x"ff",
         12310 => x"b9",
         12311 => x"2e",
         12312 => x"b9",
         12313 => x"a1",
         12314 => x"6f",
         12315 => x"57",
         12316 => x"ff",
         12317 => x"38",
         12318 => x"51",
         12319 => x"3f",
         12320 => x"08",
         12321 => x"c8",
         12322 => x"be",
         12323 => x"70",
         12324 => x"25",
         12325 => x"80",
         12326 => x"74",
         12327 => x"38",
         12328 => x"58",
         12329 => x"27",
         12330 => x"17",
         12331 => x"81",
         12332 => x"56",
         12333 => x"38",
         12334 => x"f5",
         12335 => x"b9",
         12336 => x"b9",
         12337 => x"3d",
         12338 => x"17",
         12339 => x"08",
         12340 => x"b4",
         12341 => x"2e",
         12342 => x"83",
         12343 => x"59",
         12344 => x"2e",
         12345 => x"80",
         12346 => x"54",
         12347 => x"17",
         12348 => x"33",
         12349 => x"ee",
         12350 => x"c8",
         12351 => x"85",
         12352 => x"81",
         12353 => x"18",
         12354 => x"77",
         12355 => x"19",
         12356 => x"78",
         12357 => x"83",
         12358 => x"19",
         12359 => x"fe",
         12360 => x"52",
         12361 => x"8b",
         12362 => x"b9",
         12363 => x"84",
         12364 => x"80",
         12365 => x"38",
         12366 => x"09",
         12367 => x"cd",
         12368 => x"fe",
         12369 => x"54",
         12370 => x"53",
         12371 => x"17",
         12372 => x"f2",
         12373 => x"58",
         12374 => x"08",
         12375 => x"81",
         12376 => x"38",
         12377 => x"08",
         12378 => x"b4",
         12379 => x"18",
         12380 => x"b9",
         12381 => x"55",
         12382 => x"08",
         12383 => x"38",
         12384 => x"55",
         12385 => x"09",
         12386 => x"de",
         12387 => x"b4",
         12388 => x"18",
         12389 => x"7c",
         12390 => x"33",
         12391 => x"c5",
         12392 => x"fe",
         12393 => x"55",
         12394 => x"80",
         12395 => x"52",
         12396 => x"f6",
         12397 => x"b9",
         12398 => x"84",
         12399 => x"80",
         12400 => x"38",
         12401 => x"08",
         12402 => x"e6",
         12403 => x"c8",
         12404 => x"80",
         12405 => x"53",
         12406 => x"51",
         12407 => x"3f",
         12408 => x"08",
         12409 => x"17",
         12410 => x"94",
         12411 => x"5c",
         12412 => x"27",
         12413 => x"81",
         12414 => x"0c",
         12415 => x"81",
         12416 => x"84",
         12417 => x"55",
         12418 => x"ff",
         12419 => x"56",
         12420 => x"79",
         12421 => x"39",
         12422 => x"08",
         12423 => x"39",
         12424 => x"90",
         12425 => x"0d",
         12426 => x"3d",
         12427 => x"52",
         12428 => x"ff",
         12429 => x"84",
         12430 => x"56",
         12431 => x"08",
         12432 => x"38",
         12433 => x"c8",
         12434 => x"0d",
         12435 => x"6f",
         12436 => x"70",
         12437 => x"a6",
         12438 => x"b9",
         12439 => x"84",
         12440 => x"8b",
         12441 => x"84",
         12442 => x"9f",
         12443 => x"84",
         12444 => x"84",
         12445 => x"06",
         12446 => x"80",
         12447 => x"70",
         12448 => x"06",
         12449 => x"56",
         12450 => x"38",
         12451 => x"52",
         12452 => x"52",
         12453 => x"c0",
         12454 => x"c8",
         12455 => x"5c",
         12456 => x"08",
         12457 => x"56",
         12458 => x"08",
         12459 => x"f9",
         12460 => x"c8",
         12461 => x"81",
         12462 => x"81",
         12463 => x"84",
         12464 => x"83",
         12465 => x"5a",
         12466 => x"e2",
         12467 => x"9c",
         12468 => x"05",
         12469 => x"5b",
         12470 => x"8d",
         12471 => x"22",
         12472 => x"b0",
         12473 => x"5c",
         12474 => x"18",
         12475 => x"59",
         12476 => x"57",
         12477 => x"70",
         12478 => x"34",
         12479 => x"74",
         12480 => x"58",
         12481 => x"55",
         12482 => x"81",
         12483 => x"54",
         12484 => x"78",
         12485 => x"33",
         12486 => x"c9",
         12487 => x"c8",
         12488 => x"38",
         12489 => x"dc",
         12490 => x"ff",
         12491 => x"54",
         12492 => x"53",
         12493 => x"53",
         12494 => x"52",
         12495 => x"a5",
         12496 => x"84",
         12497 => x"be",
         12498 => x"c8",
         12499 => x"34",
         12500 => x"a8",
         12501 => x"55",
         12502 => x"08",
         12503 => x"38",
         12504 => x"5b",
         12505 => x"09",
         12506 => x"e1",
         12507 => x"b4",
         12508 => x"18",
         12509 => x"77",
         12510 => x"33",
         12511 => x"e5",
         12512 => x"39",
         12513 => x"7d",
         12514 => x"81",
         12515 => x"b4",
         12516 => x"18",
         12517 => x"ac",
         12518 => x"7c",
         12519 => x"f9",
         12520 => x"c8",
         12521 => x"b9",
         12522 => x"2e",
         12523 => x"84",
         12524 => x"81",
         12525 => x"38",
         12526 => x"08",
         12527 => x"84",
         12528 => x"74",
         12529 => x"fe",
         12530 => x"84",
         12531 => x"fc",
         12532 => x"17",
         12533 => x"94",
         12534 => x"5c",
         12535 => x"27",
         12536 => x"18",
         12537 => x"84",
         12538 => x"07",
         12539 => x"18",
         12540 => x"78",
         12541 => x"a1",
         12542 => x"b9",
         12543 => x"3d",
         12544 => x"17",
         12545 => x"83",
         12546 => x"57",
         12547 => x"78",
         12548 => x"06",
         12549 => x"8b",
         12550 => x"56",
         12551 => x"70",
         12552 => x"34",
         12553 => x"75",
         12554 => x"57",
         12555 => x"18",
         12556 => x"90",
         12557 => x"19",
         12558 => x"75",
         12559 => x"34",
         12560 => x"1a",
         12561 => x"80",
         12562 => x"80",
         12563 => x"d1",
         12564 => x"7c",
         12565 => x"06",
         12566 => x"80",
         12567 => x"77",
         12568 => x"7a",
         12569 => x"34",
         12570 => x"74",
         12571 => x"cc",
         12572 => x"a0",
         12573 => x"1a",
         12574 => x"58",
         12575 => x"81",
         12576 => x"77",
         12577 => x"59",
         12578 => x"56",
         12579 => x"7d",
         12580 => x"80",
         12581 => x"64",
         12582 => x"ff",
         12583 => x"57",
         12584 => x"f2",
         12585 => x"88",
         12586 => x"80",
         12587 => x"75",
         12588 => x"83",
         12589 => x"38",
         12590 => x"0b",
         12591 => x"79",
         12592 => x"96",
         12593 => x"c8",
         12594 => x"b9",
         12595 => x"b6",
         12596 => x"84",
         12597 => x"96",
         12598 => x"b9",
         12599 => x"17",
         12600 => x"98",
         12601 => x"cc",
         12602 => x"34",
         12603 => x"5d",
         12604 => x"34",
         12605 => x"59",
         12606 => x"34",
         12607 => x"79",
         12608 => x"d9",
         12609 => x"90",
         12610 => x"34",
         12611 => x"0b",
         12612 => x"7d",
         12613 => x"80",
         12614 => x"c8",
         12615 => x"84",
         12616 => x"9f",
         12617 => x"76",
         12618 => x"74",
         12619 => x"34",
         12620 => x"57",
         12621 => x"17",
         12622 => x"39",
         12623 => x"5b",
         12624 => x"17",
         12625 => x"2a",
         12626 => x"cd",
         12627 => x"59",
         12628 => x"d8",
         12629 => x"57",
         12630 => x"a1",
         12631 => x"2a",
         12632 => x"18",
         12633 => x"2a",
         12634 => x"18",
         12635 => x"90",
         12636 => x"34",
         12637 => x"0b",
         12638 => x"7d",
         12639 => x"98",
         12640 => x"c8",
         12641 => x"96",
         12642 => x"0d",
         12643 => x"3d",
         12644 => x"5b",
         12645 => x"2e",
         12646 => x"70",
         12647 => x"33",
         12648 => x"56",
         12649 => x"2e",
         12650 => x"74",
         12651 => x"ba",
         12652 => x"38",
         12653 => x"3d",
         12654 => x"52",
         12655 => x"ff",
         12656 => x"84",
         12657 => x"56",
         12658 => x"08",
         12659 => x"38",
         12660 => x"c8",
         12661 => x"0d",
         12662 => x"3d",
         12663 => x"08",
         12664 => x"70",
         12665 => x"9f",
         12666 => x"b9",
         12667 => x"84",
         12668 => x"dc",
         12669 => x"bb",
         12670 => x"a0",
         12671 => x"56",
         12672 => x"a0",
         12673 => x"ae",
         12674 => x"58",
         12675 => x"81",
         12676 => x"77",
         12677 => x"59",
         12678 => x"55",
         12679 => x"99",
         12680 => x"78",
         12681 => x"55",
         12682 => x"05",
         12683 => x"70",
         12684 => x"34",
         12685 => x"74",
         12686 => x"3d",
         12687 => x"51",
         12688 => x"3f",
         12689 => x"08",
         12690 => x"c8",
         12691 => x"38",
         12692 => x"08",
         12693 => x"38",
         12694 => x"b9",
         12695 => x"3d",
         12696 => x"33",
         12697 => x"81",
         12698 => x"57",
         12699 => x"26",
         12700 => x"17",
         12701 => x"06",
         12702 => x"59",
         12703 => x"80",
         12704 => x"7f",
         12705 => x"b8",
         12706 => x"5d",
         12707 => x"5c",
         12708 => x"05",
         12709 => x"70",
         12710 => x"33",
         12711 => x"5a",
         12712 => x"99",
         12713 => x"e0",
         12714 => x"ff",
         12715 => x"ff",
         12716 => x"77",
         12717 => x"38",
         12718 => x"81",
         12719 => x"55",
         12720 => x"9f",
         12721 => x"75",
         12722 => x"81",
         12723 => x"77",
         12724 => x"78",
         12725 => x"30",
         12726 => x"9f",
         12727 => x"5d",
         12728 => x"80",
         12729 => x"81",
         12730 => x"5e",
         12731 => x"24",
         12732 => x"7c",
         12733 => x"5b",
         12734 => x"7b",
         12735 => x"b4",
         12736 => x"0c",
         12737 => x"3d",
         12738 => x"52",
         12739 => x"ff",
         12740 => x"84",
         12741 => x"56",
         12742 => x"08",
         12743 => x"fd",
         12744 => x"aa",
         12745 => x"09",
         12746 => x"ac",
         12747 => x"ff",
         12748 => x"84",
         12749 => x"56",
         12750 => x"08",
         12751 => x"6f",
         12752 => x"8d",
         12753 => x"05",
         12754 => x"58",
         12755 => x"70",
         12756 => x"33",
         12757 => x"05",
         12758 => x"1a",
         12759 => x"38",
         12760 => x"05",
         12761 => x"34",
         12762 => x"70",
         12763 => x"06",
         12764 => x"89",
         12765 => x"07",
         12766 => x"19",
         12767 => x"81",
         12768 => x"34",
         12769 => x"70",
         12770 => x"06",
         12771 => x"80",
         12772 => x"38",
         12773 => x"6b",
         12774 => x"38",
         12775 => x"33",
         12776 => x"71",
         12777 => x"72",
         12778 => x"5c",
         12779 => x"2e",
         12780 => x"fe",
         12781 => x"08",
         12782 => x"56",
         12783 => x"82",
         12784 => x"17",
         12785 => x"29",
         12786 => x"05",
         12787 => x"80",
         12788 => x"38",
         12789 => x"58",
         12790 => x"76",
         12791 => x"83",
         12792 => x"7e",
         12793 => x"81",
         12794 => x"b8",
         12795 => x"17",
         12796 => x"e3",
         12797 => x"b9",
         12798 => x"2e",
         12799 => x"58",
         12800 => x"b4",
         12801 => x"57",
         12802 => x"18",
         12803 => x"fb",
         12804 => x"15",
         12805 => x"ae",
         12806 => x"06",
         12807 => x"70",
         12808 => x"06",
         12809 => x"80",
         12810 => x"7b",
         12811 => x"77",
         12812 => x"34",
         12813 => x"7a",
         12814 => x"81",
         12815 => x"75",
         12816 => x"7d",
         12817 => x"34",
         12818 => x"56",
         12819 => x"18",
         12820 => x"81",
         12821 => x"34",
         12822 => x"3d",
         12823 => x"08",
         12824 => x"74",
         12825 => x"38",
         12826 => x"51",
         12827 => x"3f",
         12828 => x"08",
         12829 => x"c8",
         12830 => x"38",
         12831 => x"98",
         12832 => x"80",
         12833 => x"08",
         12834 => x"38",
         12835 => x"7a",
         12836 => x"7a",
         12837 => x"06",
         12838 => x"81",
         12839 => x"b8",
         12840 => x"16",
         12841 => x"e2",
         12842 => x"b9",
         12843 => x"2e",
         12844 => x"57",
         12845 => x"b4",
         12846 => x"55",
         12847 => x"9c",
         12848 => x"e5",
         12849 => x"0b",
         12850 => x"90",
         12851 => x"27",
         12852 => x"52",
         12853 => x"fc",
         12854 => x"b9",
         12855 => x"84",
         12856 => x"80",
         12857 => x"38",
         12858 => x"84",
         12859 => x"38",
         12860 => x"f9",
         12861 => x"51",
         12862 => x"3f",
         12863 => x"08",
         12864 => x"0c",
         12865 => x"04",
         12866 => x"b9",
         12867 => x"3d",
         12868 => x"18",
         12869 => x"33",
         12870 => x"71",
         12871 => x"78",
         12872 => x"5c",
         12873 => x"84",
         12874 => x"84",
         12875 => x"38",
         12876 => x"08",
         12877 => x"a0",
         12878 => x"b9",
         12879 => x"3d",
         12880 => x"54",
         12881 => x"53",
         12882 => x"16",
         12883 => x"e2",
         12884 => x"58",
         12885 => x"08",
         12886 => x"81",
         12887 => x"38",
         12888 => x"08",
         12889 => x"b4",
         12890 => x"17",
         12891 => x"b9",
         12892 => x"55",
         12893 => x"08",
         12894 => x"38",
         12895 => x"5d",
         12896 => x"09",
         12897 => x"93",
         12898 => x"b4",
         12899 => x"17",
         12900 => x"7b",
         12901 => x"33",
         12902 => x"c9",
         12903 => x"fd",
         12904 => x"54",
         12905 => x"53",
         12906 => x"53",
         12907 => x"52",
         12908 => x"b1",
         12909 => x"84",
         12910 => x"fc",
         12911 => x"b9",
         12912 => x"18",
         12913 => x"08",
         12914 => x"31",
         12915 => x"08",
         12916 => x"a0",
         12917 => x"fc",
         12918 => x"17",
         12919 => x"82",
         12920 => x"06",
         12921 => x"81",
         12922 => x"08",
         12923 => x"05",
         12924 => x"81",
         12925 => x"fe",
         12926 => x"79",
         12927 => x"39",
         12928 => x"02",
         12929 => x"33",
         12930 => x"80",
         12931 => x"56",
         12932 => x"96",
         12933 => x"52",
         12934 => x"ff",
         12935 => x"84",
         12936 => x"56",
         12937 => x"08",
         12938 => x"38",
         12939 => x"c8",
         12940 => x"0d",
         12941 => x"66",
         12942 => x"d0",
         12943 => x"96",
         12944 => x"b9",
         12945 => x"84",
         12946 => x"e0",
         12947 => x"cf",
         12948 => x"a0",
         12949 => x"56",
         12950 => x"74",
         12951 => x"71",
         12952 => x"33",
         12953 => x"74",
         12954 => x"56",
         12955 => x"8b",
         12956 => x"55",
         12957 => x"16",
         12958 => x"fe",
         12959 => x"84",
         12960 => x"84",
         12961 => x"96",
         12962 => x"ec",
         12963 => x"57",
         12964 => x"3d",
         12965 => x"97",
         12966 => x"a1",
         12967 => x"b9",
         12968 => x"84",
         12969 => x"80",
         12970 => x"74",
         12971 => x"0c",
         12972 => x"04",
         12973 => x"52",
         12974 => x"05",
         12975 => x"d8",
         12976 => x"c8",
         12977 => x"b9",
         12978 => x"38",
         12979 => x"05",
         12980 => x"06",
         12981 => x"75",
         12982 => x"84",
         12983 => x"19",
         12984 => x"2b",
         12985 => x"56",
         12986 => x"34",
         12987 => x"55",
         12988 => x"34",
         12989 => x"58",
         12990 => x"34",
         12991 => x"54",
         12992 => x"34",
         12993 => x"0b",
         12994 => x"78",
         12995 => x"88",
         12996 => x"c8",
         12997 => x"c8",
         12998 => x"0d",
         12999 => x"0d",
         13000 => x"5b",
         13001 => x"3d",
         13002 => x"9b",
         13003 => x"a0",
         13004 => x"b9",
         13005 => x"b9",
         13006 => x"70",
         13007 => x"08",
         13008 => x"51",
         13009 => x"80",
         13010 => x"81",
         13011 => x"5a",
         13012 => x"a4",
         13013 => x"70",
         13014 => x"25",
         13015 => x"80",
         13016 => x"38",
         13017 => x"06",
         13018 => x"80",
         13019 => x"38",
         13020 => x"08",
         13021 => x"5a",
         13022 => x"77",
         13023 => x"38",
         13024 => x"7a",
         13025 => x"7a",
         13026 => x"06",
         13027 => x"81",
         13028 => x"b8",
         13029 => x"16",
         13030 => x"dc",
         13031 => x"b9",
         13032 => x"2e",
         13033 => x"57",
         13034 => x"b4",
         13035 => x"57",
         13036 => x"7c",
         13037 => x"58",
         13038 => x"74",
         13039 => x"38",
         13040 => x"74",
         13041 => x"38",
         13042 => x"18",
         13043 => x"11",
         13044 => x"33",
         13045 => x"71",
         13046 => x"81",
         13047 => x"72",
         13048 => x"75",
         13049 => x"62",
         13050 => x"5e",
         13051 => x"76",
         13052 => x"0c",
         13053 => x"04",
         13054 => x"40",
         13055 => x"3d",
         13056 => x"fe",
         13057 => x"84",
         13058 => x"57",
         13059 => x"08",
         13060 => x"8d",
         13061 => x"2e",
         13062 => x"fe",
         13063 => x"7b",
         13064 => x"fe",
         13065 => x"54",
         13066 => x"53",
         13067 => x"53",
         13068 => x"52",
         13069 => x"ad",
         13070 => x"84",
         13071 => x"7a",
         13072 => x"06",
         13073 => x"84",
         13074 => x"83",
         13075 => x"16",
         13076 => x"08",
         13077 => x"c8",
         13078 => x"74",
         13079 => x"27",
         13080 => x"82",
         13081 => x"74",
         13082 => x"81",
         13083 => x"38",
         13084 => x"16",
         13085 => x"08",
         13086 => x"52",
         13087 => x"51",
         13088 => x"3f",
         13089 => x"54",
         13090 => x"16",
         13091 => x"33",
         13092 => x"d2",
         13093 => x"c8",
         13094 => x"fe",
         13095 => x"86",
         13096 => x"74",
         13097 => x"bb",
         13098 => x"c8",
         13099 => x"b9",
         13100 => x"e1",
         13101 => x"c8",
         13102 => x"c8",
         13103 => x"59",
         13104 => x"81",
         13105 => x"57",
         13106 => x"33",
         13107 => x"19",
         13108 => x"27",
         13109 => x"70",
         13110 => x"80",
         13111 => x"80",
         13112 => x"38",
         13113 => x"11",
         13114 => x"57",
         13115 => x"2e",
         13116 => x"e1",
         13117 => x"fd",
         13118 => x"3d",
         13119 => x"a1",
         13120 => x"05",
         13121 => x"51",
         13122 => x"3f",
         13123 => x"08",
         13124 => x"c8",
         13125 => x"38",
         13126 => x"8b",
         13127 => x"a0",
         13128 => x"05",
         13129 => x"15",
         13130 => x"38",
         13131 => x"08",
         13132 => x"81",
         13133 => x"58",
         13134 => x"78",
         13135 => x"38",
         13136 => x"3d",
         13137 => x"81",
         13138 => x"18",
         13139 => x"81",
         13140 => x"7c",
         13141 => x"ff",
         13142 => x"ff",
         13143 => x"a1",
         13144 => x"b5",
         13145 => x"c8",
         13146 => x"dc",
         13147 => x"c8",
         13148 => x"ff",
         13149 => x"80",
         13150 => x"38",
         13151 => x"0b",
         13152 => x"33",
         13153 => x"06",
         13154 => x"78",
         13155 => x"d6",
         13156 => x"78",
         13157 => x"38",
         13158 => x"33",
         13159 => x"06",
         13160 => x"74",
         13161 => x"38",
         13162 => x"09",
         13163 => x"38",
         13164 => x"06",
         13165 => x"a3",
         13166 => x"77",
         13167 => x"38",
         13168 => x"81",
         13169 => x"ff",
         13170 => x"38",
         13171 => x"55",
         13172 => x"81",
         13173 => x"81",
         13174 => x"7b",
         13175 => x"5d",
         13176 => x"a3",
         13177 => x"33",
         13178 => x"06",
         13179 => x"5a",
         13180 => x"fe",
         13181 => x"3d",
         13182 => x"56",
         13183 => x"2e",
         13184 => x"80",
         13185 => x"02",
         13186 => x"79",
         13187 => x"5c",
         13188 => x"2e",
         13189 => x"87",
         13190 => x"5a",
         13191 => x"7d",
         13192 => x"80",
         13193 => x"70",
         13194 => x"ef",
         13195 => x"b9",
         13196 => x"84",
         13197 => x"80",
         13198 => x"74",
         13199 => x"b9",
         13200 => x"3d",
         13201 => x"b5",
         13202 => x"9e",
         13203 => x"b9",
         13204 => x"ff",
         13205 => x"74",
         13206 => x"86",
         13207 => x"b9",
         13208 => x"3d",
         13209 => x"e6",
         13210 => x"fe",
         13211 => x"52",
         13212 => x"f4",
         13213 => x"b9",
         13214 => x"84",
         13215 => x"80",
         13216 => x"80",
         13217 => x"38",
         13218 => x"59",
         13219 => x"70",
         13220 => x"33",
         13221 => x"05",
         13222 => x"15",
         13223 => x"38",
         13224 => x"0b",
         13225 => x"7d",
         13226 => x"ec",
         13227 => x"c8",
         13228 => x"56",
         13229 => x"8a",
         13230 => x"8a",
         13231 => x"ff",
         13232 => x"b9",
         13233 => x"2e",
         13234 => x"fe",
         13235 => x"55",
         13236 => x"fe",
         13237 => x"08",
         13238 => x"52",
         13239 => x"b1",
         13240 => x"c8",
         13241 => x"b9",
         13242 => x"2e",
         13243 => x"81",
         13244 => x"b9",
         13245 => x"19",
         13246 => x"16",
         13247 => x"59",
         13248 => x"77",
         13249 => x"83",
         13250 => x"74",
         13251 => x"81",
         13252 => x"38",
         13253 => x"53",
         13254 => x"81",
         13255 => x"fe",
         13256 => x"84",
         13257 => x"80",
         13258 => x"ff",
         13259 => x"76",
         13260 => x"78",
         13261 => x"38",
         13262 => x"08",
         13263 => x"5a",
         13264 => x"e5",
         13265 => x"38",
         13266 => x"80",
         13267 => x"56",
         13268 => x"2e",
         13269 => x"81",
         13270 => x"81",
         13271 => x"81",
         13272 => x"fe",
         13273 => x"84",
         13274 => x"57",
         13275 => x"08",
         13276 => x"86",
         13277 => x"76",
         13278 => x"bf",
         13279 => x"76",
         13280 => x"a0",
         13281 => x"80",
         13282 => x"05",
         13283 => x"15",
         13284 => x"38",
         13285 => x"0b",
         13286 => x"8b",
         13287 => x"57",
         13288 => x"81",
         13289 => x"76",
         13290 => x"58",
         13291 => x"55",
         13292 => x"fd",
         13293 => x"70",
         13294 => x"33",
         13295 => x"05",
         13296 => x"15",
         13297 => x"38",
         13298 => x"6b",
         13299 => x"34",
         13300 => x"0b",
         13301 => x"7d",
         13302 => x"bc",
         13303 => x"c8",
         13304 => x"ce",
         13305 => x"fe",
         13306 => x"54",
         13307 => x"53",
         13308 => x"18",
         13309 => x"d4",
         13310 => x"b9",
         13311 => x"2e",
         13312 => x"80",
         13313 => x"b9",
         13314 => x"19",
         13315 => x"08",
         13316 => x"31",
         13317 => x"19",
         13318 => x"38",
         13319 => x"55",
         13320 => x"b1",
         13321 => x"c8",
         13322 => x"e8",
         13323 => x"81",
         13324 => x"fe",
         13325 => x"84",
         13326 => x"57",
         13327 => x"08",
         13328 => x"b6",
         13329 => x"39",
         13330 => x"59",
         13331 => x"fd",
         13332 => x"a1",
         13333 => x"b4",
         13334 => x"19",
         13335 => x"7a",
         13336 => x"33",
         13337 => x"fd",
         13338 => x"39",
         13339 => x"60",
         13340 => x"05",
         13341 => x"33",
         13342 => x"89",
         13343 => x"2e",
         13344 => x"08",
         13345 => x"2e",
         13346 => x"33",
         13347 => x"2e",
         13348 => x"15",
         13349 => x"22",
         13350 => x"78",
         13351 => x"38",
         13352 => x"5f",
         13353 => x"38",
         13354 => x"56",
         13355 => x"38",
         13356 => x"81",
         13357 => x"17",
         13358 => x"38",
         13359 => x"70",
         13360 => x"06",
         13361 => x"80",
         13362 => x"38",
         13363 => x"22",
         13364 => x"70",
         13365 => x"57",
         13366 => x"87",
         13367 => x"15",
         13368 => x"30",
         13369 => x"9f",
         13370 => x"c8",
         13371 => x"1c",
         13372 => x"53",
         13373 => x"81",
         13374 => x"38",
         13375 => x"78",
         13376 => x"82",
         13377 => x"56",
         13378 => x"74",
         13379 => x"fe",
         13380 => x"81",
         13381 => x"55",
         13382 => x"75",
         13383 => x"82",
         13384 => x"c8",
         13385 => x"81",
         13386 => x"b9",
         13387 => x"2e",
         13388 => x"84",
         13389 => x"81",
         13390 => x"19",
         13391 => x"2e",
         13392 => x"78",
         13393 => x"06",
         13394 => x"56",
         13395 => x"84",
         13396 => x"90",
         13397 => x"87",
         13398 => x"c8",
         13399 => x"0d",
         13400 => x"33",
         13401 => x"ac",
         13402 => x"c8",
         13403 => x"54",
         13404 => x"38",
         13405 => x"55",
         13406 => x"39",
         13407 => x"81",
         13408 => x"7d",
         13409 => x"80",
         13410 => x"81",
         13411 => x"81",
         13412 => x"38",
         13413 => x"52",
         13414 => x"dd",
         13415 => x"b9",
         13416 => x"84",
         13417 => x"ff",
         13418 => x"81",
         13419 => x"57",
         13420 => x"d7",
         13421 => x"90",
         13422 => x"7b",
         13423 => x"8c",
         13424 => x"18",
         13425 => x"18",
         13426 => x"33",
         13427 => x"5c",
         13428 => x"34",
         13429 => x"fe",
         13430 => x"08",
         13431 => x"7a",
         13432 => x"38",
         13433 => x"94",
         13434 => x"15",
         13435 => x"5d",
         13436 => x"34",
         13437 => x"d6",
         13438 => x"ff",
         13439 => x"5b",
         13440 => x"be",
         13441 => x"fe",
         13442 => x"54",
         13443 => x"ff",
         13444 => x"a1",
         13445 => x"d4",
         13446 => x"0d",
         13447 => x"a5",
         13448 => x"88",
         13449 => x"05",
         13450 => x"5f",
         13451 => x"3d",
         13452 => x"5b",
         13453 => x"2e",
         13454 => x"79",
         13455 => x"5b",
         13456 => x"26",
         13457 => x"ba",
         13458 => x"38",
         13459 => x"75",
         13460 => x"92",
         13461 => x"a4",
         13462 => x"76",
         13463 => x"38",
         13464 => x"84",
         13465 => x"70",
         13466 => x"74",
         13467 => x"38",
         13468 => x"75",
         13469 => x"bc",
         13470 => x"b9",
         13471 => x"40",
         13472 => x"52",
         13473 => x"ce",
         13474 => x"b9",
         13475 => x"ff",
         13476 => x"06",
         13477 => x"57",
         13478 => x"38",
         13479 => x"81",
         13480 => x"57",
         13481 => x"38",
         13482 => x"05",
         13483 => x"79",
         13484 => x"b0",
         13485 => x"c8",
         13486 => x"38",
         13487 => x"80",
         13488 => x"38",
         13489 => x"80",
         13490 => x"38",
         13491 => x"06",
         13492 => x"ff",
         13493 => x"2e",
         13494 => x"80",
         13495 => x"f8",
         13496 => x"80",
         13497 => x"f0",
         13498 => x"7f",
         13499 => x"83",
         13500 => x"89",
         13501 => x"08",
         13502 => x"89",
         13503 => x"4c",
         13504 => x"80",
         13505 => x"38",
         13506 => x"80",
         13507 => x"56",
         13508 => x"74",
         13509 => x"7d",
         13510 => x"df",
         13511 => x"74",
         13512 => x"79",
         13513 => x"be",
         13514 => x"84",
         13515 => x"83",
         13516 => x"83",
         13517 => x"61",
         13518 => x"33",
         13519 => x"07",
         13520 => x"57",
         13521 => x"d5",
         13522 => x"06",
         13523 => x"7d",
         13524 => x"05",
         13525 => x"33",
         13526 => x"80",
         13527 => x"38",
         13528 => x"83",
         13529 => x"12",
         13530 => x"2b",
         13531 => x"07",
         13532 => x"70",
         13533 => x"2b",
         13534 => x"07",
         13535 => x"83",
         13536 => x"12",
         13537 => x"2b",
         13538 => x"07",
         13539 => x"70",
         13540 => x"2b",
         13541 => x"07",
         13542 => x"0c",
         13543 => x"0c",
         13544 => x"44",
         13545 => x"59",
         13546 => x"4b",
         13547 => x"57",
         13548 => x"27",
         13549 => x"93",
         13550 => x"80",
         13551 => x"38",
         13552 => x"70",
         13553 => x"49",
         13554 => x"83",
         13555 => x"87",
         13556 => x"82",
         13557 => x"61",
         13558 => x"66",
         13559 => x"83",
         13560 => x"4a",
         13561 => x"58",
         13562 => x"8a",
         13563 => x"ae",
         13564 => x"2a",
         13565 => x"83",
         13566 => x"56",
         13567 => x"2e",
         13568 => x"77",
         13569 => x"83",
         13570 => x"77",
         13571 => x"70",
         13572 => x"58",
         13573 => x"86",
         13574 => x"27",
         13575 => x"52",
         13576 => x"81",
         13577 => x"b9",
         13578 => x"84",
         13579 => x"b9",
         13580 => x"f5",
         13581 => x"81",
         13582 => x"c8",
         13583 => x"b9",
         13584 => x"71",
         13585 => x"83",
         13586 => x"43",
         13587 => x"89",
         13588 => x"5c",
         13589 => x"1f",
         13590 => x"05",
         13591 => x"05",
         13592 => x"72",
         13593 => x"57",
         13594 => x"2e",
         13595 => x"74",
         13596 => x"90",
         13597 => x"60",
         13598 => x"74",
         13599 => x"f2",
         13600 => x"31",
         13601 => x"53",
         13602 => x"52",
         13603 => x"98",
         13604 => x"c8",
         13605 => x"83",
         13606 => x"38",
         13607 => x"09",
         13608 => x"dd",
         13609 => x"f5",
         13610 => x"c8",
         13611 => x"ac",
         13612 => x"f9",
         13613 => x"55",
         13614 => x"26",
         13615 => x"74",
         13616 => x"39",
         13617 => x"84",
         13618 => x"9f",
         13619 => x"b9",
         13620 => x"81",
         13621 => x"39",
         13622 => x"b9",
         13623 => x"3d",
         13624 => x"d4",
         13625 => x"33",
         13626 => x"81",
         13627 => x"57",
         13628 => x"26",
         13629 => x"1d",
         13630 => x"06",
         13631 => x"58",
         13632 => x"81",
         13633 => x"0b",
         13634 => x"5f",
         13635 => x"7d",
         13636 => x"70",
         13637 => x"33",
         13638 => x"05",
         13639 => x"9f",
         13640 => x"57",
         13641 => x"89",
         13642 => x"70",
         13643 => x"58",
         13644 => x"18",
         13645 => x"26",
         13646 => x"18",
         13647 => x"06",
         13648 => x"30",
         13649 => x"5a",
         13650 => x"2e",
         13651 => x"85",
         13652 => x"be",
         13653 => x"32",
         13654 => x"72",
         13655 => x"7b",
         13656 => x"4a",
         13657 => x"80",
         13658 => x"1c",
         13659 => x"5c",
         13660 => x"ff",
         13661 => x"56",
         13662 => x"9f",
         13663 => x"53",
         13664 => x"51",
         13665 => x"3f",
         13666 => x"b9",
         13667 => x"b6",
         13668 => x"2a",
         13669 => x"b9",
         13670 => x"56",
         13671 => x"bf",
         13672 => x"8e",
         13673 => x"26",
         13674 => x"74",
         13675 => x"fb",
         13676 => x"56",
         13677 => x"7b",
         13678 => x"ba",
         13679 => x"a3",
         13680 => x"f9",
         13681 => x"81",
         13682 => x"57",
         13683 => x"fd",
         13684 => x"6e",
         13685 => x"46",
         13686 => x"39",
         13687 => x"08",
         13688 => x"9d",
         13689 => x"38",
         13690 => x"81",
         13691 => x"fb",
         13692 => x"57",
         13693 => x"c8",
         13694 => x"0d",
         13695 => x"0c",
         13696 => x"62",
         13697 => x"99",
         13698 => x"60",
         13699 => x"74",
         13700 => x"8e",
         13701 => x"ae",
         13702 => x"61",
         13703 => x"76",
         13704 => x"58",
         13705 => x"55",
         13706 => x"8b",
         13707 => x"84",
         13708 => x"76",
         13709 => x"58",
         13710 => x"81",
         13711 => x"ff",
         13712 => x"ef",
         13713 => x"05",
         13714 => x"34",
         13715 => x"05",
         13716 => x"8d",
         13717 => x"83",
         13718 => x"4b",
         13719 => x"05",
         13720 => x"2a",
         13721 => x"8f",
         13722 => x"61",
         13723 => x"62",
         13724 => x"30",
         13725 => x"61",
         13726 => x"78",
         13727 => x"06",
         13728 => x"92",
         13729 => x"56",
         13730 => x"ff",
         13731 => x"38",
         13732 => x"ff",
         13733 => x"61",
         13734 => x"74",
         13735 => x"6b",
         13736 => x"34",
         13737 => x"05",
         13738 => x"98",
         13739 => x"61",
         13740 => x"ff",
         13741 => x"34",
         13742 => x"05",
         13743 => x"9c",
         13744 => x"88",
         13745 => x"61",
         13746 => x"7e",
         13747 => x"6b",
         13748 => x"34",
         13749 => x"84",
         13750 => x"84",
         13751 => x"61",
         13752 => x"62",
         13753 => x"f7",
         13754 => x"a7",
         13755 => x"61",
         13756 => x"a1",
         13757 => x"34",
         13758 => x"aa",
         13759 => x"83",
         13760 => x"55",
         13761 => x"05",
         13762 => x"2a",
         13763 => x"97",
         13764 => x"80",
         13765 => x"34",
         13766 => x"05",
         13767 => x"ab",
         13768 => x"90",
         13769 => x"76",
         13770 => x"58",
         13771 => x"81",
         13772 => x"ff",
         13773 => x"ef",
         13774 => x"fe",
         13775 => x"d5",
         13776 => x"83",
         13777 => x"ff",
         13778 => x"81",
         13779 => x"60",
         13780 => x"fe",
         13781 => x"81",
         13782 => x"c8",
         13783 => x"38",
         13784 => x"62",
         13785 => x"9c",
         13786 => x"57",
         13787 => x"70",
         13788 => x"34",
         13789 => x"74",
         13790 => x"75",
         13791 => x"83",
         13792 => x"38",
         13793 => x"f8",
         13794 => x"2e",
         13795 => x"57",
         13796 => x"76",
         13797 => x"45",
         13798 => x"70",
         13799 => x"34",
         13800 => x"59",
         13801 => x"81",
         13802 => x"76",
         13803 => x"75",
         13804 => x"57",
         13805 => x"66",
         13806 => x"76",
         13807 => x"7a",
         13808 => x"79",
         13809 => x"9d",
         13810 => x"c8",
         13811 => x"38",
         13812 => x"57",
         13813 => x"70",
         13814 => x"34",
         13815 => x"74",
         13816 => x"1b",
         13817 => x"58",
         13818 => x"38",
         13819 => x"40",
         13820 => x"ff",
         13821 => x"56",
         13822 => x"83",
         13823 => x"65",
         13824 => x"26",
         13825 => x"55",
         13826 => x"53",
         13827 => x"51",
         13828 => x"3f",
         13829 => x"08",
         13830 => x"74",
         13831 => x"31",
         13832 => x"db",
         13833 => x"62",
         13834 => x"38",
         13835 => x"83",
         13836 => x"8a",
         13837 => x"62",
         13838 => x"38",
         13839 => x"84",
         13840 => x"83",
         13841 => x"5e",
         13842 => x"38",
         13843 => x"56",
         13844 => x"70",
         13845 => x"34",
         13846 => x"78",
         13847 => x"d5",
         13848 => x"aa",
         13849 => x"83",
         13850 => x"78",
         13851 => x"67",
         13852 => x"81",
         13853 => x"34",
         13854 => x"05",
         13855 => x"84",
         13856 => x"43",
         13857 => x"52",
         13858 => x"fc",
         13859 => x"fe",
         13860 => x"34",
         13861 => x"08",
         13862 => x"07",
         13863 => x"86",
         13864 => x"b9",
         13865 => x"87",
         13866 => x"61",
         13867 => x"34",
         13868 => x"c7",
         13869 => x"61",
         13870 => x"34",
         13871 => x"08",
         13872 => x"05",
         13873 => x"83",
         13874 => x"62",
         13875 => x"64",
         13876 => x"05",
         13877 => x"2a",
         13878 => x"83",
         13879 => x"62",
         13880 => x"7e",
         13881 => x"05",
         13882 => x"78",
         13883 => x"79",
         13884 => x"f1",
         13885 => x"84",
         13886 => x"f7",
         13887 => x"53",
         13888 => x"51",
         13889 => x"3f",
         13890 => x"b9",
         13891 => x"b6",
         13892 => x"c8",
         13893 => x"c8",
         13894 => x"0d",
         13895 => x"0c",
         13896 => x"f9",
         13897 => x"1c",
         13898 => x"5c",
         13899 => x"7a",
         13900 => x"91",
         13901 => x"0b",
         13902 => x"22",
         13903 => x"80",
         13904 => x"74",
         13905 => x"38",
         13906 => x"56",
         13907 => x"17",
         13908 => x"57",
         13909 => x"2e",
         13910 => x"75",
         13911 => x"77",
         13912 => x"fc",
         13913 => x"84",
         13914 => x"10",
         13915 => x"05",
         13916 => x"5e",
         13917 => x"80",
         13918 => x"c8",
         13919 => x"8a",
         13920 => x"fd",
         13921 => x"77",
         13922 => x"38",
         13923 => x"e4",
         13924 => x"c8",
         13925 => x"f5",
         13926 => x"38",
         13927 => x"38",
         13928 => x"5b",
         13929 => x"38",
         13930 => x"c8",
         13931 => x"06",
         13932 => x"2e",
         13933 => x"83",
         13934 => x"39",
         13935 => x"05",
         13936 => x"2a",
         13937 => x"a1",
         13938 => x"90",
         13939 => x"61",
         13940 => x"75",
         13941 => x"76",
         13942 => x"34",
         13943 => x"80",
         13944 => x"05",
         13945 => x"80",
         13946 => x"a1",
         13947 => x"05",
         13948 => x"61",
         13949 => x"34",
         13950 => x"05",
         13951 => x"2a",
         13952 => x"a5",
         13953 => x"90",
         13954 => x"61",
         13955 => x"7c",
         13956 => x"75",
         13957 => x"34",
         13958 => x"05",
         13959 => x"ad",
         13960 => x"61",
         13961 => x"80",
         13962 => x"34",
         13963 => x"05",
         13964 => x"b1",
         13965 => x"61",
         13966 => x"80",
         13967 => x"34",
         13968 => x"80",
         13969 => x"a9",
         13970 => x"05",
         13971 => x"80",
         13972 => x"e5",
         13973 => x"55",
         13974 => x"05",
         13975 => x"70",
         13976 => x"34",
         13977 => x"74",
         13978 => x"cd",
         13979 => x"81",
         13980 => x"76",
         13981 => x"58",
         13982 => x"55",
         13983 => x"f9",
         13984 => x"54",
         13985 => x"52",
         13986 => x"be",
         13987 => x"57",
         13988 => x"08",
         13989 => x"7d",
         13990 => x"05",
         13991 => x"83",
         13992 => x"76",
         13993 => x"c8",
         13994 => x"52",
         13995 => x"bf",
         13996 => x"c3",
         13997 => x"84",
         13998 => x"9f",
         13999 => x"b9",
         14000 => x"f8",
         14001 => x"4a",
         14002 => x"81",
         14003 => x"ff",
         14004 => x"05",
         14005 => x"6a",
         14006 => x"84",
         14007 => x"61",
         14008 => x"ff",
         14009 => x"34",
         14010 => x"05",
         14011 => x"88",
         14012 => x"61",
         14013 => x"ff",
         14014 => x"34",
         14015 => x"7c",
         14016 => x"39",
         14017 => x"1f",
         14018 => x"79",
         14019 => x"d5",
         14020 => x"61",
         14021 => x"75",
         14022 => x"57",
         14023 => x"57",
         14024 => x"60",
         14025 => x"7c",
         14026 => x"5e",
         14027 => x"80",
         14028 => x"81",
         14029 => x"80",
         14030 => x"81",
         14031 => x"80",
         14032 => x"80",
         14033 => x"e4",
         14034 => x"f2",
         14035 => x"05",
         14036 => x"61",
         14037 => x"34",
         14038 => x"83",
         14039 => x"7f",
         14040 => x"7a",
         14041 => x"05",
         14042 => x"2a",
         14043 => x"83",
         14044 => x"7a",
         14045 => x"75",
         14046 => x"05",
         14047 => x"2a",
         14048 => x"83",
         14049 => x"82",
         14050 => x"05",
         14051 => x"83",
         14052 => x"76",
         14053 => x"05",
         14054 => x"83",
         14055 => x"80",
         14056 => x"ff",
         14057 => x"81",
         14058 => x"53",
         14059 => x"51",
         14060 => x"3f",
         14061 => x"1f",
         14062 => x"79",
         14063 => x"a5",
         14064 => x"57",
         14065 => x"39",
         14066 => x"7e",
         14067 => x"80",
         14068 => x"05",
         14069 => x"76",
         14070 => x"38",
         14071 => x"8e",
         14072 => x"54",
         14073 => x"52",
         14074 => x"9a",
         14075 => x"81",
         14076 => x"06",
         14077 => x"3d",
         14078 => x"8d",
         14079 => x"74",
         14080 => x"05",
         14081 => x"17",
         14082 => x"2e",
         14083 => x"77",
         14084 => x"80",
         14085 => x"55",
         14086 => x"76",
         14087 => x"b9",
         14088 => x"3d",
         14089 => x"3d",
         14090 => x"84",
         14091 => x"33",
         14092 => x"8a",
         14093 => x"38",
         14094 => x"56",
         14095 => x"9e",
         14096 => x"08",
         14097 => x"05",
         14098 => x"75",
         14099 => x"55",
         14100 => x"8e",
         14101 => x"18",
         14102 => x"88",
         14103 => x"3d",
         14104 => x"3d",
         14105 => x"74",
         14106 => x"52",
         14107 => x"ff",
         14108 => x"74",
         14109 => x"30",
         14110 => x"9f",
         14111 => x"84",
         14112 => x"1c",
         14113 => x"5a",
         14114 => x"39",
         14115 => x"51",
         14116 => x"ff",
         14117 => x"3d",
         14118 => x"ff",
         14119 => x"3d",
         14120 => x"cc",
         14121 => x"80",
         14122 => x"05",
         14123 => x"15",
         14124 => x"38",
         14125 => x"77",
         14126 => x"2e",
         14127 => x"7c",
         14128 => x"24",
         14129 => x"7d",
         14130 => x"05",
         14131 => x"75",
         14132 => x"55",
         14133 => x"b8",
         14134 => x"18",
         14135 => x"88",
         14136 => x"55",
         14137 => x"9e",
         14138 => x"ff",
         14139 => x"75",
         14140 => x"52",
         14141 => x"ff",
         14142 => x"84",
         14143 => x"86",
         14144 => x"2e",
         14145 => x"0b",
         14146 => x"0c",
         14147 => x"04",
         14148 => x"b0",
         14149 => x"54",
         14150 => x"76",
         14151 => x"9d",
         14152 => x"7b",
         14153 => x"70",
         14154 => x"2a",
         14155 => x"5a",
         14156 => x"a5",
         14157 => x"76",
         14158 => x"3f",
         14159 => x"7d",
         14160 => x"0c",
         14161 => x"04",
         14162 => x"75",
         14163 => x"9a",
         14164 => x"53",
         14165 => x"80",
         14166 => x"38",
         14167 => x"ff",
         14168 => x"84",
         14169 => x"85",
         14170 => x"83",
         14171 => x"27",
         14172 => x"b5",
         14173 => x"06",
         14174 => x"80",
         14175 => x"83",
         14176 => x"51",
         14177 => x"9c",
         14178 => x"70",
         14179 => x"06",
         14180 => x"80",
         14181 => x"38",
         14182 => x"e7",
         14183 => x"22",
         14184 => x"39",
         14185 => x"70",
         14186 => x"84",
         14187 => x"53",
         14188 => x"04",
         14189 => x"02",
         14190 => x"02",
         14191 => x"05",
         14192 => x"80",
         14193 => x"ff",
         14194 => x"70",
         14195 => x"b9",
         14196 => x"3d",
         14197 => x"83",
         14198 => x"81",
         14199 => x"70",
         14200 => x"e9",
         14201 => x"83",
         14202 => x"70",
         14203 => x"c8",
         14204 => x"3d",
         14205 => x"3d",
         14206 => x"70",
         14207 => x"26",
         14208 => x"70",
         14209 => x"06",
         14210 => x"56",
         14211 => x"ff",
         14212 => x"38",
         14213 => x"05",
         14214 => x"71",
         14215 => x"25",
         14216 => x"07",
         14217 => x"53",
         14218 => x"71",
         14219 => x"53",
         14220 => x"88",
         14221 => x"81",
         14222 => x"14",
         14223 => x"76",
         14224 => x"71",
         14225 => x"10",
         14226 => x"82",
         14227 => x"54",
         14228 => x"80",
         14229 => x"26",
         14230 => x"52",
         14231 => x"cb",
         14232 => x"70",
         14233 => x"0c",
         14234 => x"04",
         14235 => x"55",
         14236 => x"71",
         14237 => x"38",
         14238 => x"83",
         14239 => x"54",
         14240 => x"c7",
         14241 => x"83",
         14242 => x"57",
         14243 => x"d3",
         14244 => x"16",
         14245 => x"ff",
         14246 => x"f1",
         14247 => x"70",
         14248 => x"06",
         14249 => x"39",
         14250 => x"83",
         14251 => x"57",
         14252 => x"d0",
         14253 => x"ff",
         14254 => x"51",
         14255 => x"16",
         14256 => x"ff",
         14257 => x"c5",
         14258 => x"70",
         14259 => x"06",
         14260 => x"b9",
         14261 => x"31",
         14262 => x"71",
         14263 => x"ff",
         14264 => x"52",
         14265 => x"39",
         14266 => x"10",
         14267 => x"22",
         14268 => x"ef",
         14269 => x"00",
         14270 => x"ff",
         14271 => x"ff",
         14272 => x"ff",
         14273 => x"00",
         14274 => x"00",
         14275 => x"00",
         14276 => x"00",
         14277 => x"00",
         14278 => x"00",
         14279 => x"00",
         14280 => x"00",
         14281 => x"00",
         14282 => x"00",
         14283 => x"00",
         14284 => x"00",
         14285 => x"00",
         14286 => x"00",
         14287 => x"00",
         14288 => x"00",
         14289 => x"00",
         14290 => x"00",
         14291 => x"00",
         14292 => x"00",
         14293 => x"00",
         14294 => x"00",
         14295 => x"00",
         14296 => x"00",
         14297 => x"00",
         14298 => x"00",
         14299 => x"00",
         14300 => x"00",
         14301 => x"00",
         14302 => x"00",
         14303 => x"00",
         14304 => x"00",
         14305 => x"00",
         14306 => x"00",
         14307 => x"00",
         14308 => x"00",
         14309 => x"00",
         14310 => x"00",
         14311 => x"00",
         14312 => x"00",
         14313 => x"00",
         14314 => x"00",
         14315 => x"00",
         14316 => x"00",
         14317 => x"00",
         14318 => x"00",
         14319 => x"00",
         14320 => x"00",
         14321 => x"00",
         14322 => x"00",
         14323 => x"00",
         14324 => x"00",
         14325 => x"00",
         14326 => x"00",
         14327 => x"00",
         14328 => x"00",
         14329 => x"00",
         14330 => x"00",
         14331 => x"00",
         14332 => x"00",
         14333 => x"00",
         14334 => x"00",
         14335 => x"00",
         14336 => x"00",
         14337 => x"00",
         14338 => x"00",
         14339 => x"00",
         14340 => x"00",
         14341 => x"00",
         14342 => x"00",
         14343 => x"00",
         14344 => x"00",
         14345 => x"00",
         14346 => x"00",
         14347 => x"00",
         14348 => x"00",
         14349 => x"00",
         14350 => x"00",
         14351 => x"00",
         14352 => x"00",
         14353 => x"00",
         14354 => x"00",
         14355 => x"00",
         14356 => x"00",
         14357 => x"00",
         14358 => x"00",
         14359 => x"00",
         14360 => x"00",
         14361 => x"00",
         14362 => x"00",
         14363 => x"00",
         14364 => x"00",
         14365 => x"00",
         14366 => x"00",
         14367 => x"00",
         14368 => x"00",
         14369 => x"00",
         14370 => x"00",
         14371 => x"00",
         14372 => x"00",
         14373 => x"00",
         14374 => x"00",
         14375 => x"00",
         14376 => x"00",
         14377 => x"00",
         14378 => x"00",
         14379 => x"00",
         14380 => x"00",
         14381 => x"00",
         14382 => x"00",
         14383 => x"00",
         14384 => x"00",
         14385 => x"00",
         14386 => x"00",
         14387 => x"00",
         14388 => x"00",
         14389 => x"00",
         14390 => x"00",
         14391 => x"00",
         14392 => x"00",
         14393 => x"00",
         14394 => x"00",
         14395 => x"00",
         14396 => x"00",
         14397 => x"00",
         14398 => x"00",
         14399 => x"00",
         14400 => x"00",
         14401 => x"00",
         14402 => x"00",
         14403 => x"00",
         14404 => x"00",
         14405 => x"00",
         14406 => x"00",
         14407 => x"00",
         14408 => x"00",
         14409 => x"00",
         14410 => x"00",
         14411 => x"00",
         14412 => x"00",
         14413 => x"00",
         14414 => x"00",
         14415 => x"00",
         14416 => x"00",
         14417 => x"00",
         14418 => x"00",
         14419 => x"00",
         14420 => x"00",
         14421 => x"00",
         14422 => x"00",
         14423 => x"00",
         14424 => x"00",
         14425 => x"00",
         14426 => x"00",
         14427 => x"00",
         14428 => x"00",
         14429 => x"00",
         14430 => x"00",
         14431 => x"00",
         14432 => x"00",
         14433 => x"00",
         14434 => x"00",
         14435 => x"00",
         14436 => x"00",
         14437 => x"00",
         14438 => x"00",
         14439 => x"00",
         14440 => x"00",
         14441 => x"00",
         14442 => x"00",
         14443 => x"00",
         14444 => x"00",
         14445 => x"00",
         14446 => x"00",
         14447 => x"00",
         14448 => x"00",
         14449 => x"00",
         14450 => x"00",
         14451 => x"00",
         14452 => x"00",
         14453 => x"00",
         14454 => x"00",
         14455 => x"00",
         14456 => x"00",
         14457 => x"00",
         14458 => x"00",
         14459 => x"00",
         14460 => x"00",
         14461 => x"00",
         14462 => x"00",
         14463 => x"00",
         14464 => x"00",
         14465 => x"00",
         14466 => x"00",
         14467 => x"00",
         14468 => x"00",
         14469 => x"00",
         14470 => x"00",
         14471 => x"00",
         14472 => x"00",
         14473 => x"00",
         14474 => x"00",
         14475 => x"00",
         14476 => x"00",
         14477 => x"00",
         14478 => x"00",
         14479 => x"00",
         14480 => x"00",
         14481 => x"00",
         14482 => x"00",
         14483 => x"00",
         14484 => x"00",
         14485 => x"00",
         14486 => x"00",
         14487 => x"00",
         14488 => x"00",
         14489 => x"00",
         14490 => x"00",
         14491 => x"00",
         14492 => x"00",
         14493 => x"00",
         14494 => x"00",
         14495 => x"00",
         14496 => x"00",
         14497 => x"00",
         14498 => x"00",
         14499 => x"00",
         14500 => x"00",
         14501 => x"00",
         14502 => x"00",
         14503 => x"00",
         14504 => x"00",
         14505 => x"00",
         14506 => x"00",
         14507 => x"00",
         14508 => x"00",
         14509 => x"00",
         14510 => x"00",
         14511 => x"00",
         14512 => x"00",
         14513 => x"00",
         14514 => x"00",
         14515 => x"00",
         14516 => x"00",
         14517 => x"00",
         14518 => x"00",
         14519 => x"00",
         14520 => x"00",
         14521 => x"00",
         14522 => x"00",
         14523 => x"00",
         14524 => x"00",
         14525 => x"00",
         14526 => x"00",
         14527 => x"00",
         14528 => x"00",
         14529 => x"00",
         14530 => x"00",
         14531 => x"00",
         14532 => x"00",
         14533 => x"00",
         14534 => x"00",
         14535 => x"00",
         14536 => x"00",
         14537 => x"00",
         14538 => x"00",
         14539 => x"00",
         14540 => x"00",
         14541 => x"00",
         14542 => x"00",
         14543 => x"00",
         14544 => x"00",
         14545 => x"00",
         14546 => x"00",
         14547 => x"00",
         14548 => x"00",
         14549 => x"00",
         14550 => x"00",
         14551 => x"00",
         14552 => x"00",
         14553 => x"00",
         14554 => x"00",
         14555 => x"00",
         14556 => x"00",
         14557 => x"00",
         14558 => x"00",
         14559 => x"00",
         14560 => x"00",
         14561 => x"00",
         14562 => x"00",
         14563 => x"00",
         14564 => x"00",
         14565 => x"00",
         14566 => x"00",
         14567 => x"00",
         14568 => x"00",
         14569 => x"00",
         14570 => x"00",
         14571 => x"00",
         14572 => x"00",
         14573 => x"00",
         14574 => x"00",
         14575 => x"00",
         14576 => x"00",
         14577 => x"00",
         14578 => x"00",
         14579 => x"00",
         14580 => x"00",
         14581 => x"00",
         14582 => x"00",
         14583 => x"00",
         14584 => x"00",
         14585 => x"00",
         14586 => x"00",
         14587 => x"00",
         14588 => x"00",
         14589 => x"00",
         14590 => x"00",
         14591 => x"00",
         14592 => x"00",
         14593 => x"00",
         14594 => x"00",
         14595 => x"00",
         14596 => x"00",
         14597 => x"00",
         14598 => x"00",
         14599 => x"00",
         14600 => x"00",
         14601 => x"00",
         14602 => x"00",
         14603 => x"00",
         14604 => x"00",
         14605 => x"00",
         14606 => x"00",
         14607 => x"00",
         14608 => x"00",
         14609 => x"00",
         14610 => x"00",
         14611 => x"00",
         14612 => x"00",
         14613 => x"00",
         14614 => x"00",
         14615 => x"00",
         14616 => x"00",
         14617 => x"00",
         14618 => x"00",
         14619 => x"00",
         14620 => x"00",
         14621 => x"00",
         14622 => x"00",
         14623 => x"00",
         14624 => x"00",
         14625 => x"00",
         14626 => x"00",
         14627 => x"00",
         14628 => x"00",
         14629 => x"00",
         14630 => x"00",
         14631 => x"00",
         14632 => x"00",
         14633 => x"00",
         14634 => x"00",
         14635 => x"00",
         14636 => x"00",
         14637 => x"00",
         14638 => x"00",
         14639 => x"00",
         14640 => x"00",
         14641 => x"00",
         14642 => x"00",
         14643 => x"00",
         14644 => x"00",
         14645 => x"00",
         14646 => x"00",
         14647 => x"00",
         14648 => x"00",
         14649 => x"00",
         14650 => x"00",
         14651 => x"00",
         14652 => x"00",
         14653 => x"00",
         14654 => x"00",
         14655 => x"00",
         14656 => x"00",
         14657 => x"00",
         14658 => x"00",
         14659 => x"00",
         14660 => x"00",
         14661 => x"00",
         14662 => x"00",
         14663 => x"00",
         14664 => x"00",
         14665 => x"00",
         14666 => x"00",
         14667 => x"00",
         14668 => x"00",
         14669 => x"00",
         14670 => x"00",
         14671 => x"00",
         14672 => x"00",
         14673 => x"00",
         14674 => x"00",
         14675 => x"00",
         14676 => x"00",
         14677 => x"00",
         14678 => x"00",
         14679 => x"00",
         14680 => x"00",
         14681 => x"00",
         14682 => x"00",
         14683 => x"00",
         14684 => x"00",
         14685 => x"00",
         14686 => x"00",
         14687 => x"00",
         14688 => x"00",
         14689 => x"00",
         14690 => x"00",
         14691 => x"00",
         14692 => x"00",
         14693 => x"00",
         14694 => x"00",
         14695 => x"00",
         14696 => x"00",
         14697 => x"00",
         14698 => x"00",
         14699 => x"00",
         14700 => x"00",
         14701 => x"00",
         14702 => x"00",
         14703 => x"00",
         14704 => x"00",
         14705 => x"00",
         14706 => x"00",
         14707 => x"00",
         14708 => x"00",
         14709 => x"00",
         14710 => x"00",
         14711 => x"00",
         14712 => x"00",
         14713 => x"00",
         14714 => x"00",
         14715 => x"00",
         14716 => x"00",
         14717 => x"00",
         14718 => x"00",
         14719 => x"00",
         14720 => x"00",
         14721 => x"00",
         14722 => x"00",
         14723 => x"00",
         14724 => x"00",
         14725 => x"00",
         14726 => x"00",
         14727 => x"00",
         14728 => x"00",
         14729 => x"00",
         14730 => x"00",
         14731 => x"00",
         14732 => x"00",
         14733 => x"00",
         14734 => x"00",
         14735 => x"00",
         14736 => x"00",
         14737 => x"00",
         14738 => x"00",
         14739 => x"00",
         14740 => x"00",
         14741 => x"00",
         14742 => x"00",
         14743 => x"00",
         14744 => x"00",
         14745 => x"00",
         14746 => x"64",
         14747 => x"74",
         14748 => x"64",
         14749 => x"74",
         14750 => x"66",
         14751 => x"74",
         14752 => x"66",
         14753 => x"64",
         14754 => x"66",
         14755 => x"63",
         14756 => x"6d",
         14757 => x"61",
         14758 => x"6d",
         14759 => x"79",
         14760 => x"6d",
         14761 => x"66",
         14762 => x"6d",
         14763 => x"70",
         14764 => x"6d",
         14765 => x"6d",
         14766 => x"6d",
         14767 => x"68",
         14768 => x"68",
         14769 => x"68",
         14770 => x"68",
         14771 => x"63",
         14772 => x"00",
         14773 => x"6a",
         14774 => x"72",
         14775 => x"61",
         14776 => x"72",
         14777 => x"74",
         14778 => x"69",
         14779 => x"00",
         14780 => x"74",
         14781 => x"00",
         14782 => x"63",
         14783 => x"7a",
         14784 => x"74",
         14785 => x"69",
         14786 => x"6d",
         14787 => x"69",
         14788 => x"6b",
         14789 => x"00",
         14790 => x"65",
         14791 => x"55",
         14792 => x"6f",
         14793 => x"65",
         14794 => x"72",
         14795 => x"50",
         14796 => x"6d",
         14797 => x"72",
         14798 => x"6e",
         14799 => x"72",
         14800 => x"2e",
         14801 => x"54",
         14802 => x"6d",
         14803 => x"20",
         14804 => x"6e",
         14805 => x"6c",
         14806 => x"00",
         14807 => x"49",
         14808 => x"66",
         14809 => x"69",
         14810 => x"20",
         14811 => x"6f",
         14812 => x"00",
         14813 => x"46",
         14814 => x"20",
         14815 => x"6c",
         14816 => x"65",
         14817 => x"54",
         14818 => x"6f",
         14819 => x"20",
         14820 => x"72",
         14821 => x"6f",
         14822 => x"61",
         14823 => x"6c",
         14824 => x"2e",
         14825 => x"46",
         14826 => x"61",
         14827 => x"62",
         14828 => x"65",
         14829 => x"4e",
         14830 => x"6f",
         14831 => x"74",
         14832 => x"65",
         14833 => x"6c",
         14834 => x"73",
         14835 => x"20",
         14836 => x"6e",
         14837 => x"6e",
         14838 => x"73",
         14839 => x"44",
         14840 => x"20",
         14841 => x"20",
         14842 => x"62",
         14843 => x"2e",
         14844 => x"44",
         14845 => x"65",
         14846 => x"6d",
         14847 => x"20",
         14848 => x"69",
         14849 => x"6c",
         14850 => x"00",
         14851 => x"53",
         14852 => x"73",
         14853 => x"69",
         14854 => x"70",
         14855 => x"65",
         14856 => x"64",
         14857 => x"46",
         14858 => x"20",
         14859 => x"64",
         14860 => x"69",
         14861 => x"6c",
         14862 => x"00",
         14863 => x"46",
         14864 => x"20",
         14865 => x"65",
         14866 => x"20",
         14867 => x"73",
         14868 => x"00",
         14869 => x"41",
         14870 => x"73",
         14871 => x"65",
         14872 => x"64",
         14873 => x"49",
         14874 => x"6c",
         14875 => x"66",
         14876 => x"6e",
         14877 => x"2e",
         14878 => x"4e",
         14879 => x"61",
         14880 => x"66",
         14881 => x"64",
         14882 => x"4e",
         14883 => x"69",
         14884 => x"66",
         14885 => x"64",
         14886 => x"44",
         14887 => x"20",
         14888 => x"20",
         14889 => x"64",
         14890 => x"49",
         14891 => x"72",
         14892 => x"20",
         14893 => x"6f",
         14894 => x"44",
         14895 => x"20",
         14896 => x"6f",
         14897 => x"53",
         14898 => x"65",
         14899 => x"00",
         14900 => x"0a",
         14901 => x"20",
         14902 => x"65",
         14903 => x"73",
         14904 => x"20",
         14905 => x"20",
         14906 => x"65",
         14907 => x"65",
         14908 => x"00",
         14909 => x"72",
         14910 => x"00",
         14911 => x"25",
         14912 => x"58",
         14913 => x"3a",
         14914 => x"25",
         14915 => x"00",
         14916 => x"20",
         14917 => x"7c",
         14918 => x"20",
         14919 => x"25",
         14920 => x"00",
         14921 => x"20",
         14922 => x"20",
         14923 => x"00",
         14924 => x"7a",
         14925 => x"2a",
         14926 => x"73",
         14927 => x"31",
         14928 => x"34",
         14929 => x"32",
         14930 => x"76",
         14931 => x"61",
         14932 => x"20",
         14933 => x"2c",
         14934 => x"76",
         14935 => x"32",
         14936 => x"25",
         14937 => x"73",
         14938 => x"0a",
         14939 => x"4f",
         14940 => x"20",
         14941 => x"42",
         14942 => x"20",
         14943 => x"72",
         14944 => x"20",
         14945 => x"20",
         14946 => x"20",
         14947 => x"20",
         14948 => x"30",
         14949 => x"0a",
         14950 => x"20",
         14951 => x"41",
         14952 => x"41",
         14953 => x"65",
         14954 => x"20",
         14955 => x"20",
         14956 => x"20",
         14957 => x"20",
         14958 => x"30",
         14959 => x"0a",
         14960 => x"5a",
         14961 => x"49",
         14962 => x"72",
         14963 => x"74",
         14964 => x"6e",
         14965 => x"72",
         14966 => x"55",
         14967 => x"31",
         14968 => x"20",
         14969 => x"65",
         14970 => x"70",
         14971 => x"55",
         14972 => x"31",
         14973 => x"20",
         14974 => x"65",
         14975 => x"70",
         14976 => x"55",
         14977 => x"30",
         14978 => x"20",
         14979 => x"65",
         14980 => x"70",
         14981 => x"55",
         14982 => x"30",
         14983 => x"20",
         14984 => x"65",
         14985 => x"70",
         14986 => x"49",
         14987 => x"4c",
         14988 => x"20",
         14989 => x"65",
         14990 => x"70",
         14991 => x"49",
         14992 => x"4c",
         14993 => x"20",
         14994 => x"65",
         14995 => x"70",
         14996 => x"50",
         14997 => x"69",
         14998 => x"72",
         14999 => x"74",
         15000 => x"54",
         15001 => x"72",
         15002 => x"74",
         15003 => x"75",
         15004 => x"53",
         15005 => x"69",
         15006 => x"75",
         15007 => x"69",
         15008 => x"2e",
         15009 => x"45",
         15010 => x"6c",
         15011 => x"20",
         15012 => x"65",
         15013 => x"2e",
         15014 => x"61",
         15015 => x"65",
         15016 => x"2e",
         15017 => x"00",
         15018 => x"7a",
         15019 => x"7a",
         15020 => x"68",
         15021 => x"46",
         15022 => x"65",
         15023 => x"6f",
         15024 => x"69",
         15025 => x"6c",
         15026 => x"20",
         15027 => x"63",
         15028 => x"20",
         15029 => x"70",
         15030 => x"73",
         15031 => x"6e",
         15032 => x"6d",
         15033 => x"61",
         15034 => x"2e",
         15035 => x"2a",
         15036 => x"25",
         15037 => x"25",
         15038 => x"30",
         15039 => x"42",
         15040 => x"63",
         15041 => x"61",
         15042 => x"00",
         15043 => x"5a",
         15044 => x"62",
         15045 => x"25",
         15046 => x"25",
         15047 => x"73",
         15048 => x"00",
         15049 => x"43",
         15050 => x"20",
         15051 => x"6f",
         15052 => x"6e",
         15053 => x"2e",
         15054 => x"52",
         15055 => x"61",
         15056 => x"6e",
         15057 => x"70",
         15058 => x"63",
         15059 => x"6f",
         15060 => x"2e",
         15061 => x"43",
         15062 => x"69",
         15063 => x"63",
         15064 => x"20",
         15065 => x"30",
         15066 => x"20",
         15067 => x"0a",
         15068 => x"43",
         15069 => x"20",
         15070 => x"75",
         15071 => x"64",
         15072 => x"64",
         15073 => x"25",
         15074 => x"0a",
         15075 => x"45",
         15076 => x"75",
         15077 => x"67",
         15078 => x"64",
         15079 => x"20",
         15080 => x"6c",
         15081 => x"2e",
         15082 => x"25",
         15083 => x"58",
         15084 => x"38",
         15085 => x"00",
         15086 => x"25",
         15087 => x"58",
         15088 => x"34",
         15089 => x"43",
         15090 => x"61",
         15091 => x"67",
         15092 => x"00",
         15093 => x"25",
         15094 => x"78",
         15095 => x"38",
         15096 => x"3e",
         15097 => x"6c",
         15098 => x"30",
         15099 => x"0a",
         15100 => x"43",
         15101 => x"69",
         15102 => x"2e",
         15103 => x"25",
         15104 => x"58",
         15105 => x"32",
         15106 => x"43",
         15107 => x"72",
         15108 => x"2e",
         15109 => x"00",
         15110 => x"44",
         15111 => x"20",
         15112 => x"6f",
         15113 => x"0a",
         15114 => x"70",
         15115 => x"65",
         15116 => x"25",
         15117 => x"25",
         15118 => x"73",
         15119 => x"4d",
         15120 => x"72",
         15121 => x"78",
         15122 => x"73",
         15123 => x"2c",
         15124 => x"6e",
         15125 => x"20",
         15126 => x"63",
         15127 => x"20",
         15128 => x"6d",
         15129 => x"2e",
         15130 => x"3f",
         15131 => x"25",
         15132 => x"64",
         15133 => x"20",
         15134 => x"25",
         15135 => x"64",
         15136 => x"25",
         15137 => x"53",
         15138 => x"43",
         15139 => x"69",
         15140 => x"61",
         15141 => x"6e",
         15142 => x"3a",
         15143 => x"76",
         15144 => x"73",
         15145 => x"70",
         15146 => x"65",
         15147 => x"64",
         15148 => x"41",
         15149 => x"65",
         15150 => x"73",
         15151 => x"20",
         15152 => x"43",
         15153 => x"52",
         15154 => x"74",
         15155 => x"63",
         15156 => x"20",
         15157 => x"72",
         15158 => x"20",
         15159 => x"30",
         15160 => x"00",
         15161 => x"20",
         15162 => x"43",
         15163 => x"4d",
         15164 => x"72",
         15165 => x"74",
         15166 => x"20",
         15167 => x"72",
         15168 => x"20",
         15169 => x"30",
         15170 => x"00",
         15171 => x"20",
         15172 => x"53",
         15173 => x"6b",
         15174 => x"61",
         15175 => x"41",
         15176 => x"65",
         15177 => x"20",
         15178 => x"20",
         15179 => x"30",
         15180 => x"00",
         15181 => x"4d",
         15182 => x"3a",
         15183 => x"20",
         15184 => x"5a",
         15185 => x"49",
         15186 => x"20",
         15187 => x"20",
         15188 => x"20",
         15189 => x"20",
         15190 => x"20",
         15191 => x"30",
         15192 => x"00",
         15193 => x"20",
         15194 => x"53",
         15195 => x"65",
         15196 => x"6c",
         15197 => x"20",
         15198 => x"71",
         15199 => x"20",
         15200 => x"20",
         15201 => x"64",
         15202 => x"34",
         15203 => x"7a",
         15204 => x"20",
         15205 => x"57",
         15206 => x"62",
         15207 => x"20",
         15208 => x"41",
         15209 => x"6c",
         15210 => x"20",
         15211 => x"71",
         15212 => x"64",
         15213 => x"34",
         15214 => x"7a",
         15215 => x"20",
         15216 => x"53",
         15217 => x"4d",
         15218 => x"6f",
         15219 => x"46",
         15220 => x"20",
         15221 => x"20",
         15222 => x"20",
         15223 => x"64",
         15224 => x"34",
         15225 => x"7a",
         15226 => x"20",
         15227 => x"53",
         15228 => x"20",
         15229 => x"50",
         15230 => x"20",
         15231 => x"49",
         15232 => x"4c",
         15233 => x"20",
         15234 => x"57",
         15235 => x"32",
         15236 => x"20",
         15237 => x"57",
         15238 => x"42",
         15239 => x"20",
         15240 => x"00",
         15241 => x"20",
         15242 => x"49",
         15243 => x"20",
         15244 => x"4c",
         15245 => x"68",
         15246 => x"65",
         15247 => x"25",
         15248 => x"29",
         15249 => x"20",
         15250 => x"54",
         15251 => x"52",
         15252 => x"20",
         15253 => x"69",
         15254 => x"73",
         15255 => x"25",
         15256 => x"29",
         15257 => x"20",
         15258 => x"53",
         15259 => x"41",
         15260 => x"20",
         15261 => x"65",
         15262 => x"65",
         15263 => x"25",
         15264 => x"29",
         15265 => x"20",
         15266 => x"52",
         15267 => x"20",
         15268 => x"20",
         15269 => x"30",
         15270 => x"25",
         15271 => x"29",
         15272 => x"20",
         15273 => x"42",
         15274 => x"20",
         15275 => x"20",
         15276 => x"30",
         15277 => x"25",
         15278 => x"29",
         15279 => x"20",
         15280 => x"49",
         15281 => x"20",
         15282 => x"4d",
         15283 => x"30",
         15284 => x"25",
         15285 => x"29",
         15286 => x"20",
         15287 => x"53",
         15288 => x"4d",
         15289 => x"20",
         15290 => x"30",
         15291 => x"25",
         15292 => x"29",
         15293 => x"20",
         15294 => x"57",
         15295 => x"44",
         15296 => x"20",
         15297 => x"30",
         15298 => x"25",
         15299 => x"29",
         15300 => x"20",
         15301 => x"6f",
         15302 => x"6f",
         15303 => x"6f",
         15304 => x"67",
         15305 => x"55",
         15306 => x"6f",
         15307 => x"45",
         15308 => x"00",
         15309 => x"53",
         15310 => x"6c",
         15311 => x"4d",
         15312 => x"75",
         15313 => x"46",
         15314 => x"00",
         15315 => x"45",
         15316 => x"00",
         15317 => x"01",
         15318 => x"00",
         15319 => x"00",
         15320 => x"01",
         15321 => x"00",
         15322 => x"00",
         15323 => x"01",
         15324 => x"00",
         15325 => x"00",
         15326 => x"01",
         15327 => x"00",
         15328 => x"00",
         15329 => x"01",
         15330 => x"00",
         15331 => x"00",
         15332 => x"01",
         15333 => x"00",
         15334 => x"00",
         15335 => x"01",
         15336 => x"00",
         15337 => x"00",
         15338 => x"01",
         15339 => x"00",
         15340 => x"00",
         15341 => x"01",
         15342 => x"00",
         15343 => x"00",
         15344 => x"01",
         15345 => x"00",
         15346 => x"00",
         15347 => x"01",
         15348 => x"00",
         15349 => x"00",
         15350 => x"04",
         15351 => x"00",
         15352 => x"00",
         15353 => x"04",
         15354 => x"00",
         15355 => x"00",
         15356 => x"04",
         15357 => x"00",
         15358 => x"00",
         15359 => x"03",
         15360 => x"00",
         15361 => x"00",
         15362 => x"04",
         15363 => x"00",
         15364 => x"00",
         15365 => x"04",
         15366 => x"00",
         15367 => x"00",
         15368 => x"04",
         15369 => x"00",
         15370 => x"00",
         15371 => x"03",
         15372 => x"00",
         15373 => x"00",
         15374 => x"03",
         15375 => x"00",
         15376 => x"00",
         15377 => x"03",
         15378 => x"00",
         15379 => x"00",
         15380 => x"03",
         15381 => x"00",
         15382 => x"1b",
         15383 => x"1b",
         15384 => x"1b",
         15385 => x"1b",
         15386 => x"1b",
         15387 => x"1b",
         15388 => x"1b",
         15389 => x"1b",
         15390 => x"1b",
         15391 => x"1b",
         15392 => x"1b",
         15393 => x"10",
         15394 => x"0e",
         15395 => x"0d",
         15396 => x"0b",
         15397 => x"08",
         15398 => x"06",
         15399 => x"05",
         15400 => x"04",
         15401 => x"03",
         15402 => x"02",
         15403 => x"01",
         15404 => x"43",
         15405 => x"6f",
         15406 => x"70",
         15407 => x"63",
         15408 => x"74",
         15409 => x"69",
         15410 => x"72",
         15411 => x"69",
         15412 => x"20",
         15413 => x"61",
         15414 => x"6e",
         15415 => x"68",
         15416 => x"6f",
         15417 => x"68",
         15418 => x"00",
         15419 => x"21",
         15420 => x"25",
         15421 => x"75",
         15422 => x"73",
         15423 => x"46",
         15424 => x"65",
         15425 => x"6f",
         15426 => x"73",
         15427 => x"74",
         15428 => x"68",
         15429 => x"6f",
         15430 => x"66",
         15431 => x"20",
         15432 => x"45",
         15433 => x"00",
         15434 => x"3e",
         15435 => x"00",
         15436 => x"1b",
         15437 => x"00",
         15438 => x"1b",
         15439 => x"1b",
         15440 => x"1b",
         15441 => x"1b",
         15442 => x"1b",
         15443 => x"7e",
         15444 => x"1b",
         15445 => x"7e",
         15446 => x"1b",
         15447 => x"7e",
         15448 => x"1b",
         15449 => x"7e",
         15450 => x"1b",
         15451 => x"7e",
         15452 => x"1b",
         15453 => x"7e",
         15454 => x"1b",
         15455 => x"7e",
         15456 => x"1b",
         15457 => x"7e",
         15458 => x"1b",
         15459 => x"7e",
         15460 => x"1b",
         15461 => x"7e",
         15462 => x"1b",
         15463 => x"00",
         15464 => x"1b",
         15465 => x"00",
         15466 => x"1b",
         15467 => x"1b",
         15468 => x"00",
         15469 => x"1b",
         15470 => x"00",
         15471 => x"58",
         15472 => x"2c",
         15473 => x"25",
         15474 => x"64",
         15475 => x"2c",
         15476 => x"25",
         15477 => x"00",
         15478 => x"44",
         15479 => x"2d",
         15480 => x"25",
         15481 => x"63",
         15482 => x"2c",
         15483 => x"25",
         15484 => x"25",
         15485 => x"4b",
         15486 => x"3a",
         15487 => x"25",
         15488 => x"2c",
         15489 => x"25",
         15490 => x"64",
         15491 => x"52",
         15492 => x"52",
         15493 => x"72",
         15494 => x"75",
         15495 => x"72",
         15496 => x"55",
         15497 => x"30",
         15498 => x"25",
         15499 => x"00",
         15500 => x"44",
         15501 => x"30",
         15502 => x"25",
         15503 => x"00",
         15504 => x"48",
         15505 => x"30",
         15506 => x"00",
         15507 => x"4e",
         15508 => x"65",
         15509 => x"64",
         15510 => x"6e",
         15511 => x"00",
         15512 => x"53",
         15513 => x"22",
         15514 => x"3e",
         15515 => x"00",
         15516 => x"2b",
         15517 => x"5b",
         15518 => x"46",
         15519 => x"46",
         15520 => x"32",
         15521 => x"eb",
         15522 => x"53",
         15523 => x"35",
         15524 => x"4e",
         15525 => x"41",
         15526 => x"20",
         15527 => x"41",
         15528 => x"20",
         15529 => x"4e",
         15530 => x"41",
         15531 => x"20",
         15532 => x"41",
         15533 => x"20",
         15534 => x"00",
         15535 => x"00",
         15536 => x"00",
         15537 => x"00",
         15538 => x"01",
         15539 => x"09",
         15540 => x"14",
         15541 => x"1e",
         15542 => x"80",
         15543 => x"8e",
         15544 => x"45",
         15545 => x"49",
         15546 => x"90",
         15547 => x"99",
         15548 => x"59",
         15549 => x"9c",
         15550 => x"41",
         15551 => x"a5",
         15552 => x"a8",
         15553 => x"ac",
         15554 => x"b0",
         15555 => x"b4",
         15556 => x"b8",
         15557 => x"bc",
         15558 => x"c0",
         15559 => x"c4",
         15560 => x"c8",
         15561 => x"cc",
         15562 => x"d0",
         15563 => x"d4",
         15564 => x"d8",
         15565 => x"dc",
         15566 => x"e0",
         15567 => x"e4",
         15568 => x"e8",
         15569 => x"ec",
         15570 => x"f0",
         15571 => x"f4",
         15572 => x"f8",
         15573 => x"fc",
         15574 => x"2b",
         15575 => x"3d",
         15576 => x"5c",
         15577 => x"3c",
         15578 => x"7f",
         15579 => x"00",
         15580 => x"00",
         15581 => x"01",
         15582 => x"00",
         15583 => x"00",
         15584 => x"00",
         15585 => x"00",
         15586 => x"00",
         15587 => x"00",
         15588 => x"00",
         15589 => x"00",
         15590 => x"00",
         15591 => x"00",
         15592 => x"00",
         15593 => x"00",
         15594 => x"00",
         15595 => x"00",
         15596 => x"00",
         15597 => x"00",
         15598 => x"00",
         15599 => x"00",
         15600 => x"00",
         15601 => x"00",
         15602 => x"20",
         15603 => x"00",
         15604 => x"00",
         15605 => x"00",
         15606 => x"00",
         15607 => x"00",
         15608 => x"00",
         15609 => x"00",
         15610 => x"00",
         15611 => x"25",
         15612 => x"25",
         15613 => x"25",
         15614 => x"25",
         15615 => x"25",
         15616 => x"25",
         15617 => x"25",
         15618 => x"25",
         15619 => x"25",
         15620 => x"25",
         15621 => x"25",
         15622 => x"25",
         15623 => x"25",
         15624 => x"25",
         15625 => x"25",
         15626 => x"25",
         15627 => x"25",
         15628 => x"25",
         15629 => x"25",
         15630 => x"25",
         15631 => x"25",
         15632 => x"25",
         15633 => x"25",
         15634 => x"25",
         15635 => x"03",
         15636 => x"03",
         15637 => x"03",
         15638 => x"00",
         15639 => x"03",
         15640 => x"03",
         15641 => x"22",
         15642 => x"03",
         15643 => x"22",
         15644 => x"22",
         15645 => x"23",
         15646 => x"00",
         15647 => x"00",
         15648 => x"00",
         15649 => x"20",
         15650 => x"25",
         15651 => x"00",
         15652 => x"00",
         15653 => x"00",
         15654 => x"00",
         15655 => x"01",
         15656 => x"01",
         15657 => x"01",
         15658 => x"01",
         15659 => x"01",
         15660 => x"01",
         15661 => x"00",
         15662 => x"01",
         15663 => x"01",
         15664 => x"01",
         15665 => x"01",
         15666 => x"01",
         15667 => x"01",
         15668 => x"01",
         15669 => x"01",
         15670 => x"01",
         15671 => x"01",
         15672 => x"01",
         15673 => x"01",
         15674 => x"01",
         15675 => x"01",
         15676 => x"01",
         15677 => x"01",
         15678 => x"01",
         15679 => x"01",
         15680 => x"01",
         15681 => x"01",
         15682 => x"01",
         15683 => x"01",
         15684 => x"01",
         15685 => x"01",
         15686 => x"01",
         15687 => x"01",
         15688 => x"01",
         15689 => x"01",
         15690 => x"01",
         15691 => x"01",
         15692 => x"01",
         15693 => x"01",
         15694 => x"01",
         15695 => x"01",
         15696 => x"01",
         15697 => x"01",
         15698 => x"01",
         15699 => x"01",
         15700 => x"01",
         15701 => x"01",
         15702 => x"01",
         15703 => x"01",
         15704 => x"00",
         15705 => x"01",
         15706 => x"01",
         15707 => x"02",
         15708 => x"02",
         15709 => x"2c",
         15710 => x"02",
         15711 => x"2c",
         15712 => x"02",
         15713 => x"02",
         15714 => x"01",
         15715 => x"00",
         15716 => x"01",
         15717 => x"01",
         15718 => x"02",
         15719 => x"02",
         15720 => x"02",
         15721 => x"02",
         15722 => x"01",
         15723 => x"02",
         15724 => x"02",
         15725 => x"02",
         15726 => x"01",
         15727 => x"02",
         15728 => x"02",
         15729 => x"02",
         15730 => x"02",
         15731 => x"01",
         15732 => x"02",
         15733 => x"02",
         15734 => x"02",
         15735 => x"02",
         15736 => x"02",
         15737 => x"02",
         15738 => x"01",
         15739 => x"02",
         15740 => x"02",
         15741 => x"02",
         15742 => x"01",
         15743 => x"01",
         15744 => x"02",
         15745 => x"02",
         15746 => x"02",
         15747 => x"01",
         15748 => x"00",
         15749 => x"03",
         15750 => x"03",
         15751 => x"03",
         15752 => x"03",
         15753 => x"03",
         15754 => x"03",
         15755 => x"03",
         15756 => x"03",
         15757 => x"03",
         15758 => x"03",
         15759 => x"03",
         15760 => x"01",
         15761 => x"00",
         15762 => x"03",
         15763 => x"03",
         15764 => x"03",
         15765 => x"03",
         15766 => x"03",
         15767 => x"03",
         15768 => x"07",
         15769 => x"01",
         15770 => x"01",
         15771 => x"01",
         15772 => x"00",
         15773 => x"04",
         15774 => x"05",
         15775 => x"00",
         15776 => x"1d",
         15777 => x"2c",
         15778 => x"01",
         15779 => x"01",
         15780 => x"06",
         15781 => x"06",
         15782 => x"06",
         15783 => x"06",
         15784 => x"06",
         15785 => x"00",
         15786 => x"1f",
         15787 => x"1f",
         15788 => x"1f",
         15789 => x"1f",
         15790 => x"1f",
         15791 => x"1f",
         15792 => x"1f",
         15793 => x"1f",
         15794 => x"1f",
         15795 => x"1f",
         15796 => x"1f",
         15797 => x"1f",
         15798 => x"1f",
         15799 => x"1f",
         15800 => x"1f",
         15801 => x"1f",
         15802 => x"1f",
         15803 => x"1f",
         15804 => x"1f",
         15805 => x"1f",
         15806 => x"06",
         15807 => x"06",
         15808 => x"00",
         15809 => x"1f",
         15810 => x"1f",
         15811 => x"00",
         15812 => x"21",
         15813 => x"21",
         15814 => x"21",
         15815 => x"05",
         15816 => x"04",
         15817 => x"01",
         15818 => x"01",
         15819 => x"01",
         15820 => x"01",
         15821 => x"08",
         15822 => x"03",
         15823 => x"00",
         15824 => x"00",
         15825 => x"01",
         15826 => x"00",
         15827 => x"00",
         15828 => x"00",
         15829 => x"01",
         15830 => x"00",
         15831 => x"00",
         15832 => x"00",
         15833 => x"01",
         15834 => x"00",
         15835 => x"00",
         15836 => x"00",
         15837 => x"01",
         15838 => x"00",
         15839 => x"00",
         15840 => x"00",
         15841 => x"01",
         15842 => x"00",
         15843 => x"00",
         15844 => x"00",
         15845 => x"01",
         15846 => x"00",
         15847 => x"00",
         15848 => x"00",
         15849 => x"01",
         15850 => x"00",
         15851 => x"00",
         15852 => x"00",
         15853 => x"01",
         15854 => x"00",
         15855 => x"00",
         15856 => x"00",
         15857 => x"01",
         15858 => x"00",
         15859 => x"00",
         15860 => x"00",
         15861 => x"01",
         15862 => x"00",
         15863 => x"00",
         15864 => x"00",
         15865 => x"01",
         15866 => x"00",
         15867 => x"00",
         15868 => x"00",
         15869 => x"01",
         15870 => x"00",
         15871 => x"00",
         15872 => x"00",
         15873 => x"01",
         15874 => x"00",
         15875 => x"00",
         15876 => x"00",
         15877 => x"01",
         15878 => x"00",
         15879 => x"00",
         15880 => x"00",
         15881 => x"01",
         15882 => x"00",
         15883 => x"00",
         15884 => x"00",
         15885 => x"01",
         15886 => x"00",
         15887 => x"00",
         15888 => x"00",
         15889 => x"01",
         15890 => x"00",
         15891 => x"00",
         15892 => x"00",
         15893 => x"01",
         15894 => x"00",
         15895 => x"00",
         15896 => x"00",
         15897 => x"01",
         15898 => x"00",
         15899 => x"00",
         15900 => x"00",
         15901 => x"01",
         15902 => x"00",
         15903 => x"00",
         15904 => x"00",
         15905 => x"01",
         15906 => x"00",
         15907 => x"00",
         15908 => x"00",
         15909 => x"01",
         15910 => x"00",
         15911 => x"00",
         15912 => x"00",
         15913 => x"01",
         15914 => x"00",
         15915 => x"00",
         15916 => x"00",
         15917 => x"01",
         15918 => x"00",
         15919 => x"00",
         15920 => x"00",
         15921 => x"01",
         15922 => x"00",
         15923 => x"00",
         15924 => x"00",
         15925 => x"01",
         15926 => x"00",
         15927 => x"00",
         15928 => x"00",
         15929 => x"01",
         15930 => x"00",
         15931 => x"00",
         15932 => x"00",
         15933 => x"01",
         15934 => x"00",
         15935 => x"00",
         15936 => x"00",
         15937 => x"00",
         15938 => x"00",
         15939 => x"00",
         15940 => x"00",
         15941 => x"00",
         15942 => x"00",
         15943 => x"00",
         15944 => x"00",
         15945 => x"01",
         15946 => x"01",
         15947 => x"00",
         15948 => x"00",
         15949 => x"00",
         15950 => x"00",
         15951 => x"05",
         15952 => x"05",
         15953 => x"05",
         15954 => x"00",
         15955 => x"01",
         15956 => x"01",
         15957 => x"01",
         15958 => x"01",
         15959 => x"00",
         15960 => x"00",
         15961 => x"00",
         15962 => x"00",
         15963 => x"00",
         15964 => x"00",
         15965 => x"00",
         15966 => x"00",
         15967 => x"00",
         15968 => x"00",
         15969 => x"00",
         15970 => x"00",
         15971 => x"00",
         15972 => x"00",
         15973 => x"00",
         15974 => x"00",
         15975 => x"00",
         15976 => x"00",
         15977 => x"00",
         15978 => x"00",
         15979 => x"00",
         15980 => x"00",
         15981 => x"00",
         15982 => x"00",
         15983 => x"00",
         15984 => x"01",
         15985 => x"00",
         15986 => x"01",
         15987 => x"00",
         15988 => x"02",
         15989 => x"00",
         15990 => x"1b",
         15991 => x"f0",
         15992 => x"79",
         15993 => x"5d",
         15994 => x"71",
         15995 => x"75",
         15996 => x"69",
         15997 => x"6d",
         15998 => x"61",
         15999 => x"65",
         16000 => x"31",
         16001 => x"35",
         16002 => x"5c",
         16003 => x"30",
         16004 => x"f6",
         16005 => x"f1",
         16006 => x"08",
         16007 => x"f0",
         16008 => x"80",
         16009 => x"84",
         16010 => x"1b",
         16011 => x"f0",
         16012 => x"59",
         16013 => x"5d",
         16014 => x"51",
         16015 => x"55",
         16016 => x"49",
         16017 => x"4d",
         16018 => x"41",
         16019 => x"45",
         16020 => x"31",
         16021 => x"35",
         16022 => x"5c",
         16023 => x"30",
         16024 => x"f6",
         16025 => x"f1",
         16026 => x"08",
         16027 => x"f0",
         16028 => x"80",
         16029 => x"84",
         16030 => x"1b",
         16031 => x"f0",
         16032 => x"59",
         16033 => x"7d",
         16034 => x"51",
         16035 => x"55",
         16036 => x"49",
         16037 => x"4d",
         16038 => x"41",
         16039 => x"45",
         16040 => x"21",
         16041 => x"25",
         16042 => x"7c",
         16043 => x"20",
         16044 => x"f7",
         16045 => x"f9",
         16046 => x"fb",
         16047 => x"f0",
         16048 => x"85",
         16049 => x"89",
         16050 => x"1b",
         16051 => x"f0",
         16052 => x"19",
         16053 => x"1d",
         16054 => x"11",
         16055 => x"15",
         16056 => x"09",
         16057 => x"0d",
         16058 => x"01",
         16059 => x"05",
         16060 => x"f0",
         16061 => x"f0",
         16062 => x"f0",
         16063 => x"f0",
         16064 => x"f0",
         16065 => x"f0",
         16066 => x"f0",
         16067 => x"f0",
         16068 => x"80",
         16069 => x"84",
         16070 => x"bf",
         16071 => x"f0",
         16072 => x"35",
         16073 => x"b7",
         16074 => x"7c",
         16075 => x"39",
         16076 => x"3d",
         16077 => x"1d",
         16078 => x"46",
         16079 => x"74",
         16080 => x"3f",
         16081 => x"7a",
         16082 => x"d3",
         16083 => x"9d",
         16084 => x"c6",
         16085 => x"c3",
         16086 => x"f0",
         16087 => x"f0",
         16088 => x"80",
         16089 => x"84",
         16090 => x"00",
         16091 => x"00",
         16092 => x"00",
         16093 => x"00",
         16094 => x"00",
         16095 => x"00",
         16096 => x"00",
         16097 => x"00",
         16098 => x"00",
         16099 => x"00",
         16100 => x"00",
         16101 => x"00",
         16102 => x"00",
         16103 => x"00",
         16104 => x"00",
         16105 => x"00",
         16106 => x"00",
         16107 => x"00",
         16108 => x"00",
         16109 => x"00",
         16110 => x"00",
         16111 => x"00",
         16112 => x"00",
         16113 => x"00",
         16114 => x"00",
         16115 => x"00",
         16116 => x"00",
         16117 => x"f8",
         16118 => x"00",
         16119 => x"f3",
         16120 => x"00",
         16121 => x"f4",
         16122 => x"00",
         16123 => x"f1",
         16124 => x"00",
         16125 => x"f2",
         16126 => x"00",
         16127 => x"80",
         16128 => x"00",
         16129 => x"81",
         16130 => x"00",
         16131 => x"82",
         16132 => x"00",
         16133 => x"83",
         16134 => x"00",
         16135 => x"84",
         16136 => x"00",
         16137 => x"85",
         16138 => x"00",
         16139 => x"86",
         16140 => x"00",
         16141 => x"87",
         16142 => x"00",
         16143 => x"88",
         16144 => x"00",
         16145 => x"89",
         16146 => x"00",
         16147 => x"f6",
         16148 => x"00",
         16149 => x"7f",
         16150 => x"00",
         16151 => x"f9",
         16152 => x"00",
         16153 => x"e0",
         16154 => x"00",
         16155 => x"e1",
         16156 => x"00",
         16157 => x"71",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"00",
         16166 => x"00",
         16167 => x"00",
         16168 => x"00",
         16169 => x"00",
         16170 => x"00",
         16171 => x"00",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"00",
         18159 => x"50",
         18160 => x"00",
         18161 => x"cc",
         18162 => x"ce",
         18163 => x"f8",
         18164 => x"fc",
         18165 => x"e1",
         18166 => x"c4",
         18167 => x"e3",
         18168 => x"eb",
         18169 => x"00",
         18170 => x"64",
         18171 => x"68",
         18172 => x"2f",
         18173 => x"20",
         18174 => x"24",
         18175 => x"28",
         18176 => x"51",
         18177 => x"55",
         18178 => x"04",
         18179 => x"08",
         18180 => x"0c",
         18181 => x"10",
         18182 => x"14",
         18183 => x"18",
         18184 => x"59",
         18185 => x"c7",
         18186 => x"84",
         18187 => x"88",
         18188 => x"8c",
         18189 => x"90",
         18190 => x"94",
         18191 => x"98",
         18192 => x"80",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"00",
         18199 => x"00",
         18200 => x"00",
         18201 => x"00",
         18202 => x"00",
         18203 => x"00",
         18204 => x"00",
         18205 => x"00",
         18206 => x"00",
         18207 => x"00",
         18208 => x"00",
         18209 => x"00",
         18210 => x"00",
         18211 => x"00",
         18212 => x"00",
         18213 => x"00",
         18214 => x"00",
         18215 => x"00",
         18216 => x"00",
         18217 => x"00",
         18218 => x"00",
         18219 => x"00",
         18220 => x"00",
         18221 => x"00",
         18222 => x"00",
         18223 => x"00",
         18224 => x"00",
         18225 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
