---------------------------------------------------------------------------------------------------------
--
-- Name:            ChrGenRAM_DP_3208.vhd
-- Created:         Jan 2021
-- Author(s):       Philip Smart
-- Description:     Character Generator ROM/RAM for the Sharp MZ series Video Controller Core.
--                                                     
--                  This module provides a dual port inferred RAM definition (for use as ROM/RAM) for use
--                  as Character Generator ROM/RAM in the Video Controller. Port A allows 8/16/32 bit access,
--                  Port B allows for 8 bit access. The size of the RAM is declared in the generic attribute
--                  'addrbits'.
--
-- Credits:         
-- Copyright:       (c) 2018-21 Philip Smart <philip.smart@net2net.org>
--
-- History:         Jan 2021  - Initial creation.
--
---------------------------------------------------------------------------------------------------------
-- This source file is free software: you can redistribute it and-or modify
-- it under the terms of the GNU General Public License as published
-- by the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This source file is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http:--www.gnu.org-licenses->.
---------------------------------------------------------------------------------------------------------
-- Byte Addressed 32bit Port A, 8bit Port B BRAM module for the Video
-- Controller Graphics RAM implementation.
--
-- Copyright 2018-2021 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library altera;
library altera_mf;
library pkgs;
use     ieee.std_logic_1164.all;
use     ieee.std_logic_unsigned.all;
use     ieee.numeric_std.all;
use     work.VideoController_pkg.all;
use     altera.altera_syn_attributes.all;
use     altera_mf.all;

entity ChrGenRAM_DP_3208 is
    generic
    (
        addrbits             : integer := 16                                  -- Max address bit, size in bytes.
    );
    port
    (
        clkA                 : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(31 downto 0);
        memARead             : out std_logic_vector(31 downto 0);

        clkB                 : in  std_logic;
        memBAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memBWriteEnable      : in  std_logic;
        memBWrite            : in  std_logic_vector(7 downto 0);
        memBRead             : out std_logic_vector(7 downto 0)
    );
end ChrGenRAM_DP_3208;

architecture arch of ChrGenRAM_DP_3208 is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0     : ramArray :=
    (
             0 => x"00",
             1 => x"00",
             2 => x"18",
             3 => x"42",
             4 => x"7c",
             5 => x"22",
             6 => x"1c",
             7 => x"40",
             8 => x"78",
             9 => x"22",
            10 => x"7e",
            11 => x"40",
            12 => x"7e",
            13 => x"40",
            14 => x"1c",
            15 => x"42",
            16 => x"42",
            17 => x"42",
            18 => x"1c",
            19 => x"08",
            20 => x"0e",
            21 => x"04",
            22 => x"42",
            23 => x"48",
            24 => x"40",
            25 => x"40",
            26 => x"42",
            27 => x"42",
            28 => x"42",
            29 => x"46",
            30 => x"18",
            31 => x"42",
            32 => x"7c",
            33 => x"40",
            34 => x"18",
            35 => x"4a",
            36 => x"7c",
            37 => x"48",
            38 => x"3c",
            39 => x"02",
            40 => x"3e",
            41 => x"08",
            42 => x"42",
            43 => x"42",
            44 => x"42",
            45 => x"24",
            46 => x"42",
            47 => x"5a",
            48 => x"42",
            49 => x"24",
            50 => x"22",
            51 => x"08",
            52 => x"7e",
            53 => x"20",
            54 => x"0c",
            55 => x"10",
            56 => x"08",
            57 => x"0f",
            58 => x"08",
            59 => x"f8",
            60 => x"08",
            61 => x"0f",
            62 => x"08",
            63 => x"ff",
            64 => x"3c",
            65 => x"62",
            66 => x"08",
            67 => x"08",
            68 => x"3c",
            69 => x"30",
            70 => x"3c",
            71 => x"02",
            72 => x"04",
            73 => x"7e",
            74 => x"7e",
            75 => x"02",
            76 => x"1c",
            77 => x"42",
            78 => x"7e",
            79 => x"10",
            80 => x"3c",
            81 => x"42",
            82 => x"3c",
            83 => x"02",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"7e",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"10",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"40",
            99 => x"40",
           100 => x"80",
           101 => x"80",
           102 => x"01",
           103 => x"01",
           104 => x"00",
           105 => x"00",
           106 => x"10",
           107 => x"10",
           108 => x"ff",
           109 => x"00",
           110 => x"c0",
           111 => x"c0",
           112 => x"00",
           113 => x"00",
           114 => x"04",
           115 => x"04",
           116 => x"00",
           117 => x"ff",
           118 => x"0f",
           119 => x"0f",
           120 => x"00",
           121 => x"00",
           122 => x"01",
           123 => x"01",
           124 => x"00",
           125 => x"00",
           126 => x"03",
           127 => x"03",
           128 => x"10",
           129 => x"08",
           130 => x"08",
           131 => x"7f",
           132 => x"ff",
           133 => x"0f",
           134 => x"ff",
           135 => x"ff",
           136 => x"08",
           137 => x"3e",
           138 => x"00",
           139 => x"7f",
           140 => x"1c",
           141 => x"6b",
           142 => x"00",
           143 => x"7e",
           144 => x"00",
           145 => x"42",
           146 => x"3c",
           147 => x"10",
           148 => x"ff",
           149 => x"81",
           150 => x"00",
           151 => x"03",
           152 => x"00",
           153 => x"c0",
           154 => x"80",
           155 => x"f8",
           156 => x"01",
           157 => x"1f",
           158 => x"00",
           159 => x"00",
           160 => x"00",
           161 => x"08",
           162 => x"0e",
           163 => x"30",
           164 => x"3c",
           165 => x"20",
           166 => x"36",
           167 => x"3e",
           168 => x"3c",
           169 => x"04",
           170 => x"1c",
           171 => x"4c",
           172 => x"ff",
           173 => x"f0",
           174 => x"70",
           175 => x"0c",
           176 => x"00",
           177 => x"2a",
           178 => x"00",
           179 => x"08",
           180 => x"00",
           181 => x"7f",
           182 => x"f0",
           183 => x"0f",
           184 => x"00",
           185 => x"0f",
           186 => x"00",
           187 => x"f8",
           188 => x"08",
           189 => x"f8",
           190 => x"00",
           191 => x"ff",
           192 => x"00",
           193 => x"54",
           194 => x"08",
           195 => x"00",
           196 => x"24",
           197 => x"00",
           198 => x"24",
           199 => x"7e",
           200 => x"08",
           201 => x"0a",
           202 => x"00",
           203 => x"10",
           204 => x"30",
           205 => x"4a",
           206 => x"04",
           207 => x"00",
           208 => x"04",
           209 => x"10",
           210 => x"20",
           211 => x"08",
           212 => x"00",
           213 => x"08",
           214 => x"08",
           215 => x"1c",
           216 => x"0f",
           217 => x"f0",
           218 => x"81",
           219 => x"18",
           220 => x"10",
           221 => x"00",
           222 => x"08",
           223 => x"00",
           224 => x"ff",
           225 => x"00",
           226 => x"80",
           227 => x"80",
           228 => x"ff",
           229 => x"80",
           230 => x"ff",
           231 => x"01",
           232 => x"00",
           233 => x"00",
           234 => x"20",
           235 => x"20",
           236 => x"01",
           237 => x"10",
           238 => x"80",
           239 => x"08",
           240 => x"00",
           241 => x"ff",
           242 => x"08",
           243 => x"08",
           244 => x"ff",
           245 => x"00",
           246 => x"f0",
           247 => x"f0",
           248 => x"00",
           249 => x"00",
           250 => x"02",
           251 => x"02",
           252 => x"00",
           253 => x"00",
           254 => x"07",
           255 => x"07",
           256 => x"18",
           257 => x"18",
           258 => x"00",
           259 => x"3c",
           260 => x"40",
           261 => x"42",
           262 => x"00",
           263 => x"40",
           264 => x"02",
           265 => x"42",
           266 => x"00",
           267 => x"7e",
           268 => x"0c",
           269 => x"10",
           270 => x"00",
           271 => x"46",
           272 => x"40",
           273 => x"42",
           274 => x"08",
           275 => x"08",
           276 => x"04",
           277 => x"04",
           278 => x"40",
           279 => x"50",
           280 => x"18",
           281 => x"08",
           282 => x"00",
           283 => x"49",
           284 => x"00",
           285 => x"42",
           286 => x"00",
           287 => x"42",
           288 => x"00",
           289 => x"62",
           290 => x"00",
           291 => x"46",
           292 => x"00",
           293 => x"40",
           294 => x"00",
           295 => x"3c",
           296 => x"10",
           297 => x"10",
           298 => x"00",
           299 => x"42",
           300 => x"00",
           301 => x"42",
           302 => x"00",
           303 => x"49",
           304 => x"00",
           305 => x"10",
           306 => x"00",
           307 => x"46",
           308 => x"00",
           309 => x"18",
           310 => x"24",
           311 => x"3c",
           312 => x"00",
           313 => x"02",
           314 => x"03",
           315 => x"00",
           316 => x"c0",
           317 => x"00",
           318 => x"00",
           319 => x"40",
           320 => x"00",
           321 => x"c0",
           322 => x"00",
           323 => x"00",
           324 => x"44",
           325 => x"44",
           326 => x"44",
           327 => x"44",
           328 => x"20",
           329 => x"00",
           330 => x"00",
           331 => x"4c",
           332 => x"aa",
           333 => x"aa",
           334 => x"00",
           335 => x"03",
           336 => x"03",
           337 => x"00",
           338 => x"c0",
           339 => x"00",
           340 => x"38",
           341 => x"42",
           342 => x"00",
           343 => x"22",
           344 => x"00",
           345 => x"22",
           346 => x"42",
           347 => x"42",
           348 => x"42",
           349 => x"7e",
           350 => x"42",
           351 => x"42",
           352 => x"10",
           353 => x"40",
           354 => x"01",
           355 => x"20",
           356 => x"80",
           357 => x"04",
           358 => x"08",
           359 => x"02",
           360 => x"80",
           361 => x"40",
           362 => x"80",
           363 => x"20",
           364 => x"01",
           365 => x"04",
           366 => x"01",
           367 => x"02",
           368 => x"10",
           369 => x"01",
           370 => x"00",
           371 => x"80",
           372 => x"00",
           373 => x"01",
           374 => x"08",
           375 => x"80",
           376 => x"08",
           377 => x"10",
           378 => x"08",
           379 => x"ff",
           380 => x"08",
           381 => x"00",
           382 => x"00",
           383 => x"00",
           384 => x"1c",
           385 => x"08",
           386 => x"ff",
           387 => x"d5",
           388 => x"ff",
           389 => x"f7",
           390 => x"ff",
           391 => x"81",
           392 => x"ff",
           393 => x"81",
           394 => x"bd",
           395 => x"bd",
           396 => x"e3",
           397 => x"bf",
           398 => x"18",
           399 => x"5a",
           400 => x"e0",
           401 => x"42",
           402 => x"22",
           403 => x"08",
           404 => x"1c",
           405 => x"08",
           406 => x"00",
           407 => x"d2",
           408 => x"00",
           409 => x"4b",
           410 => x"22",
           411 => x"3e",
           412 => x"3c",
           413 => x"ff",
           414 => x"3c",
           415 => x"81",
           416 => x"aa",
           417 => x"aa",
           418 => x"0a",
           419 => x"0a",
           420 => x"a0",
           421 => x"a0",
           422 => x"aa",
           423 => x"00",
           424 => x"00",
           425 => x"aa",
           426 => x"aa",
           427 => x"a0",
           428 => x"aa",
           429 => x"0a",
           430 => x"80",
           431 => x"a8",
           432 => x"00",
           433 => x"0a",
           434 => x"80",
           435 => x"20",
           436 => x"08",
           437 => x"02",
           438 => x"38",
           439 => x"00",
           440 => x"00",
           441 => x"2a",
           442 => x"01",
           443 => x"04",
           444 => x"10",
           445 => x"40",
           446 => x"00",
           447 => x"54",
           448 => x"00",
           449 => x"00",
           450 => x"02",
           451 => x"02",
           452 => x"02",
           453 => x"02",
           454 => x"00",
           455 => x"88",
           456 => x"00",
           457 => x"c4",
           458 => x"11",
           459 => x"11",
           460 => x"00",
           461 => x"23",
           462 => x"00",
           463 => x"8f",
           464 => x"00",
           465 => x"f1",
           466 => x"88",
           467 => x"c0",
           468 => x"a8",
           469 => x"c0",
           470 => x"80",
           471 => x"1f",
           472 => x"00",
           473 => x"e7",
           474 => x"08",
           475 => x"00",
           476 => x"08",
           477 => x"08",
           478 => x"55",
           479 => x"55",
           480 => x"00",
           481 => x"00",
           482 => x"00",
           483 => x"00",
           484 => x"00",
           485 => x"00",
           486 => x"00",
           487 => x"00",
           488 => x"00",
           489 => x"00",
           490 => x"00",
           491 => x"00",
           492 => x"00",
           493 => x"00",
           494 => x"00",
           495 => x"00",
           496 => x"00",
           497 => x"00",
           498 => x"00",
           499 => x"00",
           500 => x"00",
           501 => x"00",
           502 => x"00",
           503 => x"00",
           504 => x"00",
           505 => x"00",
           506 => x"00",
           507 => x"00",
           508 => x"00",
           509 => x"00",
           510 => x"00",
           511 => x"00",
           512 => x"00",
           513 => x"00",
           514 => x"7c",
           515 => x"82",
           516 => x"fc",
           517 => x"ba",
           518 => x"7e",
           519 => x"a0",
           520 => x"f8",
           521 => x"aa",
           522 => x"fe",
           523 => x"88",
           524 => x"fe",
           525 => x"b8",
           526 => x"7e",
           527 => x"ae",
           528 => x"ee",
           529 => x"ba",
           530 => x"fe",
           531 => x"28",
           532 => x"1f",
           533 => x"ea",
           534 => x"e6",
           535 => x"88",
           536 => x"e0",
           537 => x"a0",
           538 => x"fe",
           539 => x"ba",
           540 => x"ee",
           541 => x"b2",
           542 => x"7c",
           543 => x"aa",
           544 => x"fc",
           545 => x"86",
           546 => x"7c",
           547 => x"aa",
           548 => x"fc",
           549 => x"84",
           550 => x"7e",
           551 => x"7a",
           552 => x"fe",
           553 => x"28",
           554 => x"ee",
           555 => x"aa",
           556 => x"ee",
           557 => x"aa",
           558 => x"ee",
           559 => x"aa",
           560 => x"c6",
           561 => x"28",
           562 => x"ee",
           563 => x"28",
           564 => x"fe",
           565 => x"28",
           566 => x"00",
           567 => x"ff",
           568 => x"00",
           569 => x"ff",
           570 => x"00",
           571 => x"38",
           572 => x"92",
           573 => x"38",
           574 => x"00",
           575 => x"fe",
           576 => x"7c",
           577 => x"aa",
           578 => x"38",
           579 => x"28",
           580 => x"7c",
           581 => x"14",
           582 => x"fc",
           583 => x"22",
           584 => x"0c",
           585 => x"b6",
           586 => x"fe",
           587 => x"7a",
           588 => x"7e",
           589 => x"82",
           590 => x"fe",
           591 => x"28",
           592 => x"7c",
           593 => x"82",
           594 => x"7c",
           595 => x"7a",
           596 => x"f8",
           597 => x"fa",
           598 => x"1f",
           599 => x"5f",
           600 => x"3c",
           601 => x"7e",
           602 => x"3c",
           603 => x"7e",
           604 => x"08",
           605 => x"77",
           606 => x"08",
           607 => x"77",
           608 => x"41",
           609 => x"7e",
           610 => x"82",
           611 => x"7e",
           612 => x"00",
           613 => x"24",
           614 => x"81",
           615 => x"18",
           616 => x"00",
           617 => x"7e",
           618 => x"24",
           619 => x"24",
           620 => x"3c",
           621 => x"d5",
           622 => x"3c",
           623 => x"d5",
           624 => x"3c",
           625 => x"99",
           626 => x"3c",
           627 => x"99",
           628 => x"42",
           629 => x"ff",
           630 => x"1c",
           631 => x"0f",
           632 => x"3c",
           633 => x"e7",
           634 => x"38",
           635 => x"f0",
           636 => x"3c",
           637 => x"ff",
           638 => x"10",
           639 => x"28",
           640 => x"00",
           641 => x"c7",
           642 => x"6b",
           643 => x"14",
           644 => x"00",
           645 => x"e3",
           646 => x"3c",
           647 => x"3c",
           648 => x"3c",
           649 => x"3c",
           650 => x"3c",
           651 => x"3c",
           652 => x"7e",
           653 => x"24",
           654 => x"7e",
           655 => x"24",
           656 => x"7e",
           657 => x"24",
           658 => x"22",
           659 => x"ff",
           660 => x"38",
           661 => x"0f",
           662 => x"3c",
           663 => x"ed",
           664 => x"1c",
           665 => x"f0",
           666 => x"3c",
           667 => x"ff",
           668 => x"3c",
           669 => x"fd",
           670 => x"1c",
           671 => x"ff",
           672 => x"38",
           673 => x"ff",
           674 => x"18",
           675 => x"3c",
           676 => x"00",
           677 => x"ff",
           678 => x"3c",
           679 => x"3c",
           680 => x"00",
           681 => x"ff",
           682 => x"20",
           683 => x"30",
           684 => x"00",
           685 => x"07",
           686 => x"3c",
           687 => x"04",
           688 => x"00",
           689 => x"e0",
           690 => x"10",
           691 => x"92",
           692 => x"00",
           693 => x"ff",
           694 => x"38",
           695 => x"7c",
           696 => x"00",
           697 => x"ff",
           698 => x"00",
           699 => x"48",
           700 => x"00",
           701 => x"50",
           702 => x"00",
           703 => x"0a",
           704 => x"00",
           705 => x"12",
           706 => x"18",
           707 => x"c3",
           708 => x"1f",
           709 => x"f0",
           710 => x"81",
           711 => x"ff",
           712 => x"f8",
           713 => x"0f",
           714 => x"bf",
           715 => x"a5",
           716 => x"ff",
           717 => x"85",
           718 => x"ff",
           719 => x"a5",
           720 => x"ff",
           721 => x"a5",
           722 => x"00",
           723 => x"00",
           724 => x"01",
           725 => x"55",
           726 => x"ff",
           727 => x"3c",
           728 => x"80",
           729 => x"aa",
           730 => x"00",
           731 => x"00",
           732 => x"00",
           733 => x"77",
           734 => x"00",
           735 => x"00",
           736 => x"00",
           737 => x"77",
           738 => x"00",
           739 => x"e7",
           740 => x"10",
           741 => x"10",
           742 => x"00",
           743 => x"ff",
           744 => x"7f",
           745 => x"08",
           746 => x"55",
           747 => x"55",
           748 => x"ff",
           749 => x"ff",
           750 => x"a5",
           751 => x"00",
           752 => x"24",
           753 => x"00",
           754 => x"ff",
           755 => x"a0",
           756 => x"ff",
           757 => x"15",
           758 => x"00",
           759 => x"a0",
           760 => x"00",
           761 => x"41",
           762 => x"a0",
           763 => x"30",
           764 => x"11",
           765 => x"0c",
           766 => x"80",
           767 => x"80",
           768 => x"01",
           769 => x"01",
           770 => x"3c",
           771 => x"10",
           772 => x"00",
           773 => x"24",
           774 => x"00",
           775 => x"42",
           776 => x"3c",
           777 => x"81",
           778 => x"00",
           779 => x"18",
           780 => x"00",
           781 => x"3c",
           782 => x"00",
           783 => x"7e",
           784 => x"3c",
           785 => x"a1",
           786 => x"ff",
           787 => x"e7",
           788 => x"ff",
           789 => x"c3",
           790 => x"ff",
           791 => x"81",
           792 => x"20",
           793 => x"ff",
           794 => x"3c",
           795 => x"ff",
           796 => x"3c",
           797 => x"99",
           798 => x"3c",
           799 => x"ff",
           800 => x"00",
           801 => x"fe",
           802 => x"0f",
           803 => x"8a",
           804 => x"f0",
           805 => x"51",
           806 => x"0f",
           807 => x"8e",
           808 => x"f0",
           809 => x"71",
           810 => x"81",
           811 => x"43",
           812 => x"81",
           813 => x"c2",
           814 => x"81",
           815 => x"40",
           816 => x"81",
           817 => x"02",
           818 => x"81",
           819 => x"43",
           820 => x"81",
           821 => x"c2",
           822 => x"81",
           823 => x"48",
           824 => x"81",
           825 => x"12",
           826 => x"08",
           827 => x"fe",
           828 => x"00",
           829 => x"30",
           830 => x"00",
           831 => x"60",
           832 => x"91",
           833 => x"c0",
           834 => x"80",
           835 => x"ff",
           836 => x"00",
           837 => x"ff",
           838 => x"00",
           839 => x"ff",
           840 => x"00",
           841 => x"fc",
           842 => x"01",
           843 => x"ff",
           844 => x"02",
           845 => x"14",
           846 => x"00",
           847 => x"10",
           848 => x"00",
           849 => x"3f",
           850 => x"00",
           851 => x"10",
           852 => x"00",
           853 => x"42",
           854 => x"00",
           855 => x"92",
           856 => x"00",
           857 => x"92",
           858 => x"00",
           859 => x"90",
           860 => x"00",
           861 => x"50",
           862 => x"00",
           863 => x"7c",
           864 => x"00",
           865 => x"55",
           866 => x"ff",
           867 => x"a3",
           868 => x"ff",
           869 => x"99",
           870 => x"00",
           871 => x"ee",
           872 => x"ff",
           873 => x"ff",
           874 => x"92",
           875 => x"10",
           876 => x"38",
           877 => x"38",
           878 => x"00",
           879 => x"ff",
           880 => x"00",
           881 => x"10",
           882 => x"7e",
           883 => x"7e",
           884 => x"00",
           885 => x"55",
           886 => x"00",
           887 => x"b0",
           888 => x"00",
           889 => x"0d",
           890 => x"00",
           891 => x"3c",
           892 => x"ff",
           893 => x"00",
           894 => x"c0",
           895 => x"f0",
           896 => x"03",
           897 => x"0f",
           898 => x"03",
           899 => x"ff",
           900 => x"c0",
           901 => x"ee",
           902 => x"0e",
           903 => x"01",
           904 => x"7a",
           905 => x"f4",
           906 => x"04",
           907 => x"6f",
           908 => x"20",
           909 => x"f6",
           910 => x"3b",
           911 => x"10",
           912 => x"dc",
           913 => x"08",
           914 => x"01",
           915 => x"0e",
           916 => x"80",
           917 => x"70",
           918 => x"1e",
           919 => x"03",
           920 => x"78",
           921 => x"c0",
           922 => x"01",
           923 => x"8c",
           924 => x"80",
           925 => x"31",
           926 => x"3f",
           927 => x"0f",
           928 => x"fc",
           929 => x"f0",
           930 => x"00",
           931 => x"02",
           932 => x"00",
           933 => x"40",
           934 => x"02",
           935 => x"1f",
           936 => x"40",
           937 => x"f8",
           938 => x"73",
           939 => x"3f",
           940 => x"ce",
           941 => x"fc",
           942 => x"0f",
           943 => x"7f",
           944 => x"f0",
           945 => x"fe",
           946 => x"f8",
           947 => x"21",
           948 => x"ff",
           949 => x"00",
           950 => x"fc",
           951 => x"81",
           952 => x"00",
           953 => x"7f",
           954 => x"00",
           955 => x"ff",
           956 => x"01",
           957 => x"ff",
           958 => x"ff",
           959 => x"80",
           960 => x"00",
           961 => x"80",
           962 => x"00",
           963 => x"f9",
           964 => x"00",
           965 => x"e9",
           966 => x"1f",
           967 => x"88",
           968 => x"40",
           969 => x"09",
           970 => x"40",
           971 => x"06",
           972 => x"40",
           973 => x"01",
           974 => x"40",
           975 => x"e1",
           976 => x"c0",
           977 => x"18",
           978 => x"01",
           979 => x"18",
           980 => x"00",
           981 => x"2a",
           982 => x"1b",
           983 => x"c9",
           984 => x"4c",
           985 => x"07",
           986 => x"7f",
           987 => x"81",
           988 => x"88",
           989 => x"88",
           990 => x"40",
           991 => x"40",
           992 => x"00",
           993 => x"ff",
           994 => x"00",
           995 => x"ff",
           996 => x"00",
           997 => x"3f",
           998 => x"00",
           999 => x"fc",
          1000 => x"10",
          1001 => x"fc",
          1002 => x"ba",
          1003 => x"38",
          1004 => x"ba",
          1005 => x"38",
          1006 => x"00",
          1007 => x"9f",
          1008 => x"00",
          1009 => x"f9",
          1010 => x"00",
          1011 => x"7f",
          1012 => x"00",
          1013 => x"fe",
          1014 => x"ff",
          1015 => x"81",
          1016 => x"e7",
          1017 => x"00",
          1018 => x"00",
          1019 => x"10",
          1020 => x"18",
          1021 => x"10",
          1022 => x"08",
          1023 => x"04",
        others => X"00"
    );

    shared variable RAM1     : ramArray :=
    (
             0 => x"00",
             1 => x"00",
             2 => x"24",
             3 => x"42",
             4 => x"22",
             5 => x"22",
             6 => x"22",
             7 => x"22",
             8 => x"24",
             9 => x"24",
            10 => x"40",
            11 => x"40",
            12 => x"40",
            13 => x"40",
            14 => x"22",
            15 => x"22",
            16 => x"42",
            17 => x"42",
            18 => x"08",
            19 => x"08",
            20 => x"04",
            21 => x"44",
            22 => x"44",
            23 => x"44",
            24 => x"40",
            25 => x"40",
            26 => x"66",
            27 => x"42",
            28 => x"62",
            29 => x"42",
            30 => x"24",
            31 => x"24",
            32 => x"42",
            33 => x"40",
            34 => x"24",
            35 => x"24",
            36 => x"42",
            37 => x"44",
            38 => x"42",
            39 => x"42",
            40 => x"08",
            41 => x"08",
            42 => x"42",
            43 => x"42",
            44 => x"42",
            45 => x"18",
            46 => x"42",
            47 => x"66",
            48 => x"42",
            49 => x"42",
            50 => x"22",
            51 => x"08",
            52 => x"02",
            53 => x"40",
            54 => x"12",
            55 => x"10",
            56 => x"08",
            57 => x"00",
            58 => x"08",
            59 => x"00",
            60 => x"08",
            61 => x"08",
            62 => x"08",
            63 => x"00",
            64 => x"42",
            65 => x"42",
            66 => x"18",
            67 => x"08",
            68 => x"42",
            69 => x"40",
            70 => x"42",
            71 => x"42",
            72 => x"0c",
            73 => x"04",
            74 => x"40",
            75 => x"44",
            76 => x"20",
            77 => x"42",
            78 => x"42",
            79 => x"10",
            80 => x"42",
            81 => x"42",
            82 => x"42",
            83 => x"04",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"08",
            90 => x"02",
            91 => x"20",
            92 => x"00",
            93 => x"18",
            94 => x"00",
            95 => x"08",
            96 => x"ff",
            97 => x"00",
            98 => x"40",
            99 => x"40",
           100 => x"80",
           101 => x"80",
           102 => x"01",
           103 => x"01",
           104 => x"00",
           105 => x"00",
           106 => x"10",
           107 => x"10",
           108 => x"ff",
           109 => x"00",
           110 => x"c0",
           111 => x"c0",
           112 => x"00",
           113 => x"ff",
           114 => x"04",
           115 => x"04",
           116 => x"00",
           117 => x"ff",
           118 => x"0f",
           119 => x"0f",
           120 => x"00",
           121 => x"00",
           122 => x"01",
           123 => x"01",
           124 => x"00",
           125 => x"00",
           126 => x"03",
           127 => x"03",
           128 => x"08",
           129 => x"08",
           130 => x"1c",
           131 => x"1c",
           132 => x"7f",
           133 => x"07",
           134 => x"ff",
           135 => x"ff",
           136 => x"1c",
           137 => x"1c",
           138 => x"00",
           139 => x"20",
           140 => x"1c",
           141 => x"08",
           142 => x"3c",
           143 => x"7e",
           144 => x"3c",
           145 => x"42",
           146 => x"42",
           147 => x"00",
           148 => x"c3",
           149 => x"81",
           150 => x"00",
           151 => x"04",
           152 => x"00",
           153 => x"20",
           154 => x"c0",
           155 => x"fc",
           156 => x"03",
           157 => x"3f",
           158 => x"00",
           159 => x"08",
           160 => x"08",
           161 => x"08",
           162 => x"18",
           163 => x"18",
           164 => x"20",
           165 => x"20",
           166 => x"7f",
           167 => x"1c",
           168 => x"04",
           169 => x"04",
           170 => x"22",
           171 => x"20",
           172 => x"fe",
           173 => x"e0",
           174 => x"18",
           175 => x"18",
           176 => x"08",
           177 => x"1c",
           178 => x"40",
           179 => x"04",
           180 => x"00",
           181 => x"02",
           182 => x"f0",
           183 => x"0f",
           184 => x"00",
           185 => x"08",
           186 => x"00",
           187 => x"08",
           188 => x"08",
           189 => x"08",
           190 => x"00",
           191 => x"08",
           192 => x"00",
           193 => x"14",
           194 => x"08",
           195 => x"00",
           196 => x"24",
           197 => x"00",
           198 => x"24",
           199 => x"24",
           200 => x"1e",
           201 => x"1c",
           202 => x"62",
           203 => x"26",
           204 => x"48",
           205 => x"44",
           206 => x"08",
           207 => x"00",
           208 => x"08",
           209 => x"08",
           210 => x"10",
           211 => x"10",
           212 => x"08",
           213 => x"08",
           214 => x"2a",
           215 => x"2a",
           216 => x"0f",
           217 => x"f0",
           218 => x"42",
           219 => x"24",
           220 => x"10",
           221 => x"00",
           222 => x"08",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"80",
           227 => x"80",
           228 => x"80",
           229 => x"80",
           230 => x"01",
           231 => x"01",
           232 => x"00",
           233 => x"00",
           234 => x"20",
           235 => x"20",
           236 => x"02",
           237 => x"20",
           238 => x"40",
           239 => x"04",
           240 => x"00",
           241 => x"00",
           242 => x"08",
           243 => x"08",
           244 => x"ff",
           245 => x"00",
           246 => x"f0",
           247 => x"f0",
           248 => x"00",
           249 => x"00",
           250 => x"02",
           251 => x"02",
           252 => x"00",
           253 => x"ff",
           254 => x"07",
           255 => x"07",
           256 => x"18",
           257 => x"18",
           258 => x"00",
           259 => x"44",
           260 => x"40",
           261 => x"62",
           262 => x"00",
           263 => x"42",
           264 => x"02",
           265 => x"46",
           266 => x"00",
           267 => x"40",
           268 => x"12",
           269 => x"10",
           270 => x"00",
           271 => x"3a",
           272 => x"40",
           273 => x"42",
           274 => x"00",
           275 => x"08",
           276 => x"00",
           277 => x"04",
           278 => x"40",
           279 => x"68",
           280 => x"08",
           281 => x"08",
           282 => x"00",
           283 => x"49",
           284 => x"00",
           285 => x"42",
           286 => x"00",
           287 => x"42",
           288 => x"00",
           289 => x"5c",
           290 => x"00",
           291 => x"3a",
           292 => x"00",
           293 => x"40",
           294 => x"00",
           295 => x"02",
           296 => x"10",
           297 => x"12",
           298 => x"00",
           299 => x"46",
           300 => x"00",
           301 => x"24",
           302 => x"00",
           303 => x"49",
           304 => x"00",
           305 => x"28",
           306 => x"00",
           307 => x"3a",
           308 => x"00",
           309 => x"20",
           310 => x"00",
           311 => x"44",
           312 => x"00",
           313 => x"04",
           314 => x"1c",
           315 => x"00",
           316 => x"38",
           317 => x"00",
           318 => x"00",
           319 => x"20",
           320 => x"00",
           321 => x"30",
           322 => x"ff",
           323 => x"ff",
           324 => x"44",
           325 => x"44",
           326 => x"ff",
           327 => x"ff",
           328 => x"10",
           329 => x"00",
           330 => x"00",
           331 => x"00",
           332 => x"44",
           333 => x"44",
           334 => x"00",
           335 => x"0c",
           336 => x"0c",
           337 => x"00",
           338 => x"30",
           339 => x"00",
           340 => x"44",
           341 => x"52",
           342 => x"22",
           343 => x"26",
           344 => x"22",
           345 => x"22",
           346 => x"00",
           347 => x"42",
           348 => x"18",
           349 => x"42",
           350 => x"18",
           351 => x"24",
           352 => x"20",
           353 => x"40",
           354 => x"06",
           355 => x"40",
           356 => x"60",
           357 => x"02",
           358 => x"04",
           359 => x"02",
           360 => x"80",
           361 => x"20",
           362 => x"40",
           363 => x"18",
           364 => x"02",
           365 => x"18",
           366 => x"01",
           367 => x"04",
           368 => x"08",
           369 => x"00",
           370 => x"00",
           371 => x"60",
           372 => x"00",
           373 => x"06",
           374 => x"10",
           375 => x"00",
           376 => x"10",
           377 => x"10",
           378 => x"08",
           379 => x"08",
           380 => x"14",
           381 => x"00",
           382 => x"00",
           383 => x"00",
           384 => x"1c",
           385 => x"00",
           386 => x"f7",
           387 => x"e3",
           388 => x"f7",
           389 => x"f7",
           390 => x"ff",
           391 => x"fb",
           392 => x"ff",
           393 => x"df",
           394 => x"bd",
           395 => x"bd",
           396 => x"dd",
           397 => x"dd",
           398 => x"24",
           399 => x"24",
           400 => x"47",
           401 => x"47",
           402 => x"3e",
           403 => x"49",
           404 => x"1c",
           405 => x"08",
           406 => x"11",
           407 => x"11",
           408 => x"88",
           409 => x"88",
           410 => x"14",
           411 => x"08",
           412 => x"7e",
           413 => x"e7",
           414 => x"42",
           415 => x"99",
           416 => x"55",
           417 => x"55",
           418 => x"05",
           419 => x"05",
           420 => x"50",
           421 => x"50",
           422 => x"55",
           423 => x"00",
           424 => x"00",
           425 => x"55",
           426 => x"54",
           427 => x"40",
           428 => x"55",
           429 => x"05",
           430 => x"40",
           431 => x"54",
           432 => x"01",
           433 => x"15",
           434 => x"80",
           435 => x"20",
           436 => x"08",
           437 => x"02",
           438 => x"28",
           439 => x"00",
           440 => x"54",
           441 => x"54",
           442 => x"01",
           443 => x"04",
           444 => x"10",
           445 => x"40",
           446 => x"c0",
           447 => x"55",
           448 => x"00",
           449 => x"02",
           450 => x"02",
           451 => x"02",
           452 => x"02",
           453 => x"02",
           454 => x"00",
           455 => x"05",
           456 => x"0e",
           457 => x"04",
           458 => x"22",
           459 => x"22",
           460 => x"70",
           461 => x"20",
           462 => x"c4",
           463 => x"94",
           464 => x"23",
           465 => x"29",
           466 => x"90",
           467 => x"a8",
           468 => x"b0",
           469 => x"a0",
           470 => x"40",
           471 => x"20",
           472 => x"00",
           473 => x"24",
           474 => x"08",
           475 => x"3e",
           476 => x"10",
           477 => x"04",
           478 => x"aa",
           479 => x"aa",
           480 => x"00",
           481 => x"00",
           482 => x"70",
           483 => x"00",
           484 => x"07",
           485 => x"00",
           486 => x"77",
           487 => x"00",
           488 => x"00",
           489 => x"70",
           490 => x"70",
           491 => x"70",
           492 => x"07",
           493 => x"70",
           494 => x"77",
           495 => x"70",
           496 => x"00",
           497 => x"07",
           498 => x"70",
           499 => x"07",
           500 => x"07",
           501 => x"07",
           502 => x"77",
           503 => x"07",
           504 => x"00",
           505 => x"77",
           506 => x"70",
           507 => x"77",
           508 => x"07",
           509 => x"77",
           510 => x"77",
           511 => x"77",
           512 => x"00",
           513 => x"00",
           514 => x"c6",
           515 => x"ba",
           516 => x"86",
           517 => x"ba",
           518 => x"c2",
           519 => x"be",
           520 => x"8c",
           521 => x"b6",
           522 => x"82",
           523 => x"be",
           524 => x"82",
           525 => x"a0",
           526 => x"82",
           527 => x"ba",
           528 => x"aa",
           529 => x"aa",
           530 => x"82",
           531 => x"ee",
           532 => x"11",
           533 => x"ba",
           534 => x"aa",
           535 => x"b4",
           536 => x"a0",
           537 => x"be",
           538 => x"82",
           539 => x"aa",
           540 => x"9a",
           541 => x"aa",
           542 => x"c6",
           543 => x"ba",
           544 => x"86",
           545 => x"bc",
           546 => x"c6",
           547 => x"b2",
           548 => x"86",
           549 => x"b4",
           550 => x"c2",
           551 => x"fa",
           552 => x"82",
           553 => x"28",
           554 => x"aa",
           555 => x"ba",
           556 => x"aa",
           557 => x"54",
           558 => x"aa",
           559 => x"aa",
           560 => x"aa",
           561 => x"54",
           562 => x"aa",
           563 => x"28",
           564 => x"82",
           565 => x"5e",
           566 => x"40",
           567 => x"7e",
           568 => x"02",
           569 => x"7e",
           570 => x"7c",
           571 => x"54",
           572 => x"54",
           573 => x"54",
           574 => x"00",
           575 => x"00",
           576 => x"82",
           577 => x"9a",
           578 => x"48",
           579 => x"6c",
           580 => x"82",
           581 => x"2e",
           582 => x"82",
           583 => x"fa",
           584 => x"14",
           585 => x"82",
           586 => x"82",
           587 => x"fa",
           588 => x"82",
           589 => x"ba",
           590 => x"82",
           591 => x"50",
           592 => x"82",
           593 => x"ba",
           594 => x"82",
           595 => x"fa",
           596 => x"88",
           597 => x"22",
           598 => x"11",
           599 => x"44",
           600 => x"5a",
           601 => x"24",
           602 => x"5a",
           603 => x"24",
           604 => x"1c",
           605 => x"3e",
           606 => x"1c",
           607 => x"3e",
           608 => x"a2",
           609 => x"ff",
           610 => x"45",
           611 => x"ff",
           612 => x"5a",
           613 => x"42",
           614 => x"a5",
           615 => x"24",
           616 => x"24",
           617 => x"24",
           618 => x"7e",
           619 => x"42",
           620 => x"5a",
           621 => x"ff",
           622 => x"5a",
           623 => x"ff",
           624 => x"42",
           625 => x"81",
           626 => x"42",
           627 => x"81",
           628 => x"42",
           629 => x"ff",
           630 => x"fe",
           631 => x"3f",
           632 => x"7e",
           633 => x"66",
           634 => x"7f",
           635 => x"fc",
           636 => x"7e",
           637 => x"ff",
           638 => x"38",
           639 => x"7c",
           640 => x"03",
           641 => x"7e",
           642 => x"7f",
           643 => x"14",
           644 => x"c0",
           645 => x"7e",
           646 => x"0c",
           647 => x"76",
           648 => x"24",
           649 => x"5a",
           650 => x"30",
           651 => x"6e",
           652 => x"7e",
           653 => x"24",
           654 => x"7e",
           655 => x"24",
           656 => x"7e",
           657 => x"24",
           658 => x"63",
           659 => x"7e",
           660 => x"6c",
           661 => x"3f",
           662 => x"3c",
           663 => x"ef",
           664 => x"36",
           665 => x"fc",
           666 => x"7e",
           667 => x"7e",
           668 => x"3c",
           669 => x"ff",
           670 => x"36",
           671 => x"ff",
           672 => x"6c",
           673 => x"ff",
           674 => x"3c",
           675 => x"18",
           676 => x"00",
           677 => x"7b",
           678 => x"3c",
           679 => x"3c",
           680 => x"00",
           681 => x"de",
           682 => x"60",
           683 => x"28",
           684 => x"40",
           685 => x"03",
           686 => x"3c",
           687 => x"04",
           688 => x"02",
           689 => x"c0",
           690 => x"10",
           691 => x"10",
           692 => x"08",
           693 => x"31",
           694 => x"10",
           695 => x"38",
           696 => x"10",
           697 => x"8c",
           698 => x"78",
           699 => x"04",
           700 => x"02",
           701 => x"60",
           702 => x"40",
           703 => x"06",
           704 => x"1e",
           705 => x"20",
           706 => x"7e",
           707 => x"81",
           708 => x"78",
           709 => x"70",
           710 => x"81",
           711 => x"7e",
           712 => x"1e",
           713 => x"0e",
           714 => x"a1",
           715 => x"bd",
           716 => x"81",
           717 => x"fd",
           718 => x"81",
           719 => x"b5",
           720 => x"80",
           721 => x"bd",
           722 => x"18",
           723 => x"7e",
           724 => x"05",
           725 => x"15",
           726 => x"00",
           727 => x"00",
           728 => x"a0",
           729 => x"a8",
           730 => x"08",
           731 => x"08",
           732 => x"00",
           733 => x"33",
           734 => x"3e",
           735 => x"3e",
           736 => x"00",
           737 => x"66",
           738 => x"00",
           739 => x"00",
           740 => x"38",
           741 => x"54",
           742 => x"00",
           743 => x"42",
           744 => x"41",
           745 => x"08",
           746 => x"55",
           747 => x"55",
           748 => x"00",
           749 => x"00",
           750 => x"42",
           751 => x"a5",
           752 => x"42",
           753 => x"81",
           754 => x"80",
           755 => x"a0",
           756 => x"01",
           757 => x"11",
           758 => x"00",
           759 => x"af",
           760 => x"00",
           761 => x"41",
           762 => x"9f",
           763 => x"30",
           764 => x"e1",
           765 => x"0c",
           766 => x"aa",
           767 => x"8f",
           768 => x"a9",
           769 => x"e1",
           770 => x"42",
           771 => x"10",
           772 => x"00",
           773 => x"18",
           774 => x"18",
           775 => x"24",
           776 => x"42",
           777 => x"81",
           778 => x"00",
           779 => x"00",
           780 => x"00",
           781 => x"3c",
           782 => x"7e",
           783 => x"7e",
           784 => x"42",
           785 => x"9d",
           786 => x"ff",
           787 => x"ff",
           788 => x"ff",
           789 => x"c3",
           790 => x"81",
           791 => x"81",
           792 => x"30",
           793 => x"7e",
           794 => x"42",
           795 => x"81",
           796 => x"5a",
           797 => x"99",
           798 => x"5a",
           799 => x"99",
           800 => x"28",
           801 => x"54",
           802 => x"30",
           803 => x"8e",
           804 => x"0c",
           805 => x"71",
           806 => x"30",
           807 => x"80",
           808 => x"0c",
           809 => x"01",
           810 => x"80",
           811 => x"40",
           812 => x"01",
           813 => x"02",
           814 => x"80",
           815 => x"40",
           816 => x"01",
           817 => x"02",
           818 => x"80",
           819 => x"40",
           820 => x"01",
           821 => x"02",
           822 => x"80",
           823 => x"40",
           824 => x"01",
           825 => x"02",
           826 => x"10",
           827 => x"fe",
           828 => x"06",
           829 => x"78",
           830 => x"52",
           831 => x"2c",
           832 => x"52",
           833 => x"00",
           834 => x"c0",
           835 => x"ff",
           836 => x"00",
           837 => x"c3",
           838 => x"00",
           839 => x"c3",
           840 => x"c0",
           841 => x"fe",
           842 => x"03",
           843 => x"ff",
           844 => x"14",
           845 => x"14",
           846 => x"fe",
           847 => x"20",
           848 => x"03",
           849 => x"7f",
           850 => x"20",
           851 => x"28",
           852 => x"3c",
           853 => x"24",
           854 => x"44",
           855 => x"6c",
           856 => x"00",
           857 => x"6c",
           858 => x"02",
           859 => x"6e",
           860 => x"1e",
           861 => x"b0",
           862 => x"00",
           863 => x"00",
           864 => x"f1",
           865 => x"51",
           866 => x"89",
           867 => x"89",
           868 => x"c3",
           869 => x"a5",
           870 => x"92",
           871 => x"38",
           872 => x"99",
           873 => x"99",
           874 => x"54",
           875 => x"10",
           876 => x"10",
           877 => x"10",
           878 => x"00",
           879 => x"aa",
           880 => x"10",
           881 => x"10",
           882 => x"42",
           883 => x"42",
           884 => x"ff",
           885 => x"55",
           886 => x"00",
           887 => x"8c",
           888 => x"00",
           889 => x"31",
           890 => x"00",
           891 => x"7e",
           892 => x"ff",
           893 => x"00",
           894 => x"e0",
           895 => x"f0",
           896 => x"07",
           897 => x"0f",
           898 => x"0c",
           899 => x"7f",
           900 => x"30",
           901 => x"f6",
           902 => x"0e",
           903 => x"01",
           904 => x"74",
           905 => x"fa",
           906 => x"4e",
           907 => x"7f",
           908 => x"72",
           909 => x"fe",
           910 => x"31",
           911 => x"1f",
           912 => x"8c",
           913 => x"f8",
           914 => x"03",
           915 => x"3e",
           916 => x"c0",
           917 => x"7c",
           918 => x"0e",
           919 => x"37",
           920 => x"70",
           921 => x"ec",
           922 => x"33",
           923 => x"df",
           924 => x"cc",
           925 => x"fb",
           926 => x"1f",
           927 => x"7f",
           928 => x"f8",
           929 => x"fe",
           930 => x"01",
           931 => x"01",
           932 => x"80",
           933 => x"80",
           934 => x"02",
           935 => x"20",
           936 => x"40",
           937 => x"04",
           938 => x"73",
           939 => x"1f",
           940 => x"ce",
           941 => x"f8",
           942 => x"0f",
           943 => x"40",
           944 => x"f0",
           945 => x"02",
           946 => x"44",
           947 => x"42",
           948 => x"05",
           949 => x"07",
           950 => x"86",
           951 => x"82",
           952 => x"00",
           953 => x"80",
           954 => x"00",
           955 => x"01",
           956 => x"01",
           957 => x"00",
           958 => x"80",
           959 => x"00",
           960 => x"00",
           961 => x"80",
           962 => x"08",
           963 => x"0a",
           964 => x"08",
           965 => x"3a",
           966 => x"28",
           967 => x"88",
           968 => x"c0",
           969 => x"02",
           970 => x"c0",
           971 => x"0a",
           972 => x"c0",
           973 => x"07",
           974 => x"a0",
           975 => x"07",
           976 => x"60",
           977 => x"60",
           978 => x"06",
           979 => x"06",
           980 => x"01",
           981 => x"2a",
           982 => x"8f",
           983 => x"a9",
           984 => x"f7",
           985 => x"02",
           986 => x"9f",
           987 => x"81",
           988 => x"02",
           989 => x"41",
           990 => x"01",
           991 => x"04",
           992 => x"30",
           993 => x"79",
           994 => x"0c",
           995 => x"9e",
           996 => x"30",
           997 => x"f9",
           998 => x"0c",
           999 => x"9f",
          1000 => x"28",
          1001 => x"78",
          1002 => x"ee",
          1003 => x"ba",
          1004 => x"fe",
          1005 => x"aa",
          1006 => x"e7",
          1007 => x"ff",
          1008 => x"e7",
          1009 => x"ff",
          1010 => x"00",
          1011 => x"63",
          1012 => x"00",
          1013 => x"c6",
          1014 => x"81",
          1015 => x"a5",
          1016 => x"81",
          1017 => x"81",
          1018 => x"04",
          1019 => x"fe",
          1020 => x"24",
          1021 => x"10",
          1022 => x"08",
          1023 => x"24",
        others => X"00"
    );

    shared variable RAM2     : ramArray :=
    (
             0 => x"00",
             1 => x"00",
             2 => x"42",
             3 => x"42",
             4 => x"22",
             5 => x"7c",
             6 => x"40",
             7 => x"1c",
             8 => x"22",
             9 => x"78",
            10 => x"40",
            11 => x"7e",
            12 => x"40",
            13 => x"40",
            14 => x"40",
            15 => x"1c",
            16 => x"42",
            17 => x"42",
            18 => x"08",
            19 => x"1c",
            20 => x"04",
            21 => x"38",
            22 => x"48",
            23 => x"42",
            24 => x"40",
            25 => x"7e",
            26 => x"5a",
            27 => x"42",
            28 => x"52",
            29 => x"42",
            30 => x"42",
            31 => x"18",
            32 => x"42",
            33 => x"40",
            34 => x"42",
            35 => x"1a",
            36 => x"42",
            37 => x"42",
            38 => x"40",
            39 => x"3c",
            40 => x"08",
            41 => x"08",
            42 => x"42",
            43 => x"3c",
            44 => x"42",
            45 => x"18",
            46 => x"42",
            47 => x"42",
            48 => x"24",
            49 => x"42",
            50 => x"22",
            51 => x"08",
            52 => x"04",
            53 => x"7e",
            54 => x"10",
            55 => x"3e",
            56 => x"08",
            57 => x"00",
            58 => x"08",
            59 => x"00",
            60 => x"08",
            61 => x"08",
            62 => x"08",
            63 => x"00",
            64 => x"46",
            65 => x"3c",
            66 => x"28",
            67 => x"3e",
            68 => x"02",
            69 => x"7e",
            70 => x"02",
            71 => x"3c",
            72 => x"14",
            73 => x"04",
            74 => x"78",
            75 => x"38",
            76 => x"40",
            77 => x"3c",
            78 => x"04",
            79 => x"10",
            80 => x"42",
            81 => x"3c",
            82 => x"42",
            83 => x"38",
            84 => x"00",
            85 => x"00",
            86 => x"7e",
            87 => x"00",
            88 => x"08",
            89 => x"08",
            90 => x"04",
            91 => x"40",
            92 => x"00",
            93 => x"18",
            94 => x"00",
            95 => x"08",
            96 => x"00",
            97 => x"00",
            98 => x"40",
            99 => x"40",
           100 => x"80",
           101 => x"80",
           102 => x"01",
           103 => x"01",
           104 => x"00",
           105 => x"00",
           106 => x"10",
           107 => x"10",
           108 => x"00",
           109 => x"00",
           110 => x"c0",
           111 => x"c0",
           112 => x"00",
           113 => x"00",
           114 => x"04",
           115 => x"04",
           116 => x"00",
           117 => x"ff",
           118 => x"0f",
           119 => x"0f",
           120 => x"00",
           121 => x"00",
           122 => x"01",
           123 => x"01",
           124 => x"00",
           125 => x"ff",
           126 => x"03",
           127 => x"03",
           128 => x"08",
           129 => x"10",
           130 => x"3e",
           131 => x"3e",
           132 => x"3f",
           133 => x"03",
           134 => x"ff",
           135 => x"ff",
           136 => x"3e",
           137 => x"08",
           138 => x"10",
           139 => x"10",
           140 => x"6b",
           141 => x"1c",
           142 => x"7e",
           143 => x"3c",
           144 => x"42",
           145 => x"3c",
           146 => x"02",
           147 => x"10",
           148 => x"81",
           149 => x"c3",
           150 => x"00",
           151 => x"08",
           152 => x"00",
           153 => x"10",
           154 => x"e0",
           155 => x"fe",
           156 => x"07",
           157 => x"7f",
           158 => x"08",
           159 => x"00",
           160 => x"1c",
           161 => x"08",
           162 => x"30",
           163 => x"0e",
           164 => x"20",
           165 => x"3c",
           166 => x"7f",
           167 => x"08",
           168 => x"04",
           169 => x"3c",
           170 => x"4a",
           171 => x"1e",
           172 => x"fc",
           173 => x"c0",
           174 => x"0c",
           175 => x"70",
           176 => x"08",
           177 => x"08",
           178 => x"20",
           179 => x"02",
           180 => x"04",
           181 => x"04",
           182 => x"f0",
           183 => x"0f",
           184 => x"00",
           185 => x"08",
           186 => x"00",
           187 => x"08",
           188 => x"08",
           189 => x"08",
           190 => x"00",
           191 => x"08",
           192 => x"01",
           193 => x"14",
           194 => x"08",
           195 => x"08",
           196 => x"24",
           197 => x"00",
           198 => x"7e",
           199 => x"24",
           200 => x"28",
           201 => x"08",
           202 => x"64",
           203 => x"46",
           204 => x"48",
           205 => x"3a",
           206 => x"10",
           207 => x"00",
           208 => x"10",
           209 => x"04",
           210 => x"08",
           211 => x"20",
           212 => x"08",
           213 => x"00",
           214 => x"1c",
           215 => x"08",
           216 => x"0f",
           217 => x"f0",
           218 => x"24",
           219 => x"42",
           220 => x"20",
           221 => x"00",
           222 => x"04",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"80",
           227 => x"80",
           228 => x"80",
           229 => x"80",
           230 => x"01",
           231 => x"01",
           232 => x"ff",
           233 => x"00",
           234 => x"20",
           235 => x"20",
           236 => x"04",
           237 => x"40",
           238 => x"20",
           239 => x"02",
           240 => x"00",
           241 => x"00",
           242 => x"08",
           243 => x"08",
           244 => x"ff",
           245 => x"00",
           246 => x"f0",
           247 => x"f0",
           248 => x"00",
           249 => x"ff",
           250 => x"02",
           251 => x"02",
           252 => x"00",
           253 => x"ff",
           254 => x"07",
           255 => x"07",
           256 => x"18",
           257 => x"18",
           258 => x"38",
           259 => x"3a",
           260 => x"5c",
           261 => x"5c",
           262 => x"3c",
           263 => x"3c",
           264 => x"3a",
           265 => x"3a",
           266 => x"3c",
           267 => x"3c",
           268 => x"10",
           269 => x"10",
           270 => x"3a",
           271 => x"02",
           272 => x"5c",
           273 => x"42",
           274 => x"18",
           275 => x"1c",
           276 => x"0c",
           277 => x"44",
           278 => x"44",
           279 => x"44",
           280 => x"08",
           281 => x"1c",
           282 => x"76",
           283 => x"49",
           284 => x"5c",
           285 => x"42",
           286 => x"3c",
           287 => x"3c",
           288 => x"5c",
           289 => x"40",
           290 => x"3a",
           291 => x"02",
           292 => x"5c",
           293 => x"40",
           294 => x"3e",
           295 => x"7c",
           296 => x"7c",
           297 => x"0c",
           298 => x"42",
           299 => x"3a",
           300 => x"42",
           301 => x"18",
           302 => x"41",
           303 => x"36",
           304 => x"44",
           305 => x"44",
           306 => x"42",
           307 => x"02",
           308 => x"7e",
           309 => x"7e",
           310 => x"38",
           311 => x"3a",
           312 => x"00",
           313 => x"08",
           314 => x"60",
           315 => x"00",
           316 => x"06",
           317 => x"00",
           318 => x"00",
           319 => x"10",
           320 => x"00",
           321 => x"0c",
           322 => x"00",
           323 => x"00",
           324 => x"44",
           325 => x"44",
           326 => x"44",
           327 => x"44",
           328 => x"08",
           329 => x"00",
           330 => x"00",
           331 => x"00",
           332 => x"aa",
           333 => x"aa",
           334 => x"00",
           335 => x"30",
           336 => x"30",
           337 => x"00",
           338 => x"0c",
           339 => x"00",
           340 => x"44",
           341 => x"4c",
           342 => x"00",
           343 => x"1a",
           344 => x"00",
           345 => x"1c",
           346 => x"42",
           347 => x"3c",
           348 => x"24",
           349 => x"42",
           350 => x"24",
           351 => x"18",
           352 => x"20",
           353 => x"80",
           354 => x"18",
           355 => x"40",
           356 => x"18",
           357 => x"02",
           358 => x"04",
           359 => x"01",
           360 => x"40",
           361 => x"20",
           362 => x"40",
           363 => x"06",
           364 => x"02",
           365 => x"60",
           366 => x"02",
           367 => x"04",
           368 => x"04",
           369 => x"00",
           370 => x"00",
           371 => x"1c",
           372 => x"00",
           373 => x"38",
           374 => x"20",
           375 => x"00",
           376 => x"10",
           377 => x"08",
           378 => x"08",
           379 => x"08",
           380 => x"22",
           381 => x"00",
           382 => x"00",
           383 => x"7e",
           384 => x"3e",
           385 => x"3e",
           386 => x"f7",
           387 => x"f7",
           388 => x"e3",
           389 => x"f7",
           390 => x"f7",
           391 => x"f7",
           392 => x"ef",
           393 => x"ef",
           394 => x"bd",
           395 => x"bd",
           396 => x"bf",
           397 => x"e3",
           398 => x"7e",
           399 => x"00",
           400 => x"42",
           401 => x"e0",
           402 => x"2a",
           403 => x"7f",
           404 => x"08",
           405 => x"14",
           406 => x"d2",
           407 => x"00",
           408 => x"4b",
           409 => x"00",
           410 => x"08",
           411 => x"1c",
           412 => x"ff",
           413 => x"7e",
           414 => x"81",
           415 => x"42",
           416 => x"aa",
           417 => x"aa",
           418 => x"0a",
           419 => x"0a",
           420 => x"a0",
           421 => x"a0",
           422 => x"aa",
           423 => x"00",
           424 => x"00",
           425 => x"aa",
           426 => x"a8",
           427 => x"80",
           428 => x"2a",
           429 => x"02",
           430 => x"a0",
           431 => x"aa",
           432 => x"02",
           433 => x"2a",
           434 => x"40",
           435 => x"10",
           436 => x"04",
           437 => x"01",
           438 => x"38",
           439 => x"00",
           440 => x"2a",
           441 => x"2a",
           442 => x"02",
           443 => x"08",
           444 => x"20",
           445 => x"80",
           446 => x"c8",
           447 => x"22",
           448 => x"00",
           449 => x"ff",
           450 => x"02",
           451 => x"07",
           452 => x"02",
           453 => x"ff",
           454 => x"20",
           455 => x"02",
           456 => x"11",
           457 => x"02",
           458 => x"44",
           459 => x"44",
           460 => x"88",
           461 => x"40",
           462 => x"a4",
           463 => x"a4",
           464 => x"25",
           465 => x"25",
           466 => x"a0",
           467 => x"98",
           468 => x"b8",
           469 => x"90",
           470 => x"20",
           471 => x"40",
           472 => x"24",
           473 => x"24",
           474 => x"3e",
           475 => x"08",
           476 => x"20",
           477 => x"02",
           478 => x"55",
           479 => x"55",
           480 => x"00",
           481 => x"00",
           482 => x"70",
           483 => x"00",
           484 => x"07",
           485 => x"00",
           486 => x"77",
           487 => x"00",
           488 => x"00",
           489 => x"70",
           490 => x"70",
           491 => x"70",
           492 => x"07",
           493 => x"70",
           494 => x"77",
           495 => x"70",
           496 => x"00",
           497 => x"07",
           498 => x"70",
           499 => x"07",
           500 => x"07",
           501 => x"07",
           502 => x"77",
           503 => x"07",
           504 => x"00",
           505 => x"77",
           506 => x"70",
           507 => x"77",
           508 => x"07",
           509 => x"77",
           510 => x"77",
           511 => x"77",
           512 => x"00",
           513 => x"00",
           514 => x"ba",
           515 => x"aa",
           516 => x"ba",
           517 => x"86",
           518 => x"be",
           519 => x"c2",
           520 => x"b6",
           521 => x"8c",
           522 => x"be",
           523 => x"82",
           524 => x"be",
           525 => x"a0",
           526 => x"be",
           527 => x"82",
           528 => x"ba",
           529 => x"aa",
           530 => x"ee",
           531 => x"82",
           532 => x"1b",
           533 => x"c6",
           534 => x"b4",
           535 => x"aa",
           536 => x"a0",
           537 => x"82",
           538 => x"aa",
           539 => x"aa",
           540 => x"8a",
           541 => x"aa",
           542 => x"ba",
           543 => x"c6",
           544 => x"ba",
           545 => x"a0",
           546 => x"ba",
           547 => x"c2",
           548 => x"ba",
           549 => x"aa",
           550 => x"be",
           551 => x"86",
           552 => x"ee",
           553 => x"28",
           554 => x"aa",
           555 => x"c6",
           556 => x"aa",
           557 => x"28",
           558 => x"aa",
           559 => x"82",
           560 => x"54",
           561 => x"aa",
           562 => x"92",
           563 => x"28",
           564 => x"fa",
           565 => x"82",
           566 => x"a0",
           567 => x"00",
           568 => x"05",
           569 => x"00",
           570 => x"d6",
           571 => x"92",
           572 => x"38",
           573 => x"92",
           574 => x"38",
           575 => x"00",
           576 => x"b2",
           577 => x"82",
           578 => x"68",
           579 => x"44",
           580 => x"ba",
           581 => x"42",
           582 => x"fa",
           583 => x"82",
           584 => x"24",
           585 => x"f6",
           586 => x"be",
           587 => x"86",
           588 => x"be",
           589 => x"82",
           590 => x"fa",
           591 => x"50",
           592 => x"ba",
           593 => x"82",
           594 => x"ba",
           595 => x"82",
           596 => x"be",
           597 => x"3e",
           598 => x"7d",
           599 => x"7c",
           600 => x"ff",
           601 => x"42",
           602 => x"ff",
           603 => x"24",
           604 => x"2a",
           605 => x"36",
           606 => x"2a",
           607 => x"36",
           608 => x"3c",
           609 => x"42",
           610 => x"3c",
           611 => x"42",
           612 => x"bd",
           613 => x"24",
           614 => x"5a",
           615 => x"c3",
           616 => x"7e",
           617 => x"24",
           618 => x"bd",
           619 => x"42",
           620 => x"ff",
           621 => x"dd",
           622 => x"ff",
           623 => x"77",
           624 => x"a5",
           625 => x"d5",
           626 => x"a5",
           627 => x"ab",
           628 => x"66",
           629 => x"7e",
           630 => x"3f",
           631 => x"fe",
           632 => x"ff",
           633 => x"42",
           634 => x"fc",
           635 => x"7f",
           636 => x"ff",
           637 => x"7e",
           638 => x"28",
           639 => x"fe",
           640 => x"07",
           641 => x"07",
           642 => x"3e",
           643 => x"1c",
           644 => x"e0",
           645 => x"e0",
           646 => x"3c",
           647 => x"76",
           648 => x"3c",
           649 => x"5a",
           650 => x"3c",
           651 => x"6e",
           652 => x"24",
           653 => x"24",
           654 => x"24",
           655 => x"24",
           656 => x"24",
           657 => x"24",
           658 => x"f7",
           659 => x"3c",
           660 => x"ff",
           661 => x"fc",
           662 => x"7e",
           663 => x"c6",
           664 => x"ff",
           665 => x"3f",
           666 => x"ff",
           667 => x"3c",
           668 => x"7e",
           669 => x"7e",
           670 => x"ff",
           671 => x"3e",
           672 => x"ff",
           673 => x"7c",
           674 => x"3c",
           675 => x"3c",
           676 => x"7b",
           677 => x"00",
           678 => x"18",
           679 => x"3c",
           680 => x"de",
           681 => x"00",
           682 => x"20",
           683 => x"3c",
           684 => x"ff",
           685 => x"00",
           686 => x"14",
           687 => x"06",
           688 => x"ff",
           689 => x"00",
           690 => x"38",
           691 => x"10",
           692 => x"10",
           693 => x"10",
           694 => x"10",
           695 => x"10",
           696 => x"08",
           697 => x"08",
           698 => x"60",
           699 => x"02",
           700 => x"04",
           701 => x"78",
           702 => x"20",
           703 => x"1e",
           704 => x"06",
           705 => x"40",
           706 => x"7e",
           707 => x"81",
           708 => x"70",
           709 => x"78",
           710 => x"81",
           711 => x"7e",
           712 => x"0e",
           713 => x"1e",
           714 => x"ad",
           715 => x"81",
           716 => x"bd",
           717 => x"01",
           718 => x"bd",
           719 => x"85",
           720 => x"bf",
           721 => x"81",
           722 => x"00",
           723 => x"00",
           724 => x"15",
           725 => x"05",
           726 => x"7e",
           727 => x"18",
           728 => x"a8",
           729 => x"a0",
           730 => x"1c",
           731 => x"1c",
           732 => x"11",
           733 => x"11",
           734 => x"1c",
           735 => x"1c",
           736 => x"44",
           737 => x"44",
           738 => x"e7",
           739 => x"00",
           740 => x"54",
           741 => x"38",
           742 => x"24",
           743 => x"24",
           744 => x"22",
           745 => x"08",
           746 => x"55",
           747 => x"55",
           748 => x"ff",
           749 => x"ff",
           750 => x"a5",
           751 => x"42",
           752 => x"81",
           753 => x"42",
           754 => x"9f",
           755 => x"a0",
           756 => x"e5",
           757 => x"15",
           758 => x"00",
           759 => x"a0",
           760 => x"00",
           761 => x"55",
           762 => x"80",
           763 => x"30",
           764 => x"01",
           765 => x"0c",
           766 => x"80",
           767 => x"80",
           768 => x"01",
           769 => x"01",
           770 => x"ab",
           771 => x"14",
           772 => x"18",
           773 => x"00",
           774 => x"24",
           775 => x"18",
           776 => x"81",
           777 => x"42",
           778 => x"00",
           779 => x"00",
           780 => x"3c",
           781 => x"00",
           782 => x"7e",
           783 => x"7e",
           784 => x"9d",
           785 => x"42",
           786 => x"ff",
           787 => x"ff",
           788 => x"c3",
           789 => x"ff",
           790 => x"81",
           791 => x"81",
           792 => x"20",
           793 => x"3c",
           794 => x"81",
           795 => x"42",
           796 => x"99",
           797 => x"5a",
           798 => x"99",
           799 => x"5a",
           800 => x"fe",
           801 => x"38",
           802 => x"40",
           803 => x"80",
           804 => x"02",
           805 => x"01",
           806 => x"40",
           807 => x"80",
           808 => x"02",
           809 => x"01",
           810 => x"88",
           811 => x"30",
           812 => x"11",
           813 => x"0c",
           814 => x"80",
           815 => x"30",
           816 => x"01",
           817 => x"0c",
           818 => x"83",
           819 => x"30",
           820 => x"c1",
           821 => x"0c",
           822 => x"87",
           823 => x"30",
           824 => x"e1",
           825 => x"0c",
           826 => x"54",
           827 => x"fe",
           828 => x"08",
           829 => x"78",
           830 => x"34",
           831 => x"4a",
           832 => x"00",
           833 => x"4a",
           834 => x"e0",
           835 => x"ff",
           836 => x"01",
           837 => x"c3",
           838 => x"80",
           839 => x"c3",
           840 => x"20",
           841 => x"ff",
           842 => x"07",
           843 => x"ff",
           844 => x"28",
           845 => x"08",
           846 => x"42",
           847 => x"42",
           848 => x"04",
           849 => x"ff",
           850 => x"10",
           851 => x"48",
           852 => x"42",
           853 => x"a5",
           854 => x"82",
           855 => x"00",
           856 => x"6c",
           857 => x"00",
           858 => x"6c",
           859 => x"00",
           860 => x"10",
           861 => x"10",
           862 => x"10",
           863 => x"10",
           864 => x"5b",
           865 => x"51",
           866 => x"91",
           867 => x"91",
           868 => x"a5",
           869 => x"c3",
           870 => x"54",
           871 => x"54",
           872 => x"99",
           873 => x"99",
           874 => x"38",
           875 => x"10",
           876 => x"38",
           877 => x"38",
           878 => x"00",
           879 => x"00",
           880 => x"10",
           881 => x"00",
           882 => x"7e",
           883 => x"7e",
           884 => x"55",
           885 => x"ff",
           886 => x"00",
           887 => x"83",
           888 => x"00",
           889 => x"c1",
           890 => x"00",
           891 => x"ff",
           892 => x"7e",
           893 => x"00",
           894 => x"f0",
           895 => x"e0",
           896 => x"0f",
           897 => x"07",
           898 => x"3f",
           899 => x"37",
           900 => x"b8",
           901 => x"fb",
           902 => x"0a",
           903 => x"03",
           904 => x"f4",
           905 => x"fd",
           906 => x"e4",
           907 => x"60",
           908 => x"27",
           909 => x"06",
           910 => x"1b",
           911 => x"0f",
           912 => x"d8",
           913 => x"f0",
           914 => x"07",
           915 => x"70",
           916 => x"e0",
           917 => x"0e",
           918 => x"06",
           919 => x"7f",
           920 => x"60",
           921 => x"fe",
           922 => x"7b",
           923 => x"7f",
           924 => x"de",
           925 => x"fe",
           926 => x"1f",
           927 => x"00",
           928 => x"f8",
           929 => x"00",
           930 => x"02",
           931 => x"1f",
           932 => x"40",
           933 => x"f8",
           934 => x"02",
           935 => x"7f",
           936 => x"40",
           937 => x"fe",
           938 => x"73",
           939 => x"0f",
           940 => x"ce",
           941 => x"f0",
           942 => x"0f",
           943 => x"7f",
           944 => x"f0",
           945 => x"fe",
           946 => x"42",
           947 => x"44",
           948 => x"07",
           949 => x"05",
           950 => x"82",
           951 => x"86",
           952 => x"80",
           953 => x"00",
           954 => x"00",
           955 => x"01",
           956 => x"01",
           957 => x"00",
           958 => x"80",
           959 => x"00",
           960 => x"00",
           961 => x"80",
           962 => x"0c",
           963 => x"0c",
           964 => x"0c",
           965 => x"0c",
           966 => x"48",
           967 => x"8f",
           968 => x"40",
           969 => x"04",
           970 => x"40",
           971 => x"1f",
           972 => x"40",
           973 => x"01",
           974 => x"20",
           975 => x"01",
           976 => x"18",
           977 => x"80",
           978 => x"18",
           979 => x"01",
           980 => x"06",
           981 => x"2a",
           982 => x"65",
           983 => x"b1",
           984 => x"f0",
           985 => x"3e",
           986 => x"31",
           987 => x"f9",
           988 => x"40",
           989 => x"00",
           990 => x"88",
           991 => x"80",
           992 => x"58",
           993 => x"30",
           994 => x"1a",
           995 => x"0c",
           996 => x"58",
           997 => x"30",
           998 => x"1a",
           999 => x"0c",
          1000 => x"68",
          1001 => x"10",
          1002 => x"aa",
          1003 => x"fe",
          1004 => x"ba",
          1005 => x"ee",
          1006 => x"42",
          1007 => x"42",
          1008 => x"42",
          1009 => x"42",
          1010 => x"fc",
          1011 => x"3e",
          1012 => x"3f",
          1013 => x"7c",
          1014 => x"a5",
          1015 => x"81",
          1016 => x"81",
          1017 => x"81",
          1018 => x"08",
          1019 => x"20",
          1020 => x"24",
          1021 => x"10",
          1022 => x"08",
          1023 => x"24",
        others => X"00"
    );

    shared variable RAM3     : ramArray :=
    (
             0 => x"00",
             1 => x"00",
             2 => x"7e",
             3 => x"00",
             4 => x"3c",
             5 => x"00",
             6 => x"40",
             7 => x"00",
             8 => x"22",
             9 => x"00",
            10 => x"78",
            11 => x"00",
            12 => x"78",
            13 => x"00",
            14 => x"4e",
            15 => x"00",
            16 => x"7e",
            17 => x"00",
            18 => x"08",
            19 => x"00",
            20 => x"04",
            21 => x"00",
            22 => x"70",
            23 => x"00",
            24 => x"40",
            25 => x"00",
            26 => x"5a",
            27 => x"00",
            28 => x"4a",
            29 => x"00",
            30 => x"42",
            31 => x"00",
            32 => x"7c",
            33 => x"00",
            34 => x"42",
            35 => x"00",
            36 => x"7c",
            37 => x"00",
            38 => x"3c",
            39 => x"00",
            40 => x"08",
            41 => x"00",
            42 => x"42",
            43 => x"00",
            44 => x"24",
            45 => x"00",
            46 => x"5a",
            47 => x"00",
            48 => x"18",
            49 => x"00",
            50 => x"1c",
            51 => x"00",
            52 => x"18",
            53 => x"00",
            54 => x"38",
            55 => x"00",
            56 => x"08",
            57 => x"00",
            58 => x"08",
            59 => x"00",
            60 => x"08",
            61 => x"08",
            62 => x"08",
            63 => x"00",
            64 => x"5a",
            65 => x"00",
            66 => x"08",
            67 => x"00",
            68 => x"0c",
            69 => x"00",
            70 => x"3c",
            71 => x"00",
            72 => x"24",
            73 => x"00",
            74 => x"04",
            75 => x"00",
            76 => x"7c",
            77 => x"00",
            78 => x"08",
            79 => x"00",
            80 => x"3c",
            81 => x"00",
            82 => x"3e",
            83 => x"00",
            84 => x"7e",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"10",
            90 => x"08",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"10",
            96 => x"00",
            97 => x"00",
            98 => x"40",
            99 => x"40",
           100 => x"80",
           101 => x"ff",
           102 => x"01",
           103 => x"ff",
           104 => x"ff",
           105 => x"00",
           106 => x"10",
           107 => x"10",
           108 => x"00",
           109 => x"00",
           110 => x"c0",
           111 => x"c0",
           112 => x"00",
           113 => x"00",
           114 => x"04",
           115 => x"04",
           116 => x"00",
           117 => x"ff",
           118 => x"0f",
           119 => x"0f",
           120 => x"00",
           121 => x"ff",
           122 => x"01",
           123 => x"01",
           124 => x"00",
           125 => x"ff",
           126 => x"03",
           127 => x"03",
           128 => x"04",
           129 => x"00",
           130 => x"7f",
           131 => x"00",
           132 => x"1f",
           133 => x"01",
           134 => x"ff",
           135 => x"ff",
           136 => x"7f",
           137 => x"00",
           138 => x"20",
           139 => x"00",
           140 => x"7f",
           141 => x"00",
           142 => x"7e",
           143 => x"00",
           144 => x"42",
           145 => x"00",
           146 => x"0c",
           147 => x"00",
           148 => x"81",
           149 => x"ff",
           150 => x"00",
           151 => x"08",
           152 => x"00",
           153 => x"10",
           154 => x"f0",
           155 => x"ff",
           156 => x"0f",
           157 => x"ff",
           158 => x"00",
           159 => x"00",
           160 => x"2a",
           161 => x"00",
           162 => x"60",
           163 => x"00",
           164 => x"20",
           165 => x"00",
           166 => x"7f",
           167 => x"00",
           168 => x"04",
           169 => x"00",
           170 => x"56",
           171 => x"00",
           172 => x"f8",
           173 => x"80",
           174 => x"06",
           175 => x"00",
           176 => x"08",
           177 => x"00",
           178 => x"10",
           179 => x"00",
           180 => x"02",
           181 => x"00",
           182 => x"f0",
           183 => x"0f",
           184 => x"00",
           185 => x"08",
           186 => x"00",
           187 => x"08",
           188 => x"08",
           189 => x"08",
           190 => x"00",
           191 => x"08",
           192 => x"3e",
           193 => x"00",
           194 => x"08",
           195 => x"00",
           196 => x"00",
           197 => x"00",
           198 => x"24",
           199 => x"00",
           200 => x"1c",
           201 => x"00",
           202 => x"08",
           203 => x"00",
           204 => x"30",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"10",
           209 => x"00",
           210 => x"08",
           211 => x"00",
           212 => x"3e",
           213 => x"00",
           214 => x"3e",
           215 => x"00",
           216 => x"0f",
           217 => x"f0",
           218 => x"18",
           219 => x"81",
           220 => x"c0",
           221 => x"00",
           222 => x"03",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"80",
           227 => x"80",
           228 => x"80",
           229 => x"80",
           230 => x"01",
           231 => x"01",
           232 => x"00",
           233 => x"00",
           234 => x"20",
           235 => x"20",
           236 => x"08",
           237 => x"80",
           238 => x"10",
           239 => x"01",
           240 => x"00",
           241 => x"00",
           242 => x"08",
           243 => x"08",
           244 => x"ff",
           245 => x"00",
           246 => x"f0",
           247 => x"f0",
           248 => x"00",
           249 => x"00",
           250 => x"02",
           251 => x"02",
           252 => x"00",
           253 => x"ff",
           254 => x"07",
           255 => x"07",
           256 => x"18",
           257 => x"00",
           258 => x"04",
           259 => x"00",
           260 => x"62",
           261 => x"00",
           262 => x"42",
           263 => x"00",
           264 => x"46",
           265 => x"00",
           266 => x"42",
           267 => x"00",
           268 => x"7c",
           269 => x"00",
           270 => x"46",
           271 => x"3c",
           272 => x"62",
           273 => x"00",
           274 => x"08",
           275 => x"00",
           276 => x"04",
           277 => x"38",
           278 => x"48",
           279 => x"00",
           280 => x"08",
           281 => x"00",
           282 => x"49",
           283 => x"00",
           284 => x"62",
           285 => x"00",
           286 => x"42",
           287 => x"00",
           288 => x"62",
           289 => x"40",
           290 => x"46",
           291 => x"02",
           292 => x"62",
           293 => x"00",
           294 => x"40",
           295 => x"00",
           296 => x"10",
           297 => x"00",
           298 => x"42",
           299 => x"00",
           300 => x"42",
           301 => x"00",
           302 => x"49",
           303 => x"00",
           304 => x"28",
           305 => x"00",
           306 => x"42",
           307 => x"3c",
           308 => x"04",
           309 => x"00",
           310 => x"04",
           311 => x"00",
           312 => x"01",
           313 => x"10",
           314 => x"80",
           315 => x"00",
           316 => x"01",
           317 => x"00",
           318 => x"80",
           319 => x"08",
           320 => x"00",
           321 => x"03",
           322 => x"00",
           323 => x"00",
           324 => x"44",
           325 => x"44",
           326 => x"44",
           327 => x"44",
           328 => x"00",
           329 => x"00",
           330 => x"32",
           331 => x"00",
           332 => x"11",
           333 => x"11",
           334 => x"00",
           335 => x"c0",
           336 => x"c0",
           337 => x"00",
           338 => x"03",
           339 => x"00",
           340 => x"4a",
           341 => x"00",
           342 => x"22",
           343 => x"00",
           344 => x"1c",
           345 => x"00",
           346 => x"42",
           347 => x"00",
           348 => x"42",
           349 => x"00",
           350 => x"42",
           351 => x"00",
           352 => x"40",
           353 => x"80",
           354 => x"20",
           355 => x"80",
           356 => x"04",
           357 => x"01",
           358 => x"02",
           359 => x"01",
           360 => x"40",
           361 => x"10",
           362 => x"20",
           363 => x"01",
           364 => x"04",
           365 => x"80",
           366 => x"02",
           367 => x"08",
           368 => x"02",
           369 => x"00",
           370 => x"00",
           371 => x"03",
           372 => x"00",
           373 => x"c0",
           374 => x"40",
           375 => x"00",
           376 => x"20",
           377 => x"00",
           378 => x"08",
           379 => x"08",
           380 => x"00",
           381 => x"00",
           382 => x"00",
           383 => x"00",
           384 => x"1c",
           385 => x"00",
           386 => x"f7",
           387 => x"ff",
           388 => x"d5",
           389 => x"ff",
           390 => x"fb",
           391 => x"ff",
           392 => x"df",
           393 => x"ff",
           394 => x"81",
           395 => x"ff",
           396 => x"bf",
           397 => x"ff",
           398 => x"ff",
           399 => x"00",
           400 => x"7e",
           401 => x"00",
           402 => x"08",
           403 => x"41",
           404 => x"3e",
           405 => x"22",
           406 => x"fc",
           407 => x"00",
           408 => x"3f",
           409 => x"00",
           410 => x"08",
           411 => x"1c",
           412 => x"db",
           413 => x"3c",
           414 => x"a5",
           415 => x"3c",
           416 => x"55",
           417 => x"55",
           418 => x"05",
           419 => x"05",
           420 => x"50",
           421 => x"50",
           422 => x"55",
           423 => x"00",
           424 => x"00",
           425 => x"55",
           426 => x"50",
           427 => x"00",
           428 => x"15",
           429 => x"01",
           430 => x"50",
           431 => x"55",
           432 => x"05",
           433 => x"55",
           434 => x"40",
           435 => x"10",
           436 => x"04",
           437 => x"01",
           438 => x"00",
           439 => x"00",
           440 => x"54",
           441 => x"00",
           442 => x"02",
           443 => x"08",
           444 => x"20",
           445 => x"80",
           446 => x"54",
           447 => x"00",
           448 => x"00",
           449 => x"02",
           450 => x"02",
           451 => x"02",
           452 => x"02",
           453 => x"02",
           454 => x"50",
           455 => x"00",
           456 => x"22",
           457 => x"01",
           458 => x"88",
           459 => x"88",
           460 => x"44",
           461 => x"80",
           462 => x"94",
           463 => x"c4",
           464 => x"29",
           465 => x"23",
           466 => x"c0",
           467 => x"b8",
           468 => x"c0",
           469 => x"88",
           470 => x"10",
           471 => x"80",
           472 => x"24",
           473 => x"00",
           474 => x"00",
           475 => x"08",
           476 => x"10",
           477 => x"04",
           478 => x"aa",
           479 => x"aa",
           480 => x"00",
           481 => x"00",
           482 => x"70",
           483 => x"00",
           484 => x"07",
           485 => x"00",
           486 => x"77",
           487 => x"00",
           488 => x"00",
           489 => x"70",
           490 => x"70",
           491 => x"70",
           492 => x"07",
           493 => x"70",
           494 => x"77",
           495 => x"70",
           496 => x"00",
           497 => x"07",
           498 => x"70",
           499 => x"07",
           500 => x"07",
           501 => x"07",
           502 => x"77",
           503 => x"07",
           504 => x"00",
           505 => x"77",
           506 => x"70",
           507 => x"77",
           508 => x"07",
           509 => x"77",
           510 => x"77",
           511 => x"77",
           512 => x"00",
           513 => x"00",
           514 => x"ba",
           515 => x"ee",
           516 => x"84",
           517 => x"fc",
           518 => x"a0",
           519 => x"7e",
           520 => x"aa",
           521 => x"f8",
           522 => x"88",
           523 => x"fe",
           524 => x"88",
           525 => x"e0",
           526 => x"a0",
           527 => x"7e",
           528 => x"82",
           529 => x"ee",
           530 => x"28",
           531 => x"fe",
           532 => x"0a",
           533 => x"7c",
           534 => x"88",
           535 => x"e6",
           536 => x"a0",
           537 => x"fe",
           538 => x"aa",
           539 => x"ee",
           540 => x"a2",
           541 => x"ee",
           542 => x"aa",
           543 => x"7c",
           544 => x"ba",
           545 => x"e0",
           546 => x"ba",
           547 => x"7c",
           548 => x"ba",
           549 => x"e6",
           550 => x"c4",
           551 => x"fc",
           552 => x"28",
           553 => x"38",
           554 => x"aa",
           555 => x"7c",
           556 => x"aa",
           557 => x"10",
           558 => x"ba",
           559 => x"fe",
           560 => x"28",
           561 => x"c6",
           562 => x"44",
           563 => x"38",
           564 => x"14",
           565 => x"fe",
           566 => x"90",
           567 => x"00",
           568 => x"09",
           569 => x"00",
           570 => x"7c",
           571 => x"00",
           572 => x"fe",
           573 => x"00",
           574 => x"54",
           575 => x"00",
           576 => x"aa",
           577 => x"7c",
           578 => x"28",
           579 => x"7c",
           580 => x"ca",
           581 => x"fe",
           582 => x"22",
           583 => x"fc",
           584 => x"54",
           585 => x"1c",
           586 => x"84",
           587 => x"fc",
           588 => x"bc",
           589 => x"7c",
           590 => x"14",
           591 => x"70",
           592 => x"7c",
           593 => x"7c",
           594 => x"82",
           595 => x"fc",
           596 => x"aa",
           597 => x"00",
           598 => x"55",
           599 => x"00",
           600 => x"e7",
           601 => x"81",
           602 => x"e7",
           603 => x"66",
           604 => x"7f",
           605 => x"63",
           606 => x"7f",
           607 => x"14",
           608 => x"5a",
           609 => x"63",
           610 => x"5a",
           611 => x"c6",
           612 => x"99",
           613 => x"00",
           614 => x"18",
           615 => x"00",
           616 => x"bd",
           617 => x"e7",
           618 => x"7e",
           619 => x"c3",
           620 => x"ab",
           621 => x"89",
           622 => x"ab",
           623 => x"22",
           624 => x"81",
           625 => x"aa",
           626 => x"81",
           627 => x"55",
           628 => x"e7",
           629 => x"3c",
           630 => x"0f",
           631 => x"1c",
           632 => x"ff",
           633 => x"42",
           634 => x"f0",
           635 => x"38",
           636 => x"ff",
           637 => x"3c",
           638 => x"28",
           639 => x"d6",
           640 => x"7e",
           641 => x"03",
           642 => x"14",
           643 => x"08",
           644 => x"7e",
           645 => x"c0",
           646 => x"18",
           647 => x"46",
           648 => x"18",
           649 => x"7e",
           650 => x"18",
           651 => x"62",
           652 => x"24",
           653 => x"6c",
           654 => x"24",
           655 => x"66",
           656 => x"24",
           657 => x"36",
           658 => x"b7",
           659 => x"3c",
           660 => x"3f",
           661 => x"38",
           662 => x"ff",
           663 => x"44",
           664 => x"fc",
           665 => x"1e",
           666 => x"bf",
           667 => x"3c",
           668 => x"ff",
           669 => x"3c",
           670 => x"ff",
           671 => x"1c",
           672 => x"ff",
           673 => x"38",
           674 => x"3c",
           675 => x"3c",
           676 => x"ff",
           677 => x"00",
           678 => x"3c",
           679 => x"18",
           680 => x"ff",
           681 => x"00",
           682 => x"20",
           683 => x"3c",
           684 => x"0b",
           685 => x"00",
           686 => x"0c",
           687 => x"04",
           688 => x"d0",
           689 => x"00",
           690 => x"7c",
           691 => x"38",
           692 => x"31",
           693 => x"08",
           694 => x"92",
           695 => x"10",
           696 => x"8c",
           697 => x"10",
           698 => x"50",
           699 => x"00",
           700 => x"48",
           701 => x"00",
           702 => x"12",
           703 => x"00",
           704 => x"0a",
           705 => x"00",
           706 => x"ff",
           707 => x"81",
           708 => x"f0",
           709 => x"1f",
           710 => x"c3",
           711 => x"18",
           712 => x"0f",
           713 => x"f8",
           714 => x"a5",
           715 => x"ff",
           716 => x"a5",
           717 => x"ff",
           718 => x"a5",
           719 => x"fd",
           720 => x"a1",
           721 => x"ff",
           722 => x"3c",
           723 => x"ff",
           724 => x"55",
           725 => x"01",
           726 => x"00",
           727 => x"00",
           728 => x"aa",
           729 => x"80",
           730 => x"3e",
           731 => x"3e",
           732 => x"33",
           733 => x"00",
           734 => x"08",
           735 => x"08",
           736 => x"66",
           737 => x"00",
           738 => x"a5",
           739 => x"00",
           740 => x"10",
           741 => x"10",
           742 => x"42",
           743 => x"00",
           744 => x"1c",
           745 => x"7f",
           746 => x"55",
           747 => x"55",
           748 => x"00",
           749 => x"00",
           750 => x"00",
           751 => x"a5",
           752 => x"00",
           753 => x"24",
           754 => x"a0",
           755 => x"a0",
           756 => x"11",
           757 => x"11",
           758 => x"ff",
           759 => x"ff",
           760 => x"ff",
           761 => x"ff",
           762 => x"ff",
           763 => x"78",
           764 => x"ff",
           765 => x"1e",
           766 => x"95",
           767 => x"ff",
           768 => x"51",
           769 => x"ff",
           770 => x"d5",
           771 => x"08",
           772 => x"24",
           773 => x"00",
           774 => x"42",
           775 => x"00",
           776 => x"81",
           777 => x"3c",
           778 => x"18",
           779 => x"00",
           780 => x"3c",
           781 => x"00",
           782 => x"7e",
           783 => x"00",
           784 => x"a1",
           785 => x"3c",
           786 => x"e7",
           787 => x"ff",
           788 => x"c3",
           789 => x"ff",
           790 => x"81",
           791 => x"ff",
           792 => x"20",
           793 => x"00",
           794 => x"ff",
           795 => x"3c",
           796 => x"99",
           797 => x"3c",
           798 => x"ff",
           799 => x"3c",
           800 => x"aa",
           801 => x"10",
           802 => x"4e",
           803 => x"81",
           804 => x"72",
           805 => x"81",
           806 => x"40",
           807 => x"81",
           808 => x"02",
           809 => x"81",
           810 => x"84",
           811 => x"0f",
           812 => x"21",
           813 => x"f0",
           814 => x"87",
           815 => x"0f",
           816 => x"e1",
           817 => x"f0",
           818 => x"84",
           819 => x"0f",
           820 => x"21",
           821 => x"f0",
           822 => x"88",
           823 => x"0f",
           824 => x"11",
           825 => x"f0",
           826 => x"fe",
           827 => x"7c",
           828 => x"10",
           829 => x"30",
           830 => x"06",
           831 => x"00",
           832 => x"03",
           833 => x"89",
           834 => x"f0",
           835 => x"ff",
           836 => x"02",
           837 => x"ff",
           838 => x"40",
           839 => x"ff",
           840 => x"10",
           841 => x"fc",
           842 => x"0f",
           843 => x"ff",
           844 => x"08",
           845 => x"00",
           846 => x"20",
           847 => x"fe",
           848 => x"08",
           849 => x"3f",
           850 => x"10",
           851 => x"86",
           852 => x"42",
           853 => x"e7",
           854 => x"82",
           855 => x"00",
           856 => x"92",
           857 => x"00",
           858 => x"90",
           859 => x"00",
           860 => x"50",
           861 => x"00",
           862 => x"00",
           863 => x"00",
           864 => x"55",
           865 => x"00",
           866 => x"c5",
           867 => x"ff",
           868 => x"99",
           869 => x"ff",
           870 => x"38",
           871 => x"92",
           872 => x"ff",
           873 => x"ff",
           874 => x"10",
           875 => x"10",
           876 => x"10",
           877 => x"10",
           878 => x"aa",
           879 => x"00",
           880 => x"7c",
           881 => x"7c",
           882 => x"42",
           883 => x"42",
           884 => x"55",
           885 => x"00",
           886 => x"c0",
           887 => x"ff",
           888 => x"03",
           889 => x"ff",
           890 => x"00",
           891 => x"ff",
           892 => x"3c",
           893 => x"00",
           894 => x"f0",
           895 => x"c0",
           896 => x"0f",
           897 => x"03",
           898 => x"3f",
           899 => x"1f",
           900 => x"dc",
           901 => x"fb",
           902 => x"04",
           903 => x"0f",
           904 => x"f4",
           905 => x"fd",
           906 => x"46",
           907 => x"3f",
           908 => x"62",
           909 => x"fc",
           910 => x"1f",
           911 => x"07",
           912 => x"f8",
           913 => x"e0",
           914 => x"06",
           915 => x"30",
           916 => x"60",
           917 => x"0c",
           918 => x"07",
           919 => x"8b",
           920 => x"e0",
           921 => x"d1",
           922 => x"59",
           923 => x"3f",
           924 => x"9a",
           925 => x"fc",
           926 => x"0f",
           927 => x"ff",
           928 => x"f0",
           929 => x"ff",
           930 => x"04",
           931 => x"1f",
           932 => x"20",
           933 => x"f8",
           934 => x"02",
           935 => x"00",
           936 => x"40",
           937 => x"00",
           938 => x"7f",
           939 => x"0f",
           940 => x"fe",
           941 => x"f0",
           942 => x"18",
           943 => x"ff",
           944 => x"18",
           945 => x"ff",
           946 => x"21",
           947 => x"f8",
           948 => x"00",
           949 => x"ff",
           950 => x"81",
           951 => x"fc",
           952 => x"40",
           953 => x"00",
           954 => x"00",
           955 => x"01",
           956 => x"01",
           957 => x"00",
           958 => x"80",
           959 => x"00",
           960 => x"00",
           961 => x"ff",
           962 => x"0a",
           963 => x"08",
           964 => x"3a",
           965 => x"08",
           966 => x"fe",
           967 => x"00",
           968 => x"e6",
           969 => x"0f",
           970 => x"e2",
           971 => x"02",
           972 => x"ef",
           973 => x"0f",
           974 => x"4f",
           975 => x"0f",
           976 => x"06",
           977 => x"fe",
           978 => x"60",
           979 => x"7f",
           980 => x"1d",
           981 => x"1f",
           982 => x"11",
           983 => x"f3",
           984 => x"18",
           985 => x"fe",
           986 => x"41",
           987 => x"fd",
           988 => x"00",
           989 => x"91",
           990 => x"00",
           991 => x"11",
           992 => x"fd",
           993 => x"00",
           994 => x"bf",
           995 => x"00",
           996 => x"fd",
           997 => x"00",
           998 => x"bf",
           999 => x"00",
          1000 => x"bc",
          1001 => x"38",
          1002 => x"38",
          1003 => x"ba",
          1004 => x"38",
          1005 => x"ba",
          1006 => x"ff",
          1007 => x"e7",
          1008 => x"ff",
          1009 => x"e7",
          1010 => x"1c",
          1011 => x"00",
          1012 => x"38",
          1013 => x"00",
          1014 => x"81",
          1015 => x"ff",
          1016 => x"00",
          1017 => x"e7",
          1018 => x"fe",
          1019 => x"40",
          1020 => x"20",
          1021 => x"10",
          1022 => x"08",
          1023 => x"18",
        others => X"00"
    );

    signal RAM0_PORTA_DO     : std_logic_vector(7 downto 0);                  -- Buffer for byte in 32bit word to be written on Port A.
    signal RAM1_PORTA_DO     : std_logic_vector(7 downto 0);                  -- Buffer for byte in 32bit word to be written on Port A.
    signal RAM2_PORTA_DO     : std_logic_vector(7 downto 0);                  -- Buffer for byte in 32bit word to be written on Port A.
    signal RAM3_PORTA_DO     : std_logic_vector(7 downto 0);                  -- Buffer for byte in 32bit word to be written on Port A.
    signal RAM_PORTA_DI      : std_logic_vector(31 downto 0);                 -- Buffer for 32bit word being read prior to assignment to external port.
    signal RAM0_PORTB_DI     : std_logic_vector(7 downto 0);                  -- Buffer for 8bit byte being read prior to assignment to external port.
    signal RAM1_PORTB_DI     : std_logic_vector(7 downto 0);                  -- Buffer for 8bit byte being read prior to assignment to external port.
    signal RAM2_PORTB_DI     : std_logic_vector(7 downto 0);                  -- Buffer for 8bit byte being read prior to assignment to external port.
    signal RAM3_PORTB_DI     : std_logic_vector(7 downto 0);                  -- Buffer for 8bit byte being read prior to assignment to external port.
    signal RAM0_PORTA_WREN   : std_logic;                                     -- Write Enable for this particular byte in 32 bit word on Port A.
    signal RAM1_PORTA_WREN   : std_logic;                                     -- Write Enable for this particular byte in 32 bit word on Port A.
    signal RAM2_PORTA_WREN   : std_logic;                                     -- Write Enable for this particular byte in 32 bit word on Port A.
    signal RAM3_PORTA_WREN   : std_logic;                                     -- Write Enable for this particular byte in 32 bit word on Port A.
    signal RAM0_PORTB_WREN   : std_logic;                                     -- Write Enable for this particular byte in 16 bit word on Port B, lowest addr = '0'.
    signal RAM1_PORTB_WREN   : std_logic;                                     -- Write Enable for this particular byte in 16 bit word on Port B, lowest addr = '0'.
    signal RAM2_PORTB_WREN   : std_logic;                                     -- Write Enable for this particular byte in 16 bit word on Port B, lowest addr = '1'.
    signal RAM3_PORTB_WREN   : std_logic;                                     -- Write Enable for this particular byte in 16 bit word on Port B, lowest addr = '1'.

begin

    -- Choose data to be written according to Byte/HWord select signals.
    RAM0_PORTA_DO   <= memAWrite(7 downto 0);
    RAM1_PORTA_DO   <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                       else
                       memAWrite(7 downto 0);
    RAM2_PORTA_DO   <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                       else
                       memAWrite(7 downto 0);
    RAM3_PORTA_DO   <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                       else
                       memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                       else
                       memAWrite(7 downto 0);

    -- Data output is according to Least significant bits. Normally, a 32bit CPU would set them to 0 so output full word when 0, it there not zero, then 
    -- process as a byte read and copy selected byte to lower 8 bits.
    memARead        <= RAM_PORTA_DI                           when memAAddr(1 downto 0) = "00"
                       else
                       X"000000" & RAM_PORTA_DI(15 downto 8)  when memAAddr(1 downto 0) = "01"
                       else
                       X"000000" & RAM_PORTA_DI(23 downto 16) when memAAddr(1 downto 0) = "10"
                       else
                       X"000000" & RAM_PORTA_DI(31 downto 24);
    memBRead        <= RAM0_PORTB_DI                          when memBAddr(1 downto 0) = "00"
                       else
                       RAM1_PORTB_DI                          when memBAddr(1 downto 0) = "01"
                       else
                       RAM2_PORTB_DI                          when memBAddr(1 downto 0) = "10"
                       else
                       RAM3_PORTB_DI;

    -- Write enable based on byte select, either write a single byte or a complete word.
    RAM0_PORTA_WREN <= '1'                                    when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                       else '0';
    RAM1_PORTA_WREN <= '1'                                    when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                       else '0';
    RAM2_PORTA_WREN <= '1'                                    when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                       else '0';
    RAM3_PORTA_WREN <= '1'                                    when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                       else '0';

    -- Port B is 16bit read and write so use the lowest address line to toggle write to a particular RAM set array.
    RAM0_PORTB_WREN <= '1'                                    when memBWriteEnable = '1' and memBAddr(1 downto 0) = "00"
                       else '0';
    RAM1_PORTB_WREN <= '1'                                    when memBWriteEnable = '1' and memBAddr(1 downto 0) = "01"
                       else '0';
    RAM2_PORTB_WREN <= '1'                                    when memBWriteEnable = '1' and memBAddr(1 downto 0) = "10"
                       else '0';
    RAM3_PORTB_WREN <= '1'                                    when memBWriteEnable = '1' and memBAddr(1 downto 0) = "11"
                       else '0';

    ---------------- PORT A - 32 bit --------------------

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clkA)
    begin
        if rising_edge(clkA) then
            if RAM0_PORTA_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_PORTA_DO;
            end if;
            RAM_PORTA_DI(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clkA)
    begin
        if rising_edge(clkA) then
            if RAM1_PORTA_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_PORTA_DO;
            end if;
            RAM_PORTA_DI(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clkA)
    begin
        if rising_edge(clkA) then
            if RAM2_PORTA_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_PORTA_DO;
            end if;
            RAM_PORTA_DI(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clkA)
    begin
        if rising_edge(clkA) then
            if RAM3_PORTA_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_PORTA_DO;
            end if;
            RAM_PORTA_DI(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
        end if;
    end process;

    ---------------- PORT B - 8 bit --------------------

        -- BRAM Byte 0 - Port B - Byte 0 - bits 7 downto 0
    process(clkB)
    begin
        if rising_edge(clkB) then
            if RAM0_PORTB_WREN = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite;
            end if;
            RAM0_PORTB_DI  <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
        end if;
    end process;

    -- BRAM Byte 1 - Port B - Byte 1 - bits 15 downto 8
    process(clkB)
    begin
        if rising_edge(clkB) then
            if RAM1_PORTB_WREN = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite;
            end if;
            RAM1_PORTB_DI  <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
        end if;
    end process;

    -- BRAM Byte 2 - Port B - Byte 2 - bits 23 downto 16
    process(clkB)
    begin
        if rising_edge(clkB) then
            if RAM2_PORTB_WREN = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite;
            end if;
            RAM2_PORTB_DI  <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
        end if;
    end process;

    -- BRAM Byte 3 - Port B - Byte 3 - bits 31 downto 24
    process(clkB)
    begin
        if rising_edge(clkB) then
            if RAM3_PORTB_WREN = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite;
            end if;
            RAM3_PORTB_DI  <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
        end if;
    end process;

end arch;
