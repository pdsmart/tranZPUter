SFL_inst : SFL PORT MAP (
		noe_in	 => noe_in_sig
	);
