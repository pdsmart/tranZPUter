//----------------------------------------------------------------------------
//  A-Z80 CPU Copyright (C) 2014,2016  Goran Devic, www.baltazarstudios.com
//
//  This program is free software; you can redistribute it and/or modify it
//  under the terms of the GNU General Public License as published by the Free
//  Software Foundation; either version 2 of the License, or (at your option)
//  any later version.
//
//  This program is distributed in the hope that it will be useful, but WITHOUT
//  ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
//  FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License for
//  more details.
//----------------------------------------------------------------------------
// Automatically generated by gencompile.py

ctl_reg_gp_we = ctl_reg_gp_we | (pla[17]&~pla[50])&(M1&T1);
ctl_reg_gp_sel_pla17npla50M1T1_2 = (pla[17]&~pla[50])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla17npla50M1T1_2,ctl_reg_gp_sel_pla17npla50M1T1_2})&(op54);
ctl_reg_gp_hilo_pla17npla50M1T1_3 = (pla[17]&~pla[50])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla17npla50M1T1_3,ctl_reg_gp_hilo_pla17npla50M1T1_3})&({~rsel3,rsel3});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[17]&~pla[50])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[17]&~pla[50])&(M1&T1);
ctl_sw_2d = ctl_sw_2d | (pla[17]&~pla[50])&(M1&T1);
ctl_sw_1d = ctl_sw_1d | (pla[17]&~pla[50])&(M1&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[17]&~pla[50])&(M1&T1);
validPLA = validPLA | (pla[17]&~pla[50])&(M1&T4);
nextM = nextM | (pla[17]&~pla[50])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[17]&~pla[50])&(M1&T4);
fMRead = fMRead | (pla[17]&~pla[50])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[17]&~pla[50])&(M2&T1);
ctl_reg_sys_hilo_pla17npla50M2T1_3 = (pla[17]&~pla[50])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla17npla50M2T1_3,ctl_reg_sys_hilo_pla17npla50M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[17]&~pla[50])&(M2&T1);
fMRead = fMRead | (pla[17]&~pla[50])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[17]&~pla[50])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[17]&~pla[50])&(M2&T2);
ctl_reg_sys_hilo_pla17npla50M2T2_4 = (pla[17]&~pla[50])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla17npla50M2T2_4,ctl_reg_sys_hilo_pla17npla50M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[17]&~pla[50])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[17]&~pla[50])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[17]&~pla[50])&(M2&T2);
fMRead = fMRead | (pla[17]&~pla[50])&(M2&T3);
setM1 = setM1 | (pla[17]&~pla[50])&(M2&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[61]&~pla[58]&~pla[59])&(M1&T1);
ctl_reg_gp_sel_pla61npla58npla59M1T1_2 = (pla[61]&~pla[58]&~pla[59])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla61npla58npla59M1T1_2,ctl_reg_gp_sel_pla61npla58npla59M1T1_2})&(op54);
ctl_reg_gp_hilo_pla61npla58npla59M1T1_3 = (pla[61]&~pla[58]&~pla[59])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla61npla58npla59M1T1_3,ctl_reg_gp_hilo_pla61npla58npla59M1T1_3})&({~rsel3,rsel3});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[61]&~pla[58]&~pla[59])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[61]&~pla[58]&~pla[59])&(M1&T1);
ctl_sw_2u = ctl_sw_2u | (pla[61]&~pla[58]&~pla[59])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[61]&~pla[58]&~pla[59])&(M1&T1);
ctl_alu_op1_oe = ctl_alu_op1_oe | (pla[61]&~pla[58]&~pla[59])&(M1&T1);
validPLA = validPLA | (pla[61]&~pla[58]&~pla[59])&(M1&T4);
setM1 = setM1 | (pla[61]&~pla[58]&~pla[59])&(M1&T4);
ctl_reg_gp_sel_pla61npla58npla59M1T4_3 = (pla[61]&~pla[58]&~pla[59])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla61npla58npla59M1T4_3,ctl_reg_gp_sel_pla61npla58npla59M1T4_3})&(op21);
ctl_reg_gp_hilo_pla61npla58npla59M1T4_4 = (pla[61]&~pla[58]&~pla[59])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla61npla58npla59M1T4_4,ctl_reg_gp_hilo_pla61npla58npla59M1T4_4})&({~rsel0,rsel0});
ctl_reg_out_hi = ctl_reg_out_hi | (pla[61]&~pla[58]&~pla[59])&(M1&T4)&(~rsel0);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[61]&~pla[58]&~pla[59])&(M1&T4)&(rsel0);
ctl_sw_2u = ctl_sw_2u | (pla[61]&~pla[58]&~pla[59])&(M1&T4)&(~rsel0);
ctl_sw_2d = ctl_sw_2d | (pla[61]&~pla[58]&~pla[59])&(M1&T4)&(rsel0);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[61]&~pla[58]&~pla[59])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[61]&~pla[58]&~pla[59])&(M1&T4);
ctl_reg_gp_we = ctl_reg_gp_we | (use_ixiy&pla[58])&(M1&T1);
ctl_reg_gp_sel_use_ixiypla58M1T1_2 = (use_ixiy&pla[58])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_use_ixiypla58M1T1_2,ctl_reg_gp_sel_use_ixiypla58M1T1_2})&(op54);
ctl_reg_gp_hilo_use_ixiypla58M1T1_3 = (use_ixiy&pla[58])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_use_ixiypla58M1T1_3,ctl_reg_gp_hilo_use_ixiypla58M1T1_3})&({~rsel3,rsel3});
ctl_reg_in_hi = ctl_reg_in_hi | (use_ixiy&pla[58])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (use_ixiy&pla[58])&(M1&T1);
ctl_sw_2d = ctl_sw_2d | (use_ixiy&pla[58])&(M1&T1);
ctl_sw_1d = ctl_sw_1d | (use_ixiy&pla[58])&(M1&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (use_ixiy&pla[58])&(M1&T1);
validPLA = validPLA | (use_ixiy&pla[58])&(M1&T4);
nextM = nextM | (use_ixiy&pla[58])&(M1&T4);
ctl_mRead = ctl_mRead | (use_ixiy&pla[58])&(M1&T4);
fMRead = fMRead | (use_ixiy&pla[58])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (use_ixiy&pla[58])&(M2&T1);
ctl_reg_sys_hilo_use_ixiypla58M2T1_3 = (use_ixiy&pla[58])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_use_ixiypla58M2T1_3,ctl_reg_sys_hilo_use_ixiypla58M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (use_ixiy&pla[58])&(M2&T1);
fMRead = fMRead | (use_ixiy&pla[58])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (use_ixiy&pla[58])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (use_ixiy&pla[58])&(M2&T2);
ctl_reg_sys_hilo_use_ixiypla58M2T2_4 = (use_ixiy&pla[58])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_use_ixiypla58M2T2_4,ctl_reg_sys_hilo_use_ixiypla58M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (use_ixiy&pla[58])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (use_ixiy&pla[58])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (use_ixiy&pla[58])&(M2&T2);
fMRead = fMRead | (use_ixiy&pla[58])&(M2&T3);
nextM = nextM | (use_ixiy&pla[58])&(M2&T3);
ixy_d = ixy_d | (use_ixiy&pla[58])&(M3&T1);
ixy_d = ixy_d | (use_ixiy&pla[58])&(M3&T2);
ixy_d = ixy_d | (use_ixiy&pla[58])&(M3&T3);
ixy_d = ixy_d | (use_ixiy&pla[58])&(M3&T4);
nextM = nextM | (use_ixiy&pla[58])&(M3&T5);
ctl_mRead = ctl_mRead | (use_ixiy&pla[58])&(M3&T5);
ixy_d = ixy_d | (use_ixiy&pla[58])&(M3&T5);
ctl_reg_gp_we = ctl_reg_gp_we | (~use_ixiy&pla[58])&(M1&T1);
ctl_reg_gp_sel_nuse_ixiypla58M1T1_2 = (~use_ixiy&pla[58])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla58M1T1_2,ctl_reg_gp_sel_nuse_ixiypla58M1T1_2})&(op54);
ctl_reg_gp_hilo_nuse_ixiypla58M1T1_3 = (~use_ixiy&pla[58])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla58M1T1_3,ctl_reg_gp_hilo_nuse_ixiypla58M1T1_3})&({~rsel3,rsel3});
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[58])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[58])&(M1&T1);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[58])&(M1&T1);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[58])&(M1&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[58])&(M1&T1);
validPLA = validPLA | (~use_ixiy&pla[58])&(M1&T4);
nextM = nextM | (~use_ixiy&pla[58])&(M1&T4);
ctl_mRead = ctl_mRead | (~use_ixiy&pla[58])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[58])&(M2&T1);
ctl_reg_gp_sel_nuse_ixiypla58M2T1_2 = (~use_ixiy&pla[58])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla58M2T1_2,ctl_reg_gp_sel_nuse_ixiypla58M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_nuse_ixiypla58M2T1_3 = (~use_ixiy&pla[58])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla58M2T1_3,ctl_reg_gp_hilo_nuse_ixiypla58M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[58])&(M2&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[58])&(M2&T1);
fMRead = fMRead | (~use_ixiy&pla[58])&(M2&T2);
fMRead = fMRead | (~use_ixiy&pla[58])&(M2&T3);
setM1 = setM1 | (~use_ixiy&pla[58])&(M2&T3);
fMRead = fMRead | (~use_ixiy&pla[58])&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[58])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[58])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[58])&(M4&T3);
setM1 = setM1 | (~use_ixiy&pla[58])&(M4&T3);
validPLA = validPLA | (use_ixiy&pla[59])&(M1&T4);
nextM = nextM | (use_ixiy&pla[59])&(M1&T4);
ctl_mRead = ctl_mRead | (use_ixiy&pla[59])&(M1&T4);
fMRead = fMRead | (use_ixiy&pla[59])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (use_ixiy&pla[59])&(M2&T1);
ctl_reg_sys_hilo_use_ixiypla59M2T1_3 = (use_ixiy&pla[59])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_use_ixiypla59M2T1_3,ctl_reg_sys_hilo_use_ixiypla59M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (use_ixiy&pla[59])&(M2&T1);
fMRead = fMRead | (use_ixiy&pla[59])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (use_ixiy&pla[59])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (use_ixiy&pla[59])&(M2&T2);
ctl_reg_sys_hilo_use_ixiypla59M2T2_4 = (use_ixiy&pla[59])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_use_ixiypla59M2T2_4,ctl_reg_sys_hilo_use_ixiypla59M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (use_ixiy&pla[59])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (use_ixiy&pla[59])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (use_ixiy&pla[59])&(M2&T2);
fMRead = fMRead | (use_ixiy&pla[59])&(M2&T3);
nextM = nextM | (use_ixiy&pla[59])&(M2&T3);
ixy_d = ixy_d | (use_ixiy&pla[59])&(M3&T1);
ixy_d = ixy_d | (use_ixiy&pla[59])&(M3&T2);
ixy_d = ixy_d | (use_ixiy&pla[59])&(M3&T3);
ixy_d = ixy_d | (use_ixiy&pla[59])&(M3&T4);
nextM = nextM | (use_ixiy&pla[59])&(M3&T5);
ctl_mWrite = ctl_mWrite | (use_ixiy&pla[59])&(M3&T5);
ixy_d = ixy_d | (use_ixiy&pla[59])&(M3&T5);
validPLA = validPLA | (~use_ixiy&pla[59])&(M1&T4);
nextM = nextM | (~use_ixiy&pla[59])&(M1&T4);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[59])&(M1&T4);
ctl_reg_gp_sel_nuse_ixiypla59M1T4_4 = (~use_ixiy&pla[59])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla59M1T4_4,ctl_reg_gp_sel_nuse_ixiypla59M1T4_4})&(op21);
ctl_reg_gp_hilo_nuse_ixiypla59M1T4_5 = (~use_ixiy&pla[59])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla59M1T4_5,ctl_reg_gp_hilo_nuse_ixiypla59M1T4_5})&({~rsel0,rsel0});
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[59])&(M1&T4)&(~rsel0);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[59])&(M1&T4)&(rsel0);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[59])&(M1&T4)&(~rsel0);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[59])&(M1&T4)&(rsel0);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[59])&(M1&T4);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[59])&(M1&T4);
fMWrite = fMWrite | (~use_ixiy&pla[59])&(M2&T1);
ctl_reg_gp_sel_nuse_ixiypla59M2T1_2 = (~use_ixiy&pla[59])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla59M2T1_2,ctl_reg_gp_sel_nuse_ixiypla59M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_nuse_ixiypla59M2T1_3 = (~use_ixiy&pla[59])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla59M2T1_3,ctl_reg_gp_hilo_nuse_ixiypla59M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[59])&(M2&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[59])&(M2&T1);
fMWrite = fMWrite | (~use_ixiy&pla[59])&(M2&T2);
fMWrite = fMWrite | (~use_ixiy&pla[59])&(M2&T3);
setM1 = setM1 | (~use_ixiy&pla[59])&(M2&T3);
fMWrite = fMWrite | (~use_ixiy&pla[59])&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[59])&(M4&T1);
ctl_reg_gp_sel_nuse_ixiypla59M4T1_3 = (~use_ixiy&pla[59])&(M4&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla59M4T1_3,ctl_reg_gp_sel_nuse_ixiypla59M4T1_3})&(op21);
ctl_reg_gp_hilo_nuse_ixiypla59M4T1_4 = (~use_ixiy&pla[59])&(M4&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla59M4T1_4,ctl_reg_gp_hilo_nuse_ixiypla59M4T1_4})&({~rsel0,rsel0});
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[59])&(M4&T1)&(~rsel0);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[59])&(M4&T1)&(rsel0);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[59])&(M4&T1)&(~rsel0);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[59])&(M4&T1)&(rsel0);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[59])&(M4&T1);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[59])&(M4&T1);
fMWrite = fMWrite | (~use_ixiy&pla[59])&(M4&T2);
fMWrite = fMWrite | (~use_ixiy&pla[59])&(M4&T3);
setM1 = setM1 | (~use_ixiy&pla[59])&(M4&T3);
validPLA = validPLA | (pla[40])&(M1&T4);
nextM = nextM | (pla[40])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[40])&(M1&T4);
fMRead = fMRead | (pla[40])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[40])&(M2&T1);
ctl_reg_sys_hilo_pla40M2T1_3 = (pla[40])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla40M2T1_3,ctl_reg_sys_hilo_pla40M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[40])&(M2&T1);
fMRead = fMRead | (pla[40])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[40])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[40])&(M2&T2);
ctl_reg_sys_hilo_pla40M2T2_4 = (pla[40])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla40M2T2_4,ctl_reg_sys_hilo_pla40M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[40])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[40])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[40])&(M2&T2);
fMRead = fMRead | (pla[40])&(M2&T3);
nextM = nextM | (pla[40])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[40])&(M2&T3);
fMRead = fMRead | (pla[40])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[40])&(M3&T1);
ctl_reg_sys_hilo_pla40M3T1_3 = (pla[40])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla40M3T1_3,ctl_reg_sys_hilo_pla40M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[40])&(M3&T1);
ixy_d = ixy_d | (pla[40])&(M3&T1);
fMRead = fMRead | (pla[40])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[40])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[40])&(M3&T2);
ctl_reg_sys_hilo_pla40M3T2_4 = (pla[40])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla40M3T2_4,ctl_reg_sys_hilo_pla40M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[40])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[40])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[40])&(M3&T2);
ixy_d = ixy_d | (pla[40])&(M3&T2);
fMRead = fMRead | (pla[40])&(M3&T3);
ixy_d = ixy_d | (pla[40])&(M3&T3);
ixy_d = ixy_d | (pla[40])&(M3&T4);
nextM = nextM | (pla[40])&(M3&T5);
ctl_mWrite = ctl_mWrite | (pla[40])&(M3&T5);
ixy_d = ixy_d | (pla[40])&(M3&T5);
validPLA = validPLA | (pla[50]&~pla[40])&(M1&T4);
nextM = nextM | (pla[50]&~pla[40])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[50]&~pla[40])&(M1&T4);
fMRead = fMRead | (pla[50]&~pla[40])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[50]&~pla[40])&(M2&T1);
ctl_reg_sys_hilo_pla50npla40M2T1_3 = (pla[50]&~pla[40])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla50npla40M2T1_3,ctl_reg_sys_hilo_pla50npla40M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[50]&~pla[40])&(M2&T1);
fMRead = fMRead | (pla[50]&~pla[40])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[50]&~pla[40])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[50]&~pla[40])&(M2&T2);
ctl_reg_sys_hilo_pla50npla40M2T2_4 = (pla[50]&~pla[40])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla50npla40M2T2_4,ctl_reg_sys_hilo_pla50npla40M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[50]&~pla[40])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[50]&~pla[40])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[50]&~pla[40])&(M2&T2);
fMRead = fMRead | (pla[50]&~pla[40])&(M2&T3);
nextM = nextM | (pla[50]&~pla[40])&(M2&T3);
ctl_mWrite = ctl_mWrite | (pla[50]&~pla[40])&(M2&T3);
fMWrite = fMWrite | (pla[50]&~pla[40])&(M3&T1);
ctl_reg_gp_sel_pla50npla40M3T1_2 = (pla[50]&~pla[40])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla50npla40M3T1_2,ctl_reg_gp_sel_pla50npla40M3T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla50npla40M3T1_3 = (pla[50]&~pla[40])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla50npla40M3T1_3,ctl_reg_gp_hilo_pla50npla40M3T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[50]&~pla[40])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[50]&~pla[40])&(M3&T1);
fMWrite = fMWrite | (pla[50]&~pla[40])&(M3&T2);
fMWrite = fMWrite | (pla[50]&~pla[40])&(M3&T3);
setM1 = setM1 | (pla[50]&~pla[40])&(M3&T3);
fMWrite = fMWrite | (pla[50]&~pla[40])&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[50]&~pla[40])&(M4&T1);
fMWrite = fMWrite | (pla[50]&~pla[40])&(M4&T2);
fMWrite = fMWrite | (pla[50]&~pla[40])&(M4&T3);
setM1 = setM1 | (pla[50]&~pla[40])&(M4&T3);
validPLA = validPLA | (pla[8]&pla[13])&(M1&T4);
nextM = nextM | (pla[8]&pla[13])&(M1&T4);
ctl_mWrite = ctl_mWrite | (pla[8]&pla[13])&(M1&T4);
ctl_reg_gp_sel_pla8pla13M1T4_4 = (pla[8]&pla[13])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla8pla13M1T4_4,ctl_reg_gp_sel_pla8pla13M1T4_4})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla8pla13M1T4_5 = (pla[8]&pla[13])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla8pla13M1T4_5,ctl_reg_gp_hilo_pla8pla13M1T4_5})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[8]&pla[13])&(M1&T4);
ctl_sw_2u = ctl_sw_2u | (pla[8]&pla[13])&(M1&T4);
ctl_sw_1u = ctl_sw_1u | (pla[8]&pla[13])&(M1&T4);
ctl_bus_db_we = ctl_bus_db_we | (pla[8]&pla[13])&(M1&T4);
fMWrite = fMWrite | (pla[8]&pla[13])&(M2&T1);
ctl_reg_gp_sel_pla8pla13M2T1_2 = (pla[8]&pla[13])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla8pla13M2T1_2,ctl_reg_gp_sel_pla8pla13M2T1_2})&(op54);
ctl_reg_gp_hilo_pla8pla13M2T1_3 = (pla[8]&pla[13])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla8pla13M2T1_3,ctl_reg_gp_hilo_pla8pla13M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[8]&pla[13])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[8]&pla[13])&(M2&T1);
fMWrite = fMWrite | (pla[8]&pla[13])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[8]&pla[13])&(M2&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[8]&pla[13])&(M2&T2);
ctl_reg_sys_hilo_pla8pla13M2T2_4 = (pla[8]&pla[13])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla8pla13M2T2_4,ctl_reg_sys_hilo_pla8pla13M2T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[8]&pla[13])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[8]&pla[13])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[8]&pla[13])&(M2&T2);
fMWrite = fMWrite | (pla[8]&pla[13])&(M2&T3);
setM1 = setM1 | (pla[8]&pla[13])&(M2&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[8]&~pla[13])&(M1&T1);
ctl_reg_gp_sel_pla8npla13M1T1_2 = (pla[8]&~pla[13])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla8npla13M1T1_2,ctl_reg_gp_sel_pla8npla13M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla8npla13M1T1_3 = (pla[8]&~pla[13])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla8npla13M1T1_3,ctl_reg_gp_hilo_pla8npla13M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[8]&~pla[13])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[8]&~pla[13])&(M1&T1);
ctl_sw_2d = ctl_sw_2d | (pla[8]&~pla[13])&(M1&T1);
ctl_sw_1d = ctl_sw_1d | (pla[8]&~pla[13])&(M1&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[8]&~pla[13])&(M1&T1);
validPLA = validPLA | (pla[8]&~pla[13])&(M1&T4);
nextM = nextM | (pla[8]&~pla[13])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[8]&~pla[13])&(M1&T4);
fMRead = fMRead | (pla[8]&~pla[13])&(M2&T1);
ctl_reg_gp_sel_pla8npla13M2T1_2 = (pla[8]&~pla[13])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla8npla13M2T1_2,ctl_reg_gp_sel_pla8npla13M2T1_2})&(op54);
ctl_reg_gp_hilo_pla8npla13M2T1_3 = (pla[8]&~pla[13])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla8npla13M2T1_3,ctl_reg_gp_hilo_pla8npla13M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[8]&~pla[13])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[8]&~pla[13])&(M2&T1);
fMRead = fMRead | (pla[8]&~pla[13])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[8]&~pla[13])&(M2&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[8]&~pla[13])&(M2&T2);
ctl_reg_sys_hilo_pla8npla13M2T2_4 = (pla[8]&~pla[13])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla8npla13M2T2_4,ctl_reg_sys_hilo_pla8npla13M2T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[8]&~pla[13])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[8]&~pla[13])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[8]&~pla[13])&(M2&T2);
fMRead = fMRead | (pla[8]&~pla[13])&(M2&T3);
setM1 = setM1 | (pla[8]&~pla[13])&(M2&T3);
validPLA = validPLA | (pla[38]&pla[13])&(M1&T4);
nextM = nextM | (pla[38]&pla[13])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[38]&pla[13])&(M1&T4);
fMRead = fMRead | (pla[38]&pla[13])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[38]&pla[13])&(M2&T1);
ctl_reg_sys_hilo_pla38pla13M2T1_3 = (pla[38]&pla[13])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38pla13M2T1_3,ctl_reg_sys_hilo_pla38pla13M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[38]&pla[13])&(M2&T1);
fMRead = fMRead | (pla[38]&pla[13])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[38]&pla[13])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[38]&pla[13])&(M2&T2);
ctl_reg_sys_hilo_pla38pla13M2T2_4 = (pla[38]&pla[13])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38pla13M2T2_4,ctl_reg_sys_hilo_pla38pla13M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[38]&pla[13])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[38]&pla[13])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[38]&pla[13])&(M2&T2);
fMRead = fMRead | (pla[38]&pla[13])&(M2&T3);
nextM = nextM | (pla[38]&pla[13])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[38]&pla[13])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[38]&pla[13])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[38]&pla[13])&(M2&T3);
ctl_reg_sys_hilo_pla38pla13M2T3_6 = (pla[38]&pla[13])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38pla13M2T3_6,ctl_reg_sys_hilo_pla38pla13M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[38]&pla[13])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[38]&pla[13])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[38]&pla[13])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[38]&pla[13])&(M2&T3);
fMRead = fMRead | (pla[38]&pla[13])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[38]&pla[13])&(M3&T1);
ctl_reg_sys_hilo_pla38pla13M3T1_3 = (pla[38]&pla[13])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38pla13M3T1_3,ctl_reg_sys_hilo_pla38pla13M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[38]&pla[13])&(M3&T1);
fMRead = fMRead | (pla[38]&pla[13])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[38]&pla[13])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[38]&pla[13])&(M3&T2);
ctl_reg_sys_hilo_pla38pla13M3T2_4 = (pla[38]&pla[13])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38pla13M3T2_4,ctl_reg_sys_hilo_pla38pla13M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[38]&pla[13])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[38]&pla[13])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[38]&pla[13])&(M3&T2);
fMRead = fMRead | (pla[38]&pla[13])&(M3&T3);
nextM = nextM | (pla[38]&pla[13])&(M3&T3);
ctl_mWrite = ctl_mWrite | (pla[38]&pla[13])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[38]&pla[13])&(M3&T3);
ctl_reg_sys_hilo_pla38pla13M3T3_5 = (pla[38]&pla[13])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38pla13M3T3_5,ctl_reg_sys_hilo_pla38pla13M3T3_5})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[38]&pla[13])&(M3&T3);
ctl_al_we = ctl_al_we | (pla[38]&pla[13])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[38]&pla[13])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[38]&pla[13])&(M3&T3);
ctl_reg_sys_hilo_pla38pla13M3T3_10 = (pla[38]&pla[13])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38pla13M3T3_10,ctl_reg_sys_hilo_pla38pla13M3T3_10})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[38]&pla[13])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[38]&pla[13])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[38]&pla[13])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[38]&pla[13])&(M3&T3);
fMWrite = fMWrite | (pla[38]&pla[13])&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[38]&pla[13])&(M4&T1);
ctl_reg_gp_sel_pla38pla13M4T1_3 = (pla[38]&pla[13])&(M4&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla38pla13M4T1_3,ctl_reg_gp_sel_pla38pla13M4T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla38pla13M4T1_4 = (pla[38]&pla[13])&(M4&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla38pla13M4T1_4,ctl_reg_gp_hilo_pla38pla13M4T1_4})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[38]&pla[13])&(M4&T1);
ctl_sw_2u = ctl_sw_2u | (pla[38]&pla[13])&(M4&T1);
ctl_sw_1u = ctl_sw_1u | (pla[38]&pla[13])&(M4&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[38]&pla[13])&(M4&T1);
fMWrite = fMWrite | (pla[38]&pla[13])&(M4&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[38]&pla[13])&(M4&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[38]&pla[13])&(M4&T2);
ctl_reg_sys_hilo_pla38pla13M4T2_4 = (pla[38]&pla[13])&(M4&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38pla13M4T2_4,ctl_reg_sys_hilo_pla38pla13M4T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[38]&pla[13])&(M4&T2);
ctl_inc_cy = ctl_inc_cy | (pla[38]&pla[13])&(M4&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[38]&pla[13])&(M4&T2);
fMWrite = fMWrite | (pla[38]&pla[13])&(M4&T3);
setM1 = setM1 | (pla[38]&pla[13])&(M4&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[38]&~pla[13])&(M1&T1);
ctl_reg_gp_sel_pla38npla13M1T1_2 = (pla[38]&~pla[13])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla38npla13M1T1_2,ctl_reg_gp_sel_pla38npla13M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla38npla13M1T1_3 = (pla[38]&~pla[13])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla38npla13M1T1_3,ctl_reg_gp_hilo_pla38npla13M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[38]&~pla[13])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[38]&~pla[13])&(M1&T1);
ctl_sw_2d = ctl_sw_2d | (pla[38]&~pla[13])&(M1&T1);
ctl_sw_1d = ctl_sw_1d | (pla[38]&~pla[13])&(M1&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[38]&~pla[13])&(M1&T1);
validPLA = validPLA | (pla[38]&~pla[13])&(M1&T4);
nextM = nextM | (pla[38]&~pla[13])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[38]&~pla[13])&(M1&T4);
fMRead = fMRead | (pla[38]&~pla[13])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[38]&~pla[13])&(M2&T1);
ctl_reg_sys_hilo_pla38npla13M2T1_3 = (pla[38]&~pla[13])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38npla13M2T1_3,ctl_reg_sys_hilo_pla38npla13M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[38]&~pla[13])&(M2&T1);
fMRead = fMRead | (pla[38]&~pla[13])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[38]&~pla[13])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[38]&~pla[13])&(M2&T2);
ctl_reg_sys_hilo_pla38npla13M2T2_4 = (pla[38]&~pla[13])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38npla13M2T2_4,ctl_reg_sys_hilo_pla38npla13M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[38]&~pla[13])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[38]&~pla[13])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[38]&~pla[13])&(M2&T2);
fMRead = fMRead | (pla[38]&~pla[13])&(M2&T3);
nextM = nextM | (pla[38]&~pla[13])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[38]&~pla[13])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[38]&~pla[13])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[38]&~pla[13])&(M2&T3);
ctl_reg_sys_hilo_pla38npla13M2T3_6 = (pla[38]&~pla[13])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38npla13M2T3_6,ctl_reg_sys_hilo_pla38npla13M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[38]&~pla[13])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[38]&~pla[13])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[38]&~pla[13])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[38]&~pla[13])&(M2&T3);
fMRead = fMRead | (pla[38]&~pla[13])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[38]&~pla[13])&(M3&T1);
ctl_reg_sys_hilo_pla38npla13M3T1_3 = (pla[38]&~pla[13])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38npla13M3T1_3,ctl_reg_sys_hilo_pla38npla13M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[38]&~pla[13])&(M3&T1);
fMRead = fMRead | (pla[38]&~pla[13])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[38]&~pla[13])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[38]&~pla[13])&(M3&T2);
ctl_reg_sys_hilo_pla38npla13M3T2_4 = (pla[38]&~pla[13])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38npla13M3T2_4,ctl_reg_sys_hilo_pla38npla13M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[38]&~pla[13])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[38]&~pla[13])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[38]&~pla[13])&(M3&T2);
fMRead = fMRead | (pla[38]&~pla[13])&(M3&T3);
nextM = nextM | (pla[38]&~pla[13])&(M3&T3);
ctl_mRead = ctl_mRead | (pla[38]&~pla[13])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[38]&~pla[13])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[38]&~pla[13])&(M3&T3);
ctl_reg_sys_hilo_pla38npla13M3T3_6 = (pla[38]&~pla[13])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38npla13M3T3_6,ctl_reg_sys_hilo_pla38npla13M3T3_6})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[38]&~pla[13])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[38]&~pla[13])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[38]&~pla[13])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[38]&~pla[13])&(M3&T3);
fMRead = fMRead | (pla[38]&~pla[13])&(M4&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[38]&~pla[13])&(M4&T1);
ctl_reg_sys_hilo_pla38npla13M4T1_3 = (pla[38]&~pla[13])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38npla13M4T1_3,ctl_reg_sys_hilo_pla38npla13M4T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[38]&~pla[13])&(M4&T1);
ctl_al_we = ctl_al_we | (pla[38]&~pla[13])&(M4&T1);
fMRead = fMRead | (pla[38]&~pla[13])&(M4&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[38]&~pla[13])&(M4&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[38]&~pla[13])&(M4&T2);
ctl_reg_sys_hilo_pla38npla13M4T2_4 = (pla[38]&~pla[13])&(M4&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla38npla13M4T2_4,ctl_reg_sys_hilo_pla38npla13M4T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[38]&~pla[13])&(M4&T2);
ctl_inc_cy = ctl_inc_cy | (pla[38]&~pla[13])&(M4&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[38]&~pla[13])&(M4&T2);
fMRead = fMRead | (pla[38]&~pla[13])&(M4&T3);
setM1 = setM1 | (pla[38]&~pla[13])&(M4&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[83])&(M1&T1);
ctl_reg_gp_sel_pla83M1T1_2 = (pla[83])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla83M1T1_2,ctl_reg_gp_sel_pla83M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla83M1T1_3 = (pla[83])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla83M1T1_3,ctl_reg_gp_hilo_pla83M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[83])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[83])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[83])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[83])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[83])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[83])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[83])&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (pla[83])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (pla[83])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[83])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[83])&(M1&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[83])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[83])&(M1&T1);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[83])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[83])&(M1&T1);
ctl_pf_sel_pla83M1T1_19 = (pla[83])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla83M1T1_19,ctl_pf_sel_pla83M1T1_19})&(`PFSEL_IFF2);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[83])&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[83])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[83])&(M1&T2);
ctl_reg_gp_sel_pla83M1T2_2 = (pla[83])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla83M1T2_2,ctl_reg_gp_sel_pla83M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla83M1T2_3 = (pla[83])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla83M1T2_3,ctl_reg_gp_hilo_pla83M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[83])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[83])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[83])&(M1&T2);
ctl_reg_gp_sel_pla83M1T3_1 = (pla[83])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla83M1T3_1,ctl_reg_gp_sel_pla83M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla83M1T3_2 = (pla[83])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla83M1T3_2,ctl_reg_gp_hilo_pla83M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[83])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[83])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[83])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[83])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[83])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[83])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[83])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[83])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[83])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[83])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[83])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[83])&(M1&T3);
validPLA = validPLA | (pla[83])&(M1&T4);
ctl_reg_sel_ir = ctl_reg_sel_ir | (pla[83])&(M1&T4);
ctl_reg_sys_hilo_pla83M1T4_3 = (pla[83])&(M1&T4);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla83M1T4_3,ctl_reg_sys_hilo_pla83M1T4_3})&({~op3,op3});
ctl_sw_4u = ctl_sw_4u | (pla[83])&(M1&T4);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[83])&(M1&T4)&(~rsel3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[83])&(M1&T4)&(rsel3);
ctl_sw_2u = ctl_sw_2u | (pla[83])&(M1&T4)&(~rsel3);
ctl_sw_2d = ctl_sw_2d | (pla[83])&(M1&T4)&(rsel3);
ctl_flags_alu = ctl_flags_alu | (pla[83])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[83])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[83])&(M1&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[83])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[83])&(M1&T4);
ctl_alu_core_R = ctl_alu_core_R | (pla[83])&(M1&T4);
ctl_alu_core_V = ctl_alu_core_V | (pla[83])&(M1&T4);
ctl_alu_core_S = ctl_alu_core_S | (pla[83])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[83])&(M1&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[83])&(M1&T4);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[83])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[83])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[83])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[83])&(M1&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[83])&(M1&T4);
setM1 = setM1 | (pla[83])&(M1&T5);
ctl_reg_gp_sel_pla57M1T3_1 = (pla[57])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla57M1T3_1,ctl_reg_gp_sel_pla57M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla57M1T3_2 = (pla[57])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla57M1T3_2,ctl_reg_gp_hilo_pla57M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[57])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[57])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[57])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[57])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[57])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[57])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[57])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[57])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[57])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[57])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[57])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[57])&(M1&T3);
validPLA = validPLA | (pla[57])&(M1&T4);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[57])&(M1&T4);
ctl_reg_sel_ir = ctl_reg_sel_ir | (pla[57])&(M1&T4);
ctl_reg_sys_hilo_pla57M1T4_4 = (pla[57])&(M1&T4);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla57M1T4_4,ctl_reg_sys_hilo_pla57M1T4_4})&({~op3,op3});
ctl_sw_4d = ctl_sw_4d | (pla[57])&(M1&T4);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[57])&(M1&T4);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[57])&(M1&T4);
ctl_sw_2u = ctl_sw_2u | (pla[57])&(M1&T4);
ctl_alu_oe = ctl_alu_oe | (pla[57])&(M1&T4);
ctl_alu_op1_oe = ctl_alu_op1_oe | (pla[57])&(M1&T4);
setM1 = setM1 | (pla[57])&(M1&T5);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[7])&(M1&T1);
ctl_reg_gp_sel_pla7M1T1_2 = (pla[7])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla7M1T1_2,ctl_reg_gp_sel_pla7M1T1_2})&(op54);
ctl_reg_gp_hilo_pla7M1T1_3 = (pla[7])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla7M1T1_3,ctl_reg_gp_hilo_pla7M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[7])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[7])&(M1&T1);
ctl_sw_2d = ctl_sw_2d | (pla[7])&(M1&T1);
ctl_sw_1d = ctl_sw_1d | (pla[7])&(M1&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[7])&(M1&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[7])&(M1&T1);
validPLA = validPLA | (pla[7])&(M1&T4);
nextM = nextM | (pla[7])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[7])&(M1&T4);
fMRead = fMRead | (pla[7])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[7])&(M2&T1);
ctl_reg_sys_hilo_pla7M2T1_3 = (pla[7])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla7M2T1_3,ctl_reg_sys_hilo_pla7M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[7])&(M2&T1);
fMRead = fMRead | (pla[7])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[7])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[7])&(M2&T2);
ctl_reg_sys_hilo_pla7M2T2_4 = (pla[7])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla7M2T2_4,ctl_reg_sys_hilo_pla7M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[7])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[7])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[7])&(M2&T2);
fMRead = fMRead | (pla[7])&(M2&T3);
nextM = nextM | (pla[7])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[7])&(M2&T3);
fMRead = fMRead | (pla[7])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[7])&(M3&T1);
ctl_reg_sys_hilo_pla7M3T1_3 = (pla[7])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla7M3T1_3,ctl_reg_sys_hilo_pla7M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[7])&(M3&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[7])&(M3&T1);
ctl_reg_gp_sel_pla7M3T1_6 = (pla[7])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla7M3T1_6,ctl_reg_gp_sel_pla7M3T1_6})&(op54);
ctl_reg_gp_hilo_pla7M3T1_7 = (pla[7])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla7M3T1_7,ctl_reg_gp_hilo_pla7M3T1_7})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[7])&(M3&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[7])&(M3&T1);
ctl_sw_2d = ctl_sw_2d | (pla[7])&(M3&T1);
ctl_sw_1d = ctl_sw_1d | (pla[7])&(M3&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[7])&(M3&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[7])&(M3&T1);
fMRead = fMRead | (pla[7])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[7])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[7])&(M3&T2);
ctl_reg_sys_hilo_pla7M3T2_4 = (pla[7])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla7M3T2_4,ctl_reg_sys_hilo_pla7M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[7])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[7])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[7])&(M3&T2);
fMRead = fMRead | (pla[7])&(M3&T3);
setM1 = setM1 | (pla[7])&(M3&T3);
validPLA = validPLA | (pla[30]&pla[13])&(M1&T4);
nextM = nextM | (pla[30]&pla[13])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[30]&pla[13])&(M1&T4);
fMRead = fMRead | (pla[30]&pla[13])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[30]&pla[13])&(M2&T1);
ctl_reg_sys_hilo_pla30pla13M2T1_3 = (pla[30]&pla[13])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30pla13M2T1_3,ctl_reg_sys_hilo_pla30pla13M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[30]&pla[13])&(M2&T1);
fMRead = fMRead | (pla[30]&pla[13])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[30]&pla[13])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[30]&pla[13])&(M2&T2);
ctl_reg_sys_hilo_pla30pla13M2T2_4 = (pla[30]&pla[13])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30pla13M2T2_4,ctl_reg_sys_hilo_pla30pla13M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[30]&pla[13])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[30]&pla[13])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[30]&pla[13])&(M2&T2);
fMRead = fMRead | (pla[30]&pla[13])&(M2&T3);
nextM = nextM | (pla[30]&pla[13])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[30]&pla[13])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[30]&pla[13])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&pla[13])&(M2&T3);
ctl_reg_sys_hilo_pla30pla13M2T3_6 = (pla[30]&pla[13])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30pla13M2T3_6,ctl_reg_sys_hilo_pla30pla13M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[30]&pla[13])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[30]&pla[13])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[30]&pla[13])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[30]&pla[13])&(M2&T3);
fMRead = fMRead | (pla[30]&pla[13])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[30]&pla[13])&(M3&T1);
ctl_reg_sys_hilo_pla30pla13M3T1_3 = (pla[30]&pla[13])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30pla13M3T1_3,ctl_reg_sys_hilo_pla30pla13M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[30]&pla[13])&(M3&T1);
fMRead = fMRead | (pla[30]&pla[13])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[30]&pla[13])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[30]&pla[13])&(M3&T2);
ctl_reg_sys_hilo_pla30pla13M3T2_4 = (pla[30]&pla[13])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30pla13M3T2_4,ctl_reg_sys_hilo_pla30pla13M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[30]&pla[13])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[30]&pla[13])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[30]&pla[13])&(M3&T2);
fMRead = fMRead | (pla[30]&pla[13])&(M3&T3);
nextM = nextM | (pla[30]&pla[13])&(M3&T3);
ctl_mWrite = ctl_mWrite | (pla[30]&pla[13])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&pla[13])&(M3&T3);
ctl_reg_sys_hilo_pla30pla13M3T3_5 = (pla[30]&pla[13])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30pla13M3T3_5,ctl_reg_sys_hilo_pla30pla13M3T3_5})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[30]&pla[13])&(M3&T3);
ctl_al_we = ctl_al_we | (pla[30]&pla[13])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[30]&pla[13])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&pla[13])&(M3&T3);
ctl_reg_sys_hilo_pla30pla13M3T3_10 = (pla[30]&pla[13])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30pla13M3T3_10,ctl_reg_sys_hilo_pla30pla13M3T3_10})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[30]&pla[13])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[30]&pla[13])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[30]&pla[13])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[30]&pla[13])&(M3&T3);
fMWrite = fMWrite | (pla[30]&pla[13])&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[30]&pla[13])&(M4&T1);
ctl_reg_gp_sel_pla30pla13M4T1_3 = (pla[30]&pla[13])&(M4&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla30pla13M4T1_3,ctl_reg_gp_sel_pla30pla13M4T1_3})&(op54);
ctl_reg_gp_hilo_pla30pla13M4T1_4 = (pla[30]&pla[13])&(M4&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla30pla13M4T1_4,ctl_reg_gp_hilo_pla30pla13M4T1_4})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[30]&pla[13])&(M4&T1);
ctl_sw_1u = ctl_sw_1u | (pla[30]&pla[13])&(M4&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[30]&pla[13])&(M4&T1);
fMWrite = fMWrite | (pla[30]&pla[13])&(M4&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[30]&pla[13])&(M4&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&pla[13])&(M4&T2);
ctl_reg_sys_hilo_pla30pla13M4T2_4 = (pla[30]&pla[13])&(M4&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30pla13M4T2_4,ctl_reg_sys_hilo_pla30pla13M4T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[30]&pla[13])&(M4&T2);
ctl_inc_cy = ctl_inc_cy | (pla[30]&pla[13])&(M4&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[30]&pla[13])&(M4&T2);
fMWrite = fMWrite | (pla[30]&pla[13])&(M4&T3);
nextM = nextM | (pla[30]&pla[13])&(M4&T3);
ctl_mWrite = ctl_mWrite | (pla[30]&pla[13])&(M4&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&pla[13])&(M4&T3);
ctl_reg_sys_hilo_pla30pla13M4T3_5 = (pla[30]&pla[13])&(M4&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30pla13M4T3_5,ctl_reg_sys_hilo_pla30pla13M4T3_5})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[30]&pla[13])&(M4&T3);
ctl_al_we = ctl_al_we | (pla[30]&pla[13])&(M4&T3);
fMWrite = fMWrite | (pla[30]&pla[13])&(M5&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[30]&pla[13])&(M5&T1);
ctl_reg_gp_sel_pla30pla13M5T1_3 = (pla[30]&pla[13])&(M5&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla30pla13M5T1_3,ctl_reg_gp_sel_pla30pla13M5T1_3})&(op54);
ctl_reg_gp_hilo_pla30pla13M5T1_4 = (pla[30]&pla[13])&(M5&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla30pla13M5T1_4,ctl_reg_gp_hilo_pla30pla13M5T1_4})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[30]&pla[13])&(M5&T1);
ctl_sw_2u = ctl_sw_2u | (pla[30]&pla[13])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (pla[30]&pla[13])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[30]&pla[13])&(M5&T1);
fMWrite = fMWrite | (pla[30]&pla[13])&(M5&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[30]&pla[13])&(M5&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&pla[13])&(M5&T2);
ctl_reg_sys_hilo_pla30pla13M5T2_4 = (pla[30]&pla[13])&(M5&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30pla13M5T2_4,ctl_reg_sys_hilo_pla30pla13M5T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[30]&pla[13])&(M5&T2);
ctl_inc_cy = ctl_inc_cy | (pla[30]&pla[13])&(M5&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[30]&pla[13])&(M5&T2);
fMWrite = fMWrite | (pla[30]&pla[13])&(M5&T3);
setM1 = setM1 | (pla[30]&pla[13])&(M5&T3);
validPLA = validPLA | (pla[30]&~pla[13])&(M1&T4);
nextM = nextM | (pla[30]&~pla[13])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[30]&~pla[13])&(M1&T4);
fMRead = fMRead | (pla[30]&~pla[13])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[30]&~pla[13])&(M2&T1);
ctl_reg_sys_hilo_pla30npla13M2T1_3 = (pla[30]&~pla[13])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30npla13M2T1_3,ctl_reg_sys_hilo_pla30npla13M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[30]&~pla[13])&(M2&T1);
fMRead = fMRead | (pla[30]&~pla[13])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[30]&~pla[13])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[30]&~pla[13])&(M2&T2);
ctl_reg_sys_hilo_pla30npla13M2T2_4 = (pla[30]&~pla[13])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30npla13M2T2_4,ctl_reg_sys_hilo_pla30npla13M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[30]&~pla[13])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[30]&~pla[13])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[30]&~pla[13])&(M2&T2);
fMRead = fMRead | (pla[30]&~pla[13])&(M2&T3);
nextM = nextM | (pla[30]&~pla[13])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[30]&~pla[13])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[30]&~pla[13])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&~pla[13])&(M2&T3);
ctl_reg_sys_hilo_pla30npla13M2T3_6 = (pla[30]&~pla[13])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30npla13M2T3_6,ctl_reg_sys_hilo_pla30npla13M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[30]&~pla[13])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[30]&~pla[13])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[30]&~pla[13])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[30]&~pla[13])&(M2&T3);
fMRead = fMRead | (pla[30]&~pla[13])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[30]&~pla[13])&(M3&T1);
ctl_reg_sys_hilo_pla30npla13M3T1_3 = (pla[30]&~pla[13])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30npla13M3T1_3,ctl_reg_sys_hilo_pla30npla13M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[30]&~pla[13])&(M3&T1);
fMRead = fMRead | (pla[30]&~pla[13])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[30]&~pla[13])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[30]&~pla[13])&(M3&T2);
ctl_reg_sys_hilo_pla30npla13M3T2_4 = (pla[30]&~pla[13])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30npla13M3T2_4,ctl_reg_sys_hilo_pla30npla13M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[30]&~pla[13])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[30]&~pla[13])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[30]&~pla[13])&(M3&T2);
fMRead = fMRead | (pla[30]&~pla[13])&(M3&T3);
nextM = nextM | (pla[30]&~pla[13])&(M3&T3);
ctl_mRead = ctl_mRead | (pla[30]&~pla[13])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[30]&~pla[13])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&~pla[13])&(M3&T3);
ctl_reg_sys_hilo_pla30npla13M3T3_6 = (pla[30]&~pla[13])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30npla13M3T3_6,ctl_reg_sys_hilo_pla30npla13M3T3_6})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[30]&~pla[13])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[30]&~pla[13])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[30]&~pla[13])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[30]&~pla[13])&(M3&T3);
fMRead = fMRead | (pla[30]&~pla[13])&(M4&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&~pla[13])&(M4&T1);
ctl_reg_sys_hilo_pla30npla13M4T1_3 = (pla[30]&~pla[13])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30npla13M4T1_3,ctl_reg_sys_hilo_pla30npla13M4T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[30]&~pla[13])&(M4&T1);
ctl_al_we = ctl_al_we | (pla[30]&~pla[13])&(M4&T1);
fMRead = fMRead | (pla[30]&~pla[13])&(M4&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[30]&~pla[13])&(M4&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&~pla[13])&(M4&T2);
ctl_reg_sys_hilo_pla30npla13M4T2_4 = (pla[30]&~pla[13])&(M4&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30npla13M4T2_4,ctl_reg_sys_hilo_pla30npla13M4T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[30]&~pla[13])&(M4&T2);
ctl_inc_cy = ctl_inc_cy | (pla[30]&~pla[13])&(M4&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[30]&~pla[13])&(M4&T2);
fMRead = fMRead | (pla[30]&~pla[13])&(M4&T3);
nextM = nextM | (pla[30]&~pla[13])&(M4&T3);
ctl_mRead = ctl_mRead | (pla[30]&~pla[13])&(M4&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[30]&~pla[13])&(M4&T3);
ctl_reg_gp_sel_pla30npla13M4T3_5 = (pla[30]&~pla[13])&(M4&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla30npla13M4T3_5,ctl_reg_gp_sel_pla30npla13M4T3_5})&(op54);
ctl_reg_gp_hilo_pla30npla13M4T3_6 = (pla[30]&~pla[13])&(M4&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla30npla13M4T3_6,ctl_reg_gp_hilo_pla30npla13M4T3_6})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[30]&~pla[13])&(M4&T3);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[30]&~pla[13])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (pla[30]&~pla[13])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (pla[30]&~pla[13])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[30]&~pla[13])&(M4&T3);
fMRead = fMRead | (pla[30]&~pla[13])&(M5&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&~pla[13])&(M5&T1);
ctl_reg_sys_hilo_pla30npla13M5T1_3 = (pla[30]&~pla[13])&(M5&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30npla13M5T1_3,ctl_reg_sys_hilo_pla30npla13M5T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[30]&~pla[13])&(M5&T1);
ctl_al_we = ctl_al_we | (pla[30]&~pla[13])&(M5&T1);
fMRead = fMRead | (pla[30]&~pla[13])&(M5&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[30]&~pla[13])&(M5&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[30]&~pla[13])&(M5&T2);
ctl_reg_sys_hilo_pla30npla13M5T2_4 = (pla[30]&~pla[13])&(M5&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla30npla13M5T2_4,ctl_reg_sys_hilo_pla30npla13M5T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[30]&~pla[13])&(M5&T2);
ctl_inc_cy = ctl_inc_cy | (pla[30]&~pla[13])&(M5&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[30]&~pla[13])&(M5&T2);
fMRead = fMRead | (pla[30]&~pla[13])&(M5&T3);
setM1 = setM1 | (pla[30]&~pla[13])&(M5&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[30]&~pla[13])&(M5&T3);
ctl_reg_gp_sel_pla30npla13M5T3_4 = (pla[30]&~pla[13])&(M5&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla30npla13M5T3_4,ctl_reg_gp_sel_pla30npla13M5T3_4})&(op54);
ctl_reg_gp_hilo_pla30npla13M5T3_5 = (pla[30]&~pla[13])&(M5&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla30npla13M5T3_5,ctl_reg_gp_hilo_pla30npla13M5T3_5})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[30]&~pla[13])&(M5&T3);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[30]&~pla[13])&(M5&T3);
ctl_sw_2d = ctl_sw_2d | (pla[30]&~pla[13])&(M5&T3);
ctl_sw_1d = ctl_sw_1d | (pla[30]&~pla[13])&(M5&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[30]&~pla[13])&(M5&T3);
validPLA = validPLA | (pla[31]&pla[33])&(M1&T4);
nextM = nextM | (pla[31]&pla[33])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[31]&pla[33])&(M1&T4);
fMRead = fMRead | (pla[31]&pla[33])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[31]&pla[33])&(M2&T1);
ctl_reg_sys_hilo_pla31pla33M2T1_3 = (pla[31]&pla[33])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31pla33M2T1_3,ctl_reg_sys_hilo_pla31pla33M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[31]&pla[33])&(M2&T1);
fMRead = fMRead | (pla[31]&pla[33])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[31]&pla[33])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[31]&pla[33])&(M2&T2);
ctl_reg_sys_hilo_pla31pla33M2T2_4 = (pla[31]&pla[33])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31pla33M2T2_4,ctl_reg_sys_hilo_pla31pla33M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[31]&pla[33])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[31]&pla[33])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[31]&pla[33])&(M2&T2);
fMRead = fMRead | (pla[31]&pla[33])&(M2&T3);
nextM = nextM | (pla[31]&pla[33])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[31]&pla[33])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[31]&pla[33])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&pla[33])&(M2&T3);
ctl_reg_sys_hilo_pla31pla33M2T3_6 = (pla[31]&pla[33])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31pla33M2T3_6,ctl_reg_sys_hilo_pla31pla33M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[31]&pla[33])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[31]&pla[33])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[31]&pla[33])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[31]&pla[33])&(M2&T3);
fMRead = fMRead | (pla[31]&pla[33])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[31]&pla[33])&(M3&T1);
ctl_reg_sys_hilo_pla31pla33M3T1_3 = (pla[31]&pla[33])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31pla33M3T1_3,ctl_reg_sys_hilo_pla31pla33M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[31]&pla[33])&(M3&T1);
fMRead = fMRead | (pla[31]&pla[33])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[31]&pla[33])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[31]&pla[33])&(M3&T2);
ctl_reg_sys_hilo_pla31pla33M3T2_4 = (pla[31]&pla[33])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31pla33M3T2_4,ctl_reg_sys_hilo_pla31pla33M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[31]&pla[33])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[31]&pla[33])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[31]&pla[33])&(M3&T2);
fMRead = fMRead | (pla[31]&pla[33])&(M3&T3);
nextM = nextM | (pla[31]&pla[33])&(M3&T3);
ctl_mWrite = ctl_mWrite | (pla[31]&pla[33])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&pla[33])&(M3&T3);
ctl_reg_sys_hilo_pla31pla33M3T3_5 = (pla[31]&pla[33])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31pla33M3T3_5,ctl_reg_sys_hilo_pla31pla33M3T3_5})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[31]&pla[33])&(M3&T3);
ctl_al_we = ctl_al_we | (pla[31]&pla[33])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[31]&pla[33])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&pla[33])&(M3&T3);
ctl_reg_sys_hilo_pla31pla33M3T3_10 = (pla[31]&pla[33])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31pla33M3T3_10,ctl_reg_sys_hilo_pla31pla33M3T3_10})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[31]&pla[33])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[31]&pla[33])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[31]&pla[33])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[31]&pla[33])&(M3&T3);
fMWrite = fMWrite | (pla[31]&pla[33])&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[31]&pla[33])&(M4&T1);
ctl_reg_gp_sel_pla31pla33M4T1_3 = (pla[31]&pla[33])&(M4&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla31pla33M4T1_3,ctl_reg_gp_sel_pla31pla33M4T1_3})&(op54);
ctl_reg_gp_hilo_pla31pla33M4T1_4 = (pla[31]&pla[33])&(M4&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla31pla33M4T1_4,ctl_reg_gp_hilo_pla31pla33M4T1_4})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[31]&pla[33])&(M4&T1);
ctl_sw_1u = ctl_sw_1u | (pla[31]&pla[33])&(M4&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[31]&pla[33])&(M4&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[31]&pla[33])&(M4&T1);
fMWrite = fMWrite | (pla[31]&pla[33])&(M4&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[31]&pla[33])&(M4&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&pla[33])&(M4&T2);
ctl_reg_sys_hilo_pla31pla33M4T2_4 = (pla[31]&pla[33])&(M4&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31pla33M4T2_4,ctl_reg_sys_hilo_pla31pla33M4T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[31]&pla[33])&(M4&T2);
ctl_inc_cy = ctl_inc_cy | (pla[31]&pla[33])&(M4&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[31]&pla[33])&(M4&T2);
fMWrite = fMWrite | (pla[31]&pla[33])&(M4&T3);
nextM = nextM | (pla[31]&pla[33])&(M4&T3);
ctl_mWrite = ctl_mWrite | (pla[31]&pla[33])&(M4&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&pla[33])&(M4&T3);
ctl_reg_sys_hilo_pla31pla33M4T3_5 = (pla[31]&pla[33])&(M4&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31pla33M4T3_5,ctl_reg_sys_hilo_pla31pla33M4T3_5})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[31]&pla[33])&(M4&T3);
ctl_al_we = ctl_al_we | (pla[31]&pla[33])&(M4&T3);
fMWrite = fMWrite | (pla[31]&pla[33])&(M5&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[31]&pla[33])&(M5&T1);
ctl_reg_gp_sel_pla31pla33M5T1_3 = (pla[31]&pla[33])&(M5&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla31pla33M5T1_3,ctl_reg_gp_sel_pla31pla33M5T1_3})&(op54);
ctl_reg_gp_hilo_pla31pla33M5T1_4 = (pla[31]&pla[33])&(M5&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla31pla33M5T1_4,ctl_reg_gp_hilo_pla31pla33M5T1_4})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[31]&pla[33])&(M5&T1);
ctl_sw_2u = ctl_sw_2u | (pla[31]&pla[33])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (pla[31]&pla[33])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[31]&pla[33])&(M5&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[31]&pla[33])&(M5&T1);
fMWrite = fMWrite | (pla[31]&pla[33])&(M5&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[31]&pla[33])&(M5&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&pla[33])&(M5&T2);
ctl_reg_sys_hilo_pla31pla33M5T2_4 = (pla[31]&pla[33])&(M5&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31pla33M5T2_4,ctl_reg_sys_hilo_pla31pla33M5T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[31]&pla[33])&(M5&T2);
ctl_inc_cy = ctl_inc_cy | (pla[31]&pla[33])&(M5&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[31]&pla[33])&(M5&T2);
fMWrite = fMWrite | (pla[31]&pla[33])&(M5&T3);
setM1 = setM1 | (pla[31]&pla[33])&(M5&T3);
validPLA = validPLA | (pla[31]&~pla[33])&(M1&T4);
nextM = nextM | (pla[31]&~pla[33])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[31]&~pla[33])&(M1&T4);
fMRead = fMRead | (pla[31]&~pla[33])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[31]&~pla[33])&(M2&T1);
ctl_reg_sys_hilo_pla31npla33M2T1_3 = (pla[31]&~pla[33])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31npla33M2T1_3,ctl_reg_sys_hilo_pla31npla33M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[31]&~pla[33])&(M2&T1);
fMRead = fMRead | (pla[31]&~pla[33])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[31]&~pla[33])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[31]&~pla[33])&(M2&T2);
ctl_reg_sys_hilo_pla31npla33M2T2_4 = (pla[31]&~pla[33])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31npla33M2T2_4,ctl_reg_sys_hilo_pla31npla33M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[31]&~pla[33])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[31]&~pla[33])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[31]&~pla[33])&(M2&T2);
fMRead = fMRead | (pla[31]&~pla[33])&(M2&T3);
nextM = nextM | (pla[31]&~pla[33])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[31]&~pla[33])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[31]&~pla[33])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&~pla[33])&(M2&T3);
ctl_reg_sys_hilo_pla31npla33M2T3_6 = (pla[31]&~pla[33])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31npla33M2T3_6,ctl_reg_sys_hilo_pla31npla33M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[31]&~pla[33])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[31]&~pla[33])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[31]&~pla[33])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[31]&~pla[33])&(M2&T3);
fMRead = fMRead | (pla[31]&~pla[33])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[31]&~pla[33])&(M3&T1);
ctl_reg_sys_hilo_pla31npla33M3T1_3 = (pla[31]&~pla[33])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31npla33M3T1_3,ctl_reg_sys_hilo_pla31npla33M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[31]&~pla[33])&(M3&T1);
fMRead = fMRead | (pla[31]&~pla[33])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[31]&~pla[33])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[31]&~pla[33])&(M3&T2);
ctl_reg_sys_hilo_pla31npla33M3T2_4 = (pla[31]&~pla[33])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31npla33M3T2_4,ctl_reg_sys_hilo_pla31npla33M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[31]&~pla[33])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[31]&~pla[33])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[31]&~pla[33])&(M3&T2);
fMRead = fMRead | (pla[31]&~pla[33])&(M3&T3);
nextM = nextM | (pla[31]&~pla[33])&(M3&T3);
ctl_mRead = ctl_mRead | (pla[31]&~pla[33])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[31]&~pla[33])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&~pla[33])&(M3&T3);
ctl_reg_sys_hilo_pla31npla33M3T3_6 = (pla[31]&~pla[33])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31npla33M3T3_6,ctl_reg_sys_hilo_pla31npla33M3T3_6})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[31]&~pla[33])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[31]&~pla[33])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[31]&~pla[33])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[31]&~pla[33])&(M3&T3);
fMRead = fMRead | (pla[31]&~pla[33])&(M4&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&~pla[33])&(M4&T1);
ctl_reg_sys_hilo_pla31npla33M4T1_3 = (pla[31]&~pla[33])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31npla33M4T1_3,ctl_reg_sys_hilo_pla31npla33M4T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[31]&~pla[33])&(M4&T1);
ctl_al_we = ctl_al_we | (pla[31]&~pla[33])&(M4&T1);
fMRead = fMRead | (pla[31]&~pla[33])&(M4&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[31]&~pla[33])&(M4&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&~pla[33])&(M4&T2);
ctl_reg_sys_hilo_pla31npla33M4T2_4 = (pla[31]&~pla[33])&(M4&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31npla33M4T2_4,ctl_reg_sys_hilo_pla31npla33M4T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[31]&~pla[33])&(M4&T2);
ctl_inc_cy = ctl_inc_cy | (pla[31]&~pla[33])&(M4&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[31]&~pla[33])&(M4&T2);
fMRead = fMRead | (pla[31]&~pla[33])&(M4&T3);
nextM = nextM | (pla[31]&~pla[33])&(M4&T3);
ctl_mRead = ctl_mRead | (pla[31]&~pla[33])&(M4&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[31]&~pla[33])&(M4&T3);
ctl_reg_gp_sel_pla31npla33M4T3_5 = (pla[31]&~pla[33])&(M4&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla31npla33M4T3_5,ctl_reg_gp_sel_pla31npla33M4T3_5})&(op54);
ctl_reg_gp_hilo_pla31npla33M4T3_6 = (pla[31]&~pla[33])&(M4&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla31npla33M4T3_6,ctl_reg_gp_hilo_pla31npla33M4T3_6})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[31]&~pla[33])&(M4&T3);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[31]&~pla[33])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (pla[31]&~pla[33])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (pla[31]&~pla[33])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[31]&~pla[33])&(M4&T3);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[31]&~pla[33])&(M4&T3);
fMRead = fMRead | (pla[31]&~pla[33])&(M5&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&~pla[33])&(M5&T1);
ctl_reg_sys_hilo_pla31npla33M5T1_3 = (pla[31]&~pla[33])&(M5&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31npla33M5T1_3,ctl_reg_sys_hilo_pla31npla33M5T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[31]&~pla[33])&(M5&T1);
ctl_al_we = ctl_al_we | (pla[31]&~pla[33])&(M5&T1);
fMRead = fMRead | (pla[31]&~pla[33])&(M5&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[31]&~pla[33])&(M5&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[31]&~pla[33])&(M5&T2);
ctl_reg_sys_hilo_pla31npla33M5T2_4 = (pla[31]&~pla[33])&(M5&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla31npla33M5T2_4,ctl_reg_sys_hilo_pla31npla33M5T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[31]&~pla[33])&(M5&T2);
ctl_inc_cy = ctl_inc_cy | (pla[31]&~pla[33])&(M5&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[31]&~pla[33])&(M5&T2);
fMRead = fMRead | (pla[31]&~pla[33])&(M5&T3);
setM1 = setM1 | (pla[31]&~pla[33])&(M5&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[31]&~pla[33])&(M5&T3);
ctl_reg_gp_sel_pla31npla33M5T3_4 = (pla[31]&~pla[33])&(M5&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla31npla33M5T3_4,ctl_reg_gp_sel_pla31npla33M5T3_4})&(op54);
ctl_reg_gp_hilo_pla31npla33M5T3_5 = (pla[31]&~pla[33])&(M5&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla31npla33M5T3_5,ctl_reg_gp_hilo_pla31npla33M5T3_5})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[31]&~pla[33])&(M5&T3);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[31]&~pla[33])&(M5&T3);
ctl_sw_2d = ctl_sw_2d | (pla[31]&~pla[33])&(M5&T3);
ctl_sw_1d = ctl_sw_1d | (pla[31]&~pla[33])&(M5&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[31]&~pla[33])&(M5&T3);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[31]&~pla[33])&(M5&T3);
validPLA = validPLA | (pla[5])&(M1&T4);
ctl_reg_gp_sel_pla5M1T4_2 = (pla[5])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla5M1T4_2,ctl_reg_gp_sel_pla5M1T4_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla5M1T4_3 = (pla[5])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla5M1T4_3,ctl_reg_gp_hilo_pla5M1T4_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[5])&(M1&T4);
ctl_al_we = ctl_al_we | (pla[5])&(M1&T4);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[5])&(M1&T5);
ctl_reg_gp_sel_pla5M1T5_2 = (pla[5])&(M1&T5);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla5M1T5_2,ctl_reg_gp_sel_pla5M1T5_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla5M1T5_3 = (pla[5])&(M1&T5);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla5M1T5_3,ctl_reg_gp_hilo_pla5M1T5_3})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[5])&(M1&T5);
ctl_sw_4u = ctl_sw_4u | (pla[5])&(M1&T5);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[5])&(M1&T5);
setM1 = setM1 | (pla[5])&(M1&T6);
validPLA = validPLA | (pla[23]&pla[16])&(M1&T4);
nextM = nextM | (pla[23]&pla[16])&(M1&T5);
ctl_mWrite = ctl_mWrite | (pla[23]&pla[16])&(M1&T5);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[23]&pla[16])&(M1&T5);
ctl_reg_gp_sel_pla23pla16M1T5_4 = (pla[23]&pla[16])&(M1&T5);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23pla16M1T5_4,ctl_reg_gp_sel_pla23pla16M1T5_4})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla23pla16M1T5_5 = (pla[23]&pla[16])&(M1&T5);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23pla16M1T5_5,ctl_reg_gp_hilo_pla23pla16M1T5_5})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[23]&pla[16])&(M1&T5);
ctl_inc_cy = ctl_inc_cy | (pla[23]&pla[16])&(M1&T5)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[23]&pla[16])&(M1&T5);
ctl_al_we = ctl_al_we | (pla[23]&pla[16])&(M1&T5);
fMWrite = fMWrite | (pla[23]&pla[16])&(M2&T1);
ctl_inc_cy = ctl_inc_cy | (pla[23]&pla[16])&(M2&T1)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[23]&pla[16])&(M2&T1);
ctl_apin_mux = ctl_apin_mux | (pla[23]&pla[16])&(M2&T1);
ctl_reg_gp_sel_pla23pla16M2T1_5 = (pla[23]&pla[16])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23pla16M2T1_5,ctl_reg_gp_sel_pla23pla16M2T1_5})&(op54);
ctl_reg_gp_hilo_pla23pla16M2T1_6 = (pla[23]&pla[16])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23pla16M2T1_6,ctl_reg_gp_hilo_pla23pla16M2T1_6})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[23]&pla[16])&(M2&T1);
ctl_sw_2u = ctl_sw_2u | (pla[23]&pla[16])&(M2&T1);
ctl_sw_1u = ctl_sw_1u | (pla[23]&pla[16])&(M2&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[23]&pla[16])&(M2&T1);
fMWrite = fMWrite | (pla[23]&pla[16])&(M2&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[23]&pla[16])&(M2&T2);
ctl_reg_gp_sel_pla23pla16M2T2_3 = (pla[23]&pla[16])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23pla16M2T2_3,ctl_reg_gp_sel_pla23pla16M2T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla23pla16M2T2_4 = (pla[23]&pla[16])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23pla16M2T2_4,ctl_reg_gp_hilo_pla23pla16M2T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[23]&pla[16])&(M2&T2);
ctl_sw_4u = ctl_sw_4u | (pla[23]&pla[16])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[23]&pla[16])&(M2&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[23]&pla[16])&(M2&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[23]&pla[16])&(M2&T2);
fMWrite = fMWrite | (pla[23]&pla[16])&(M2&T3);
nextM = nextM | (pla[23]&pla[16])&(M2&T3);
ctl_mWrite = ctl_mWrite | (pla[23]&pla[16])&(M2&T3);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[23]&pla[16])&(M2&T3);
ctl_reg_gp_sel_pla23pla16M2T3_5 = (pla[23]&pla[16])&(M2&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23pla16M2T3_5,ctl_reg_gp_sel_pla23pla16M2T3_5})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla23pla16M2T3_6 = (pla[23]&pla[16])&(M2&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23pla16M2T3_6,ctl_reg_gp_hilo_pla23pla16M2T3_6})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[23]&pla[16])&(M2&T3);
ctl_inc_cy = ctl_inc_cy | (pla[23]&pla[16])&(M2&T3)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[23]&pla[16])&(M2&T3);
ctl_al_we = ctl_al_we | (pla[23]&pla[16])&(M2&T3);
fMWrite = fMWrite | (pla[23]&pla[16])&(M3&T1);
ctl_inc_cy = ctl_inc_cy | (pla[23]&pla[16])&(M3&T1)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[23]&pla[16])&(M3&T1);
ctl_apin_mux = ctl_apin_mux | (pla[23]&pla[16])&(M3&T1);
ctl_reg_gp_sel_pla23pla16M3T1_5 = (pla[23]&pla[16])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23pla16M3T1_5,ctl_reg_gp_sel_pla23pla16M3T1_5})&(op54);
ctl_reg_gp_hilo_pla23pla16M3T1_6 = (pla[23]&pla[16])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23pla16M3T1_6,ctl_reg_gp_hilo_pla23pla16M3T1_6})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[23]&pla[16])&(M3&T1);
ctl_sw_1u = ctl_sw_1u | (pla[23]&pla[16])&(M3&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[23]&pla[16])&(M3&T1);
fMWrite = fMWrite | (pla[23]&pla[16])&(M3&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[23]&pla[16])&(M3&T2);
ctl_reg_gp_sel_pla23pla16M3T2_3 = (pla[23]&pla[16])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23pla16M3T2_3,ctl_reg_gp_sel_pla23pla16M3T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla23pla16M3T2_4 = (pla[23]&pla[16])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23pla16M3T2_4,ctl_reg_gp_hilo_pla23pla16M3T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[23]&pla[16])&(M3&T2);
ctl_sw_4u = ctl_sw_4u | (pla[23]&pla[16])&(M3&T2);
ctl_inc_cy = ctl_inc_cy | (pla[23]&pla[16])&(M3&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[23]&pla[16])&(M3&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[23]&pla[16])&(M3&T2);
fMWrite = fMWrite | (pla[23]&pla[16])&(M3&T3);
setM1 = setM1 | (pla[23]&pla[16])&(M3&T3);
validPLA = validPLA | (pla[23]&~pla[16])&(M1&T4);
nextM = nextM | (pla[23]&~pla[16])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[23]&~pla[16])&(M1&T4);
fMRead = fMRead | (pla[23]&~pla[16])&(M2&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[23]&~pla[16])&(M2&T1);
ctl_reg_gp_sel_pla23npla16M2T1_3 = (pla[23]&~pla[16])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23npla16M2T1_3,ctl_reg_gp_sel_pla23npla16M2T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla23npla16M2T1_4 = (pla[23]&~pla[16])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23npla16M2T1_4,ctl_reg_gp_hilo_pla23npla16M2T1_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[23]&~pla[16])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[23]&~pla[16])&(M2&T1);
fMRead = fMRead | (pla[23]&~pla[16])&(M2&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[23]&~pla[16])&(M2&T2);
ctl_reg_gp_sel_pla23npla16M2T2_3 = (pla[23]&~pla[16])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23npla16M2T2_3,ctl_reg_gp_sel_pla23npla16M2T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla23npla16M2T2_4 = (pla[23]&~pla[16])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23npla16M2T2_4,ctl_reg_gp_hilo_pla23npla16M2T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[23]&~pla[16])&(M2&T2);
ctl_sw_4u = ctl_sw_4u | (pla[23]&~pla[16])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[23]&~pla[16])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[23]&~pla[16])&(M2&T2);
fMRead = fMRead | (pla[23]&~pla[16])&(M2&T3);
nextM = nextM | (pla[23]&~pla[16])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[23]&~pla[16])&(M2&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[23]&~pla[16])&(M2&T3);
ctl_reg_gp_sel_pla23npla16M2T3_5 = (pla[23]&~pla[16])&(M2&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23npla16M2T3_5,ctl_reg_gp_sel_pla23npla16M2T3_5})&(op54);
ctl_reg_gp_hilo_pla23npla16M2T3_6 = (pla[23]&~pla[16])&(M2&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23npla16M2T3_6,ctl_reg_gp_hilo_pla23npla16M2T3_6})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[23]&~pla[16])&(M2&T3);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[23]&~pla[16])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[23]&~pla[16])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[23]&~pla[16])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[23]&~pla[16])&(M2&T3);
fMRead = fMRead | (pla[23]&~pla[16])&(M3&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[23]&~pla[16])&(M3&T1);
ctl_reg_gp_sel_pla23npla16M3T1_3 = (pla[23]&~pla[16])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23npla16M3T1_3,ctl_reg_gp_sel_pla23npla16M3T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla23npla16M3T1_4 = (pla[23]&~pla[16])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23npla16M3T1_4,ctl_reg_gp_hilo_pla23npla16M3T1_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[23]&~pla[16])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[23]&~pla[16])&(M3&T1);
fMRead = fMRead | (pla[23]&~pla[16])&(M3&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[23]&~pla[16])&(M3&T2);
ctl_reg_gp_sel_pla23npla16M3T2_3 = (pla[23]&~pla[16])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23npla16M3T2_3,ctl_reg_gp_sel_pla23npla16M3T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla23npla16M3T2_4 = (pla[23]&~pla[16])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23npla16M3T2_4,ctl_reg_gp_hilo_pla23npla16M3T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[23]&~pla[16])&(M3&T2);
ctl_sw_4u = ctl_sw_4u | (pla[23]&~pla[16])&(M3&T2);
ctl_inc_cy = ctl_inc_cy | (pla[23]&~pla[16])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[23]&~pla[16])&(M3&T2);
fMRead = fMRead | (pla[23]&~pla[16])&(M3&T3);
setM1 = setM1 | (pla[23]&~pla[16])&(M3&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[23]&~pla[16])&(M3&T3);
ctl_reg_gp_sel_pla23npla16M3T3_4 = (pla[23]&~pla[16])&(M3&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla23npla16M3T3_4,ctl_reg_gp_sel_pla23npla16M3T3_4})&(op54);
ctl_reg_gp_hilo_pla23npla16M3T3_5 = (pla[23]&~pla[16])&(M3&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla23npla16M3T3_5,ctl_reg_gp_hilo_pla23npla16M3T3_5})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[23]&~pla[16])&(M3&T3);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[23]&~pla[16])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[23]&~pla[16])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[23]&~pla[16])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[23]&~pla[16])&(M3&T3);
ctl_reg_ex_de_hl = ctl_reg_ex_de_hl | (pla[2])&(M1&T2);
validPLA = validPLA | (pla[2])&(M1&T4);
setM1 = setM1 | (pla[2])&(M1&T4);
ctl_reg_ex_af = ctl_reg_ex_af | (pla[39])&(M1&T2);
validPLA = validPLA | (pla[39])&(M1&T4);
setM1 = setM1 | (pla[39])&(M1&T4);
ctl_reg_exx = ctl_reg_exx | (pla[1])&(M1&T2);
validPLA = validPLA | (pla[1])&(M1&T4);
setM1 = setM1 | (pla[1])&(M1&T4);
validPLA = validPLA | (pla[10])&(M1&T4);
nextM = nextM | (pla[10])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[10])&(M1&T4);
fMRead = fMRead | (pla[10])&(M2&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[10])&(M2&T1);
ctl_reg_gp_sel_pla10M2T1_3 = (pla[10])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M2T1_3,ctl_reg_gp_sel_pla10M2T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla10M2T1_4 = (pla[10])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M2T1_4,ctl_reg_gp_hilo_pla10M2T1_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[10])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[10])&(M2&T1);
fMRead = fMRead | (pla[10])&(M2&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[10])&(M2&T2);
ctl_reg_gp_sel_pla10M2T2_3 = (pla[10])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M2T2_3,ctl_reg_gp_sel_pla10M2T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla10M2T2_4 = (pla[10])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M2T2_4,ctl_reg_gp_hilo_pla10M2T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[10])&(M2&T2);
ctl_sw_4u = ctl_sw_4u | (pla[10])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[10])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[10])&(M2&T2);
fMRead = fMRead | (pla[10])&(M2&T3);
nextM = nextM | (pla[10])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[10])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[10])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[10])&(M2&T3);
ctl_reg_sys_hilo_pla10M2T3_6 = (pla[10])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla10M2T3_6,ctl_reg_sys_hilo_pla10M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[10])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[10])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[10])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[10])&(M2&T3);
fMRead = fMRead | (pla[10])&(M3&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[10])&(M3&T1);
ctl_reg_gp_sel_pla10M3T1_3 = (pla[10])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M3T1_3,ctl_reg_gp_sel_pla10M3T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla10M3T1_4 = (pla[10])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M3T1_4,ctl_reg_gp_hilo_pla10M3T1_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[10])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[10])&(M3&T1);
fMRead = fMRead | (pla[10])&(M3&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[10])&(M3&T2);
ctl_reg_gp_sel_pla10M3T2_3 = (pla[10])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M3T2_3,ctl_reg_gp_sel_pla10M3T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla10M3T2_4 = (pla[10])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M3T2_4,ctl_reg_gp_hilo_pla10M3T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[10])&(M3&T2);
ctl_sw_4u = ctl_sw_4u | (pla[10])&(M3&T2);
ctl_inc_cy = ctl_inc_cy | (pla[10])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[10])&(M3&T2);
fMRead = fMRead | (pla[10])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[10])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[10])&(M3&T3);
ctl_reg_sys_hilo_pla10M3T3_4 = (pla[10])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla10M3T3_4,ctl_reg_sys_hilo_pla10M3T3_4})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[10])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[10])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[10])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[10])&(M3&T3);
nextM = nextM | (pla[10])&(M3&T4);
ctl_mWrite = ctl_mWrite | (pla[10])&(M3&T4);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[10])&(M3&T4);
ctl_reg_gp_sel_pla10M3T4_4 = (pla[10])&(M3&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M3T4_4,ctl_reg_gp_sel_pla10M3T4_4})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla10M3T4_5 = (pla[10])&(M3&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M3T4_5,ctl_reg_gp_hilo_pla10M3T4_5})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[10])&(M3&T4);
ctl_inc_cy = ctl_inc_cy | (pla[10])&(M3&T4)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[10])&(M3&T4);
ctl_al_we = ctl_al_we | (pla[10])&(M3&T4);
fMWrite = fMWrite | (pla[10])&(M4&T1);
ctl_inc_cy = ctl_inc_cy | (pla[10])&(M4&T1)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[10])&(M4&T1);
ctl_apin_mux = ctl_apin_mux | (pla[10])&(M4&T1);
ctl_reg_gp_sel_pla10M4T1_5 = (pla[10])&(M4&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M4T1_5,ctl_reg_gp_sel_pla10M4T1_5})&(op54);
ctl_reg_gp_hilo_pla10M4T1_6 = (pla[10])&(M4&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M4T1_6,ctl_reg_gp_hilo_pla10M4T1_6})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[10])&(M4&T1);
ctl_sw_2u = ctl_sw_2u | (pla[10])&(M4&T1);
ctl_sw_1u = ctl_sw_1u | (pla[10])&(M4&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[10])&(M4&T1);
fMWrite = fMWrite | (pla[10])&(M4&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[10])&(M4&T2);
ctl_reg_gp_sel_pla10M4T2_3 = (pla[10])&(M4&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M4T2_3,ctl_reg_gp_sel_pla10M4T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla10M4T2_4 = (pla[10])&(M4&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M4T2_4,ctl_reg_gp_hilo_pla10M4T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[10])&(M4&T2);
ctl_sw_4u = ctl_sw_4u | (pla[10])&(M4&T2);
ctl_inc_cy = ctl_inc_cy | (pla[10])&(M4&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[10])&(M4&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[10])&(M4&T2);
fMWrite = fMWrite | (pla[10])&(M4&T3);
nextM = nextM | (pla[10])&(M4&T3);
ctl_mWrite = ctl_mWrite | (pla[10])&(M4&T3);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[10])&(M4&T3);
ctl_reg_gp_sel_pla10M4T3_5 = (pla[10])&(M4&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M4T3_5,ctl_reg_gp_sel_pla10M4T3_5})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla10M4T3_6 = (pla[10])&(M4&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M4T3_6,ctl_reg_gp_hilo_pla10M4T3_6})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[10])&(M4&T3);
ctl_inc_cy = ctl_inc_cy | (pla[10])&(M4&T3)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[10])&(M4&T3);
ctl_al_we = ctl_al_we | (pla[10])&(M4&T3);
fMWrite = fMWrite | (pla[10])&(M5&T1);
ctl_inc_cy = ctl_inc_cy | (pla[10])&(M5&T1)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[10])&(M5&T1);
ctl_apin_mux = ctl_apin_mux | (pla[10])&(M5&T1);
ctl_reg_gp_sel_pla10M5T1_5 = (pla[10])&(M5&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M5T1_5,ctl_reg_gp_sel_pla10M5T1_5})&(op54);
ctl_reg_gp_hilo_pla10M5T1_6 = (pla[10])&(M5&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M5T1_6,ctl_reg_gp_hilo_pla10M5T1_6})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[10])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (pla[10])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[10])&(M5&T1);
fMWrite = fMWrite | (pla[10])&(M5&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[10])&(M5&T2);
ctl_reg_gp_sel_pla10M5T2_3 = (pla[10])&(M5&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M5T2_3,ctl_reg_gp_sel_pla10M5T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla10M5T2_4 = (pla[10])&(M5&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M5T2_4,ctl_reg_gp_hilo_pla10M5T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[10])&(M5&T2);
ctl_sw_4u = ctl_sw_4u | (pla[10])&(M5&T2);
ctl_inc_cy = ctl_inc_cy | (pla[10])&(M5&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[10])&(M5&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[10])&(M5&T2);
fMWrite = fMWrite | (pla[10])&(M5&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[10])&(M5&T3);
ctl_reg_sys_hilo_pla10M5T3_3 = (pla[10])&(M5&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla10M5T3_3,ctl_reg_sys_hilo_pla10M5T3_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[10])&(M5&T3);
ctl_al_we = ctl_al_we | (pla[10])&(M5&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[10])&(M5&T4);
ctl_reg_gp_sel_pla10M5T4_2 = (pla[10])&(M5&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla10M5T4_2,ctl_reg_gp_sel_pla10M5T4_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla10M5T4_3 = (pla[10])&(M5&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla10M5T4_3,ctl_reg_gp_hilo_pla10M5T4_3})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[10])&(M5&T4);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[10])&(M5&T4);
setM1 = setM1 | (pla[10])&(M5&T5);
nonRep = nonRep | (pla[0]);
ctl_flags_alu = ctl_flags_alu | (pla[12])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[12])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[12])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[12])&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (pla[12])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (pla[12])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[12])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[12])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[12])&(M1&T1);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[12])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[12])&(M1&T1);
ctl_pf_sel_pla12M1T1_12 = (pla[12])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla12M1T1_12,ctl_pf_sel_pla12M1T1_12})&(`PFSEL_REP);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[12])&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[12])&(M1&T1);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (pla[12])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[12])&(M1&T2);
ctl_reg_gp_sel_pla12M1T2_2 = (pla[12])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla12M1T2_2,ctl_reg_gp_sel_pla12M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla12M1T2_3 = (pla[12])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla12M1T2_3,ctl_reg_gp_hilo_pla12M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[12])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[12])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[12])&(M1&T2);
ctl_reg_gp_sel_pla12M1T3_1 = (pla[12])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla12M1T3_1,ctl_reg_gp_sel_pla12M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla12M1T3_2 = (pla[12])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla12M1T3_2,ctl_reg_gp_hilo_pla12M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[12])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[12])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[12])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[12])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[12])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[12])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[12])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[12])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[12])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[12])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[12])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[12])&(M1&T3);
validPLA = validPLA | (pla[12])&(M1&T4);
nextM = nextM | (pla[12])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[12])&(M1&T4);
fMRead = fMRead | (pla[12])&(M2&T1);
ctl_reg_gp_sel_pla12M2T1_2 = (pla[12])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla12M2T1_2,ctl_reg_gp_sel_pla12M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla12M2T1_3 = (pla[12])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla12M2T1_3,ctl_reg_gp_hilo_pla12M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[12])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[12])&(M2&T1);
fMRead = fMRead | (pla[12])&(M2&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[12])&(M2&T2);
ctl_reg_gp_sel_pla12M2T2_3 = (pla[12])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla12M2T2_3,ctl_reg_gp_sel_pla12M2T2_3})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla12M2T2_4 = (pla[12])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla12M2T2_4,ctl_reg_gp_hilo_pla12M2T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[12])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[12])&(M2&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[12])&(M2&T2)&(op3);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[12])&(M2&T2);
fMRead = fMRead | (pla[12])&(M2&T3);
nextM = nextM | (pla[12])&(M2&T3);
ctl_mWrite = ctl_mWrite | (pla[12])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[12])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[12])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[12])&(M2&T3);
ctl_flags_alu = ctl_flags_alu | (pla[12])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[12])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[12])&(M2&T3);
ctl_alu_op_low = ctl_alu_op_low | (pla[12])&(M2&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[12])&(M2&T3)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[12])&(M2&T3)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[12])&(M2&T3)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[12])&(M2&T3);
ctl_flags_cf2_we = ctl_flags_cf2_we | (pla[12])&(M2&T3);
fMWrite = fMWrite | (pla[12])&(M3&T1);
ctl_reg_gp_sel_pla12M3T1_2 = (pla[12])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla12M3T1_2,ctl_reg_gp_sel_pla12M3T1_2})&(`GP_REG_DE);
ctl_reg_gp_hilo_pla12M3T1_3 = (pla[12])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla12M3T1_3,ctl_reg_gp_hilo_pla12M3T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[12])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[12])&(M3&T1);
ctl_flags_alu = ctl_flags_alu | (pla[12])&(M3&T1);
ctl_alu_oe = ctl_alu_oe | (pla[12])&(M3&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[12])&(M3&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[12])&(M3&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[12])&(M3&T1)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[12])&(M3&T1)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[12])&(M3&T1)&(~ctl_alu_op_low);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (pla[12])&(M3&T1);
fMWrite = fMWrite | (pla[12])&(M3&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[12])&(M3&T2);
ctl_reg_gp_sel_pla12M3T2_3 = (pla[12])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla12M3T2_3,ctl_reg_gp_sel_pla12M3T2_3})&(`GP_REG_DE);
ctl_reg_gp_hilo_pla12M3T2_4 = (pla[12])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla12M3T2_4,ctl_reg_gp_hilo_pla12M3T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[12])&(M3&T2);
ctl_inc_cy = ctl_inc_cy | (pla[12])&(M3&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[12])&(M3&T2)&(op3);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[12])&(M3&T2);
fMWrite = fMWrite | (pla[12])&(M3&T3);
ctl_reg_gp_sel_pla12M3T3_2 = (pla[12])&(M3&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla12M3T3_2,ctl_reg_gp_sel_pla12M3T3_2})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla12M3T3_3 = (pla[12])&(M3&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla12M3T3_3,ctl_reg_gp_hilo_pla12M3T3_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[12])&(M3&T3);
ctl_al_we = ctl_al_we | (pla[12])&(M3&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[12])&(M3&T4);
ctl_reg_gp_sel_pla12M3T4_2 = (pla[12])&(M3&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla12M3T4_2,ctl_reg_gp_sel_pla12M3T4_2})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla12M3T4_3 = (pla[12])&(M3&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla12M3T4_3,ctl_reg_gp_hilo_pla12M3T4_3})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[12])&(M3&T4);
ctl_inc_cy = ctl_inc_cy | (pla[12])&(M3&T4)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[12])&(M3&T4);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[12])&(M3&T4);
ctl_repeat_we = ctl_repeat_we | (pla[12])&(M3&T4);
nextM = nextM | (pla[12])&(M3&T5);
setM1 = setM1 | (pla[12])&(M3&T5)&(nonRep|~repeat_en);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[12])&(M4&T1);
ctl_reg_sys_hilo_pla12M4T1_2 = (pla[12])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla12M4T1_2,ctl_reg_sys_hilo_pla12M4T1_2})&(2'b11);
ctl_al_we = ctl_al_we | (pla[12])&(M4&T1);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[12])&(M4&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[12])&(M4&T2);
ctl_reg_sys_hilo_pla12M4T2_3 = (pla[12])&(M4&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla12M4T2_3,ctl_reg_sys_hilo_pla12M4T2_3})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[12])&(M4&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[12])&(M4&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[12])&(M4&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[12])&(M4&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[12])&(M4&T3);
ctl_reg_sys_hilo_pla12M4T3_2 = (pla[12])&(M4&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla12M4T3_2,ctl_reg_sys_hilo_pla12M4T3_2})&(2'b11);
ctl_al_we = ctl_al_we | (pla[12])&(M4&T3);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[12])&(M4&T4);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[12])&(M4&T4);
ctl_reg_sys_hilo_pla12M4T4_3 = (pla[12])&(M4&T4);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla12M4T4_3,ctl_reg_sys_hilo_pla12M4T4_3})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[12])&(M4&T4)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[12])&(M4&T4)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[12])&(M4&T4);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[12])&(M4&T4);
setM1 = setM1 | (pla[12])&(M4&T5);
ctl_flags_alu = ctl_flags_alu | (pla[11])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[11])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[11])&(M1&T1);
ctl_alu_op1_sel_zero = ctl_alu_op1_sel_zero | (pla[11])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[11])&(M1&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[11])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[11])&(M1&T1)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[11])&(M1&T1)&(~ctl_alu_op_low);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[11])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[11])&(M1&T1);
ctl_pf_sel_pla11M1T1_11 = (pla[11])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla11M1T1_11,ctl_pf_sel_pla11M1T1_11})&(`PFSEL_REP);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[11])&(M1&T1);
ctl_flags_nf_set = ctl_flags_nf_set | (pla[11])&(M1&T1);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (pla[11])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[11])&(M1&T2);
ctl_reg_gp_sel_pla11M1T2_2 = (pla[11])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla11M1T2_2,ctl_reg_gp_sel_pla11M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla11M1T2_3 = (pla[11])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla11M1T2_3,ctl_reg_gp_hilo_pla11M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[11])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[11])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[11])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (pla[11])&(M1&T2)&(flags_nf);
ctl_reg_gp_sel_pla11M1T3_1 = (pla[11])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla11M1T3_1,ctl_reg_gp_sel_pla11M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla11M1T3_2 = (pla[11])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla11M1T3_2,ctl_reg_gp_hilo_pla11M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[11])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[11])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[11])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[11])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[11])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[11])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[11])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[11])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[11])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[11])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[11])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[11])&(M1&T3);
validPLA = validPLA | (pla[11])&(M1&T4);
nextM = nextM | (pla[11])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[11])&(M1&T4);
fMRead = fMRead | (pla[11])&(M2&T1);
ctl_reg_gp_sel_pla11M2T1_2 = (pla[11])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla11M2T1_2,ctl_reg_gp_sel_pla11M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla11M2T1_3 = (pla[11])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla11M2T1_3,ctl_reg_gp_hilo_pla11M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[11])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[11])&(M2&T1);
fMRead = fMRead | (pla[11])&(M2&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[11])&(M2&T2);
ctl_reg_gp_sel_pla11M2T2_3 = (pla[11])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla11M2T2_3,ctl_reg_gp_sel_pla11M2T2_3})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla11M2T2_4 = (pla[11])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla11M2T2_4,ctl_reg_gp_hilo_pla11M2T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[11])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[11])&(M2&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[11])&(M2&T2)&(op3);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[11])&(M2&T2);
fMRead = fMRead | (pla[11])&(M2&T3);
nextM = nextM | (pla[11])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[11])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[11])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[11])&(M2&T3);
ctl_flags_alu = ctl_flags_alu | (pla[11])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[11])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[11])&(M2&T3);
ctl_alu_op_low = ctl_alu_op_low | (pla[11])&(M2&T3);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[11])&(M2&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[11])&(M2&T3)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[11])&(M2&T3)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[11])&(M2&T3);
ctl_flags_cf2_we = ctl_flags_cf2_we | (pla[11])&(M2&T3);
ctl_flags_alu = ctl_flags_alu | (pla[11])&(M3&T1);
ctl_alu_oe = ctl_alu_oe | (pla[11])&(M3&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[11])&(M3&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[11])&(M3&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[11])&(M3&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[11])&(M3&T1)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[11])&(M3&T1)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[11])&(M3&T1);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (pla[11])&(M3&T1);
ctl_reg_gp_sel_pla11M3T3_1 = (pla[11])&(M3&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla11M3T3_1,ctl_reg_gp_sel_pla11M3T3_1})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla11M3T3_2 = (pla[11])&(M3&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla11M3T3_2,ctl_reg_gp_hilo_pla11M3T3_2})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[11])&(M3&T3);
ctl_al_we = ctl_al_we | (pla[11])&(M3&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[11])&(M3&T4);
ctl_reg_gp_sel_pla11M3T4_2 = (pla[11])&(M3&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla11M3T4_2,ctl_reg_gp_sel_pla11M3T4_2})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla11M3T4_3 = (pla[11])&(M3&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla11M3T4_3,ctl_reg_gp_hilo_pla11M3T4_3})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[11])&(M3&T4);
ctl_inc_cy = ctl_inc_cy | (pla[11])&(M3&T4)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[11])&(M3&T4);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[11])&(M3&T4);
ctl_repeat_we = ctl_repeat_we | (pla[11])&(M3&T4);
nextM = nextM | (pla[11])&(M3&T5);
setM1 = setM1 | (pla[11])&(M3&T5)&(nonRep|~repeat_en|flags_zf);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[11])&(M4&T1);
ctl_reg_sys_hilo_pla11M4T1_2 = (pla[11])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla11M4T1_2,ctl_reg_sys_hilo_pla11M4T1_2})&(2'b11);
ctl_al_we = ctl_al_we | (pla[11])&(M4&T1);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[11])&(M4&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[11])&(M4&T2);
ctl_reg_sys_hilo_pla11M4T2_3 = (pla[11])&(M4&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla11M4T2_3,ctl_reg_sys_hilo_pla11M4T2_3})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[11])&(M4&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[11])&(M4&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[11])&(M4&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[11])&(M4&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[11])&(M4&T3);
ctl_reg_sys_hilo_pla11M4T3_2 = (pla[11])&(M4&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla11M4T3_2,ctl_reg_sys_hilo_pla11M4T3_2})&(2'b11);
ctl_al_we = ctl_al_we | (pla[11])&(M4&T3);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[11])&(M4&T4);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[11])&(M4&T4);
ctl_reg_sys_hilo_pla11M4T4_3 = (pla[11])&(M4&T4);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla11M4T4_3,ctl_reg_sys_hilo_pla11M4T4_3})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[11])&(M4&T4)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[11])&(M4&T4)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[11])&(M4&T4);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[11])&(M4&T4);
setM1 = setM1 | (pla[11])&(M4&T5);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[65]&~pla[52])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[65]&~pla[52])&(M1&T1);
ctl_sw_2u = ctl_sw_2u | (pla[65]&~pla[52])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[65]&~pla[52])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[65]&~pla[52])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[65]&~pla[52])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[65]&~pla[52])&(M1&T1);
ctl_state_alu = ctl_state_alu | (pla[65]&~pla[52])&(M1&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[65]&~pla[52])&(M1&T1);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[65]&~pla[52])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[65]&~pla[52])&(M1&T2);
ctl_reg_gp_sel_pla65npla52M1T2_2 = (pla[65]&~pla[52])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla65npla52M1T2_2,ctl_reg_gp_sel_pla65npla52M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla65npla52M1T2_3 = (pla[65]&~pla[52])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla65npla52M1T2_3,ctl_reg_gp_hilo_pla65npla52M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[65]&~pla[52])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[65]&~pla[52])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[65]&~pla[52])&(M1&T2);
ctl_state_alu = ctl_state_alu | (pla[65]&~pla[52])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (pla[65]&~pla[52])&(M1&T2)&(flags_nf);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[65]&~pla[52])&(M1&T2)&(flags_nf);
ctl_reg_gp_sel_pla65npla52M1T3_1 = (pla[65]&~pla[52])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla65npla52M1T3_1,ctl_reg_gp_sel_pla65npla52M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla65npla52M1T3_2 = (pla[65]&~pla[52])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla65npla52M1T3_2,ctl_reg_gp_hilo_pla65npla52M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[65]&~pla[52])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[65]&~pla[52])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[65]&~pla[52])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[65]&~pla[52])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[65]&~pla[52])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[65]&~pla[52])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[65]&~pla[52])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[65]&~pla[52])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[65]&~pla[52])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[65]&~pla[52])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[65]&~pla[52])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[65]&~pla[52])&(M1&T3);
validPLA = validPLA | (pla[65]&~pla[52])&(M1&T4);
setM1 = setM1 | (pla[65]&~pla[52])&(M1&T4);
ctl_reg_gp_sel_pla65npla52M1T4_3 = (pla[65]&~pla[52])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla65npla52M1T4_3,ctl_reg_gp_sel_pla65npla52M1T4_3})&(op21);
ctl_reg_gp_hilo_pla65npla52M1T4_4 = (pla[65]&~pla[52])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla65npla52M1T4_4,ctl_reg_gp_hilo_pla65npla52M1T4_4})&({~rsel0,rsel0});
ctl_reg_out_hi = ctl_reg_out_hi | (pla[65]&~pla[52])&(M1&T4)&(~rsel0);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[65]&~pla[52])&(M1&T4)&(rsel0);
ctl_sw_2u = ctl_sw_2u | (pla[65]&~pla[52])&(M1&T4)&(~rsel0);
ctl_sw_2d = ctl_sw_2d | (pla[65]&~pla[52])&(M1&T4)&(rsel0);
ctl_flags_alu = ctl_flags_alu | (pla[65]&~pla[52])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[65]&~pla[52])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[65]&~pla[52])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[65]&~pla[52])&(M1&T4);
ctl_state_alu = ctl_state_alu | (pla[65]&~pla[52])&(M1&T4);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[65]&~pla[52])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[65]&~pla[52])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[65]&~pla[52])&(M1&T4);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[64])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[64])&(M1&T1);
ctl_sw_2u = ctl_sw_2u | (pla[64])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[64])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[64])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[64])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[64])&(M1&T1);
ctl_state_alu = ctl_state_alu | (pla[64])&(M1&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[64])&(M1&T1);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[64])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[64])&(M1&T2);
ctl_reg_gp_sel_pla64M1T2_2 = (pla[64])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla64M1T2_2,ctl_reg_gp_sel_pla64M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla64M1T2_3 = (pla[64])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla64M1T2_3,ctl_reg_gp_hilo_pla64M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[64])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[64])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[64])&(M1&T2);
ctl_state_alu = ctl_state_alu | (pla[64])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (pla[64])&(M1&T2)&(flags_nf);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[64])&(M1&T2)&(flags_nf);
ctl_reg_gp_sel_pla64M1T3_1 = (pla[64])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla64M1T3_1,ctl_reg_gp_sel_pla64M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla64M1T3_2 = (pla[64])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla64M1T3_2,ctl_reg_gp_hilo_pla64M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[64])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[64])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[64])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[64])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[64])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[64])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[64])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[64])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[64])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[64])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[64])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[64])&(M1&T3);
validPLA = validPLA | (pla[64])&(M1&T4);
nextM = nextM | (pla[64])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[64])&(M1&T4);
ctl_reg_gp_sel_pla64M1T4_4 = (pla[64])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla64M1T4_4,ctl_reg_gp_sel_pla64M1T4_4})&(op21);
ctl_reg_gp_hilo_pla64M1T4_5 = (pla[64])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla64M1T4_5,ctl_reg_gp_hilo_pla64M1T4_5})&({~rsel0,rsel0});
ctl_reg_out_hi = ctl_reg_out_hi | (pla[64])&(M1&T4)&(~rsel0);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[64])&(M1&T4)&(rsel0);
ctl_sw_2u = ctl_sw_2u | (pla[64])&(M1&T4)&(~rsel0);
ctl_sw_2d = ctl_sw_2d | (pla[64])&(M1&T4)&(rsel0);
ctl_flags_alu = ctl_flags_alu | (pla[64])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[64])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[64])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[64])&(M1&T4);
ctl_state_alu = ctl_state_alu | (pla[64])&(M1&T4);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[64])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[64])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[64])&(M1&T4);
fMRead = fMRead | (pla[64])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[64])&(M2&T1);
ctl_reg_sys_hilo_pla64M2T1_3 = (pla[64])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla64M2T1_3,ctl_reg_sys_hilo_pla64M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[64])&(M2&T1);
ctl_state_alu = ctl_state_alu | (pla[64])&(M2&T1);
fMRead = fMRead | (pla[64])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[64])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[64])&(M2&T2);
ctl_reg_sys_hilo_pla64M2T2_4 = (pla[64])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla64M2T2_4,ctl_reg_sys_hilo_pla64M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[64])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[64])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[64])&(M2&T2);
fMRead = fMRead | (pla[64])&(M2&T3);
setM1 = setM1 | (pla[64])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[64])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[64])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[64])&(M2&T3);
ctl_flags_alu = ctl_flags_alu | (pla[64])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[64])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[64])&(M2&T3);
ctl_alu_op_low = ctl_alu_op_low | (pla[64])&(M2&T3);
ctl_state_alu = ctl_state_alu | (pla[64])&(M2&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[64])&(M2&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[64])&(M2&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[64])&(M2&T3);
ctl_reg_gp_sel_use_ixiypla52M1T3_1 = (use_ixiy&pla[52])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_use_ixiypla52M1T3_1,ctl_reg_gp_sel_use_ixiypla52M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_use_ixiypla52M1T3_2 = (use_ixiy&pla[52])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_use_ixiypla52M1T3_2,ctl_reg_gp_hilo_use_ixiypla52M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (use_ixiy&pla[52])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (use_ixiy&pla[52])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (use_ixiy&pla[52])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (use_ixiy&pla[52])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (use_ixiy&pla[52])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (use_ixiy&pla[52])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (use_ixiy&pla[52])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (use_ixiy&pla[52])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (use_ixiy&pla[52])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (use_ixiy&pla[52])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (use_ixiy&pla[52])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (use_ixiy&pla[52])&(M1&T3);
validPLA = validPLA | (use_ixiy&pla[52])&(M1&T4);
nextM = nextM | (use_ixiy&pla[52])&(M1&T4);
ctl_mRead = ctl_mRead | (use_ixiy&pla[52])&(M1&T4);
fMRead = fMRead | (use_ixiy&pla[52])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (use_ixiy&pla[52])&(M2&T1);
ctl_reg_sys_hilo_use_ixiypla52M2T1_3 = (use_ixiy&pla[52])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_use_ixiypla52M2T1_3,ctl_reg_sys_hilo_use_ixiypla52M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (use_ixiy&pla[52])&(M2&T1);
fMRead = fMRead | (use_ixiy&pla[52])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (use_ixiy&pla[52])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (use_ixiy&pla[52])&(M2&T2);
ctl_reg_sys_hilo_use_ixiypla52M2T2_4 = (use_ixiy&pla[52])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_use_ixiypla52M2T2_4,ctl_reg_sys_hilo_use_ixiypla52M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (use_ixiy&pla[52])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (use_ixiy&pla[52])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (use_ixiy&pla[52])&(M2&T2);
fMRead = fMRead | (use_ixiy&pla[52])&(M2&T3);
nextM = nextM | (use_ixiy&pla[52])&(M2&T3);
ixy_d = ixy_d | (use_ixiy&pla[52])&(M3&T1);
ixy_d = ixy_d | (use_ixiy&pla[52])&(M3&T2);
ixy_d = ixy_d | (use_ixiy&pla[52])&(M3&T3);
ixy_d = ixy_d | (use_ixiy&pla[52])&(M3&T4);
nextM = nextM | (use_ixiy&pla[52])&(M3&T5);
ctl_mRead = ctl_mRead | (use_ixiy&pla[52])&(M3&T5);
ixy_d = ixy_d | (use_ixiy&pla[52])&(M3&T5);
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[52])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[52])&(M1&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[52])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[52])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[52])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[52])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[52])&(M1&T1);
ctl_state_alu = ctl_state_alu | (~use_ixiy&pla[52])&(M1&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[52])&(M1&T1);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[52])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (~use_ixiy&pla[52])&(M1&T2);
ctl_reg_gp_sel_nuse_ixiypla52M1T2_2 = (~use_ixiy&pla[52])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla52M1T2_2,ctl_reg_gp_sel_nuse_ixiypla52M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla52M1T2_3 = (~use_ixiy&pla[52])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla52M1T2_3,ctl_reg_gp_hilo_nuse_ixiypla52M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[52])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[52])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (~use_ixiy&pla[52])&(M1&T2);
ctl_state_alu = ctl_state_alu | (~use_ixiy&pla[52])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (~use_ixiy&pla[52])&(M1&T2)&(flags_nf);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[52])&(M1&T2)&(flags_nf);
ctl_reg_gp_sel_nuse_ixiypla52M1T3_1 = (~use_ixiy&pla[52])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla52M1T3_1,ctl_reg_gp_sel_nuse_ixiypla52M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla52M1T3_2 = (~use_ixiy&pla[52])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla52M1T3_2,ctl_reg_gp_hilo_nuse_ixiypla52M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[52])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[52])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[52])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[52])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[52])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[52])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[52])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[52])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[52])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[52])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[52])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[52])&(M1&T3);
validPLA = validPLA | (~use_ixiy&pla[52])&(M1&T4);
nextM = nextM | (~use_ixiy&pla[52])&(M1&T4);
ctl_mRead = ctl_mRead | (~use_ixiy&pla[52])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[52])&(M2&T1);
ctl_reg_gp_sel_nuse_ixiypla52M2T1_2 = (~use_ixiy&pla[52])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla52M2T1_2,ctl_reg_gp_sel_nuse_ixiypla52M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_nuse_ixiypla52M2T1_3 = (~use_ixiy&pla[52])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla52M2T1_3,ctl_reg_gp_hilo_nuse_ixiypla52M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[52])&(M2&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[52])&(M2&T1);
fMRead = fMRead | (~use_ixiy&pla[52])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (~use_ixiy&pla[52])&(M2&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~use_ixiy&pla[52])&(M2&T2);
ctl_reg_sys_hilo_nuse_ixiypla52M2T2_4 = (~use_ixiy&pla[52])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nuse_ixiypla52M2T2_4,ctl_reg_sys_hilo_nuse_ixiypla52M2T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (~use_ixiy&pla[52])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (~use_ixiy&pla[52])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[52])&(M2&T2);
fMRead = fMRead | (~use_ixiy&pla[52])&(M2&T3);
setM1 = setM1 | (~use_ixiy&pla[52])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[52])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[52])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[52])&(M2&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[52])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[52])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[52])&(M2&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[52])&(M2&T3);
ctl_state_alu = ctl_state_alu | (~use_ixiy&pla[52])&(M2&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[52])&(M2&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[52])&(M2&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[52])&(M2&T3);
fMRead = fMRead | (~use_ixiy&pla[52])&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[52])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[52])&(M4&T2);
ctl_reg_gp_sel_nuse_ixiypla52M4T2_2 = (~use_ixiy&pla[52])&(M4&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla52M4T2_2,ctl_reg_gp_sel_nuse_ixiypla52M4T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla52M4T2_3 = (~use_ixiy&pla[52])&(M4&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla52M4T2_3,ctl_reg_gp_hilo_nuse_ixiypla52M4T2_3})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[52])&(M4&T2);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[52])&(M4&T2);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[52])&(M4&T2);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[52])&(M4&T2)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[52])&(M4&T2);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[52])&(M4&T2);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[52])&(M4&T2);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[52])&(M4&T2);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[52])&(M4&T2);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[52])&(M4&T2);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[52])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[52])&(M4&T3);
setM1 = setM1 | (~use_ixiy&pla[52])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[52])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[52])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[52])&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[52])&(M4&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[52])&(M4&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[52])&(M4&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[52])&(M4&T3);
ctl_state_alu = ctl_state_alu | (~use_ixiy&pla[52])&(M4&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[52])&(M4&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[52])&(M4&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[52])&(M4&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[66]&~pla[53])&(M1&T1);
ctl_reg_gp_sel_pla66npla53M1T1_2 = (pla[66]&~pla[53])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla66npla53M1T1_2,ctl_reg_gp_sel_pla66npla53M1T1_2})&(op54);
ctl_reg_gp_hilo_pla66npla53M1T1_3 = (pla[66]&~pla[53])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla66npla53M1T1_3,ctl_reg_gp_hilo_pla66npla53M1T1_3})&({~rsel3,rsel3});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[66]&~pla[53])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[66]&~pla[53])&(M1&T1);
ctl_sw_2u = ctl_sw_2u | (pla[66]&~pla[53])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[66]&~pla[53])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[66]&~pla[53])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[66]&~pla[53])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[66]&~pla[53])&(M1&T1);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[66]&~pla[53])&(M1&T1)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[66]&~pla[53])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[66]&~pla[53])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[66]&~pla[53])&(M1&T1);
ctl_pf_sel_pla66npla53M1T1_15 = (pla[66]&~pla[53])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla66npla53M1T1_15,ctl_pf_sel_pla66npla53M1T1_15})&(`PFSEL_V);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (pla[66]&~pla[53])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[66]&~pla[53])&(M1&T2);
ctl_reg_gp_sel_pla66npla53M1T2_2 = (pla[66]&~pla[53])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla66npla53M1T2_2,ctl_reg_gp_sel_pla66npla53M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla66npla53M1T2_3 = (pla[66]&~pla[53])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla66npla53M1T2_3,ctl_reg_gp_hilo_pla66npla53M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[66]&~pla[53])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[66]&~pla[53])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[66]&~pla[53])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (pla[66]&~pla[53])&(M1&T2)&(flags_nf);
ctl_reg_gp_sel_pla66npla53M1T3_1 = (pla[66]&~pla[53])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla66npla53M1T3_1,ctl_reg_gp_sel_pla66npla53M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla66npla53M1T3_2 = (pla[66]&~pla[53])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla66npla53M1T3_2,ctl_reg_gp_hilo_pla66npla53M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[66]&~pla[53])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[66]&~pla[53])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[66]&~pla[53])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[66]&~pla[53])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[66]&~pla[53])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[66]&~pla[53])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[66]&~pla[53])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[66]&~pla[53])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[66]&~pla[53])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[66]&~pla[53])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[66]&~pla[53])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[66]&~pla[53])&(M1&T3);
validPLA = validPLA | (pla[66]&~pla[53])&(M1&T4);
setM1 = setM1 | (pla[66]&~pla[53])&(M1&T4);
ctl_bus_zero_oe = ctl_bus_zero_oe | (pla[66]&~pla[53])&(M1&T4)&(op4&op5&~op3);
ctl_reg_gp_sel_pla66npla53M1T4nop4op5nop3_1 = (pla[66]&~pla[53])&(M1&T4)&(~(op4&op5&~op3));
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla66npla53M1T4nop4op5nop3_1,ctl_reg_gp_sel_pla66npla53M1T4nop4op5nop3_1})&(op54);
ctl_reg_gp_hilo_pla66npla53M1T4nop4op5nop3_2 = (pla[66]&~pla[53])&(M1&T4)&(~(op4&op5&~op3));
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla66npla53M1T4nop4op5nop3_2,ctl_reg_gp_hilo_pla66npla53M1T4nop4op5nop3_2})&({~rsel3,rsel3});
ctl_reg_out_hi = ctl_reg_out_hi | (pla[66]&~pla[53])&(M1&T4)&(~rsel3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[66]&~pla[53])&(M1&T4)&(rsel3);
ctl_sw_2u = ctl_sw_2u | (pla[66]&~pla[53])&(M1&T4)&(~rsel3);
ctl_sw_2d = ctl_sw_2d | (pla[66]&~pla[53])&(M1&T4)&(rsel3);
ctl_flags_alu = ctl_flags_alu | (pla[66]&~pla[53])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[66]&~pla[53])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_zero = ctl_alu_op2_sel_zero | (pla[66]&~pla[53])&(M1&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[66]&~pla[53])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[66]&~pla[53])&(M1&T4);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[66]&~pla[53])&(M1&T4)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[66]&~pla[53])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[66]&~pla[53])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[66]&~pla[53])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[66]&~pla[53])&(M1&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[66]&~pla[53])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[66]&~pla[53])&(M1&T4);
ctl_flags_cf2_we = ctl_flags_cf2_we | (pla[66]&~pla[53])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[75])&(M1&T1);
ctl_flags_nf_set = ctl_flags_nf_set | (pla[75])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[75])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[75])&(M1&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[75])&(M1&T1);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[75])&(M1&T4);
ctl_flags_nf_set = ctl_flags_nf_set | (pla[75])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[75])&(M1&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[75])&(M1&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[75])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | ((M2|M4)&pla[75]);
ctl_flags_nf_set = ctl_flags_nf_set | ((M2|M4)&pla[75]);
ctl_flags_cf_set = ctl_flags_cf_set | ((M2|M4)&pla[75]);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | ((M2|M4)&pla[75]);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | ((M2|M4)&pla[75]);
ctl_reg_gp_sel_use_ixiypla53M1T3_1 = (use_ixiy&pla[53])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_use_ixiypla53M1T3_1,ctl_reg_gp_sel_use_ixiypla53M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_use_ixiypla53M1T3_2 = (use_ixiy&pla[53])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_use_ixiypla53M1T3_2,ctl_reg_gp_hilo_use_ixiypla53M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (use_ixiy&pla[53])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (use_ixiy&pla[53])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (use_ixiy&pla[53])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (use_ixiy&pla[53])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (use_ixiy&pla[53])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (use_ixiy&pla[53])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (use_ixiy&pla[53])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (use_ixiy&pla[53])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (use_ixiy&pla[53])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (use_ixiy&pla[53])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (use_ixiy&pla[53])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (use_ixiy&pla[53])&(M1&T3);
validPLA = validPLA | (use_ixiy&pla[53])&(M1&T4);
nextM = nextM | (use_ixiy&pla[53])&(M1&T4);
ctl_mRead = ctl_mRead | (use_ixiy&pla[53])&(M1&T4);
fMRead = fMRead | (use_ixiy&pla[53])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (use_ixiy&pla[53])&(M2&T1);
ctl_reg_sys_hilo_use_ixiypla53M2T1_3 = (use_ixiy&pla[53])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_use_ixiypla53M2T1_3,ctl_reg_sys_hilo_use_ixiypla53M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (use_ixiy&pla[53])&(M2&T1);
fMRead = fMRead | (use_ixiy&pla[53])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (use_ixiy&pla[53])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (use_ixiy&pla[53])&(M2&T2);
ctl_reg_sys_hilo_use_ixiypla53M2T2_4 = (use_ixiy&pla[53])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_use_ixiypla53M2T2_4,ctl_reg_sys_hilo_use_ixiypla53M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (use_ixiy&pla[53])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (use_ixiy&pla[53])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (use_ixiy&pla[53])&(M2&T2);
fMRead = fMRead | (use_ixiy&pla[53])&(M2&T3);
nextM = nextM | (use_ixiy&pla[53])&(M2&T3);
ixy_d = ixy_d | (use_ixiy&pla[53])&(M3&T1);
ixy_d = ixy_d | (use_ixiy&pla[53])&(M3&T2);
ixy_d = ixy_d | (use_ixiy&pla[53])&(M3&T3);
ixy_d = ixy_d | (use_ixiy&pla[53])&(M3&T4);
nextM = nextM | (use_ixiy&pla[53])&(M3&T5);
ctl_mRead = ctl_mRead | (use_ixiy&pla[53])&(M3&T5);
ixy_d = ixy_d | (use_ixiy&pla[53])&(M3&T5);
ctl_reg_gp_we = ctl_reg_gp_we | (~use_ixiy&pla[53])&(M1&T2);
ctl_reg_gp_sel_nuse_ixiypla53M1T2_2 = (~use_ixiy&pla[53])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla53M1T2_2,ctl_reg_gp_sel_nuse_ixiypla53M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla53M1T2_3 = (~use_ixiy&pla[53])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla53M1T2_3,ctl_reg_gp_hilo_nuse_ixiypla53M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[53])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[53])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (~use_ixiy&pla[53])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (~use_ixiy&pla[53])&(M1&T2)&(flags_nf);
ctl_reg_gp_sel_nuse_ixiypla53M1T3_1 = (~use_ixiy&pla[53])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla53M1T3_1,ctl_reg_gp_sel_nuse_ixiypla53M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla53M1T3_2 = (~use_ixiy&pla[53])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla53M1T3_2,ctl_reg_gp_hilo_nuse_ixiypla53M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[53])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[53])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[53])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[53])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[53])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[53])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[53])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[53])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[53])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[53])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[53])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[53])&(M1&T3);
validPLA = validPLA | (~use_ixiy&pla[53])&(M1&T4);
nextM = nextM | (~use_ixiy&pla[53])&(M1&T4);
ctl_mRead = ctl_mRead | (~use_ixiy&pla[53])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[53])&(M2&T1);
ctl_reg_gp_sel_nuse_ixiypla53M2T1_2 = (~use_ixiy&pla[53])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla53M2T1_2,ctl_reg_gp_sel_nuse_ixiypla53M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_nuse_ixiypla53M2T1_3 = (~use_ixiy&pla[53])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla53M2T1_3,ctl_reg_gp_hilo_nuse_ixiypla53M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[53])&(M2&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[53])&(M2&T1);
fMRead = fMRead | (~use_ixiy&pla[53])&(M2&T2);
fMRead = fMRead | (~use_ixiy&pla[53])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[53])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[53])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[53])&(M2&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[53])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[53])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_zero = ctl_alu_op2_sel_zero | (~use_ixiy&pla[53])&(M2&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[53])&(M2&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[53])&(M2&T3);
ctl_alu_core_hf = ctl_alu_core_hf | (~use_ixiy&pla[53])&(M2&T3)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[53])&(M2&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[53])&(M2&T3);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[53])&(M2&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[53])&(M2&T3);
ctl_flags_cf2_we = ctl_flags_cf2_we | (~use_ixiy&pla[53])&(M2&T3);
nextM = nextM | (~use_ixiy&pla[53])&(M2&T4);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[53])&(M2&T4);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[53])&(M2&T4);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[53])&(M2&T4);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[53])&(M2&T4);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[53])&(M2&T4);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[53])&(M2&T4);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[53])&(M2&T4);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[53])&(M2&T4);
ctl_alu_core_hf = ctl_alu_core_hf | (~use_ixiy&pla[53])&(M2&T4)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[53])&(M2&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[53])&(M2&T4);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[53])&(M2&T4);
ctl_pf_sel_nuse_ixiypla53M2T4_14 = (~use_ixiy&pla[53])&(M2&T4);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_nuse_ixiypla53M2T4_14,ctl_pf_sel_nuse_ixiypla53M2T4_14})&(`PFSEL_V);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (~use_ixiy&pla[53])&(M2&T4);
fMWrite = fMWrite | (~use_ixiy&pla[53])&(M3&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[53])&(M3&T1);
fMWrite = fMWrite | (~use_ixiy&pla[53])&(M3&T2);
fMWrite = fMWrite | (~use_ixiy&pla[53])&(M3&T3);
setM1 = setM1 | (~use_ixiy&pla[53])&(M3&T3);
fMRead = fMRead | (~use_ixiy&pla[53])&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[53])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[53])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[53])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[53])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[53])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[53])&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[53])&(M4&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[53])&(M4&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_zero = ctl_alu_op2_sel_zero | (~use_ixiy&pla[53])&(M4&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[53])&(M4&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[53])&(M4&T3);
ctl_alu_core_hf = ctl_alu_core_hf | (~use_ixiy&pla[53])&(M4&T3)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[53])&(M4&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[53])&(M4&T3);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[53])&(M4&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[53])&(M4&T3);
ctl_flags_cf2_we = ctl_flags_cf2_we | (~use_ixiy&pla[53])&(M4&T3);
nextM = nextM | (~use_ixiy&pla[53])&(M4&T4);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[53])&(M4&T4);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[53])&(M4&T4);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[53])&(M4&T4);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[53])&(M4&T4);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[53])&(M4&T4);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[53])&(M4&T4);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[53])&(M4&T4);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[53])&(M4&T4);
ctl_alu_core_hf = ctl_alu_core_hf | (~use_ixiy&pla[53])&(M4&T4)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[53])&(M4&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[53])&(M4&T4);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[53])&(M4&T4);
ctl_pf_sel_nuse_ixiypla53M4T4_14 = (~use_ixiy&pla[53])&(M4&T4);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_nuse_ixiypla53M4T4_14,ctl_pf_sel_nuse_ixiypla53M4T4_14})&(`PFSEL_V);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (~use_ixiy&pla[53])&(M4&T4);
fMWrite = fMWrite | (~use_ixiy&pla[53])&(M5&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[53])&(M5&T1);
fMWrite = fMWrite | (~use_ixiy&pla[53])&(M5&T2);
fMWrite = fMWrite | (~use_ixiy&pla[53])&(M5&T3);
setM1 = setM1 | (~use_ixiy&pla[53])&(M5&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[69])&(M1&T2);
ctl_reg_gp_sel_pla69M1T2_2 = (pla[69])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla69M1T2_2,ctl_reg_gp_sel_pla69M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla69M1T2_3 = (pla[69])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla69M1T2_3,ctl_reg_gp_hilo_pla69M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[69])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[69])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[69])&(M1&T2);
ctl_reg_gp_sel_pla69M1T3_1 = (pla[69])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla69M1T3_1,ctl_reg_gp_sel_pla69M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla69M1T3_2 = (pla[69])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla69M1T3_2,ctl_reg_gp_hilo_pla69M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[69])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[69])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[69])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[69])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[69])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[69])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[69])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[69])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[69])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[69])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[69])&(M1&T3);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[69])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[69])&(M1&T3);
validPLA = validPLA | (pla[69])&(M1&T4);
nextM = nextM | (pla[69])&(M1&T4);
ctl_reg_gp_sel_pla69M1T4_3 = (pla[69])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla69M1T4_3,ctl_reg_gp_sel_pla69M1T4_3})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla69M1T4_4 = (pla[69])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla69M1T4_4,ctl_reg_gp_hilo_pla69M1T4_4})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[69])&(M1&T4);
ctl_sw_2d = ctl_sw_2d | (pla[69])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[69])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[69])&(M1&T4);
ctl_reg_gp_sel_pla69M2T1_1 = (pla[69])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla69M2T1_1,ctl_reg_gp_sel_pla69M2T1_1})&(op54);
ctl_reg_gp_hilo_pla69M2T1_2 = (pla[69])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla69M2T1_2,ctl_reg_gp_hilo_pla69M2T1_2})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[69])&(M2&T1);
ctl_sw_2d = ctl_sw_2d | (pla[69])&(M2&T1);
ctl_flags_alu = ctl_flags_alu | (pla[69])&(M2&T1);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[69])&(M2&T1)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[69])&(M2&T1);
ctl_alu_op_low = ctl_alu_op_low | (pla[69])&(M2&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[69])&(M2&T1)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[69])&(M2&T1)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[69])&(M2&T1)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[69])&(M2&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[69])&(M2&T1);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[69])&(M2&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[69])&(M2&T2);
ctl_reg_sys_hilo_pla69M2T2_3 = (pla[69])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla69M2T2_3,ctl_reg_sys_hilo_pla69M2T2_3})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[69])&(M2&T2);
ctl_sw_2u = ctl_sw_2u | (pla[69])&(M2&T2);
ctl_flags_alu = ctl_flags_alu | (pla[69])&(M2&T2);
ctl_alu_oe = ctl_alu_oe | (pla[69])&(M2&T2);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[69])&(M2&T2);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[69])&(M2&T2);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[69])&(M2&T2)&(~ctl_alu_op_low);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[69])&(M2&T2);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[69])&(M2&T2);
ctl_reg_gp_sel_pla69M2T3_1 = (pla[69])&(M2&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla69M2T3_1,ctl_reg_gp_sel_pla69M2T3_1})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla69M2T3_2 = (pla[69])&(M2&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla69M2T3_2,ctl_reg_gp_hilo_pla69M2T3_2})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[69])&(M2&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[69])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[69])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[69])&(M2&T3);
nextM = nextM | (pla[69])&(M2&T4);
ctl_reg_gp_sel_pla69M2T4_2 = (pla[69])&(M2&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla69M2T4_2,ctl_reg_gp_sel_pla69M2T4_2})&(op54);
ctl_reg_gp_hilo_pla69M2T4_3 = (pla[69])&(M2&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla69M2T4_3,ctl_reg_gp_hilo_pla69M2T4_3})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[69])&(M2&T4);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[69])&(M2&T4);
ctl_flags_alu = ctl_flags_alu | (pla[69])&(M2&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[69])&(M2&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[69])&(M2&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[69])&(M2&T4);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[69])&(M2&T4)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[69])&(M2&T4);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[69])&(M2&T4);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[69])&(M3&T1);
ctl_reg_sys_hilo_pla69M3T1_2 = (pla[69])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla69M3T1_2,ctl_reg_sys_hilo_pla69M3T1_2})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[69])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[69])&(M3&T1);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[69])&(M3&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[69])&(M3&T1);
ctl_reg_sys_hilo_pla69M3T1_7 = (pla[69])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla69M3T1_7,ctl_reg_sys_hilo_pla69M3T1_7})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[69])&(M3&T1);
ctl_sw_2u = ctl_sw_2u | (pla[69])&(M3&T1);
ctl_flags_alu = ctl_flags_alu | (pla[69])&(M3&T1);
ctl_alu_oe = ctl_alu_oe | (pla[69])&(M3&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[69])&(M3&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[69])&(M3&T1);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[69])&(M3&T1)&(~ctl_alu_op_low);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[69])&(M3&T1);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[69])&(M3&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[69])&(M3&T2);
ctl_reg_gp_sel_pla69M3T2_2 = (pla[69])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla69M3T2_2,ctl_reg_gp_sel_pla69M3T2_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla69M3T2_3 = (pla[69])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla69M3T2_3,ctl_reg_gp_hilo_pla69M3T2_3})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[69])&(M3&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[69])&(M3&T2);
setM1 = setM1 | (pla[69])&(M3&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (op3&pla[68])&(M1&T2);
ctl_reg_gp_sel_op3pla68M1T2_2 = (op3&pla[68])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_op3pla68M1T2_2,ctl_reg_gp_sel_op3pla68M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_op3pla68M1T2_3 = (op3&pla[68])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_op3pla68M1T2_3,ctl_reg_gp_hilo_op3pla68M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (op3&pla[68])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (op3&pla[68])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (op3&pla[68])&(M1&T2);
ctl_reg_gp_sel_op3pla68M1T3_1 = (op3&pla[68])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_op3pla68M1T3_1,ctl_reg_gp_sel_op3pla68M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_op3pla68M1T3_2 = (op3&pla[68])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_op3pla68M1T3_2,ctl_reg_gp_hilo_op3pla68M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (op3&pla[68])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (op3&pla[68])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (op3&pla[68])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (op3&pla[68])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (op3&pla[68])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (op3&pla[68])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (op3&pla[68])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (op3&pla[68])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (op3&pla[68])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (op3&pla[68])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (op3&pla[68])&(M1&T3);
ctl_flags_nf_clr = ctl_flags_nf_clr | (op3&pla[68])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (op3&pla[68])&(M1&T3);
validPLA = validPLA | (op3&pla[68])&(M1&T4);
nextM = nextM | (op3&pla[68])&(M1&T4);
ctl_reg_gp_sel_op3pla68M1T4_3 = (op3&pla[68])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_op3pla68M1T4_3,ctl_reg_gp_sel_op3pla68M1T4_3})&(`GP_REG_HL);
ctl_reg_gp_hilo_op3pla68M1T4_4 = (op3&pla[68])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_op3pla68M1T4_4,ctl_reg_gp_hilo_op3pla68M1T4_4})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (op3&pla[68])&(M1&T4);
ctl_sw_2d = ctl_sw_2d | (op3&pla[68])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (op3&pla[68])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (op3&pla[68])&(M1&T4);
ctl_reg_gp_sel_op3pla68M2T1_1 = (op3&pla[68])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_op3pla68M2T1_1,ctl_reg_gp_sel_op3pla68M2T1_1})&(op54);
ctl_reg_gp_hilo_op3pla68M2T1_2 = (op3&pla[68])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_op3pla68M2T1_2,ctl_reg_gp_hilo_op3pla68M2T1_2})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (op3&pla[68])&(M2&T1);
ctl_sw_2d = ctl_sw_2d | (op3&pla[68])&(M2&T1);
ctl_flags_alu = ctl_flags_alu | (op3&pla[68])&(M2&T1);
ctl_alu_shift_oe = ctl_alu_shift_oe | (op3&pla[68])&(M2&T1)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (op3&pla[68])&(M2&T1);
ctl_alu_op_low = ctl_alu_op_low | (op3&pla[68])&(M2&T1);
ctl_alu_core_hf = ctl_alu_core_hf | (op3&pla[68])&(M2&T1)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (op3&pla[68])&(M2&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (op3&pla[68])&(M2&T1);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (op3&pla[68])&(M2&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (op3&pla[68])&(M2&T2);
ctl_reg_sys_hilo_op3pla68M2T2_3 = (op3&pla[68])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_op3pla68M2T2_3,ctl_reg_sys_hilo_op3pla68M2T2_3})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (op3&pla[68])&(M2&T2);
ctl_sw_2u = ctl_sw_2u | (op3&pla[68])&(M2&T2);
ctl_flags_alu = ctl_flags_alu | (op3&pla[68])&(M2&T2);
ctl_alu_oe = ctl_alu_oe | (op3&pla[68])&(M2&T2);
ctl_alu_res_oe = ctl_alu_res_oe | (op3&pla[68])&(M2&T2);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (op3&pla[68])&(M2&T2);
ctl_alu_core_hf = ctl_alu_core_hf | (op3&pla[68])&(M2&T2)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (op3&pla[68])&(M2&T2);
ctl_flags_xy_we = ctl_flags_xy_we | (op3&pla[68])&(M2&T2);
ctl_flags_cf_we = ctl_flags_cf_we | (op3&pla[68])&(M2&T2);
ctl_reg_gp_sel_op3pla68M2T3_1 = (op3&pla[68])&(M2&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_op3pla68M2T3_1,ctl_reg_gp_sel_op3pla68M2T3_1})&(`GP_REG_HL);
ctl_reg_gp_hilo_op3pla68M2T3_2 = (op3&pla[68])&(M2&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_op3pla68M2T3_2,ctl_reg_gp_hilo_op3pla68M2T3_2})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (op3&pla[68])&(M2&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (op3&pla[68])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (op3&pla[68])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (op3&pla[68])&(M2&T3);
nextM = nextM | (op3&pla[68])&(M2&T4);
ctl_reg_gp_sel_op3pla68M2T4_2 = (op3&pla[68])&(M2&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_op3pla68M2T4_2,ctl_reg_gp_sel_op3pla68M2T4_2})&(op54);
ctl_reg_gp_hilo_op3pla68M2T4_3 = (op3&pla[68])&(M2&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_op3pla68M2T4_3,ctl_reg_gp_hilo_op3pla68M2T4_3})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (op3&pla[68])&(M2&T4);
ctl_reg_out_lo = ctl_reg_out_lo | (op3&pla[68])&(M2&T4);
ctl_flags_alu = ctl_flags_alu | (op3&pla[68])&(M2&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (op3&pla[68])&(M2&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (op3&pla[68])&(M2&T4);
ctl_alu_op_low = ctl_alu_op_low | (op3&pla[68])&(M2&T4);
ctl_alu_core_hf = ctl_alu_core_hf | (op3&pla[68])&(M2&T4)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (op3&pla[68])&(M2&T4);
ctl_reg_use_sp = ctl_reg_use_sp | (op3&pla[68])&(M2&T4);
ctl_reg_sel_wz = ctl_reg_sel_wz | (op3&pla[68])&(M3&T1);
ctl_reg_sys_hilo_op3pla68M3T1_2 = (op3&pla[68])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_op3pla68M3T1_2,ctl_reg_sys_hilo_op3pla68M3T1_2})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (op3&pla[68])&(M3&T1);
ctl_al_we = ctl_al_we | (op3&pla[68])&(M3&T1);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (op3&pla[68])&(M3&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (op3&pla[68])&(M3&T1);
ctl_reg_sys_hilo_op3pla68M3T1_7 = (op3&pla[68])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_op3pla68M3T1_7,ctl_reg_sys_hilo_op3pla68M3T1_7})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (op3&pla[68])&(M3&T1);
ctl_sw_2u = ctl_sw_2u | (op3&pla[68])&(M3&T1);
ctl_flags_alu = ctl_flags_alu | (op3&pla[68])&(M3&T1);
ctl_alu_oe = ctl_alu_oe | (op3&pla[68])&(M3&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (op3&pla[68])&(M3&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (op3&pla[68])&(M3&T1);
ctl_alu_core_hf = ctl_alu_core_hf | (op3&pla[68])&(M3&T1)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (op3&pla[68])&(M3&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (op3&pla[68])&(M3&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (op3&pla[68])&(M3&T1);
ctl_pf_sel_op3pla68M3T1_18 = (op3&pla[68])&(M3&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_op3pla68M3T1_18,ctl_pf_sel_op3pla68M3T1_18})&(`PFSEL_V);
ctl_flags_cf_we = ctl_flags_cf_we | (op3&pla[68])&(M3&T1);
ctl_alu_zero_16bit = ctl_alu_zero_16bit | (op3&pla[68])&(M3&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (op3&pla[68])&(M3&T2);
ctl_reg_gp_sel_op3pla68M3T2_2 = (op3&pla[68])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_op3pla68M3T2_2,ctl_reg_gp_sel_op3pla68M3T2_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_op3pla68M3T2_3 = (op3&pla[68])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_op3pla68M3T2_3,ctl_reg_gp_hilo_op3pla68M3T2_3})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (op3&pla[68])&(M3&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (op3&pla[68])&(M3&T2);
setM1 = setM1 | (op3&pla[68])&(M3&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (~op3&pla[68])&(M1&T2);
ctl_reg_gp_sel_nop3pla68M1T2_2 = (~op3&pla[68])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nop3pla68M1T2_2,ctl_reg_gp_sel_nop3pla68M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_nop3pla68M1T2_3 = (~op3&pla[68])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nop3pla68M1T2_3,ctl_reg_gp_hilo_nop3pla68M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (~op3&pla[68])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (~op3&pla[68])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (~op3&pla[68])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (~op3&pla[68])&(M1&T2)&(flags_nf);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~op3&pla[68])&(M1&T2)&(flags_nf);
ctl_reg_gp_sel_nop3pla68M1T3_1 = (~op3&pla[68])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nop3pla68M1T3_1,ctl_reg_gp_sel_nop3pla68M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nop3pla68M1T3_2 = (~op3&pla[68])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nop3pla68M1T3_2,ctl_reg_gp_hilo_nop3pla68M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~op3&pla[68])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~op3&pla[68])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~op3&pla[68])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~op3&pla[68])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~op3&pla[68])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~op3&pla[68])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~op3&pla[68])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~op3&pla[68])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~op3&pla[68])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~op3&pla[68])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~op3&pla[68])&(M1&T3);
ctl_flags_nf_set = ctl_flags_nf_set | (~op3&pla[68])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~op3&pla[68])&(M1&T3);
validPLA = validPLA | (~op3&pla[68])&(M1&T4);
nextM = nextM | (~op3&pla[68])&(M1&T4);
ctl_reg_gp_sel_nop3pla68M1T4_3 = (~op3&pla[68])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nop3pla68M1T4_3,ctl_reg_gp_sel_nop3pla68M1T4_3})&(`GP_REG_HL);
ctl_reg_gp_hilo_nop3pla68M1T4_4 = (~op3&pla[68])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nop3pla68M1T4_4,ctl_reg_gp_hilo_nop3pla68M1T4_4})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (~op3&pla[68])&(M1&T4);
ctl_sw_2d = ctl_sw_2d | (~op3&pla[68])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~op3&pla[68])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~op3&pla[68])&(M1&T4);
ctl_reg_gp_sel_nop3pla68M2T1_1 = (~op3&pla[68])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nop3pla68M2T1_1,ctl_reg_gp_sel_nop3pla68M2T1_1})&(op54);
ctl_reg_gp_hilo_nop3pla68M2T1_2 = (~op3&pla[68])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nop3pla68M2T1_2,ctl_reg_gp_hilo_nop3pla68M2T1_2})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (~op3&pla[68])&(M2&T1);
ctl_sw_2d = ctl_sw_2d | (~op3&pla[68])&(M2&T1);
ctl_flags_alu = ctl_flags_alu | (~op3&pla[68])&(M2&T1);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~op3&pla[68])&(M2&T1)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~op3&pla[68])&(M2&T1);
ctl_alu_op_low = ctl_alu_op_low | (~op3&pla[68])&(M2&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~op3&pla[68])&(M2&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~op3&pla[68])&(M2&T1)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (~op3&pla[68])&(M2&T1)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (~op3&pla[68])&(M2&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (~op3&pla[68])&(M2&T1);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (~op3&pla[68])&(M2&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~op3&pla[68])&(M2&T2);
ctl_reg_sys_hilo_nop3pla68M2T2_3 = (~op3&pla[68])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nop3pla68M2T2_3,ctl_reg_sys_hilo_nop3pla68M2T2_3})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (~op3&pla[68])&(M2&T2);
ctl_sw_2u = ctl_sw_2u | (~op3&pla[68])&(M2&T2);
ctl_flags_alu = ctl_flags_alu | (~op3&pla[68])&(M2&T2);
ctl_alu_oe = ctl_alu_oe | (~op3&pla[68])&(M2&T2);
ctl_alu_res_oe = ctl_alu_res_oe | (~op3&pla[68])&(M2&T2);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~op3&pla[68])&(M2&T2);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~op3&pla[68])&(M2&T2);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~op3&pla[68])&(M2&T2)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (~op3&pla[68])&(M2&T2)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (~op3&pla[68])&(M2&T2);
ctl_flags_xy_we = ctl_flags_xy_we | (~op3&pla[68])&(M2&T2);
ctl_flags_cf_we = ctl_flags_cf_we | (~op3&pla[68])&(M2&T2);
ctl_reg_gp_sel_nop3pla68M2T3_1 = (~op3&pla[68])&(M2&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nop3pla68M2T3_1,ctl_reg_gp_sel_nop3pla68M2T3_1})&(`GP_REG_HL);
ctl_reg_gp_hilo_nop3pla68M2T3_2 = (~op3&pla[68])&(M2&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nop3pla68M2T3_2,ctl_reg_gp_hilo_nop3pla68M2T3_2})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (~op3&pla[68])&(M2&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~op3&pla[68])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~op3&pla[68])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~op3&pla[68])&(M2&T3);
nextM = nextM | (~op3&pla[68])&(M2&T4);
ctl_reg_gp_sel_nop3pla68M2T4_2 = (~op3&pla[68])&(M2&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nop3pla68M2T4_2,ctl_reg_gp_sel_nop3pla68M2T4_2})&(op54);
ctl_reg_gp_hilo_nop3pla68M2T4_3 = (~op3&pla[68])&(M2&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nop3pla68M2T4_3,ctl_reg_gp_hilo_nop3pla68M2T4_3})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (~op3&pla[68])&(M2&T4);
ctl_reg_out_lo = ctl_reg_out_lo | (~op3&pla[68])&(M2&T4);
ctl_flags_alu = ctl_flags_alu | (~op3&pla[68])&(M2&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~op3&pla[68])&(M2&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~op3&pla[68])&(M2&T4);
ctl_alu_op_low = ctl_alu_op_low | (~op3&pla[68])&(M2&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~op3&pla[68])&(M2&T4);
ctl_alu_core_hf = ctl_alu_core_hf | (~op3&pla[68])&(M2&T4)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (~op3&pla[68])&(M2&T4);
ctl_reg_use_sp = ctl_reg_use_sp | (~op3&pla[68])&(M2&T4);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~op3&pla[68])&(M3&T1);
ctl_reg_sys_hilo_nop3pla68M3T1_2 = (~op3&pla[68])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nop3pla68M3T1_2,ctl_reg_sys_hilo_nop3pla68M3T1_2})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~op3&pla[68])&(M3&T1);
ctl_al_we = ctl_al_we | (~op3&pla[68])&(M3&T1);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (~op3&pla[68])&(M3&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~op3&pla[68])&(M3&T1);
ctl_reg_sys_hilo_nop3pla68M3T1_7 = (~op3&pla[68])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nop3pla68M3T1_7,ctl_reg_sys_hilo_nop3pla68M3T1_7})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (~op3&pla[68])&(M3&T1);
ctl_sw_2u = ctl_sw_2u | (~op3&pla[68])&(M3&T1);
ctl_flags_alu = ctl_flags_alu | (~op3&pla[68])&(M3&T1);
ctl_alu_oe = ctl_alu_oe | (~op3&pla[68])&(M3&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~op3&pla[68])&(M3&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~op3&pla[68])&(M3&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~op3&pla[68])&(M3&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~op3&pla[68])&(M3&T1)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (~op3&pla[68])&(M3&T1)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (~op3&pla[68])&(M3&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (~op3&pla[68])&(M3&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (~op3&pla[68])&(M3&T1);
ctl_pf_sel_nop3pla68M3T1_20 = (~op3&pla[68])&(M3&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_nop3pla68M3T1_20,ctl_pf_sel_nop3pla68M3T1_20})&(`PFSEL_V);
ctl_flags_cf_we = ctl_flags_cf_we | (~op3&pla[68])&(M3&T1);
ctl_alu_zero_16bit = ctl_alu_zero_16bit | (~op3&pla[68])&(M3&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (~op3&pla[68])&(M3&T2);
ctl_reg_gp_sel_nop3pla68M3T2_2 = (~op3&pla[68])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nop3pla68M3T2_2,ctl_reg_gp_sel_nop3pla68M3T2_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_nop3pla68M3T2_3 = (~op3&pla[68])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nop3pla68M3T2_3,ctl_reg_gp_hilo_nop3pla68M3T2_3})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (~op3&pla[68])&(M3&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~op3&pla[68])&(M3&T2);
setM1 = setM1 | (~op3&pla[68])&(M3&T3);
validPLA = validPLA | (pla[9])&(M1&T4);
ctl_reg_gp_sel_pla9M1T4_2 = (pla[9])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla9M1T4_2,ctl_reg_gp_sel_pla9M1T4_2})&(op54);
ctl_reg_gp_hilo_pla9M1T4_3 = (pla[9])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla9M1T4_3,ctl_reg_gp_hilo_pla9M1T4_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[9])&(M1&T4);
ctl_al_we = ctl_al_we | (pla[9])&(M1&T4);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[9])&(M1&T4);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[9])&(M1&T5);
ctl_reg_gp_sel_pla9M1T5_2 = (pla[9])&(M1&T5);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla9M1T5_2,ctl_reg_gp_sel_pla9M1T5_2})&(op54);
ctl_reg_gp_hilo_pla9M1T5_3 = (pla[9])&(M1&T5);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla9M1T5_3,ctl_reg_gp_hilo_pla9M1T5_3})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[9])&(M1&T5);
ctl_inc_cy = ctl_inc_cy | (pla[9])&(M1&T5)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[9])&(M1&T5)&(op3);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[9])&(M1&T5);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[9])&(M1&T5);
setM1 = setM1 | (pla[9])&(M1&T6);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[77])&(M1&T1);
ctl_reg_gp_sel_pla77M1T1_2 = (pla[77])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla77M1T1_2,ctl_reg_gp_sel_pla77M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla77M1T1_3 = (pla[77])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla77M1T1_3,ctl_reg_gp_hilo_pla77M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[77])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[77])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[77])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[77])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[77])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[77])&(M1&T1);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[77])&(M1&T1)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[77])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[77])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[77])&(M1&T1);
ctl_pf_sel_pla77M1T1_14 = (pla[77])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla77M1T1_14,ctl_pf_sel_pla77M1T1_14})&(`PFSEL_P);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[77])&(M1&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[77])&(M1&T1)&(flags_nf);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[77])&(M1&T1)&(~flags_nf);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[77])&(M1&T2);
ctl_reg_gp_sel_pla77M1T2_2 = (pla[77])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla77M1T2_2,ctl_reg_gp_sel_pla77M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla77M1T2_3 = (pla[77])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla77M1T2_3,ctl_reg_gp_hilo_pla77M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[77])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[77])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[77])&(M1&T2);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (pla[77])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (pla[77])&(M1&T2)&(flags_nf);
ctl_reg_gp_sel_pla77M1T3_1 = (pla[77])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla77M1T3_1,ctl_reg_gp_sel_pla77M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla77M1T3_2 = (pla[77])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla77M1T3_2,ctl_reg_gp_hilo_pla77M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[77])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[77])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[77])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[77])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[77])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[77])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[77])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[77])&(M1&T3);
ctl_flags_hf2_we = ctl_flags_hf2_we | (pla[77])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[77])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[77])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[77])&(M1&T3);
validPLA = validPLA | (pla[77])&(M1&T4);
setM1 = setM1 | (pla[77])&(M1&T4);
ctl_sw_2d = ctl_sw_2d | (pla[77])&(M1&T4);
ctl_flags_alu = ctl_flags_alu | (pla[77])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[77])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[77])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[77])&(M1&T4);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[77])&(M1&T4)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[77])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[77])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[77])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[77])&(M1&T4);
ctl_flags_cf2_we = ctl_flags_cf2_we | (pla[77])&(M1&T4);
ctl_flags_cf2_sel_daa = ctl_flags_cf2_sel_daa | (pla[77])&(M1&T4);
ctl_daa_oe = ctl_daa_oe | (pla[77])&(M1&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[77])&(M1&T4)&(flags_nf);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[77])&(M1&T4)&(~flags_nf);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[81])&(M1&T1);
ctl_reg_gp_sel_pla81M1T1_2 = (pla[81])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla81M1T1_2,ctl_reg_gp_sel_pla81M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla81M1T1_3 = (pla[81])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla81M1T1_3,ctl_reg_gp_hilo_pla81M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[81])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[81])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[81])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[81])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[81])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[81])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[81])&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (pla[81])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (pla[81])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[81])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[81])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[81])&(M1&T1);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[81])&(M1&T1);
ctl_flags_nf_set = ctl_flags_nf_set | (pla[81])&(M1&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[81])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[81])&(M1&T2);
ctl_reg_gp_sel_pla81M1T2_2 = (pla[81])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla81M1T2_2,ctl_reg_gp_sel_pla81M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla81M1T2_3 = (pla[81])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla81M1T2_3,ctl_reg_gp_hilo_pla81M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[81])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[81])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[81])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (pla[81])&(M1&T2)&(flags_nf);
ctl_reg_gp_sel_pla81M1T3_1 = (pla[81])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla81M1T3_1,ctl_reg_gp_sel_pla81M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla81M1T3_2 = (pla[81])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla81M1T3_2,ctl_reg_gp_hilo_pla81M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[81])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[81])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[81])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[81])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[81])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[81])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[81])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[81])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[81])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[81])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[81])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[81])&(M1&T3);
validPLA = validPLA | (pla[81])&(M1&T4);
setM1 = setM1 | (pla[81])&(M1&T4);
ctl_flags_alu = ctl_flags_alu | (pla[81])&(M1&T4);
ctl_alu_op1_sel_zero = ctl_alu_op1_sel_zero | (pla[81])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[81])&(M1&T4);
ctl_alu_core_R = ctl_alu_core_R | (pla[81])&(M1&T4);
ctl_alu_core_V = ctl_alu_core_V | (pla[81])&(M1&T4);
ctl_alu_core_S = ctl_alu_core_S | (pla[81])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[81])&(M1&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[81])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[81])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[81])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[81])&(M1&T4);
ctl_flags_nf_set = ctl_flags_nf_set | (pla[81])&(M1&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[81])&(M1&T4);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[82])&(M1&T1);
ctl_reg_gp_sel_pla82M1T1_2 = (pla[82])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla82M1T1_2,ctl_reg_gp_sel_pla82M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla82M1T1_3 = (pla[82])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla82M1T1_3,ctl_reg_gp_hilo_pla82M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[82])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[82])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[82])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[82])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[82])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[82])&(M1&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[82])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[82])&(M1&T1)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[82])&(M1&T1)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[82])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[82])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[82])&(M1&T1);
ctl_pf_sel_pla82M1T1_16 = (pla[82])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla82M1T1_16,ctl_pf_sel_pla82M1T1_16})&(`PFSEL_V);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[82])&(M1&T1);
ctl_flags_nf_set = ctl_flags_nf_set | (pla[82])&(M1&T1);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[82])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[82])&(M1&T2);
ctl_reg_gp_sel_pla82M1T2_2 = (pla[82])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla82M1T2_2,ctl_reg_gp_sel_pla82M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla82M1T2_3 = (pla[82])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla82M1T2_3,ctl_reg_gp_hilo_pla82M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[82])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[82])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[82])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (pla[82])&(M1&T2)&(flags_nf);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[82])&(M1&T2)&(flags_nf);
ctl_reg_gp_sel_pla82M1T3_1 = (pla[82])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla82M1T3_1,ctl_reg_gp_sel_pla82M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla82M1T3_2 = (pla[82])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla82M1T3_2,ctl_reg_gp_hilo_pla82M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[82])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[82])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[82])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[82])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[82])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[82])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[82])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[82])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[82])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[82])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[82])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[82])&(M1&T3);
validPLA = validPLA | (pla[82])&(M1&T4);
setM1 = setM1 | (pla[82])&(M1&T4);
ctl_flags_alu = ctl_flags_alu | (pla[82])&(M1&T4);
ctl_alu_op1_sel_zero = ctl_alu_op1_sel_zero | (pla[82])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[82])&(M1&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[82])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[82])&(M1&T4)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[82])&(M1&T4)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[82])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[82])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[82])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[82])&(M1&T4);
ctl_flags_nf_set = ctl_flags_nf_set | (pla[82])&(M1&T4);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[82])&(M1&T4);
ctl_flags_alu = ctl_flags_alu | (pla[89])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[89])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[89])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[89])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[89])&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (pla[89])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (pla[89])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[89])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[89])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[89])&(M1&T1);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[89])&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[89])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[89])&(M1&T2);
ctl_reg_gp_sel_pla89M1T2_2 = (pla[89])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla89M1T2_2,ctl_reg_gp_sel_pla89M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla89M1T2_3 = (pla[89])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla89M1T2_3,ctl_reg_gp_hilo_pla89M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[89])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[89])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[89])&(M1&T2);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[89])&(M1&T2);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[89])&(M1&T2);
ctl_flags_hf_cpl = ctl_flags_hf_cpl | (pla[89])&(M1&T2)&(~flags_cf);
ctl_reg_gp_sel_pla89M1T3_1 = (pla[89])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla89M1T3_1,ctl_reg_gp_sel_pla89M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla89M1T3_2 = (pla[89])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla89M1T3_2,ctl_reg_gp_hilo_pla89M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[89])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[89])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[89])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[89])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[89])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[89])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[89])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[89])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[89])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[89])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[89])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[89])&(M1&T3);
validPLA = validPLA | (pla[89])&(M1&T4);
setM1 = setM1 | (pla[89])&(M1&T4);
ctl_flags_alu = ctl_flags_alu | (pla[89])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[89])&(M1&T4);
ctl_alu_core_R = ctl_alu_core_R | (pla[89])&(M1&T4);
ctl_alu_core_V = ctl_alu_core_V | (pla[89])&(M1&T4);
ctl_alu_core_S = ctl_alu_core_S | (pla[89])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[89])&(M1&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[89])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[89])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[89])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[89])&(M1&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[89])&(M1&T4);
ctl_flags_alu = ctl_flags_alu | (pla[92])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[92])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[92])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[92])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[92])&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (pla[92])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (pla[92])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[92])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[92])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[92])&(M1&T1);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[92])&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[92])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[92])&(M1&T2);
ctl_reg_gp_sel_pla92M1T2_2 = (pla[92])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla92M1T2_2,ctl_reg_gp_sel_pla92M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla92M1T2_3 = (pla[92])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla92M1T2_3,ctl_reg_gp_hilo_pla92M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[92])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[92])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[92])&(M1&T2);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[92])&(M1&T2);
ctl_reg_gp_sel_pla92M1T3_1 = (pla[92])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla92M1T3_1,ctl_reg_gp_sel_pla92M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla92M1T3_2 = (pla[92])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla92M1T3_2,ctl_reg_gp_hilo_pla92M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[92])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[92])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[92])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[92])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[92])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[92])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[92])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[92])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[92])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[92])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[92])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[92])&(M1&T3);
validPLA = validPLA | (pla[92])&(M1&T4);
setM1 = setM1 | (pla[92])&(M1&T4);
ctl_flags_alu = ctl_flags_alu | (pla[92])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[92])&(M1&T4);
ctl_alu_core_R = ctl_alu_core_R | (pla[92])&(M1&T4);
ctl_alu_core_V = ctl_alu_core_V | (pla[92])&(M1&T4);
ctl_alu_core_S = ctl_alu_core_S | (pla[92])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[92])&(M1&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[92])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[92])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[92])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[92])&(M1&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[92])&(M1&T4);
ctl_state_halt_set = ctl_state_halt_set | (pla[95])&(M1&T3);
validPLA = validPLA | (pla[95])&(M1&T4);
setM1 = setM1 | (pla[95])&(M1&T4);
ctl_iffx_bit = ctl_iffx_bit | (pla[97])&(M1&T3)&(op3);
ctl_iffx_we = ctl_iffx_we | (pla[97])&(M1&T3);
validPLA = validPLA | (pla[97])&(M1&T4);
setM1 = setM1 | (pla[97])&(M1&T4);
ctl_no_ints = ctl_no_ints | (pla[97])&(M1&T4);
ctl_sw_1d = ctl_sw_1d | (pla[96])&(M1&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[96])&(M1&T3);
ctl_im_we = ctl_im_we | (pla[96])&(M1&T3);
validPLA = validPLA | (pla[96])&(M1&T4);
setM1 = setM1 | (pla[96])&(M1&T4);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[25])&(M1&T1);
ctl_reg_gp_sel_pla25M1T1_2 = (pla[25])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla25M1T1_2,ctl_reg_gp_sel_pla25M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla25M1T1_3 = (pla[25])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla25M1T1_3,ctl_reg_gp_hilo_pla25M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[25])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[25])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[25])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[25])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[25])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[25])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[25])&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (pla[25])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (pla[25])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[25])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[25])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[25])&(M1&T1);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[25])&(M1&T1);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[25])&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[25])&(M1&T1);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[25])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[25])&(M1&T2);
ctl_reg_gp_sel_pla25M1T2_2 = (pla[25])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla25M1T2_2,ctl_reg_gp_sel_pla25M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla25M1T2_3 = (pla[25])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla25M1T2_3,ctl_reg_gp_hilo_pla25M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[25])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[25])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[25])&(M1&T2);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (pla[25])&(M1&T2);
ctl_reg_gp_sel_pla25M1T3_1 = (pla[25])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla25M1T3_1,ctl_reg_gp_sel_pla25M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla25M1T3_2 = (pla[25])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla25M1T3_2,ctl_reg_gp_hilo_pla25M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[25])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[25])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[25])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[25])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[25])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[25])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[25])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[25])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[25])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[25])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[25])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[25])&(M1&T3);
validPLA = validPLA | (pla[25])&(M1&T4);
setM1 = setM1 | (pla[25])&(M1&T4);
ctl_reg_gp_sel_pla25M1T4_3 = (pla[25])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla25M1T4_3,ctl_reg_gp_sel_pla25M1T4_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla25M1T4_4 = (pla[25])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla25M1T4_4,ctl_reg_gp_hilo_pla25M1T4_4})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[25])&(M1&T4);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[25])&(M1&T4);
ctl_flags_alu = ctl_flags_alu | (pla[25])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[25])&(M1&T4);
ctl_shift_en = ctl_shift_en | (pla[25])&(M1&T4);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[25])&(M1&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[25])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[25])&(M1&T4);
ctl_alu_core_R = ctl_alu_core_R | (pla[25])&(M1&T4);
ctl_alu_core_V = ctl_alu_core_V | (pla[25])&(M1&T4);
ctl_alu_core_S = ctl_alu_core_S | (pla[25])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[25])&(M1&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[25])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[25])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[25])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[25])&(M1&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[25])&(M1&T4);
ctl_flags_cf2_we = ctl_flags_cf2_we | (pla[25])&(M1&T4);
ctl_flags_cf2_sel_shift = ctl_flags_cf2_sel_shift | (pla[25])&(M1&T4);
ctl_reg_gp_we = ctl_reg_gp_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_reg_gp_sel_nuse_ixiypla70npla55M1T1_2 = (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla70npla55M1T1_2,ctl_reg_gp_sel_nuse_ixiypla70npla55M1T1_2})&(op21);
ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T1_3 = (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T1_3,ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T1_3})&({~rsel0,rsel0});
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_pf_sel_nuse_ixiypla70npla55M1T1_20 = (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_nuse_ixiypla70npla55M1T1_20,ctl_pf_sel_nuse_ixiypla70npla55M1T1_20})&(`PFSEL_P);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T2);
ctl_reg_gp_sel_nuse_ixiypla70npla55M1T2_2 = (~use_ixiy&pla[70]&~pla[55])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla70npla55M1T2_2,ctl_reg_gp_sel_nuse_ixiypla70npla55M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T2_3 = (~use_ixiy&pla[70]&~pla[55])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T2_3,ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[70]&~pla[55])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[70]&~pla[55])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (~use_ixiy&pla[70]&~pla[55])&(M1&T2);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (~use_ixiy&pla[70]&~pla[55])&(M1&T2);
ctl_reg_gp_sel_nuse_ixiypla70npla55M1T3_1 = (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla70npla55M1T3_1,ctl_reg_gp_sel_nuse_ixiypla70npla55M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T3_2 = (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T3_2,ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[70]&~pla[55])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T3);
validPLA = validPLA | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
setM1 = setM1 | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_reg_gp_sel_nuse_ixiypla70npla55M1T4_3 = (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla70npla55M1T4_3,ctl_reg_gp_sel_nuse_ixiypla70npla55M1T4_3})&(op21);
ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T4_4 = (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T4_4,ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T4_4})&({~rsel0,rsel0});
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[70]&~pla[55])&(M1&T4)&(~rsel0);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[70]&~pla[55])&(M1&T4)&(rsel0);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[70]&~pla[55])&(M1&T4)&(~rsel0);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[70]&~pla[55])&(M1&T4)&(rsel0);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_shift_en = ctl_shift_en | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_flags_cf2_we = ctl_flags_cf2_we | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
ctl_flags_cf2_sel_shift = ctl_flags_cf2_sel_shift | (~use_ixiy&pla[70]&~pla[55])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[70]&~pla[55])&(M4&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~use_ixiy&pla[70]&~pla[55])&(M4&T1);
ctl_reg_sys_hilo_nuse_ixiypla70npla55M4T1_3 = (~use_ixiy&pla[70]&~pla[55])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nuse_ixiypla70npla55M4T1_3,ctl_reg_sys_hilo_nuse_ixiypla70npla55M4T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[70]&~pla[55])&(M4&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[70]&~pla[55])&(M4&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[70]&~pla[55])&(M4&T1);
ctl_ir_we = ctl_ir_we | (~use_ixiy&pla[70]&~pla[55])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[70]&~pla[55])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
nextM = nextM | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_shift_en = ctl_shift_en | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_flags_cf2_we = ctl_flags_cf2_we | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
ctl_flags_cf2_sel_shift = ctl_flags_cf2_sel_shift | (~use_ixiy&pla[70]&~pla[55])&(M4&T3);
fMWrite = fMWrite | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_pf_sel_nuse_ixiypla70npla55M5T1_19 = (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_nuse_ixiypla70npla55M5T1_19,ctl_pf_sel_nuse_ixiypla70npla55M5T1_19})&(`PFSEL_P);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[70]&~pla[55])&(M5&T1);
fMWrite = fMWrite | (~use_ixiy&pla[70]&~pla[55])&(M5&T2);
fMWrite = fMWrite | (~use_ixiy&pla[70]&~pla[55])&(M5&T3);
setM1 = setM1 | (~use_ixiy&pla[70]&~pla[55])&(M5&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (~use_ixiy&pla[70]&pla[55])&(M1&T2);
ctl_reg_gp_sel_nuse_ixiypla70pla55M1T2_2 = (~use_ixiy&pla[70]&pla[55])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla70pla55M1T2_2,ctl_reg_gp_sel_nuse_ixiypla70pla55M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla70pla55M1T2_3 = (~use_ixiy&pla[70]&pla[55])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla70pla55M1T2_3,ctl_reg_gp_hilo_nuse_ixiypla70pla55M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[70]&pla[55])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[70]&pla[55])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (~use_ixiy&pla[70]&pla[55])&(M1&T2);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (~use_ixiy&pla[70]&pla[55])&(M1&T2);
ctl_reg_gp_sel_nuse_ixiypla70pla55M1T3_1 = (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla70pla55M1T3_1,ctl_reg_gp_sel_nuse_ixiypla70pla55M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla70pla55M1T3_2 = (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla70pla55M1T3_2,ctl_reg_gp_hilo_nuse_ixiypla70pla55M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[70]&pla[55])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[70]&pla[55])&(M1&T3);
validPLA = validPLA | (~use_ixiy&pla[70]&pla[55])&(M1&T4);
nextM = nextM | (~use_ixiy&pla[70]&pla[55])&(M1&T4);
ctl_mRead = ctl_mRead | (~use_ixiy&pla[70]&pla[55])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[70]&pla[55])&(M2&T1);
ctl_reg_gp_sel_nuse_ixiypla70pla55M2T1_2 = (~use_ixiy&pla[70]&pla[55])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla70pla55M2T1_2,ctl_reg_gp_sel_nuse_ixiypla70pla55M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_nuse_ixiypla70pla55M2T1_3 = (~use_ixiy&pla[70]&pla[55])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla70pla55M2T1_3,ctl_reg_gp_hilo_nuse_ixiypla70pla55M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[70]&pla[55])&(M2&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[70]&pla[55])&(M2&T1);
fMRead = fMRead | (~use_ixiy&pla[70]&pla[55])&(M2&T2);
fMRead = fMRead | (~use_ixiy&pla[70]&pla[55])&(M2&T3);
nextM = nextM | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_shift_en = ctl_shift_en | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_flags_cf2_we = ctl_flags_cf2_we | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
ctl_flags_cf2_sel_shift = ctl_flags_cf2_sel_shift | (~use_ixiy&pla[70]&pla[55])&(M2&T4);
fMWrite = fMWrite | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_pf_sel_nuse_ixiypla70pla55M3T1_19 = (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_nuse_ixiypla70pla55M3T1_19,ctl_pf_sel_nuse_ixiypla70pla55M3T1_19})&(`PFSEL_P);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[70]&pla[55])&(M3&T1);
fMWrite = fMWrite | (~use_ixiy&pla[70]&pla[55])&(M3&T2);
fMWrite = fMWrite | (~use_ixiy&pla[70]&pla[55])&(M3&T3);
setM1 = setM1 | (~use_ixiy&pla[70]&pla[55])&(M3&T3);
fMRead = fMRead | (~use_ixiy&pla[70]&pla[55])&(M4&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~use_ixiy&pla[70]&pla[55])&(M4&T1);
ctl_reg_sys_hilo_nuse_ixiypla70pla55M4T1_3 = (~use_ixiy&pla[70]&pla[55])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nuse_ixiypla70pla55M4T1_3,ctl_reg_sys_hilo_nuse_ixiypla70pla55M4T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[70]&pla[55])&(M4&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[70]&pla[55])&(M4&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[70]&pla[55])&(M4&T1);
ctl_ir_we = ctl_ir_we | (~use_ixiy&pla[70]&pla[55])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[70]&pla[55])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
nextM = nextM | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_shift_en = ctl_shift_en | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_flags_cf2_we = ctl_flags_cf2_we | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
ctl_flags_cf2_sel_shift = ctl_flags_cf2_sel_shift | (~use_ixiy&pla[70]&pla[55])&(M4&T3);
fMWrite = fMWrite | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_pf_sel_nuse_ixiypla70pla55M5T1_19 = (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_nuse_ixiypla70pla55M5T1_19,ctl_pf_sel_nuse_ixiypla70pla55M5T1_19})&(`PFSEL_P);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[70]&pla[55])&(M5&T1);
fMWrite = fMWrite | (~use_ixiy&pla[70]&pla[55])&(M5&T2);
fMWrite = fMWrite | (~use_ixiy&pla[70]&pla[55])&(M5&T3);
setM1 = setM1 | (~use_ixiy&pla[70]&pla[55])&(M5&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[15]&op3)&(M1&T1);
ctl_reg_gp_sel_pla15op3M1T1_2 = (pla[15]&op3)&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla15op3M1T1_2,ctl_reg_gp_sel_pla15op3M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla15op3M1T1_3 = (pla[15]&op3)&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla15op3M1T1_3,ctl_reg_gp_hilo_pla15op3M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[15]&op3)&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[15]&op3)&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[15]&op3)&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[15]&op3)&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[15]&op3)&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[15]&op3)&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[15]&op3)&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (pla[15]&op3)&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (pla[15]&op3)&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[15]&op3)&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[15]&op3)&(M1&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[15]&op3)&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[15]&op3)&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[15]&op3)&(M1&T1);
ctl_pf_sel_pla15op3M1T1_18 = (pla[15]&op3)&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla15op3M1T1_18,ctl_pf_sel_pla15op3M1T1_18})&(`PFSEL_P);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[15]&op3)&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[15]&op3)&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[15]&op3)&(M1&T2);
ctl_reg_gp_sel_pla15op3M1T2_2 = (pla[15]&op3)&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla15op3M1T2_2,ctl_reg_gp_sel_pla15op3M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla15op3M1T2_3 = (pla[15]&op3)&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla15op3M1T2_3,ctl_reg_gp_hilo_pla15op3M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[15]&op3)&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[15]&op3)&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[15]&op3)&(M1&T2);
ctl_reg_gp_sel_pla15op3M1T3_1 = (pla[15]&op3)&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla15op3M1T3_1,ctl_reg_gp_sel_pla15op3M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla15op3M1T3_2 = (pla[15]&op3)&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla15op3M1T3_2,ctl_reg_gp_hilo_pla15op3M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[15]&op3)&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[15]&op3)&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[15]&op3)&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[15]&op3)&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[15]&op3)&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[15]&op3)&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[15]&op3)&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[15]&op3)&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[15]&op3)&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[15]&op3)&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[15]&op3)&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[15]&op3)&(M1&T3);
validPLA = validPLA | (pla[15]&op3)&(M1&T4);
nextM = nextM | (pla[15]&op3)&(M1&T4);
ctl_mRead = ctl_mRead | (pla[15]&op3)&(M1&T4);
fMRead = fMRead | (pla[15]&op3)&(M2&T1);
ctl_reg_gp_sel_pla15op3M2T1_2 = (pla[15]&op3)&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla15op3M2T1_2,ctl_reg_gp_sel_pla15op3M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla15op3M2T1_3 = (pla[15]&op3)&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla15op3M2T1_3,ctl_reg_gp_hilo_pla15op3M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[15]&op3)&(M2&T1);
ctl_al_we = ctl_al_we | (pla[15]&op3)&(M2&T1);
fMRead = fMRead | (pla[15]&op3)&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[15]&op3)&(M2&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[15]&op3)&(M2&T2);
ctl_reg_sys_hilo_pla15op3M2T2_4 = (pla[15]&op3)&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla15op3M2T2_4,ctl_reg_sys_hilo_pla15op3M2T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[15]&op3)&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[15]&op3)&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[15]&op3)&(M2&T2);
fMRead = fMRead | (pla[15]&op3)&(M2&T3);
nextM = nextM | (pla[15]&op3)&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[15]&op3)&(M3&T1);
ctl_sw_1d = ctl_sw_1d | (pla[15]&op3)&(M3&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[15]&op3)&(M3&T1);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[15]&op3)&(M3&T1)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_lq = ctl_alu_op2_sel_lq | (pla[15]&op3)&(M3&T1);
ctl_alu_op_low = ctl_alu_op_low | (pla[15]&op3)&(M3&T1);
nextM = nextM | (pla[15]&op3)&(M3&T4);
ctl_mWrite = ctl_mWrite | (pla[15]&op3)&(M3&T4);
ctl_sw_2d = ctl_sw_2d | (pla[15]&op3)&(M3&T4);
ctl_sw_1d = ctl_sw_1d | (pla[15]&op3)&(M3&T4);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[15]&op3)&(M3&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[15]&op3)&(M3&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_low = ctl_alu_op1_sel_low | (pla[15]&op3)&(M3&T4);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[15]&op3)&(M3&T4);
fMWrite = fMWrite | (pla[15]&op3)&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[15]&op3)&(M4&T1);
ctl_sw_2u = ctl_sw_2u | (pla[15]&op3)&(M4&T1);
ctl_sw_1u = ctl_sw_1u | (pla[15]&op3)&(M4&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[15]&op3)&(M4&T1);
ctl_alu_oe = ctl_alu_oe | (pla[15]&op3)&(M4&T1);
ctl_alu_op2_oe = ctl_alu_op2_oe | (pla[15]&op3)&(M4&T1);
fMWrite = fMWrite | (pla[15]&op3)&(M4&T2);
ctl_alu_op1_oe = ctl_alu_op1_oe | (pla[15]&op3)&(M4&T2);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[15]&op3)&(M4&T2);
fMWrite = fMWrite | (pla[15]&op3)&(M4&T3);
setM1 = setM1 | (pla[15]&op3)&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (pla[15]&op3)&(M4&T3);
ctl_alu_op_low = ctl_alu_op_low | (pla[15]&op3)&(M4&T3);
ctl_alu_core_R = ctl_alu_core_R | (pla[15]&op3)&(M4&T3);
ctl_alu_core_V = ctl_alu_core_V | (pla[15]&op3)&(M4&T3);
ctl_alu_core_S = ctl_alu_core_S | (pla[15]&op3)&(M4&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[15]&op3)&(M4&T3);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[15]&op3)&(M4&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[15]&op3)&(M4&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[15]&op3)&(M4&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[15]&op3)&(M4&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[15]&op3)&(M4&T3);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[15]&op3)&(M4&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[15]&~op3)&(M1&T1);
ctl_reg_gp_sel_pla15nop3M1T1_2 = (pla[15]&~op3)&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla15nop3M1T1_2,ctl_reg_gp_sel_pla15nop3M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla15nop3M1T1_3 = (pla[15]&~op3)&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla15nop3M1T1_3,ctl_reg_gp_hilo_pla15nop3M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[15]&~op3)&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[15]&~op3)&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[15]&~op3)&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[15]&~op3)&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[15]&~op3)&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[15]&~op3)&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[15]&~op3)&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (pla[15]&~op3)&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (pla[15]&~op3)&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[15]&~op3)&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[15]&~op3)&(M1&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[15]&~op3)&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[15]&~op3)&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[15]&~op3)&(M1&T1);
ctl_pf_sel_pla15nop3M1T1_18 = (pla[15]&~op3)&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla15nop3M1T1_18,ctl_pf_sel_pla15nop3M1T1_18})&(`PFSEL_P);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[15]&~op3)&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[15]&~op3)&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[15]&~op3)&(M1&T2);
ctl_reg_gp_sel_pla15nop3M1T2_2 = (pla[15]&~op3)&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla15nop3M1T2_2,ctl_reg_gp_sel_pla15nop3M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla15nop3M1T2_3 = (pla[15]&~op3)&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla15nop3M1T2_3,ctl_reg_gp_hilo_pla15nop3M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[15]&~op3)&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[15]&~op3)&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[15]&~op3)&(M1&T2);
ctl_reg_gp_sel_pla15nop3M1T3_1 = (pla[15]&~op3)&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla15nop3M1T3_1,ctl_reg_gp_sel_pla15nop3M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla15nop3M1T3_2 = (pla[15]&~op3)&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla15nop3M1T3_2,ctl_reg_gp_hilo_pla15nop3M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[15]&~op3)&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[15]&~op3)&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[15]&~op3)&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[15]&~op3)&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[15]&~op3)&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[15]&~op3)&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[15]&~op3)&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[15]&~op3)&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[15]&~op3)&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[15]&~op3)&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[15]&~op3)&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[15]&~op3)&(M1&T3);
validPLA = validPLA | (pla[15]&~op3)&(M1&T4);
nextM = nextM | (pla[15]&~op3)&(M1&T4);
ctl_mRead = ctl_mRead | (pla[15]&~op3)&(M1&T4);
fMRead = fMRead | (pla[15]&~op3)&(M2&T1);
ctl_reg_gp_sel_pla15nop3M2T1_2 = (pla[15]&~op3)&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla15nop3M2T1_2,ctl_reg_gp_sel_pla15nop3M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla15nop3M2T1_3 = (pla[15]&~op3)&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla15nop3M2T1_3,ctl_reg_gp_hilo_pla15nop3M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[15]&~op3)&(M2&T1);
ctl_al_we = ctl_al_we | (pla[15]&~op3)&(M2&T1);
fMRead = fMRead | (pla[15]&~op3)&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[15]&~op3)&(M2&T2);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[15]&~op3)&(M2&T2);
ctl_reg_sys_hilo_pla15nop3M2T2_4 = (pla[15]&~op3)&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla15nop3M2T2_4,ctl_reg_sys_hilo_pla15nop3M2T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[15]&~op3)&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[15]&~op3)&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[15]&~op3)&(M2&T2);
fMRead = fMRead | (pla[15]&~op3)&(M2&T3);
nextM = nextM | (pla[15]&~op3)&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[15]&~op3)&(M3&T1);
ctl_sw_1d = ctl_sw_1d | (pla[15]&~op3)&(M3&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[15]&~op3)&(M3&T1);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[15]&~op3)&(M3&T1)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_lq = ctl_alu_op2_sel_lq | (pla[15]&~op3)&(M3&T1);
ctl_alu_op1_sel_low = ctl_alu_op1_sel_low | (pla[15]&~op3)&(M3&T1);
ctl_alu_op_low = ctl_alu_op_low | (pla[15]&~op3)&(M3&T1);
ctl_sw_2u = ctl_sw_2u | (pla[15]&~op3)&(M3&T2);
ctl_sw_1u = ctl_sw_1u | (pla[15]&~op3)&(M3&T2);
ctl_bus_db_we = ctl_bus_db_we | (pla[15]&~op3)&(M3&T2);
ctl_alu_oe = ctl_alu_oe | (pla[15]&~op3)&(M3&T2);
ctl_alu_op2_oe = ctl_alu_op2_oe | (pla[15]&~op3)&(M3&T2);
ctl_reg_gp_sel_pla15nop3M3T3_1 = (pla[15]&~op3)&(M3&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla15nop3M3T3_1,ctl_reg_gp_sel_pla15nop3M3T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla15nop3M3T3_2 = (pla[15]&~op3)&(M3&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla15nop3M3T3_2,ctl_reg_gp_hilo_pla15nop3M3T3_2})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[15]&~op3)&(M3&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[15]&~op3)&(M3&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[15]&~op3)&(M3&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_lq = ctl_alu_op2_sel_lq | (pla[15]&~op3)&(M3&T3);
ctl_alu_op_low = ctl_alu_op_low | (pla[15]&~op3)&(M3&T3);
nextM = nextM | (pla[15]&~op3)&(M3&T4);
ctl_mWrite = ctl_mWrite | (pla[15]&~op3)&(M3&T4);
ctl_sw_2d = ctl_sw_2d | (pla[15]&~op3)&(M3&T4);
ctl_sw_1d = ctl_sw_1d | (pla[15]&~op3)&(M3&T4);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[15]&~op3)&(M3&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[15]&~op3)&(M3&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_low = ctl_alu_op1_sel_low | (pla[15]&~op3)&(M3&T4);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[15]&~op3)&(M3&T4);
fMWrite = fMWrite | (pla[15]&~op3)&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[15]&~op3)&(M4&T1);
ctl_sw_2u = ctl_sw_2u | (pla[15]&~op3)&(M4&T1);
ctl_sw_1u = ctl_sw_1u | (pla[15]&~op3)&(M4&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[15]&~op3)&(M4&T1);
ctl_alu_oe = ctl_alu_oe | (pla[15]&~op3)&(M4&T1);
ctl_alu_op2_oe = ctl_alu_op2_oe | (pla[15]&~op3)&(M4&T1);
fMWrite = fMWrite | (pla[15]&~op3)&(M4&T2);
ctl_alu_op1_oe = ctl_alu_op1_oe | (pla[15]&~op3)&(M4&T2);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[15]&~op3)&(M4&T2);
fMWrite = fMWrite | (pla[15]&~op3)&(M4&T3);
setM1 = setM1 | (pla[15]&~op3)&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (pla[15]&~op3)&(M4&T3);
ctl_alu_op_low = ctl_alu_op_low | (pla[15]&~op3)&(M4&T3);
ctl_alu_core_R = ctl_alu_core_R | (pla[15]&~op3)&(M4&T3);
ctl_alu_core_V = ctl_alu_core_V | (pla[15]&~op3)&(M4&T3);
ctl_alu_core_S = ctl_alu_core_S | (pla[15]&~op3)&(M4&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[15]&~op3)&(M4&T3);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[15]&~op3)&(M4&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[15]&~op3)&(M4&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[15]&~op3)&(M4&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[15]&~op3)&(M4&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[15]&~op3)&(M4&T3);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[15]&~op3)&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_pf_sel_nuse_ixiypla72npla55M1T1_10 = (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_nuse_ixiypla72npla55M1T1_10,ctl_pf_sel_nuse_ixiypla72npla55M1T1_10})&(`PFSEL_P);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[72]&~pla[55])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T2);
ctl_reg_gp_sel_nuse_ixiypla72npla55M1T2_2 = (~use_ixiy&pla[72]&~pla[55])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla72npla55M1T2_2,ctl_reg_gp_sel_nuse_ixiypla72npla55M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T2_3 = (~use_ixiy&pla[72]&~pla[55])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T2_3,ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[72]&~pla[55])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[72]&~pla[55])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (~use_ixiy&pla[72]&~pla[55])&(M1&T2);
ctl_reg_gp_sel_nuse_ixiypla72npla55M1T3_1 = (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla72npla55M1T3_1,ctl_reg_gp_sel_nuse_ixiypla72npla55M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T3_2 = (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T3_2,ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T3);
validPLA = validPLA | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
setM1 = setM1 | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_reg_gp_sel_nuse_ixiypla72npla55M1T4_3 = (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla72npla55M1T4_3,ctl_reg_gp_sel_nuse_ixiypla72npla55M1T4_3})&(op21);
ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T4_4 = (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T4_4,ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T4_4})&({~rsel0,rsel0});
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[72]&~pla[55])&(M1&T4)&(~rsel0);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[72]&~pla[55])&(M1&T4)&(rsel0);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[72]&~pla[55])&(M1&T4)&(~rsel0);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[72]&~pla[55])&(M1&T4)&(rsel0);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[72]&~pla[55])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[72]&~pla[55])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[72]&~pla[55])&(M4&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[72]&~pla[55])&(M4&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[72]&~pla[55])&(M4&T1);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[72]&~pla[55])&(M4&T1);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[72]&~pla[55])&(M4&T1);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[72]&~pla[55])&(M4&T1);
ctl_ir_we = ctl_ir_we | (~use_ixiy&pla[72]&~pla[55])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[72]&~pla[55])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[72]&~pla[55])&(M4&T3);
setM1 = setM1 | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[72]&~pla[55])&(M4&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[72]&~pla[55])&(M4&T4);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_pf_sel_nuse_ixiypla72pla55M1T1_10 = (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_nuse_ixiypla72pla55M1T1_10,ctl_pf_sel_nuse_ixiypla72pla55M1T1_10})&(`PFSEL_P);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[72]&pla[55])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (~use_ixiy&pla[72]&pla[55])&(M1&T2);
ctl_reg_gp_sel_nuse_ixiypla72pla55M1T2_2 = (~use_ixiy&pla[72]&pla[55])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla72pla55M1T2_2,ctl_reg_gp_sel_nuse_ixiypla72pla55M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla72pla55M1T2_3 = (~use_ixiy&pla[72]&pla[55])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla72pla55M1T2_3,ctl_reg_gp_hilo_nuse_ixiypla72pla55M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[72]&pla[55])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[72]&pla[55])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (~use_ixiy&pla[72]&pla[55])&(M1&T2);
ctl_reg_gp_sel_nuse_ixiypla72pla55M1T3_1 = (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla72pla55M1T3_1,ctl_reg_gp_sel_nuse_ixiypla72pla55M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla72pla55M1T3_2 = (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla72pla55M1T3_2,ctl_reg_gp_hilo_nuse_ixiypla72pla55M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[72]&pla[55])&(M1&T3);
validPLA = validPLA | (~use_ixiy&pla[72]&pla[55])&(M1&T4);
nextM = nextM | (~use_ixiy&pla[72]&pla[55])&(M1&T4);
ctl_mRead = ctl_mRead | (~use_ixiy&pla[72]&pla[55])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[72]&pla[55])&(M2&T1);
ctl_reg_gp_sel_nuse_ixiypla72pla55M2T1_2 = (~use_ixiy&pla[72]&pla[55])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla72pla55M2T1_2,ctl_reg_gp_sel_nuse_ixiypla72pla55M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_nuse_ixiypla72pla55M2T1_3 = (~use_ixiy&pla[72]&pla[55])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla72pla55M2T1_3,ctl_reg_gp_hilo_nuse_ixiypla72pla55M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[72]&pla[55])&(M2&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[72]&pla[55])&(M2&T1);
fMRead = fMRead | (~use_ixiy&pla[72]&pla[55])&(M2&T2);
fMRead = fMRead | (~use_ixiy&pla[72]&pla[55])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~use_ixiy&pla[72]&pla[55])&(M2&T3);
ctl_reg_sys_hilo_nuse_ixiypla72pla55M2T3_3 = (~use_ixiy&pla[72]&pla[55])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nuse_ixiypla72pla55M2T3_3,ctl_reg_sys_hilo_nuse_ixiypla72pla55M2T3_3})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (~use_ixiy&pla[72]&pla[55])&(M2&T3);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[72]&pla[55])&(M2&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[72]&pla[55])&(M2&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[72]&pla[55])&(M2&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[72]&pla[55])&(M2&T3);
setM1 = setM1 | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[72]&pla[55])&(M2&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[72]&pla[55])&(M2&T4);
fMRead = fMRead | (~use_ixiy&pla[72]&pla[55])&(M4&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~use_ixiy&pla[72]&pla[55])&(M4&T1);
ctl_reg_sys_hilo_nuse_ixiypla72pla55M4T1_3 = (~use_ixiy&pla[72]&pla[55])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nuse_ixiypla72pla55M4T1_3,ctl_reg_sys_hilo_nuse_ixiypla72pla55M4T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[72]&pla[55])&(M4&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[72]&pla[55])&(M4&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[72]&pla[55])&(M4&T1);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[72]&pla[55])&(M4&T1);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[72]&pla[55])&(M4&T1);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[72]&pla[55])&(M4&T1);
ctl_ir_we = ctl_ir_we | (~use_ixiy&pla[72]&pla[55])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[72]&pla[55])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[72]&pla[55])&(M4&T3);
setM1 = setM1 | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[72]&pla[55])&(M4&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (~use_ixiy&pla[72]&pla[55])&(M4&T4);
ctl_reg_gp_we = ctl_reg_gp_we | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_reg_gp_sel_nuse_ixiypla74npla55M1T1_2 = (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla74npla55M1T1_2,ctl_reg_gp_sel_nuse_ixiypla74npla55M1T1_2})&(op21);
ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T1_3 = (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T1_3,ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T1_3})&({~rsel0,rsel0});
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[74]&~pla[55])&(M1&T1);
ctl_reg_gp_sel_nuse_ixiypla74npla55M1T3_1 = (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla74npla55M1T3_1,ctl_reg_gp_sel_nuse_ixiypla74npla55M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T3_2 = (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T3_2,ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[74]&~pla[55])&(M1&T3);
validPLA = validPLA | (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
setM1 = setM1 | (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
ctl_reg_gp_sel_nuse_ixiypla74npla55M1T4_3 = (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla74npla55M1T4_3,ctl_reg_gp_sel_nuse_ixiypla74npla55M1T4_3})&(op21);
ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T4_4 = (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T4_4,ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T4_4})&({~rsel0,rsel0});
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[74]&~pla[55])&(M1&T4)&(~rsel0);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[74]&~pla[55])&(M1&T4)&(rsel0);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[74]&~pla[55])&(M1&T4)&(~rsel0);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[74]&~pla[55])&(M1&T4)&(rsel0);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[74]&~pla[55])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[74]&~pla[55])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[74]&~pla[55])&(M4&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~use_ixiy&pla[74]&~pla[55])&(M4&T1);
ctl_reg_sys_hilo_nuse_ixiypla74npla55M4T1_3 = (~use_ixiy&pla[74]&~pla[55])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nuse_ixiypla74npla55M4T1_3,ctl_reg_sys_hilo_nuse_ixiypla74npla55M4T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[74]&~pla[55])&(M4&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[74]&~pla[55])&(M4&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[74]&~pla[55])&(M4&T1);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[74]&~pla[55])&(M4&T1);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[74]&~pla[55])&(M4&T1);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[74]&~pla[55])&(M4&T1);
ctl_ir_we = ctl_ir_we | (~use_ixiy&pla[74]&~pla[55])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[74]&~pla[55])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
nextM = nextM | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[74]&~pla[55])&(M4&T3)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[74]&~pla[55])&(M4&T3);
fMWrite = fMWrite | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[74]&~pla[55])&(M5&T1);
fMWrite = fMWrite | (~use_ixiy&pla[74]&~pla[55])&(M5&T2);
fMWrite = fMWrite | (~use_ixiy&pla[74]&~pla[55])&(M5&T3);
setM1 = setM1 | (~use_ixiy&pla[74]&~pla[55])&(M5&T3);
ctl_reg_gp_sel_nuse_ixiypla74pla55M1T3_1 = (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla74pla55M1T3_1,ctl_reg_gp_sel_nuse_ixiypla74pla55M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla74pla55M1T3_2 = (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla74pla55M1T3_2,ctl_reg_gp_hilo_nuse_ixiypla74pla55M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[74]&pla[55])&(M1&T3);
validPLA = validPLA | (~use_ixiy&pla[74]&pla[55])&(M1&T4);
nextM = nextM | (~use_ixiy&pla[74]&pla[55])&(M1&T4);
ctl_mRead = ctl_mRead | (~use_ixiy&pla[74]&pla[55])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[74]&pla[55])&(M2&T1);
ctl_reg_gp_sel_nuse_ixiypla74pla55M2T1_2 = (~use_ixiy&pla[74]&pla[55])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla74pla55M2T1_2,ctl_reg_gp_sel_nuse_ixiypla74pla55M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_nuse_ixiypla74pla55M2T1_3 = (~use_ixiy&pla[74]&pla[55])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla74pla55M2T1_3,ctl_reg_gp_hilo_nuse_ixiypla74pla55M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[74]&pla[55])&(M2&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[74]&pla[55])&(M2&T1);
fMRead = fMRead | (~use_ixiy&pla[74]&pla[55])&(M2&T2);
fMRead = fMRead | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[74]&pla[55])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[74]&pla[55])&(M2&T3);
nextM = nextM | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[74]&pla[55])&(M2&T4);
fMWrite = fMWrite | (~use_ixiy&pla[74]&pla[55])&(M3&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[74]&pla[55])&(M3&T1);
fMWrite = fMWrite | (~use_ixiy&pla[74]&pla[55])&(M3&T2);
fMWrite = fMWrite | (~use_ixiy&pla[74]&pla[55])&(M3&T3);
setM1 = setM1 | (~use_ixiy&pla[74]&pla[55])&(M3&T3);
fMRead = fMRead | (~use_ixiy&pla[74]&pla[55])&(M4&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~use_ixiy&pla[74]&pla[55])&(M4&T1);
ctl_reg_sys_hilo_nuse_ixiypla74pla55M4T1_3 = (~use_ixiy&pla[74]&pla[55])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nuse_ixiypla74pla55M4T1_3,ctl_reg_sys_hilo_nuse_ixiypla74pla55M4T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[74]&pla[55])&(M4&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[74]&pla[55])&(M4&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[74]&pla[55])&(M4&T1);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[74]&pla[55])&(M4&T1);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[74]&pla[55])&(M4&T1);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[74]&pla[55])&(M4&T1);
ctl_ir_we = ctl_ir_we | (~use_ixiy&pla[74]&pla[55])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[74]&pla[55])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
nextM = nextM | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[74]&pla[55])&(M4&T3)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[74]&pla[55])&(M4&T3);
fMWrite = fMWrite | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_alu_core_R = ctl_alu_core_R | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_alu_core_V = ctl_alu_core_V | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (~use_ixiy&pla[74]&pla[55])&(M5&T1);
fMWrite = fMWrite | (~use_ixiy&pla[74]&pla[55])&(M5&T2);
fMWrite = fMWrite | (~use_ixiy&pla[74]&pla[55])&(M5&T3);
setM1 = setM1 | (~use_ixiy&pla[74]&pla[55])&(M5&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_reg_gp_sel_nuse_ixiypla73npla55M1T1_2 = (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla73npla55M1T1_2,ctl_reg_gp_sel_nuse_ixiypla73npla55M1T1_2})&(op21);
ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T1_3 = (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T1_3,ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T1_3})&({~rsel0,rsel0});
ctl_reg_in_hi = ctl_reg_in_hi | (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~use_ixiy&pla[73]&~pla[55])&(M1&T1);
ctl_reg_gp_sel_nuse_ixiypla73npla55M1T3_1 = (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla73npla55M1T3_1,ctl_reg_gp_sel_nuse_ixiypla73npla55M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T3_2 = (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T3_2,ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[73]&~pla[55])&(M1&T3);
validPLA = validPLA | (~use_ixiy&pla[73]&~pla[55])&(M1&T4);
setM1 = setM1 | (~use_ixiy&pla[73]&~pla[55])&(M1&T4);
ctl_reg_gp_sel_nuse_ixiypla73npla55M1T4_3 = (~use_ixiy&pla[73]&~pla[55])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla73npla55M1T4_3,ctl_reg_gp_sel_nuse_ixiypla73npla55M1T4_3})&(op21);
ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T4_4 = (~use_ixiy&pla[73]&~pla[55])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T4_4,ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T4_4})&({~rsel0,rsel0});
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[73]&~pla[55])&(M1&T4)&(~rsel0);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[73]&~pla[55])&(M1&T4)&(rsel0);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[73]&~pla[55])&(M1&T4)&(~rsel0);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[73]&~pla[55])&(M1&T4)&(rsel0);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[73]&~pla[55])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[73]&~pla[55])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[73]&~pla[55])&(M1&T4);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[73]&~pla[55])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[73]&~pla[55])&(M1&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~use_ixiy&pla[73]&~pla[55])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[73]&~pla[55])&(M4&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~use_ixiy&pla[73]&~pla[55])&(M4&T1);
ctl_reg_sys_hilo_nuse_ixiypla73npla55M4T1_3 = (~use_ixiy&pla[73]&~pla[55])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nuse_ixiypla73npla55M4T1_3,ctl_reg_sys_hilo_nuse_ixiypla73npla55M4T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[73]&~pla[55])&(M4&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[73]&~pla[55])&(M4&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[73]&~pla[55])&(M4&T1);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[73]&~pla[55])&(M4&T1);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[73]&~pla[55])&(M4&T1);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[73]&~pla[55])&(M4&T1);
ctl_ir_we = ctl_ir_we | (~use_ixiy&pla[73]&~pla[55])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[73]&~pla[55])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
nextM = nextM | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[73]&~pla[55])&(M4&T3)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~use_ixiy&pla[73]&~pla[55])&(M4&T3);
fMWrite = fMWrite | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~use_ixiy&pla[73]&~pla[55])&(M5&T1);
fMWrite = fMWrite | (~use_ixiy&pla[73]&~pla[55])&(M5&T2);
fMWrite = fMWrite | (~use_ixiy&pla[73]&~pla[55])&(M5&T3);
setM1 = setM1 | (~use_ixiy&pla[73]&~pla[55])&(M5&T3);
ctl_reg_gp_sel_nuse_ixiypla73pla55M1T3_1 = (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla73pla55M1T3_1,ctl_reg_gp_sel_nuse_ixiypla73pla55M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_nuse_ixiypla73pla55M1T3_2 = (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla73pla55M1T3_2,ctl_reg_gp_hilo_nuse_ixiypla73pla55M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (~use_ixiy&pla[73]&pla[55])&(M1&T3);
validPLA = validPLA | (~use_ixiy&pla[73]&pla[55])&(M1&T4);
nextM = nextM | (~use_ixiy&pla[73]&pla[55])&(M1&T4);
ctl_mRead = ctl_mRead | (~use_ixiy&pla[73]&pla[55])&(M1&T4);
fMRead = fMRead | (~use_ixiy&pla[73]&pla[55])&(M2&T1);
ctl_reg_gp_sel_nuse_ixiypla73pla55M2T1_2 = (~use_ixiy&pla[73]&pla[55])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_nuse_ixiypla73pla55M2T1_2,ctl_reg_gp_sel_nuse_ixiypla73pla55M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_nuse_ixiypla73pla55M2T1_3 = (~use_ixiy&pla[73]&pla[55])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_nuse_ixiypla73pla55M2T1_3,ctl_reg_gp_hilo_nuse_ixiypla73pla55M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[73]&pla[55])&(M2&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[73]&pla[55])&(M2&T1);
fMRead = fMRead | (~use_ixiy&pla[73]&pla[55])&(M2&T2);
fMRead = fMRead | (~use_ixiy&pla[73]&pla[55])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[73]&pla[55])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[73]&pla[55])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[73]&pla[55])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[73]&pla[55])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[73]&pla[55])&(M2&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[73]&pla[55])&(M2&T3);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[73]&pla[55])&(M2&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[73]&pla[55])&(M2&T3);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~use_ixiy&pla[73]&pla[55])&(M2&T3);
nextM = nextM | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~use_ixiy&pla[73]&pla[55])&(M2&T4);
fMWrite = fMWrite | (~use_ixiy&pla[73]&pla[55])&(M3&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[73]&pla[55])&(M3&T1);
fMWrite = fMWrite | (~use_ixiy&pla[73]&pla[55])&(M3&T2);
fMWrite = fMWrite | (~use_ixiy&pla[73]&pla[55])&(M3&T3);
setM1 = setM1 | (~use_ixiy&pla[73]&pla[55])&(M3&T3);
fMRead = fMRead | (~use_ixiy&pla[73]&pla[55])&(M4&T1);
ctl_reg_sel_wz = ctl_reg_sel_wz | (~use_ixiy&pla[73]&pla[55])&(M4&T1);
ctl_reg_sys_hilo_nuse_ixiypla73pla55M4T1_3 = (~use_ixiy&pla[73]&pla[55])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_nuse_ixiypla73pla55M4T1_3,ctl_reg_sys_hilo_nuse_ixiypla73pla55M4T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (~use_ixiy&pla[73]&pla[55])&(M4&T1);
ctl_al_we = ctl_al_we | (~use_ixiy&pla[73]&pla[55])&(M4&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[73]&pla[55])&(M4&T1);
ctl_alu_bs_oe = ctl_alu_bs_oe | (~use_ixiy&pla[73]&pla[55])&(M4&T1);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (~use_ixiy&pla[73]&pla[55])&(M4&T1);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[73]&pla[55])&(M4&T1);
ctl_ir_we = ctl_ir_we | (~use_ixiy&pla[73]&pla[55])&(M4&T1);
fMRead = fMRead | (~use_ixiy&pla[73]&pla[55])&(M4&T2);
fMRead = fMRead | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
nextM = nextM | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
ctl_mWrite = ctl_mWrite | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
ctl_flags_alu = ctl_flags_alu | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (~use_ixiy&pla[73]&pla[55])&(M4&T3)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
ctl_alu_op_low = ctl_alu_op_low | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~use_ixiy&pla[73]&pla[55])&(M4&T3);
fMWrite = fMWrite | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
ctl_sw_2u = ctl_sw_2u | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
ctl_alu_oe = ctl_alu_oe | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
ctl_alu_core_S = ctl_alu_core_S | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (~use_ixiy&pla[73]&pla[55])&(M5&T1);
fMWrite = fMWrite | (~use_ixiy&pla[73]&pla[55])&(M5&T2);
fMWrite = fMWrite | (~use_ixiy&pla[73]&pla[55])&(M5&T3);
setM1 = setM1 | (~use_ixiy&pla[73]&pla[55])&(M5&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[37]&~pla[28])&(M1&T1);
ctl_reg_gp_sel_pla37npla28M1T1_2 = (pla[37]&~pla[28])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla37npla28M1T1_2,ctl_reg_gp_sel_pla37npla28M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla37npla28M1T1_3 = (pla[37]&~pla[28])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla37npla28M1T1_3,ctl_reg_gp_hilo_pla37npla28M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[37]&~pla[28])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[37]&~pla[28])&(M1&T1);
ctl_sw_2d = ctl_sw_2d | (pla[37]&~pla[28])&(M1&T1);
ctl_sw_1d = ctl_sw_1d | (pla[37]&~pla[28])&(M1&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[37]&~pla[28])&(M1&T1);
validPLA = validPLA | (pla[37]&~pla[28])&(M1&T4);
nextM = nextM | (pla[37]&~pla[28])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[37]&~pla[28])&(M1&T4);
fMRead = fMRead | (pla[37]&~pla[28])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[37]&~pla[28])&(M2&T1);
ctl_reg_sys_hilo_pla37npla28M2T1_3 = (pla[37]&~pla[28])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla37npla28M2T1_3,ctl_reg_sys_hilo_pla37npla28M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[37]&~pla[28])&(M2&T1);
fMRead = fMRead | (pla[37]&~pla[28])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[37]&~pla[28])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[37]&~pla[28])&(M2&T2);
ctl_reg_sys_hilo_pla37npla28M2T2_4 = (pla[37]&~pla[28])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla37npla28M2T2_4,ctl_reg_sys_hilo_pla37npla28M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[37]&~pla[28])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[37]&~pla[28])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[37]&~pla[28])&(M2&T2);
fMRead = fMRead | (pla[37]&~pla[28])&(M2&T3);
nextM = nextM | (pla[37]&~pla[28])&(M2&T3);
ctl_iorw = ctl_iorw | (pla[37]&~pla[28])&(M2&T3);
fIORead = fIORead | (pla[37]&~pla[28])&(M3&T1);
ctl_reg_gp_sel_pla37npla28M3T1_2 = (pla[37]&~pla[28])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla37npla28M3T1_2,ctl_reg_gp_sel_pla37npla28M3T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla37npla28M3T1_3 = (pla[37]&~pla[28])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla37npla28M3T1_3,ctl_reg_gp_hilo_pla37npla28M3T1_3})&(2'b10);
ctl_sw_4d = ctl_sw_4d | (pla[37]&~pla[28])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[37]&~pla[28])&(M3&T1);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[37]&~pla[28])&(M3&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[37]&~pla[28])&(M3&T1);
ctl_sw_1d = ctl_sw_1d | (pla[37]&~pla[28])&(M3&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[37]&~pla[28])&(M3&T1);
fIORead = fIORead | (pla[37]&~pla[28])&(M3&T2);
fIORead = fIORead | (pla[37]&~pla[28])&(M3&T3);
fIORead = fIORead | (pla[37]&~pla[28])&(M3&T4);
setM1 = setM1 | (pla[37]&~pla[28])&(M3&T4);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[27]&~pla[34])&(M1&T1);
ctl_reg_gp_sel_pla27npla34M1T1_2 = (pla[27]&~pla[34])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla27npla34M1T1_2,ctl_reg_gp_sel_pla27npla34M1T1_2})&(op54);
ctl_reg_gp_hilo_pla27npla34M1T1_3 = (pla[27]&~pla[34])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla27npla34M1T1_3,ctl_reg_gp_hilo_pla27npla34M1T1_3})&({~rsel3,rsel3});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[27]&~pla[34])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[27]&~pla[34])&(M1&T1);
ctl_sw_2d = ctl_sw_2d | (pla[27]&~pla[34])&(M1&T1);
ctl_sw_1d = ctl_sw_1d | (pla[27]&~pla[34])&(M1&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[27]&~pla[34])&(M1&T1);
ctl_flags_alu = ctl_flags_alu | (pla[27]&~pla[34])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[27]&~pla[34])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[27]&~pla[34])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[27]&~pla[34])&(M1&T1);
ctl_alu_core_V = ctl_alu_core_V | (pla[27]&~pla[34])&(M1&T1);
ctl_alu_core_S = ctl_alu_core_S | (pla[27]&~pla[34])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[27]&~pla[34])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[27]&~pla[34])&(M1&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[27]&~pla[34])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[27]&~pla[34])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[27]&~pla[34])&(M1&T1);
ctl_pf_sel_pla27npla34M1T1_20 = (pla[27]&~pla[34])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla27npla34M1T1_20,ctl_pf_sel_pla27npla34M1T1_20})&(`PFSEL_P);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[27]&~pla[34])&(M1&T1);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[27]&~pla[34])&(M1&T1);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[27]&~pla[34])&(M1&T2);
ctl_reg_gp_sel_pla27npla34M1T2_2 = (pla[27]&~pla[34])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla27npla34M1T2_2,ctl_reg_gp_sel_pla27npla34M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla27npla34M1T2_3 = (pla[27]&~pla[34])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla27npla34M1T2_3,ctl_reg_gp_hilo_pla27npla34M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[27]&~pla[34])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[27]&~pla[34])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[27]&~pla[34])&(M1&T2);
ctl_reg_gp_sel_pla27npla34M1T3_1 = (pla[27]&~pla[34])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla27npla34M1T3_1,ctl_reg_gp_sel_pla27npla34M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla27npla34M1T3_2 = (pla[27]&~pla[34])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla27npla34M1T3_2,ctl_reg_gp_hilo_pla27npla34M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[27]&~pla[34])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[27]&~pla[34])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[27]&~pla[34])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[27]&~pla[34])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[27]&~pla[34])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[27]&~pla[34])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[27]&~pla[34])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[27]&~pla[34])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[27]&~pla[34])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[27]&~pla[34])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[27]&~pla[34])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[27]&~pla[34])&(M1&T3);
validPLA = validPLA | (pla[27]&~pla[34])&(M1&T4);
nextM = nextM | (pla[27]&~pla[34])&(M1&T4);
ctl_iorw = ctl_iorw | (pla[27]&~pla[34])&(M1&T4);
fIORead = fIORead | (pla[27]&~pla[34])&(M2&T1);
ctl_reg_gp_sel_pla27npla34M2T1_2 = (pla[27]&~pla[34])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla27npla34M2T1_2,ctl_reg_gp_sel_pla27npla34M2T1_2})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla27npla34M2T1_3 = (pla[27]&~pla[34])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla27npla34M2T1_3,ctl_reg_gp_hilo_pla27npla34M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[27]&~pla[34])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[27]&~pla[34])&(M2&T1);
fIORead = fIORead | (pla[27]&~pla[34])&(M2&T2);
fIORead = fIORead | (pla[27]&~pla[34])&(M2&T3);
fIORead = fIORead | (pla[27]&~pla[34])&(M2&T4);
setM1 = setM1 | (pla[27]&~pla[34])&(M2&T4);
ctl_sw_2d = ctl_sw_2d | (pla[27]&~pla[34])&(M2&T4);
ctl_sw_1d = ctl_sw_1d | (pla[27]&~pla[34])&(M2&T4);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[27]&~pla[34])&(M2&T4);
ctl_flags_alu = ctl_flags_alu | (pla[27]&~pla[34])&(M2&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[27]&~pla[34])&(M2&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[27]&~pla[34])&(M2&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[27]&~pla[34])&(M2&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[27]&~pla[34])&(M2&T4);
ctl_alu_core_R = ctl_alu_core_R | (pla[27]&~pla[34])&(M2&T4);
ctl_alu_core_V = ctl_alu_core_V | (pla[27]&~pla[34])&(M2&T4);
ctl_alu_core_S = ctl_alu_core_S | (pla[27]&~pla[34])&(M2&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[27]&~pla[34])&(M2&T4);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[27]&~pla[34])&(M2&T4);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[27]&~pla[34])&(M2&T4);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[27]&~pla[34])&(M2&T4);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[27]&~pla[34])&(M2&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[27]&~pla[34])&(M2&T4);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[27]&~pla[34])&(M2&T4);
validPLA = validPLA | (pla[37]&pla[28])&(M1&T4);
nextM = nextM | (pla[37]&pla[28])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[37]&pla[28])&(M1&T4);
fMRead = fMRead | (pla[37]&pla[28])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[37]&pla[28])&(M2&T1);
ctl_reg_sys_hilo_pla37pla28M2T1_3 = (pla[37]&pla[28])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla37pla28M2T1_3,ctl_reg_sys_hilo_pla37pla28M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[37]&pla[28])&(M2&T1);
fMRead = fMRead | (pla[37]&pla[28])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[37]&pla[28])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[37]&pla[28])&(M2&T2);
ctl_reg_sys_hilo_pla37pla28M2T2_4 = (pla[37]&pla[28])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla37pla28M2T2_4,ctl_reg_sys_hilo_pla37pla28M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[37]&pla[28])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[37]&pla[28])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[37]&pla[28])&(M2&T2);
fMRead = fMRead | (pla[37]&pla[28])&(M2&T3);
nextM = nextM | (pla[37]&pla[28])&(M2&T3);
ctl_iorw = ctl_iorw | (pla[37]&pla[28])&(M2&T3);
ctl_reg_gp_sel_pla37pla28M2T3_4 = (pla[37]&pla[28])&(M2&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla37pla28M2T3_4,ctl_reg_gp_sel_pla37pla28M2T3_4})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla37pla28M2T3_5 = (pla[37]&pla[28])&(M2&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla37pla28M2T3_5,ctl_reg_gp_hilo_pla37pla28M2T3_5})&(2'b10);
ctl_sw_4d = ctl_sw_4d | (pla[37]&pla[28])&(M2&T3);
ctl_al_we = ctl_al_we | (pla[37]&pla[28])&(M2&T3);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[37]&pla[28])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[37]&pla[28])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[37]&pla[28])&(M2&T3);
fIOWrite = fIOWrite | (pla[37]&pla[28])&(M3&T1);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[37]&pla[28])&(M3&T1);
ctl_reg_gp_sel_pla37pla28M3T1_3 = (pla[37]&pla[28])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla37pla28M3T1_3,ctl_reg_gp_sel_pla37pla28M3T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla37pla28M3T1_4 = (pla[37]&pla[28])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla37pla28M3T1_4,ctl_reg_gp_hilo_pla37pla28M3T1_4})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[37]&pla[28])&(M3&T1);
ctl_sw_2u = ctl_sw_2u | (pla[37]&pla[28])&(M3&T1);
ctl_sw_1u = ctl_sw_1u | (pla[37]&pla[28])&(M3&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[37]&pla[28])&(M3&T1);
fIOWrite = fIOWrite | (pla[37]&pla[28])&(M3&T2);
fIOWrite = fIOWrite | (pla[37]&pla[28])&(M3&T3);
fIOWrite = fIOWrite | (pla[37]&pla[28])&(M3&T4);
setM1 = setM1 | (pla[37]&pla[28])&(M3&T4);
validPLA = validPLA | (pla[27]&pla[34])&(M1&T4);
nextM = nextM | (pla[27]&pla[34])&(M1&T4);
ctl_iorw = ctl_iorw | (pla[27]&pla[34])&(M1&T4);
ctl_bus_zero_oe = ctl_bus_zero_oe | (pla[27]&pla[34])&(M1&T4)&(op4&op5&~op3);
ctl_reg_gp_sel_pla27pla34M1T4nop4op5nop3_1 = (pla[27]&pla[34])&(M1&T4)&(~(op4&op5&~op3));
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla27pla34M1T4nop4op5nop3_1,ctl_reg_gp_sel_pla27pla34M1T4nop4op5nop3_1})&(op54);
ctl_reg_gp_hilo_pla27pla34M1T4nop4op5nop3_2 = (pla[27]&pla[34])&(M1&T4)&(~(op4&op5&~op3));
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla27pla34M1T4nop4op5nop3_2,ctl_reg_gp_hilo_pla27pla34M1T4nop4op5nop3_2})&({~rsel3,rsel3});
ctl_reg_out_hi = ctl_reg_out_hi | (pla[27]&pla[34])&(M1&T4)&(~rsel3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[27]&pla[34])&(M1&T4)&(rsel3);
ctl_sw_2u = ctl_sw_2u | (pla[27]&pla[34])&(M1&T4)&(~rsel3);
ctl_sw_2d = ctl_sw_2d | (pla[27]&pla[34])&(M1&T4)&(rsel3);
ctl_sw_1u = ctl_sw_1u | (pla[27]&pla[34])&(M1&T4);
ctl_bus_db_we = ctl_bus_db_we | (pla[27]&pla[34])&(M1&T4);
fIOWrite = fIOWrite | (pla[27]&pla[34])&(M2&T1);
ctl_reg_gp_sel_pla27pla34M2T1_2 = (pla[27]&pla[34])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla27pla34M2T1_2,ctl_reg_gp_sel_pla27pla34M2T1_2})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla27pla34M2T1_3 = (pla[27]&pla[34])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla27pla34M2T1_3,ctl_reg_gp_hilo_pla27pla34M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[27]&pla[34])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[27]&pla[34])&(M2&T1);
fIOWrite = fIOWrite | (pla[27]&pla[34])&(M2&T2);
fIOWrite = fIOWrite | (pla[27]&pla[34])&(M2&T3);
fIOWrite = fIOWrite | (pla[27]&pla[34])&(M2&T4);
setM1 = setM1 | (pla[27]&pla[34])&(M2&T4);
ctl_alu_oe = ctl_alu_oe | (pla[91]&pla[21])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[91]&pla[21])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[91]&pla[21])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[91]&pla[21])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[91]&pla[21])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[91]&pla[21])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[91]&pla[21])&(M1&T1);
ctl_pf_sel_pla91pla21M1T1_8 = (pla[91]&pla[21])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla91pla21M1T1_8,ctl_pf_sel_pla91pla21M1T1_8})&(`PFSEL_P);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[91]&pla[21])&(M1&T2);
ctl_reg_gp_sel_pla91pla21M1T2_2 = (pla[91]&pla[21])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla21M1T2_2,ctl_reg_gp_sel_pla91pla21M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla91pla21M1T2_3 = (pla[91]&pla[21])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla21M1T2_3,ctl_reg_gp_hilo_pla91pla21M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[91]&pla[21])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[91]&pla[21])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[91]&pla[21])&(M1&T2);
ctl_reg_gp_sel_pla91pla21M1T3_1 = (pla[91]&pla[21])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla21M1T3_1,ctl_reg_gp_sel_pla91pla21M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla91pla21M1T3_2 = (pla[91]&pla[21])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla21M1T3_2,ctl_reg_gp_hilo_pla91pla21M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[91]&pla[21])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[91]&pla[21])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[91]&pla[21])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[91]&pla[21])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[91]&pla[21])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[91]&pla[21])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[91]&pla[21])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[91]&pla[21])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[91]&pla[21])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[91]&pla[21])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[91]&pla[21])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[91]&pla[21])&(M1&T3);
validPLA = validPLA | (pla[91]&pla[21])&(M1&T4);
nextM = nextM | (pla[91]&pla[21])&(M1&T5);
ctl_iorw = ctl_iorw | (pla[91]&pla[21])&(M1&T5);
fIORead = fIORead | (pla[91]&pla[21])&(M2&T1);
ctl_reg_gp_sel_pla91pla21M2T1_2 = (pla[91]&pla[21])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla21M2T1_2,ctl_reg_gp_sel_pla91pla21M2T1_2})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla91pla21M2T1_3 = (pla[91]&pla[21])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla21M2T1_3,ctl_reg_gp_hilo_pla91pla21M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[91]&pla[21])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[91]&pla[21])&(M2&T1);
fIORead = fIORead | (pla[91]&pla[21])&(M2&T2);
ctl_reg_gp_sel_pla91pla21M2T2_2 = (pla[91]&pla[21])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla21M2T2_2,ctl_reg_gp_sel_pla91pla21M2T2_2})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla91pla21M2T2_3 = (pla[91]&pla[21])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla21M2T2_3,ctl_reg_gp_hilo_pla91pla21M2T2_3})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[91]&pla[21])&(M2&T2);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[91]&pla[21])&(M2&T2);
ctl_flags_alu = ctl_flags_alu | (pla[91]&pla[21])&(M2&T2);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[91]&pla[21])&(M2&T2)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_zero = ctl_alu_op2_sel_zero | (pla[91]&pla[21])&(M2&T2);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[91]&pla[21])&(M2&T2);
ctl_alu_op_low = ctl_alu_op_low | (pla[91]&pla[21])&(M2&T2);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[91]&pla[21])&(M2&T2)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[91]&pla[21])&(M2&T2)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[91]&pla[21])&(M2&T2)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[91]&pla[21])&(M2&T2);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[91]&pla[21])&(M2&T2);
fIORead = fIORead | (pla[91]&pla[21])&(M2&T3);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[91]&pla[21])&(M2&T3);
ctl_reg_gp_sel_pla91pla21M2T3_3 = (pla[91]&pla[21])&(M2&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla21M2T3_3,ctl_reg_gp_sel_pla91pla21M2T3_3})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla91pla21M2T3_4 = (pla[91]&pla[21])&(M2&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla21M2T3_4,ctl_reg_gp_hilo_pla91pla21M2T3_4})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[91]&pla[21])&(M2&T3);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[91]&pla[21])&(M2&T3);
ctl_flags_alu = ctl_flags_alu | (pla[91]&pla[21])&(M2&T3);
ctl_alu_oe = ctl_alu_oe | (pla[91]&pla[21])&(M2&T3);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[91]&pla[21])&(M2&T3);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[91]&pla[21])&(M2&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[91]&pla[21])&(M2&T3)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[91]&pla[21])&(M2&T3)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[91]&pla[21])&(M2&T3)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[91]&pla[21])&(M2&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[91]&pla[21])&(M2&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[91]&pla[21])&(M2&T3);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[91]&pla[21])&(M2&T3);
fIORead = fIORead | (pla[91]&pla[21])&(M2&T4);
nextM = nextM | (pla[91]&pla[21])&(M2&T4);
ctl_mWrite = ctl_mWrite | (pla[91]&pla[21])&(M2&T4);
ctl_sw_2d = ctl_sw_2d | (pla[91]&pla[21])&(M2&T4);
ctl_sw_1d = ctl_sw_1d | (pla[91]&pla[21])&(M2&T4);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[91]&pla[21])&(M2&T4);
ctl_flags_alu = ctl_flags_alu | (pla[91]&pla[21])&(M2&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[91]&pla[21])&(M2&T4)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[91]&pla[21])&(M2&T4);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[91]&pla[21])&(M2&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[91]&pla[21])&(M2&T4);
fMWrite = fMWrite | (pla[91]&pla[21])&(M3&T1);
ctl_reg_gp_sel_pla91pla21M3T1_2 = (pla[91]&pla[21])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla21M3T1_2,ctl_reg_gp_sel_pla91pla21M3T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla91pla21M3T1_3 = (pla[91]&pla[21])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla21M3T1_3,ctl_reg_gp_hilo_pla91pla21M3T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[91]&pla[21])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[91]&pla[21])&(M3&T1);
fMWrite = fMWrite | (pla[91]&pla[21])&(M3&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[91]&pla[21])&(M3&T2);
ctl_reg_gp_sel_pla91pla21M3T2_3 = (pla[91]&pla[21])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla21M3T2_3,ctl_reg_gp_sel_pla91pla21M3T2_3})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla91pla21M3T2_4 = (pla[91]&pla[21])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla21M3T2_4,ctl_reg_gp_hilo_pla91pla21M3T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[91]&pla[21])&(M3&T2);
ctl_inc_cy = ctl_inc_cy | (pla[91]&pla[21])&(M3&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[91]&pla[21])&(M3&T2)&(op3);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[91]&pla[21])&(M3&T2);
fMWrite = fMWrite | (pla[91]&pla[21])&(M3&T3);
nextM = nextM | (pla[91]&pla[21])&(M3&T3);
setM1 = setM1 | (pla[91]&pla[21])&(M3&T3)&(nonRep|flags_zf);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[91]&pla[21])&(M4&T1);
ctl_reg_sys_hilo_pla91pla21M4T1_2 = (pla[91]&pla[21])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla91pla21M4T1_2,ctl_reg_sys_hilo_pla91pla21M4T1_2})&(2'b11);
ctl_al_we = ctl_al_we | (pla[91]&pla[21])&(M4&T1);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[91]&pla[21])&(M4&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[91]&pla[21])&(M4&T2);
ctl_reg_sys_hilo_pla91pla21M4T2_3 = (pla[91]&pla[21])&(M4&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla91pla21M4T2_3,ctl_reg_sys_hilo_pla91pla21M4T2_3})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[91]&pla[21])&(M4&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[91]&pla[21])&(M4&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[91]&pla[21])&(M4&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[91]&pla[21])&(M4&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[91]&pla[21])&(M4&T3);
ctl_reg_sys_hilo_pla91pla21M4T3_2 = (pla[91]&pla[21])&(M4&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla91pla21M4T3_2,ctl_reg_sys_hilo_pla91pla21M4T3_2})&(2'b11);
ctl_al_we = ctl_al_we | (pla[91]&pla[21])&(M4&T3);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[91]&pla[21])&(M4&T4);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[91]&pla[21])&(M4&T4);
ctl_reg_sys_hilo_pla91pla21M4T4_3 = (pla[91]&pla[21])&(M4&T4);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla91pla21M4T4_3,ctl_reg_sys_hilo_pla91pla21M4T4_3})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[91]&pla[21])&(M4&T4)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[91]&pla[21])&(M4&T4)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[91]&pla[21])&(M4&T4);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[91]&pla[21])&(M4&T4);
setM1 = setM1 | (pla[91]&pla[21])&(M4&T5);
ctl_flags_alu = ctl_flags_alu | (pla[91]&pla[20])&(M1&T1);
ctl_alu_oe = ctl_alu_oe | (pla[91]&pla[20])&(M1&T1);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[91]&pla[20])&(M1&T1);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[91]&pla[20])&(M1&T1);
ctl_alu_core_R = ctl_alu_core_R | (pla[91]&pla[20])&(M1&T1);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[91]&pla[20])&(M1&T1);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[91]&pla[20])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[91]&pla[20])&(M1&T1);
ctl_pf_sel_pla91pla20M1T1_9 = (pla[91]&pla[20])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla91pla20M1T1_9,ctl_pf_sel_pla91pla20M1T1_9})&(`PFSEL_P);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[91]&pla[20])&(M1&T2);
ctl_reg_gp_sel_pla91pla20M1T2_2 = (pla[91]&pla[20])&(M1&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla20M1T2_2,ctl_reg_gp_sel_pla91pla20M1T2_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla91pla20M1T2_3 = (pla[91]&pla[20])&(M1&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla20M1T2_3,ctl_reg_gp_hilo_pla91pla20M1T2_3})&(2'b01);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[91]&pla[20])&(M1&T2);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[91]&pla[20])&(M1&T2);
ctl_flags_oe = ctl_flags_oe | (pla[91]&pla[20])&(M1&T2);
ctl_reg_gp_sel_pla91pla20M1T3_1 = (pla[91]&pla[20])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla20M1T3_1,ctl_reg_gp_sel_pla91pla20M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla91pla20M1T3_2 = (pla[91]&pla[20])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla20M1T3_2,ctl_reg_gp_hilo_pla91pla20M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[91]&pla[20])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[91]&pla[20])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[91]&pla[20])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[91]&pla[20])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[91]&pla[20])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[91]&pla[20])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[91]&pla[20])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[91]&pla[20])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[91]&pla[20])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[91]&pla[20])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[91]&pla[20])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[91]&pla[20])&(M1&T3);
validPLA = validPLA | (pla[91]&pla[20])&(M1&T4);
ctl_reg_gp_sel_pla91pla20M1T4_2 = (pla[91]&pla[20])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla20M1T4_2,ctl_reg_gp_sel_pla91pla20M1T4_2})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla91pla20M1T4_3 = (pla[91]&pla[20])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla20M1T4_3,ctl_reg_gp_hilo_pla91pla20M1T4_3})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[91]&pla[20])&(M1&T4);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[91]&pla[20])&(M1&T4);
ctl_flags_alu = ctl_flags_alu | (pla[91]&pla[20])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[91]&pla[20])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_zero = ctl_alu_op2_sel_zero | (pla[91]&pla[20])&(M1&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[91]&pla[20])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[91]&pla[20])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[91]&pla[20])&(M1&T4)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[91]&pla[20])&(M1&T4)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[91]&pla[20])&(M1&T4)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[91]&pla[20])&(M1&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[91]&pla[20])&(M1&T4);
nextM = nextM | (pla[91]&pla[20])&(M1&T5);
ctl_mRead = ctl_mRead | (pla[91]&pla[20])&(M1&T5);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[91]&pla[20])&(M1&T5);
ctl_reg_gp_sel_pla91pla20M1T5_4 = (pla[91]&pla[20])&(M1&T5);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla20M1T5_4,ctl_reg_gp_sel_pla91pla20M1T5_4})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla91pla20M1T5_5 = (pla[91]&pla[20])&(M1&T5);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla20M1T5_5,ctl_reg_gp_hilo_pla91pla20M1T5_5})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[91]&pla[20])&(M1&T5);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[91]&pla[20])&(M1&T5);
ctl_flags_alu = ctl_flags_alu | (pla[91]&pla[20])&(M1&T5);
ctl_alu_oe = ctl_alu_oe | (pla[91]&pla[20])&(M1&T5);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[91]&pla[20])&(M1&T5);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[91]&pla[20])&(M1&T5);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[91]&pla[20])&(M1&T5)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[91]&pla[20])&(M1&T5)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[91]&pla[20])&(M1&T5)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[91]&pla[20])&(M1&T5);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[91]&pla[20])&(M1&T5);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[91]&pla[20])&(M1&T5);
fMRead = fMRead | (pla[91]&pla[20])&(M2&T1);
ctl_reg_gp_sel_pla91pla20M2T1_2 = (pla[91]&pla[20])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla20M2T1_2,ctl_reg_gp_sel_pla91pla20M2T1_2})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla91pla20M2T1_3 = (pla[91]&pla[20])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla20M2T1_3,ctl_reg_gp_hilo_pla91pla20M2T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[91]&pla[20])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[91]&pla[20])&(M2&T1);
fMRead = fMRead | (pla[91]&pla[20])&(M2&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[91]&pla[20])&(M2&T2);
ctl_reg_gp_sel_pla91pla20M2T2_3 = (pla[91]&pla[20])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla20M2T2_3,ctl_reg_gp_sel_pla91pla20M2T2_3})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla91pla20M2T2_4 = (pla[91]&pla[20])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla20M2T2_4,ctl_reg_gp_hilo_pla91pla20M2T2_4})&(2'b11);
ctl_sw_4u = ctl_sw_4u | (pla[91]&pla[20])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[91]&pla[20])&(M2&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[91]&pla[20])&(M2&T2)&(op3);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[91]&pla[20])&(M2&T2);
fMRead = fMRead | (pla[91]&pla[20])&(M2&T3);
nextM = nextM | (pla[91]&pla[20])&(M2&T3);
ctl_iorw = ctl_iorw | (pla[91]&pla[20])&(M2&T3);
ctl_reg_gp_sel_pla91pla20M2T3_4 = (pla[91]&pla[20])&(M2&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla20M2T3_4,ctl_reg_gp_sel_pla91pla20M2T3_4})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla91pla20M2T3_5 = (pla[91]&pla[20])&(M2&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla20M2T3_5,ctl_reg_gp_hilo_pla91pla20M2T3_5})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[91]&pla[20])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[91]&pla[20])&(M2&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[91]&pla[20])&(M2&T3)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[91]&pla[20])&(M2&T3);
fIOWrite = fIOWrite | (pla[91]&pla[20])&(M3&T1);
ctl_reg_gp_sel_pla91pla20M3T1_2 = (pla[91]&pla[20])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla91pla20M3T1_2,ctl_reg_gp_sel_pla91pla20M3T1_2})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla91pla20M3T1_3 = (pla[91]&pla[20])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla91pla20M3T1_3,ctl_reg_gp_hilo_pla91pla20M3T1_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[91]&pla[20])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[91]&pla[20])&(M3&T1);
fIOWrite = fIOWrite | (pla[91]&pla[20])&(M3&T2);
ctl_sw_2d = ctl_sw_2d | (pla[91]&pla[20])&(M3&T2);
ctl_sw_1d = ctl_sw_1d | (pla[91]&pla[20])&(M3&T2);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[91]&pla[20])&(M3&T2);
ctl_flags_alu = ctl_flags_alu | (pla[91]&pla[20])&(M3&T2);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[91]&pla[20])&(M3&T2)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[91]&pla[20])&(M3&T2);
ctl_alu_op_low = ctl_alu_op_low | (pla[91]&pla[20])&(M3&T2);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[91]&pla[20])&(M3&T2)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[91]&pla[20])&(M3&T2)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[91]&pla[20])&(M3&T2)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[91]&pla[20])&(M3&T2);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[91]&pla[20])&(M3&T2);
fIOWrite = fIOWrite | (pla[91]&pla[20])&(M3&T3);
ctl_flags_alu = ctl_flags_alu | (pla[91]&pla[20])&(M3&T3);
ctl_alu_oe = ctl_alu_oe | (pla[91]&pla[20])&(M3&T3);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[91]&pla[20])&(M3&T3);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[91]&pla[20])&(M3&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[91]&pla[20])&(M3&T3)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[91]&pla[20])&(M3&T3)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[91]&pla[20])&(M3&T3)&(~ctl_alu_op_low);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[91]&pla[20])&(M3&T3);
fIOWrite = fIOWrite | (pla[91]&pla[20])&(M3&T4);
nextM = nextM | (pla[91]&pla[20])&(M3&T4);
setM1 = setM1 | (pla[91]&pla[20])&(M3&T4)&(nonRep|flags_zf);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[91]&pla[20])&(M4&T1);
ctl_reg_sys_hilo_pla91pla20M4T1_2 = (pla[91]&pla[20])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla91pla20M4T1_2,ctl_reg_sys_hilo_pla91pla20M4T1_2})&(2'b11);
ctl_al_we = ctl_al_we | (pla[91]&pla[20])&(M4&T1);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[91]&pla[20])&(M4&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[91]&pla[20])&(M4&T2);
ctl_reg_sys_hilo_pla91pla20M4T2_3 = (pla[91]&pla[20])&(M4&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla91pla20M4T2_3,ctl_reg_sys_hilo_pla91pla20M4T2_3})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[91]&pla[20])&(M4&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[91]&pla[20])&(M4&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[91]&pla[20])&(M4&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[91]&pla[20])&(M4&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[91]&pla[20])&(M4&T3);
ctl_reg_sys_hilo_pla91pla20M4T3_2 = (pla[91]&pla[20])&(M4&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla91pla20M4T3_2,ctl_reg_sys_hilo_pla91pla20M4T3_2})&(2'b11);
ctl_al_we = ctl_al_we | (pla[91]&pla[20])&(M4&T3);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[91]&pla[20])&(M4&T4);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[91]&pla[20])&(M4&T4);
ctl_reg_sys_hilo_pla91pla20M4T4_3 = (pla[91]&pla[20])&(M4&T4);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla91pla20M4T4_3,ctl_reg_sys_hilo_pla91pla20M4T4_3})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[91]&pla[20])&(M4&T4)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[91]&pla[20])&(M4&T4)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[91]&pla[20])&(M4&T4);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[91]&pla[20])&(M4&T4);
setM1 = setM1 | (pla[91]&pla[20])&(M4&T5);
validPLA = validPLA | (pla[29])&(M1&T4);
nextM = nextM | (pla[29])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[29])&(M1&T4);
fMRead = fMRead | (pla[29])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[29])&(M2&T1);
ctl_reg_sys_hilo_pla29M2T1_3 = (pla[29])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla29M2T1_3,ctl_reg_sys_hilo_pla29M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[29])&(M2&T1);
fMRead = fMRead | (pla[29])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[29])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[29])&(M2&T2);
ctl_reg_sys_hilo_pla29M2T2_4 = (pla[29])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla29M2T2_4,ctl_reg_sys_hilo_pla29M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[29])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[29])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[29])&(M2&T2);
fMRead = fMRead | (pla[29])&(M2&T3);
nextM = nextM | (pla[29])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[29])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[29])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[29])&(M2&T3);
ctl_reg_sys_hilo_pla29M2T3_6 = (pla[29])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla29M2T3_6,ctl_reg_sys_hilo_pla29M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[29])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[29])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[29])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[29])&(M2&T3);
fMRead = fMRead | (pla[29])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[29])&(M3&T1);
ctl_reg_sys_hilo_pla29M3T1_3 = (pla[29])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla29M3T1_3,ctl_reg_sys_hilo_pla29M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[29])&(M3&T1);
fMRead = fMRead | (pla[29])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[29])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[29])&(M3&T2);
ctl_reg_sys_hilo_pla29M3T2_4 = (pla[29])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla29M3T2_4,ctl_reg_sys_hilo_pla29M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[29])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[29])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[29])&(M3&T2);
fMRead = fMRead | (pla[29])&(M3&T3);
setM1 = setM1 | (pla[29])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[29])&(M3&T3);
ctl_reg_sys_hilo_pla29M3T3_4 = (pla[29])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla29M3T3_4,ctl_reg_sys_hilo_pla29M3T3_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[29])&(M3&T3);
ctl_al_we = ctl_al_we | (pla[29])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[29])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[29])&(M3&T3);
ctl_reg_sys_hilo_pla29M3T3_9 = (pla[29])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla29M3T3_9,ctl_reg_sys_hilo_pla29M3T3_9})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[29])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[29])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[29])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[29])&(M3&T3);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[29])&(M3&T3);
ctl_reg_gp_sel_pla43M1T3_1 = (pla[43])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla43M1T3_1,ctl_reg_gp_sel_pla43M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla43M1T3_2 = (pla[43])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla43M1T3_2,ctl_reg_gp_hilo_pla43M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[43])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[43])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[43])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[43])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[43])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[43])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[43])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[43])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[43])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[43])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[43])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[43])&(M1&T3);
validPLA = validPLA | (pla[43])&(M1&T4);
nextM = nextM | (pla[43])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[43])&(M1&T4);
fMRead = fMRead | (pla[43])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[43])&(M2&T1);
ctl_reg_sys_hilo_pla43M2T1_3 = (pla[43])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla43M2T1_3,ctl_reg_sys_hilo_pla43M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[43])&(M2&T1);
fMRead = fMRead | (pla[43])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[43])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[43])&(M2&T2);
ctl_reg_sys_hilo_pla43M2T2_4 = (pla[43])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla43M2T2_4,ctl_reg_sys_hilo_pla43M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[43])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[43])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[43])&(M2&T2);
fMRead = fMRead | (pla[43])&(M2&T3);
nextM = nextM | (pla[43])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[43])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[43])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[43])&(M2&T3);
ctl_reg_sys_hilo_pla43M2T3_6 = (pla[43])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla43M2T3_6,ctl_reg_sys_hilo_pla43M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[43])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[43])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[43])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[43])&(M2&T3);
fMRead = fMRead | (pla[43])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[43])&(M3&T1);
ctl_reg_sys_hilo_pla43M3T1_3 = (pla[43])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla43M3T1_3,ctl_reg_sys_hilo_pla43M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[43])&(M3&T1);
fMRead = fMRead | (pla[43])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[43])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[43])&(M3&T2);
ctl_reg_sys_hilo_pla43M3T2_4 = (pla[43])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla43M3T2_4,ctl_reg_sys_hilo_pla43M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[43])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[43])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[43])&(M3&T2);
fMRead = fMRead | (pla[43])&(M3&T3);
setM1 = setM1 | (pla[43])&(M3&T3);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[43])&(M3&T3)&(flags_cond_true);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[43])&(M3&T3)&(flags_cond_true);
ctl_reg_sys_hilo_pla43M3T3_5 = (pla[43])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla43M3T3_5,ctl_reg_sys_hilo_pla43M3T3_5})&({flags_cond_true,flags_cond_true});
ctl_sw_4d = ctl_sw_4d | (pla[43])&(M3&T3)&(flags_cond_true);
ctl_al_we = ctl_al_we | (pla[43])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[43])&(M3&T3)&(flags_cond_true);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[43])&(M3&T3)&(flags_cond_true);
ctl_reg_sys_hilo_pla43M3T3_10 = (pla[43])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla43M3T3_10,ctl_reg_sys_hilo_pla43M3T3_10})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[43])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[43])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[43])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[43])&(M3&T3);
ctl_reg_gp_sel_pla47M1T3_1 = (pla[47])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla47M1T3_1,ctl_reg_gp_sel_pla47M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla47M1T3_2 = (pla[47])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla47M1T3_2,ctl_reg_gp_hilo_pla47M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[47])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[47])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[47])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[47])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[47])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[47])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[47])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[47])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[47])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[47])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[47])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[47])&(M1&T3);
validPLA = validPLA | (pla[47])&(M1&T4);
nextM = nextM | (pla[47])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[47])&(M1&T4);
fMRead = fMRead | (pla[47])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[47])&(M2&T1);
ctl_reg_sys_hilo_pla47M2T1_3 = (pla[47])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla47M2T1_3,ctl_reg_sys_hilo_pla47M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[47])&(M2&T1);
fMRead = fMRead | (pla[47])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[47])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[47])&(M2&T2);
ctl_reg_sys_hilo_pla47M2T2_4 = (pla[47])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla47M2T2_4,ctl_reg_sys_hilo_pla47M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[47])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[47])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[47])&(M2&T2);
fMRead = fMRead | (pla[47])&(M2&T3);
nextM = nextM | (pla[47])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[47])&(M3&T1);
ctl_sw_1d = ctl_sw_1d | (pla[47])&(M3&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[47])&(M3&T1);
ctl_flags_alu = ctl_flags_alu | (pla[47])&(M3&T1);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[47])&(M3&T1)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[47])&(M3&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[47])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[47])&(M3&T2);
ctl_reg_sys_hilo_pla47M3T2_2 = (pla[47])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla47M3T2_2,ctl_reg_sys_hilo_pla47M3T2_2})&(2'b01);
ctl_sw_4u = ctl_sw_4u | (pla[47])&(M3&T2);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[47])&(M3&T2);
ctl_sw_2d = ctl_sw_2d | (pla[47])&(M3&T2);
ctl_flags_alu = ctl_flags_alu | (pla[47])&(M3&T2);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[47])&(M3&T2)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[47])&(M3&T2);
ctl_alu_op_low = ctl_alu_op_low | (pla[47])&(M3&T2);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[47])&(M3&T2)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[47])&(M3&T2)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[47])&(M3&T2)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[47])&(M3&T2);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[47])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[47])&(M3&T3);
ctl_reg_sys_hilo_pla47M3T3_3 = (pla[47])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla47M3T3_3,ctl_reg_sys_hilo_pla47M3T3_3})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[47])&(M3&T3);
ctl_sw_2u = ctl_sw_2u | (pla[47])&(M3&T3);
ctl_flags_alu = ctl_flags_alu | (pla[47])&(M3&T3);
ctl_alu_oe = ctl_alu_oe | (pla[47])&(M3&T3);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[47])&(M3&T3);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[47])&(M3&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[47])&(M3&T3)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[47])&(M3&T3)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[47])&(M3&T3)&(~ctl_alu_op_low);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[47])&(M3&T3);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[47])&(M3&T4);
ctl_reg_sys_hilo_pla47M3T4_2 = (pla[47])&(M3&T4);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla47M3T4_2,ctl_reg_sys_hilo_pla47M3T4_2})&(2'b10);
ctl_sw_4u = ctl_sw_4u | (pla[47])&(M3&T4);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[47])&(M3&T4);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[47])&(M3&T4);
ctl_flags_alu = ctl_flags_alu | (pla[47])&(M3&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[47])&(M3&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_zero = ctl_alu_op2_sel_zero | (pla[47])&(M3&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[47])&(M3&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[47])&(M3&T4);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[47])&(M3&T4)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[47])&(M3&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[47])&(M3&T4)&(flags_sf);
setM1 = setM1 | (pla[47])&(M3&T5);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[47])&(M3&T5);
ctl_reg_sys_hilo_pla47M3T5_3 = (pla[47])&(M3&T5);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla47M3T5_3,ctl_reg_sys_hilo_pla47M3T5_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[47])&(M3&T5);
ctl_al_we = ctl_al_we | (pla[47])&(M3&T5);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[47])&(M3&T5);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[47])&(M3&T5);
ctl_reg_sys_hilo_pla47M3T5_8 = (pla[47])&(M3&T5);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla47M3T5_8,ctl_reg_sys_hilo_pla47M3T5_8})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[47])&(M3&T5);
ctl_flags_alu = ctl_flags_alu | (pla[47])&(M3&T5);
ctl_alu_oe = ctl_alu_oe | (pla[47])&(M3&T5);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[47])&(M3&T5);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[47])&(M3&T5);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[47])&(M3&T5)&(~ctl_alu_op_low);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[47])&(M3&T5)&(flags_sf);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[47])&(M3&T5);
ctl_reg_gp_sel_pla48M1T3_1 = (pla[48])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla48M1T3_1,ctl_reg_gp_sel_pla48M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla48M1T3_2 = (pla[48])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla48M1T3_2,ctl_reg_gp_hilo_pla48M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[48])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[48])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[48])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[48])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[48])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[48])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[48])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[48])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[48])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[48])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[48])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[48])&(M1&T3);
validPLA = validPLA | (pla[48])&(M1&T4);
nextM = nextM | (pla[48])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[48])&(M1&T4);
ctl_cond_short = ctl_cond_short | (pla[48])&(M1&T4);
fMRead = fMRead | (pla[48])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[48])&(M2&T1);
ctl_reg_sys_hilo_pla48M2T1_3 = (pla[48])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla48M2T1_3,ctl_reg_sys_hilo_pla48M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[48])&(M2&T1);
fMRead = fMRead | (pla[48])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[48])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[48])&(M2&T2);
ctl_reg_sys_hilo_pla48M2T2_4 = (pla[48])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla48M2T2_4,ctl_reg_sys_hilo_pla48M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[48])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[48])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[48])&(M2&T2);
fMRead = fMRead | (pla[48])&(M2&T3);
nextM = nextM | (pla[48])&(M2&T3);
setM1 = setM1 | (pla[48])&(M2&T3)&(~flags_cond_true);
ctl_sw_2d = ctl_sw_2d | (pla[48])&(M3&T1);
ctl_sw_1d = ctl_sw_1d | (pla[48])&(M3&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[48])&(M3&T1);
ctl_flags_alu = ctl_flags_alu | (pla[48])&(M3&T1);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[48])&(M3&T1)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[48])&(M3&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[48])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[48])&(M3&T2);
ctl_reg_sys_hilo_pla48M3T2_2 = (pla[48])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla48M3T2_2,ctl_reg_sys_hilo_pla48M3T2_2})&(2'b01);
ctl_sw_4u = ctl_sw_4u | (pla[48])&(M3&T2);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[48])&(M3&T2);
ctl_sw_2d = ctl_sw_2d | (pla[48])&(M3&T2);
ctl_flags_alu = ctl_flags_alu | (pla[48])&(M3&T2);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[48])&(M3&T2)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[48])&(M3&T2);
ctl_alu_op_low = ctl_alu_op_low | (pla[48])&(M3&T2);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[48])&(M3&T2)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[48])&(M3&T2)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[48])&(M3&T2)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[48])&(M3&T2);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[48])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[48])&(M3&T3);
ctl_reg_sys_hilo_pla48M3T3_3 = (pla[48])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla48M3T3_3,ctl_reg_sys_hilo_pla48M3T3_3})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[48])&(M3&T3);
ctl_sw_2u = ctl_sw_2u | (pla[48])&(M3&T3);
ctl_flags_alu = ctl_flags_alu | (pla[48])&(M3&T3);
ctl_alu_oe = ctl_alu_oe | (pla[48])&(M3&T3);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[48])&(M3&T3);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[48])&(M3&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[48])&(M3&T3)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[48])&(M3&T3)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[48])&(M3&T3)&(~ctl_alu_op_low);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[48])&(M3&T3);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[48])&(M3&T4);
ctl_reg_sys_hilo_pla48M3T4_2 = (pla[48])&(M3&T4);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla48M3T4_2,ctl_reg_sys_hilo_pla48M3T4_2})&(2'b10);
ctl_sw_4u = ctl_sw_4u | (pla[48])&(M3&T4);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[48])&(M3&T4);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[48])&(M3&T4);
ctl_flags_alu = ctl_flags_alu | (pla[48])&(M3&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[48])&(M3&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_zero = ctl_alu_op2_sel_zero | (pla[48])&(M3&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[48])&(M3&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[48])&(M3&T4);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[48])&(M3&T4)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[48])&(M3&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[48])&(M3&T4)&(flags_sf);
setM1 = setM1 | (pla[48])&(M3&T5);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[48])&(M3&T5);
ctl_reg_sys_hilo_pla48M3T5_3 = (pla[48])&(M3&T5);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla48M3T5_3,ctl_reg_sys_hilo_pla48M3T5_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[48])&(M3&T5);
ctl_al_we = ctl_al_we | (pla[48])&(M3&T5);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[48])&(M3&T5);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[48])&(M3&T5);
ctl_reg_sys_hilo_pla48M3T5_8 = (pla[48])&(M3&T5);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla48M3T5_8,ctl_reg_sys_hilo_pla48M3T5_8})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[48])&(M3&T5);
ctl_flags_alu = ctl_flags_alu | (pla[48])&(M3&T5);
ctl_alu_oe = ctl_alu_oe | (pla[48])&(M3&T5);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[48])&(M3&T5);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[48])&(M3&T5);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[48])&(M3&T5)&(~ctl_alu_op_low);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[48])&(M3&T5)&(flags_sf);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[48])&(M3&T5);
validPLA = validPLA | (pla[6])&(M1&T4);
setM1 = setM1 | (pla[6])&(M1&T4);
ctl_reg_gp_sel_pla6M1T4_3 = (pla[6])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla6M1T4_3,ctl_reg_gp_sel_pla6M1T4_3})&(`GP_REG_HL);
ctl_reg_gp_hilo_pla6M1T4_4 = (pla[6])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla6M1T4_4,ctl_reg_gp_hilo_pla6M1T4_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[6])&(M1&T4);
ctl_al_we = ctl_al_we | (pla[6])&(M1&T4);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[6])&(M1&T4);
ctl_reg_gp_sel_pla26M1T3_1 = (pla[26])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla26M1T3_1,ctl_reg_gp_sel_pla26M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla26M1T3_2 = (pla[26])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla26M1T3_2,ctl_reg_gp_hilo_pla26M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[26])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[26])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[26])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[26])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[26])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[26])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[26])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[26])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[26])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[26])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[26])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[26])&(M1&T3);
validPLA = validPLA | (pla[26])&(M1&T4);
ctl_reg_gp_sel_pla26M1T4_2 = (pla[26])&(M1&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla26M1T4_2,ctl_reg_gp_sel_pla26M1T4_2})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla26M1T4_3 = (pla[26])&(M1&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla26M1T4_3,ctl_reg_gp_hilo_pla26M1T4_3})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[26])&(M1&T4);
ctl_flags_alu = ctl_flags_alu | (pla[26])&(M1&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[26])&(M1&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_zero = ctl_alu_op2_sel_zero | (pla[26])&(M1&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[26])&(M1&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[26])&(M1&T4);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[26])&(M1&T4)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[26])&(M1&T4)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[26])&(M1&T4)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[26])&(M1&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[26])&(M1&T4);
nextM = nextM | (pla[26])&(M1&T5);
ctl_mRead = ctl_mRead | (pla[26])&(M1&T5);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[26])&(M1&T5);
ctl_reg_gp_sel_pla26M1T5_4 = (pla[26])&(M1&T5);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla26M1T5_4,ctl_reg_gp_sel_pla26M1T5_4})&(`GP_REG_BC);
ctl_reg_gp_hilo_pla26M1T5_5 = (pla[26])&(M1&T5);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla26M1T5_5,ctl_reg_gp_hilo_pla26M1T5_5})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[26])&(M1&T5);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[26])&(M1&T5);
ctl_flags_alu = ctl_flags_alu | (pla[26])&(M1&T5);
ctl_alu_oe = ctl_alu_oe | (pla[26])&(M1&T5);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[26])&(M1&T5);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[26])&(M1&T5);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[26])&(M1&T5)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[26])&(M1&T5)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[26])&(M1&T5)&(~ctl_alu_op_low);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[26])&(M1&T5);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[26])&(M1&T5);
fMRead = fMRead | (pla[26])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[26])&(M2&T1);
ctl_reg_sys_hilo_pla26M2T1_3 = (pla[26])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla26M2T1_3,ctl_reg_sys_hilo_pla26M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[26])&(M2&T1);
fMRead = fMRead | (pla[26])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[26])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[26])&(M2&T2);
ctl_reg_sys_hilo_pla26M2T2_4 = (pla[26])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla26M2T2_4,ctl_reg_sys_hilo_pla26M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[26])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[26])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[26])&(M2&T2);
fMRead = fMRead | (pla[26])&(M2&T3);
nextM = nextM | (pla[26])&(M2&T3);
setM1 = setM1 | (pla[26])&(M2&T3)&(flags_zf);
ctl_sw_2d = ctl_sw_2d | (pla[26])&(M3&T1);
ctl_sw_1d = ctl_sw_1d | (pla[26])&(M3&T1);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[26])&(M3&T1);
ctl_flags_alu = ctl_flags_alu | (pla[26])&(M3&T1);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[26])&(M3&T1)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[26])&(M3&T1);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[26])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[26])&(M3&T2);
ctl_reg_sys_hilo_pla26M3T2_2 = (pla[26])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla26M3T2_2,ctl_reg_sys_hilo_pla26M3T2_2})&(2'b01);
ctl_sw_4u = ctl_sw_4u | (pla[26])&(M3&T2);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[26])&(M3&T2);
ctl_sw_2d = ctl_sw_2d | (pla[26])&(M3&T2);
ctl_flags_alu = ctl_flags_alu | (pla[26])&(M3&T2);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[26])&(M3&T2)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[26])&(M3&T2);
ctl_alu_op_low = ctl_alu_op_low | (pla[26])&(M3&T2);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[26])&(M3&T2)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[26])&(M3&T2)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[26])&(M3&T2)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[26])&(M3&T2);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[26])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[26])&(M3&T3);
ctl_reg_sys_hilo_pla26M3T3_3 = (pla[26])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla26M3T3_3,ctl_reg_sys_hilo_pla26M3T3_3})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[26])&(M3&T3);
ctl_sw_2u = ctl_sw_2u | (pla[26])&(M3&T3);
ctl_flags_alu = ctl_flags_alu | (pla[26])&(M3&T3);
ctl_alu_oe = ctl_alu_oe | (pla[26])&(M3&T3);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[26])&(M3&T3);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[26])&(M3&T3);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[26])&(M3&T3)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[26])&(M3&T3)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[26])&(M3&T3)&(~ctl_alu_op_low);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[26])&(M3&T3);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[26])&(M3&T4);
ctl_reg_sys_hilo_pla26M3T4_2 = (pla[26])&(M3&T4);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla26M3T4_2,ctl_reg_sys_hilo_pla26M3T4_2})&(2'b10);
ctl_sw_4u = ctl_sw_4u | (pla[26])&(M3&T4);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[26])&(M3&T4);
ctl_flags_alu = ctl_flags_alu | (pla[26])&(M3&T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[26])&(M3&T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_zero = ctl_alu_op2_sel_zero | (pla[26])&(M3&T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[26])&(M3&T4);
ctl_alu_op_low = ctl_alu_op_low | (pla[26])&(M3&T4);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[26])&(M3&T4)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[26])&(M3&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[26])&(M3&T4)&(flags_sf);
setM1 = setM1 | (pla[26])&(M3&T5);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[26])&(M3&T5);
ctl_reg_sys_hilo_pla26M3T5_3 = (pla[26])&(M3&T5);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla26M3T5_3,ctl_reg_sys_hilo_pla26M3T5_3})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[26])&(M3&T5);
ctl_al_we = ctl_al_we | (pla[26])&(M3&T5);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[26])&(M3&T5);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[26])&(M3&T5);
ctl_reg_sys_hilo_pla26M3T5_8 = (pla[26])&(M3&T5);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla26M3T5_8,ctl_reg_sys_hilo_pla26M3T5_8})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[26])&(M3&T5);
ctl_flags_alu = ctl_flags_alu | (pla[26])&(M3&T5);
ctl_alu_oe = ctl_alu_oe | (pla[26])&(M3&T5);
ctl_alu_res_oe = ctl_alu_res_oe | (pla[26])&(M3&T5);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (pla[26])&(M3&T5);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[26])&(M3&T5)&(~ctl_alu_op_low);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[26])&(M3&T5)&(flags_sf);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[26])&(M3&T5);
validPLA = validPLA | (pla[24])&(M1&T4);
nextM = nextM | (pla[24])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[24])&(M1&T4);
fMRead = fMRead | (pla[24])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[24])&(M2&T1);
ctl_reg_sys_hilo_pla24M2T1_3 = (pla[24])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla24M2T1_3,ctl_reg_sys_hilo_pla24M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[24])&(M2&T1);
fMRead = fMRead | (pla[24])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[24])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[24])&(M2&T2);
ctl_reg_sys_hilo_pla24M2T2_4 = (pla[24])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla24M2T2_4,ctl_reg_sys_hilo_pla24M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[24])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[24])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[24])&(M2&T2);
fMRead = fMRead | (pla[24])&(M2&T3);
nextM = nextM | (pla[24])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[24])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[24])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[24])&(M2&T3);
ctl_reg_sys_hilo_pla24M2T3_6 = (pla[24])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla24M2T3_6,ctl_reg_sys_hilo_pla24M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[24])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[24])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[24])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[24])&(M2&T3);
fMRead = fMRead | (pla[24])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[24])&(M3&T1);
ctl_reg_sys_hilo_pla24M3T1_3 = (pla[24])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla24M3T1_3,ctl_reg_sys_hilo_pla24M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[24])&(M3&T1);
fMRead = fMRead | (pla[24])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[24])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[24])&(M3&T2);
ctl_reg_sys_hilo_pla24M3T2_4 = (pla[24])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla24M3T2_4,ctl_reg_sys_hilo_pla24M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[24])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[24])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[24])&(M3&T2);
fMRead = fMRead | (pla[24])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[24])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[24])&(M3&T3);
ctl_reg_sys_hilo_pla24M3T3_4 = (pla[24])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla24M3T3_4,ctl_reg_sys_hilo_pla24M3T3_4})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[24])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[24])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[24])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[24])&(M3&T3);
nextM = nextM | (pla[24])&(M3&T4);
ctl_mWrite = ctl_mWrite | (pla[24])&(M3&T4);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[24])&(M3&T4);
ctl_reg_gp_sel_pla24M3T4_4 = (pla[24])&(M3&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla24M3T4_4,ctl_reg_gp_sel_pla24M3T4_4})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla24M3T4_5 = (pla[24])&(M3&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla24M3T4_5,ctl_reg_gp_hilo_pla24M3T4_5})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[24])&(M3&T4);
ctl_inc_cy = ctl_inc_cy | (pla[24])&(M3&T4)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[24])&(M3&T4);
ctl_al_we = ctl_al_we | (pla[24])&(M3&T4);
fMWrite = fMWrite | (pla[24])&(M4&T1);
ctl_inc_cy = ctl_inc_cy | (pla[24])&(M4&T1)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[24])&(M4&T1);
ctl_apin_mux = ctl_apin_mux | (pla[24])&(M4&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[24])&(M4&T1);
ctl_reg_sys_hilo_pla24M4T1_6 = (pla[24])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla24M4T1_6,ctl_reg_sys_hilo_pla24M4T1_6})&(2'b10);
ctl_sw_4u = ctl_sw_4u | (pla[24])&(M4&T1);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[24])&(M4&T1);
ctl_sw_2u = ctl_sw_2u | (pla[24])&(M4&T1);
ctl_sw_1u = ctl_sw_1u | (pla[24])&(M4&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[24])&(M4&T1);
fMWrite = fMWrite | (pla[24])&(M4&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[24])&(M4&T2);
ctl_reg_gp_sel_pla24M4T2_3 = (pla[24])&(M4&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla24M4T2_3,ctl_reg_gp_sel_pla24M4T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla24M4T2_4 = (pla[24])&(M4&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla24M4T2_4,ctl_reg_gp_hilo_pla24M4T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[24])&(M4&T2);
ctl_sw_4u = ctl_sw_4u | (pla[24])&(M4&T2);
ctl_inc_cy = ctl_inc_cy | (pla[24])&(M4&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[24])&(M4&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[24])&(M4&T2);
fMWrite = fMWrite | (pla[24])&(M4&T3);
nextM = nextM | (pla[24])&(M4&T3);
ctl_mWrite = ctl_mWrite | (pla[24])&(M4&T3);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[24])&(M4&T3);
ctl_reg_gp_sel_pla24M4T3_5 = (pla[24])&(M4&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla24M4T3_5,ctl_reg_gp_sel_pla24M4T3_5})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla24M4T3_6 = (pla[24])&(M4&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla24M4T3_6,ctl_reg_gp_hilo_pla24M4T3_6})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[24])&(M4&T3);
ctl_inc_cy = ctl_inc_cy | (pla[24])&(M4&T3)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[24])&(M4&T3);
ctl_al_we = ctl_al_we | (pla[24])&(M4&T3);
fMWrite = fMWrite | (pla[24])&(M5&T1);
ctl_inc_cy = ctl_inc_cy | (pla[24])&(M5&T1)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[24])&(M5&T1);
ctl_apin_mux = ctl_apin_mux | (pla[24])&(M5&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[24])&(M5&T1);
ctl_reg_sys_hilo_pla24M5T1_6 = (pla[24])&(M5&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla24M5T1_6,ctl_reg_sys_hilo_pla24M5T1_6})&(2'b01);
ctl_sw_4u = ctl_sw_4u | (pla[24])&(M5&T1);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[24])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (pla[24])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[24])&(M5&T1);
fMWrite = fMWrite | (pla[24])&(M5&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[24])&(M5&T2);
ctl_reg_gp_sel_pla24M5T2_3 = (pla[24])&(M5&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla24M5T2_3,ctl_reg_gp_sel_pla24M5T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla24M5T2_4 = (pla[24])&(M5&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla24M5T2_4,ctl_reg_gp_hilo_pla24M5T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[24])&(M5&T2);
ctl_sw_4u = ctl_sw_4u | (pla[24])&(M5&T2);
ctl_inc_cy = ctl_inc_cy | (pla[24])&(M5&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[24])&(M5&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[24])&(M5&T2);
fMWrite = fMWrite | (pla[24])&(M5&T3);
setM1 = setM1 | (pla[24])&(M5&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[24])&(M5&T3);
ctl_reg_sys_hilo_pla24M5T3_4 = (pla[24])&(M5&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla24M5T3_4,ctl_reg_sys_hilo_pla24M5T3_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[24])&(M5&T3);
ctl_al_we = ctl_al_we | (pla[24])&(M5&T3);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[24])&(M5&T3);
ctl_reg_gp_sel_pla42M1T3_1 = (pla[42])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla42M1T3_1,ctl_reg_gp_sel_pla42M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla42M1T3_2 = (pla[42])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla42M1T3_2,ctl_reg_gp_hilo_pla42M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[42])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[42])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[42])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[42])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[42])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[42])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[42])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[42])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[42])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[42])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[42])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[42])&(M1&T3);
validPLA = validPLA | (pla[42])&(M1&T4);
nextM = nextM | (pla[42])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[42])&(M1&T4);
fMRead = fMRead | (pla[42])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[42])&(M2&T1);
ctl_reg_sys_hilo_pla42M2T1_3 = (pla[42])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla42M2T1_3,ctl_reg_sys_hilo_pla42M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[42])&(M2&T1);
fMRead = fMRead | (pla[42])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[42])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[42])&(M2&T2);
ctl_reg_sys_hilo_pla42M2T2_4 = (pla[42])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla42M2T2_4,ctl_reg_sys_hilo_pla42M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[42])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[42])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[42])&(M2&T2);
fMRead = fMRead | (pla[42])&(M2&T3);
nextM = nextM | (pla[42])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[42])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[42])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[42])&(M2&T3);
ctl_reg_sys_hilo_pla42M2T3_6 = (pla[42])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla42M2T3_6,ctl_reg_sys_hilo_pla42M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[42])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[42])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[42])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[42])&(M2&T3);
fMRead = fMRead | (pla[42])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[42])&(M3&T1);
ctl_reg_sys_hilo_pla42M3T1_3 = (pla[42])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla42M3T1_3,ctl_reg_sys_hilo_pla42M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[42])&(M3&T1);
fMRead = fMRead | (pla[42])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[42])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[42])&(M3&T2);
ctl_reg_sys_hilo_pla42M3T2_4 = (pla[42])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla42M3T2_4,ctl_reg_sys_hilo_pla42M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[42])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[42])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[42])&(M3&T2);
fMRead = fMRead | (pla[42])&(M3&T3);
nextM = nextM | (pla[42])&(M3&T3)&(~flags_cond_true);
setM1 = setM1 | (pla[42])&(M3&T3)&(~flags_cond_true);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[42])&(M3&T3)&(flags_cond_true);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[42])&(M3&T3)&(flags_cond_true);
ctl_reg_sys_hilo_pla42M3T3_6 = (pla[42])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla42M3T3_6,ctl_reg_sys_hilo_pla42M3T3_6})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[42])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[42])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[42])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[42])&(M3&T3);
nextM = nextM | (pla[42])&(M3&T4);
ctl_mWrite = ctl_mWrite | (pla[42])&(M3&T4);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[42])&(M3&T4);
ctl_reg_gp_sel_pla42M3T4_4 = (pla[42])&(M3&T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla42M3T4_4,ctl_reg_gp_sel_pla42M3T4_4})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla42M3T4_5 = (pla[42])&(M3&T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla42M3T4_5,ctl_reg_gp_hilo_pla42M3T4_5})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[42])&(M3&T4);
ctl_inc_cy = ctl_inc_cy | (pla[42])&(M3&T4)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[42])&(M3&T4);
ctl_al_we = ctl_al_we | (pla[42])&(M3&T4);
fMWrite = fMWrite | (pla[42])&(M4&T1);
ctl_inc_cy = ctl_inc_cy | (pla[42])&(M4&T1)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[42])&(M4&T1);
ctl_apin_mux = ctl_apin_mux | (pla[42])&(M4&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[42])&(M4&T1);
ctl_reg_sys_hilo_pla42M4T1_6 = (pla[42])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla42M4T1_6,ctl_reg_sys_hilo_pla42M4T1_6})&(2'b10);
ctl_sw_4u = ctl_sw_4u | (pla[42])&(M4&T1);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[42])&(M4&T1);
ctl_sw_2u = ctl_sw_2u | (pla[42])&(M4&T1);
ctl_sw_1u = ctl_sw_1u | (pla[42])&(M4&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[42])&(M4&T1);
fMWrite = fMWrite | (pla[42])&(M4&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[42])&(M4&T2);
ctl_reg_gp_sel_pla42M4T2_3 = (pla[42])&(M4&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla42M4T2_3,ctl_reg_gp_sel_pla42M4T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla42M4T2_4 = (pla[42])&(M4&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla42M4T2_4,ctl_reg_gp_hilo_pla42M4T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[42])&(M4&T2);
ctl_sw_4u = ctl_sw_4u | (pla[42])&(M4&T2);
ctl_inc_cy = ctl_inc_cy | (pla[42])&(M4&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[42])&(M4&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[42])&(M4&T2);
fMWrite = fMWrite | (pla[42])&(M4&T3);
nextM = nextM | (pla[42])&(M4&T3);
ctl_mWrite = ctl_mWrite | (pla[42])&(M4&T3);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[42])&(M4&T3);
ctl_reg_gp_sel_pla42M4T3_5 = (pla[42])&(M4&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla42M4T3_5,ctl_reg_gp_sel_pla42M4T3_5})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla42M4T3_6 = (pla[42])&(M4&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla42M4T3_6,ctl_reg_gp_hilo_pla42M4T3_6})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[42])&(M4&T3);
ctl_inc_cy = ctl_inc_cy | (pla[42])&(M4&T3)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[42])&(M4&T3);
ctl_al_we = ctl_al_we | (pla[42])&(M4&T3);
fMWrite = fMWrite | (pla[42])&(M5&T1);
ctl_inc_cy = ctl_inc_cy | (pla[42])&(M5&T1)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[42])&(M5&T1);
ctl_apin_mux = ctl_apin_mux | (pla[42])&(M5&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[42])&(M5&T1);
ctl_reg_sys_hilo_pla42M5T1_6 = (pla[42])&(M5&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla42M5T1_6,ctl_reg_sys_hilo_pla42M5T1_6})&(2'b01);
ctl_sw_4u = ctl_sw_4u | (pla[42])&(M5&T1);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[42])&(M5&T1);
ctl_sw_1u = ctl_sw_1u | (pla[42])&(M5&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[42])&(M5&T1);
fMWrite = fMWrite | (pla[42])&(M5&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[42])&(M5&T2);
ctl_reg_gp_sel_pla42M5T2_3 = (pla[42])&(M5&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla42M5T2_3,ctl_reg_gp_sel_pla42M5T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla42M5T2_4 = (pla[42])&(M5&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla42M5T2_4,ctl_reg_gp_hilo_pla42M5T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[42])&(M5&T2);
ctl_sw_4u = ctl_sw_4u | (pla[42])&(M5&T2);
ctl_inc_cy = ctl_inc_cy | (pla[42])&(M5&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[42])&(M5&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[42])&(M5&T2);
fMWrite = fMWrite | (pla[42])&(M5&T3);
setM1 = setM1 | (pla[42])&(M5&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[42])&(M5&T3);
ctl_reg_sys_hilo_pla42M5T3_4 = (pla[42])&(M5&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla42M5T3_4,ctl_reg_sys_hilo_pla42M5T3_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[42])&(M5&T3);
ctl_al_we = ctl_al_we | (pla[42])&(M5&T3);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[42])&(M5&T3);
validPLA = validPLA | (pla[35])&(M1&T4);
nextM = nextM | (pla[35])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[35])&(M1&T4);
fMRead = fMRead | (pla[35])&(M2&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[35])&(M2&T1);
ctl_reg_gp_sel_pla35M2T1_3 = (pla[35])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla35M2T1_3,ctl_reg_gp_sel_pla35M2T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla35M2T1_4 = (pla[35])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla35M2T1_4,ctl_reg_gp_hilo_pla35M2T1_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[35])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[35])&(M2&T1);
fMRead = fMRead | (pla[35])&(M2&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[35])&(M2&T2);
ctl_reg_gp_sel_pla35M2T2_3 = (pla[35])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla35M2T2_3,ctl_reg_gp_sel_pla35M2T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla35M2T2_4 = (pla[35])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla35M2T2_4,ctl_reg_gp_hilo_pla35M2T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[35])&(M2&T2);
ctl_sw_4u = ctl_sw_4u | (pla[35])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[35])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[35])&(M2&T2);
fMRead = fMRead | (pla[35])&(M2&T3);
nextM = nextM | (pla[35])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[35])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[35])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[35])&(M2&T3);
ctl_reg_sys_hilo_pla35M2T3_6 = (pla[35])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla35M2T3_6,ctl_reg_sys_hilo_pla35M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[35])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[35])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[35])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[35])&(M2&T3);
fMRead = fMRead | (pla[35])&(M3&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[35])&(M3&T1);
ctl_reg_gp_sel_pla35M3T1_3 = (pla[35])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla35M3T1_3,ctl_reg_gp_sel_pla35M3T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla35M3T1_4 = (pla[35])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla35M3T1_4,ctl_reg_gp_hilo_pla35M3T1_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[35])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[35])&(M3&T1);
fMRead = fMRead | (pla[35])&(M3&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[35])&(M3&T2);
ctl_reg_gp_sel_pla35M3T2_3 = (pla[35])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla35M3T2_3,ctl_reg_gp_sel_pla35M3T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla35M3T2_4 = (pla[35])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla35M3T2_4,ctl_reg_gp_hilo_pla35M3T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[35])&(M3&T2);
ctl_sw_4u = ctl_sw_4u | (pla[35])&(M3&T2);
ctl_inc_cy = ctl_inc_cy | (pla[35])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[35])&(M3&T2);
fMRead = fMRead | (pla[35])&(M3&T3);
setM1 = setM1 | (pla[35])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[35])&(M3&T3);
ctl_reg_sys_hilo_pla35M3T3_4 = (pla[35])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla35M3T3_4,ctl_reg_sys_hilo_pla35M3T3_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[35])&(M3&T3);
ctl_al_we = ctl_al_we | (pla[35])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[35])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[35])&(M3&T3);
ctl_reg_sys_hilo_pla35M3T3_9 = (pla[35])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla35M3T3_9,ctl_reg_sys_hilo_pla35M3T3_9})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[35])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[35])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[35])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[35])&(M3&T3);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[35])&(M3&T3);
ctl_reg_gp_sel_pla45M1T3_1 = (pla[45])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla45M1T3_1,ctl_reg_gp_sel_pla45M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla45M1T3_2 = (pla[45])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla45M1T3_2,ctl_reg_gp_hilo_pla45M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[45])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[45])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[45])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[45])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[45])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[45])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[45])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[45])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[45])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[45])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[45])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[45])&(M1&T3);
validPLA = validPLA | (pla[45])&(M1&T4);
nextM = nextM | (pla[45])&(M1&T5);
ctl_mRead = ctl_mRead | (pla[45])&(M1&T5);
setM1 = setM1 | (pla[45])&(M1&T5)&(~flags_cond_true);
fMRead = fMRead | (pla[45])&(M2&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[45])&(M2&T1);
ctl_reg_gp_sel_pla45M2T1_3 = (pla[45])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla45M2T1_3,ctl_reg_gp_sel_pla45M2T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla45M2T1_4 = (pla[45])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla45M2T1_4,ctl_reg_gp_hilo_pla45M2T1_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[45])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[45])&(M2&T1);
fMRead = fMRead | (pla[45])&(M2&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[45])&(M2&T2);
ctl_reg_gp_sel_pla45M2T2_3 = (pla[45])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla45M2T2_3,ctl_reg_gp_sel_pla45M2T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla45M2T2_4 = (pla[45])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla45M2T2_4,ctl_reg_gp_hilo_pla45M2T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[45])&(M2&T2);
ctl_sw_4u = ctl_sw_4u | (pla[45])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[45])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[45])&(M2&T2);
fMRead = fMRead | (pla[45])&(M2&T3);
nextM = nextM | (pla[45])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[45])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[45])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[45])&(M2&T3);
ctl_reg_sys_hilo_pla45M2T3_6 = (pla[45])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla45M2T3_6,ctl_reg_sys_hilo_pla45M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[45])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[45])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[45])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[45])&(M2&T3);
fMRead = fMRead | (pla[45])&(M3&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[45])&(M3&T1);
ctl_reg_gp_sel_pla45M3T1_3 = (pla[45])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla45M3T1_3,ctl_reg_gp_sel_pla45M3T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla45M3T1_4 = (pla[45])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla45M3T1_4,ctl_reg_gp_hilo_pla45M3T1_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[45])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[45])&(M3&T1);
fMRead = fMRead | (pla[45])&(M3&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[45])&(M3&T2);
ctl_reg_gp_sel_pla45M3T2_3 = (pla[45])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla45M3T2_3,ctl_reg_gp_sel_pla45M3T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla45M3T2_4 = (pla[45])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla45M3T2_4,ctl_reg_gp_hilo_pla45M3T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[45])&(M3&T2);
ctl_sw_4u = ctl_sw_4u | (pla[45])&(M3&T2);
ctl_inc_cy = ctl_inc_cy | (pla[45])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[45])&(M3&T2);
fMRead = fMRead | (pla[45])&(M3&T3);
setM1 = setM1 | (pla[45])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[45])&(M3&T3);
ctl_reg_sys_hilo_pla45M3T3_4 = (pla[45])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla45M3T3_4,ctl_reg_sys_hilo_pla45M3T3_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[45])&(M3&T3);
ctl_al_we = ctl_al_we | (pla[45])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[45])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[45])&(M3&T3);
ctl_reg_sys_hilo_pla45M3T3_9 = (pla[45])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla45M3T3_9,ctl_reg_sys_hilo_pla45M3T3_9})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[45])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[45])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[45])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[45])&(M3&T3);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[45])&(M3&T3);
validPLA = validPLA | (pla[46])&(M1&T4);
nextM = nextM | (pla[46])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[46])&(M1&T4);
ctl_iff1_iff2 = ctl_iff1_iff2 | (pla[46])&(M1&T4);
fMRead = fMRead | (pla[46])&(M2&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[46])&(M2&T1);
ctl_reg_gp_sel_pla46M2T1_3 = (pla[46])&(M2&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla46M2T1_3,ctl_reg_gp_sel_pla46M2T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla46M2T1_4 = (pla[46])&(M2&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla46M2T1_4,ctl_reg_gp_hilo_pla46M2T1_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[46])&(M2&T1);
ctl_al_we = ctl_al_we | (pla[46])&(M2&T1);
fMRead = fMRead | (pla[46])&(M2&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[46])&(M2&T2);
ctl_reg_gp_sel_pla46M2T2_3 = (pla[46])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla46M2T2_3,ctl_reg_gp_sel_pla46M2T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla46M2T2_4 = (pla[46])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla46M2T2_4,ctl_reg_gp_hilo_pla46M2T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[46])&(M2&T2);
ctl_sw_4u = ctl_sw_4u | (pla[46])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[46])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[46])&(M2&T2);
fMRead = fMRead | (pla[46])&(M2&T3);
nextM = nextM | (pla[46])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[46])&(M2&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[46])&(M2&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[46])&(M2&T3);
ctl_reg_sys_hilo_pla46M2T3_6 = (pla[46])&(M2&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla46M2T3_6,ctl_reg_sys_hilo_pla46M2T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[46])&(M2&T3);
ctl_sw_2d = ctl_sw_2d | (pla[46])&(M2&T3);
ctl_sw_1d = ctl_sw_1d | (pla[46])&(M2&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[46])&(M2&T3);
fMRead = fMRead | (pla[46])&(M3&T1);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[46])&(M3&T1);
ctl_reg_gp_sel_pla46M3T1_3 = (pla[46])&(M3&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla46M3T1_3,ctl_reg_gp_sel_pla46M3T1_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla46M3T1_4 = (pla[46])&(M3&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla46M3T1_4,ctl_reg_gp_hilo_pla46M3T1_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[46])&(M3&T1);
ctl_al_we = ctl_al_we | (pla[46])&(M3&T1);
fMRead = fMRead | (pla[46])&(M3&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[46])&(M3&T2);
ctl_reg_gp_sel_pla46M3T2_3 = (pla[46])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla46M3T2_3,ctl_reg_gp_sel_pla46M3T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla46M3T2_4 = (pla[46])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla46M3T2_4,ctl_reg_gp_hilo_pla46M3T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[46])&(M3&T2);
ctl_sw_4u = ctl_sw_4u | (pla[46])&(M3&T2);
ctl_inc_cy = ctl_inc_cy | (pla[46])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[46])&(M3&T2);
fMRead = fMRead | (pla[46])&(M3&T3);
setM1 = setM1 | (pla[46])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[46])&(M3&T3);
ctl_reg_sys_hilo_pla46M3T3_4 = (pla[46])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla46M3T3_4,ctl_reg_sys_hilo_pla46M3T3_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[46])&(M3&T3);
ctl_al_we = ctl_al_we | (pla[46])&(M3&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[46])&(M3&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[46])&(M3&T3);
ctl_reg_sys_hilo_pla46M3T3_9 = (pla[46])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla46M3T3_9,ctl_reg_sys_hilo_pla46M3T3_9})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[46])&(M3&T3);
ctl_sw_2d = ctl_sw_2d | (pla[46])&(M3&T3);
ctl_sw_1d = ctl_sw_1d | (pla[46])&(M3&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[46])&(M3&T3);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[46])&(M3&T3);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[56])&(M1&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[56])&(M1&T3);
ctl_reg_sys_hilo_pla56M1T3_3 = (pla[56])&(M1&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla56M1T3_3,ctl_reg_sys_hilo_pla56M1T3_3})&(2'b11);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[56])&(M1&T3);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[56])&(M1&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[56])&(M1&T3);
ctl_alu_oe = ctl_alu_oe | (pla[56])&(M1&T3);
ctl_alu_op1_oe = ctl_alu_op1_oe | (pla[56])&(M1&T3);
ctl_alu_op1_sel_zero = ctl_alu_op1_sel_zero | (pla[56])&(M1&T3);
ctl_sw_mask543_en = ctl_sw_mask543_en | (pla[56])&(M1&T3)&(~((in_intr&im2)|in_nmi));
ctl_sw_1d = ctl_sw_1d | (pla[56])&(M1&T3)&(~in_nmi);
ctl_66_oe = ctl_66_oe | (pla[56])&(M1&T3)&(in_nmi);
ctl_bus_ff_oe = ctl_bus_ff_oe | (pla[56])&(M1&T3)&(in_intr&im1);
validPLA = validPLA | (pla[56])&(M1&T4);
nextM = nextM | (pla[56])&(M1&T5);
ctl_mWrite = ctl_mWrite | (pla[56])&(M1&T5);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[56])&(M1&T5);
ctl_reg_gp_sel_pla56M1T5_4 = (pla[56])&(M1&T5);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla56M1T5_4,ctl_reg_gp_sel_pla56M1T5_4})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla56M1T5_5 = (pla[56])&(M1&T5);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla56M1T5_5,ctl_reg_gp_hilo_pla56M1T5_5})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[56])&(M1&T5);
ctl_inc_cy = ctl_inc_cy | (pla[56])&(M1&T5)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[56])&(M1&T5);
ctl_al_we = ctl_al_we | (pla[56])&(M1&T5);
ctl_sw_2d = ctl_sw_2d | (pla[56])&(M1&T5);
ctl_sw_1d = ctl_sw_1d | (pla[56])&(M1&T5);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[56])&(M1&T5);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[56])&(M1&T5)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[56])&(M1&T5);
fMWrite = fMWrite | (pla[56])&(M2&T1);
ctl_inc_cy = ctl_inc_cy | (pla[56])&(M2&T1)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[56])&(M2&T1);
ctl_apin_mux = ctl_apin_mux | (pla[56])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[56])&(M2&T1);
ctl_reg_sys_hilo_pla56M2T1_6 = (pla[56])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla56M2T1_6,ctl_reg_sys_hilo_pla56M2T1_6})&(2'b10);
ctl_sw_4u = ctl_sw_4u | (pla[56])&(M2&T1);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[56])&(M2&T1);
ctl_sw_2u = ctl_sw_2u | (pla[56])&(M2&T1);
ctl_sw_1u = ctl_sw_1u | (pla[56])&(M2&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[56])&(M2&T1);
fMWrite = fMWrite | (pla[56])&(M2&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[56])&(M2&T2);
ctl_reg_gp_sel_pla56M2T2_3 = (pla[56])&(M2&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla56M2T2_3,ctl_reg_gp_sel_pla56M2T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla56M2T2_4 = (pla[56])&(M2&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla56M2T2_4,ctl_reg_gp_hilo_pla56M2T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[56])&(M2&T2);
ctl_sw_4u = ctl_sw_4u | (pla[56])&(M2&T2);
ctl_inc_cy = ctl_inc_cy | (pla[56])&(M2&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[56])&(M2&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[56])&(M2&T2);
fMWrite = fMWrite | (pla[56])&(M2&T3);
nextM = nextM | (pla[56])&(M2&T3);
ctl_mWrite = ctl_mWrite | (pla[56])&(M2&T3);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[56])&(M2&T3);
ctl_reg_gp_sel_pla56M2T3_5 = (pla[56])&(M2&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla56M2T3_5,ctl_reg_gp_sel_pla56M2T3_5})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla56M2T3_6 = (pla[56])&(M2&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla56M2T3_6,ctl_reg_gp_hilo_pla56M2T3_6})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[56])&(M2&T3);
ctl_inc_cy = ctl_inc_cy | (pla[56])&(M2&T3)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[56])&(M2&T3);
ctl_al_we = ctl_al_we | (pla[56])&(M2&T3);
fMWrite = fMWrite | (pla[56])&(M3&T1);
ctl_inc_cy = ctl_inc_cy | (pla[56])&(M3&T1)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[56])&(M3&T1);
ctl_apin_mux = ctl_apin_mux | (pla[56])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[56])&(M3&T1);
ctl_reg_sys_hilo_pla56M3T1_6 = (pla[56])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla56M3T1_6,ctl_reg_sys_hilo_pla56M3T1_6})&(2'b01);
ctl_sw_4u = ctl_sw_4u | (pla[56])&(M3&T1);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[56])&(M3&T1);
ctl_sw_1u = ctl_sw_1u | (pla[56])&(M3&T1);
ctl_bus_db_we = ctl_bus_db_we | (pla[56])&(M3&T1);
fMWrite = fMWrite | (pla[56])&(M3&T2);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[56])&(M3&T2);
ctl_reg_gp_sel_pla56M3T2_3 = (pla[56])&(M3&T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla56M3T2_3,ctl_reg_gp_sel_pla56M3T2_3})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla56M3T2_4 = (pla[56])&(M3&T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla56M3T2_4,ctl_reg_gp_hilo_pla56M3T2_4})&(2'b11);
ctl_reg_use_sp = ctl_reg_use_sp | (pla[56])&(M3&T2);
ctl_sw_4u = ctl_sw_4u | (pla[56])&(M3&T2);
ctl_inc_cy = ctl_inc_cy | (pla[56])&(M3&T2)&(~pc_inc_hold);
ctl_inc_dec = ctl_inc_dec | (pla[56])&(M3&T2);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[56])&(M3&T2);
fMWrite = fMWrite | (pla[56])&(M3&T3);
nextM = nextM | (pla[56])&(M3&T3);
ctl_mRead = ctl_mRead | (pla[56])&(M3&T3)&(in_intr&im2);
setM1 = setM1 | (pla[56])&(M3&T3)&(~(in_intr&im2));
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[56])&(M3&T3);
ctl_reg_sys_hilo_pla56M3T3_6 = (pla[56])&(M3&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla56M3T3_6,ctl_reg_sys_hilo_pla56M3T3_6})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[56])&(M3&T3);
ctl_al_we = ctl_al_we | (pla[56])&(M3&T3);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[56])&(M3&T3);
fMRead = fMRead | (pla[56])&(M4&T1);
ctl_reg_sel_ir = ctl_reg_sel_ir | (pla[56])&(M4&T1);
ctl_reg_sys_hilo_pla56M4T1_3 = (pla[56])&(M4&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla56M4T1_3,ctl_reg_sys_hilo_pla56M4T1_3})&(2'b10);
ctl_sw_4d = ctl_sw_4d | (pla[56])&(M4&T1);
ctl_al_we = ctl_al_we | (pla[56])&(M4&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[56])&(M4&T1);
ctl_sw_2u = ctl_sw_2u | (pla[56])&(M4&T1);
ctl_alu_oe = ctl_alu_oe | (pla[56])&(M4&T1);
ctl_alu_op1_oe = ctl_alu_op1_oe | (pla[56])&(M4&T1);
fMRead = fMRead | (pla[56])&(M4&T2);
ctl_sw_4u = ctl_sw_4u | (pla[56])&(M4&T2);
ctl_inc_cy = ctl_inc_cy | (pla[56])&(M4&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[56])&(M4&T2);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[56])&(M4&T2);
ctl_sw_2d = ctl_sw_2d | (pla[56])&(M4&T2);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[56])&(M4&T2)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[56])&(M4&T2);
fMRead = fMRead | (pla[56])&(M4&T3);
nextM = nextM | (pla[56])&(M4&T3);
ctl_mRead = ctl_mRead | (pla[56])&(M4&T3);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (pla[56])&(M4&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[56])&(M4&T3);
ctl_reg_sys_hilo_pla56M4T3_6 = (pla[56])&(M4&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla56M4T3_6,ctl_reg_sys_hilo_pla56M4T3_6})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (pla[56])&(M4&T3);
ctl_sw_2d = ctl_sw_2d | (pla[56])&(M4&T3);
ctl_sw_1d = ctl_sw_1d | (pla[56])&(M4&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[56])&(M4&T3);
fMRead = fMRead | (pla[56])&(M5&T1);
ctl_reg_sel_ir = ctl_reg_sel_ir | (pla[56])&(M5&T1);
ctl_reg_sys_hilo_pla56M5T1_3 = (pla[56])&(M5&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla56M5T1_3,ctl_reg_sys_hilo_pla56M5T1_3})&(2'b10);
ctl_sw_4d = ctl_sw_4d | (pla[56])&(M5&T1);
ctl_al_we = ctl_al_we | (pla[56])&(M5&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[56])&(M5&T1);
ctl_sw_2u = ctl_sw_2u | (pla[56])&(M5&T1);
ctl_alu_oe = ctl_alu_oe | (pla[56])&(M5&T1);
ctl_alu_op1_oe = ctl_alu_op1_oe | (pla[56])&(M5&T1);
fMRead = fMRead | (pla[56])&(M5&T2);
ctl_inc_cy = ctl_inc_cy | (pla[56])&(M5&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[56])&(M5&T2);
fMRead = fMRead | (pla[56])&(M5&T3);
setM1 = setM1 | (pla[56])&(M5&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[56])&(M5&T3);
ctl_reg_sys_hilo_pla56M5T3_4 = (pla[56])&(M5&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla56M5T3_4,ctl_reg_sys_hilo_pla56M5T3_4})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (pla[56])&(M5&T3);
ctl_al_we = ctl_al_we | (pla[56])&(M5&T3);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (pla[56])&(M5&T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (pla[56])&(M5&T3);
ctl_reg_sys_hilo_pla56M5T3_9 = (pla[56])&(M5&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla56M5T3_9,ctl_reg_sys_hilo_pla56M5T3_9})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (pla[56])&(M5&T3);
ctl_sw_2d = ctl_sw_2d | (pla[56])&(M5&T3);
ctl_sw_1d = ctl_sw_1d | (pla[56])&(M5&T3);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[56])&(M5&T3);
ctl_reg_not_pc = ctl_reg_not_pc | (pla[56])&(M5&T3);
ctl_reg_gp_sel_pla49M1T3_1 = (pla[49])&(M1&T3);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla49M1T3_1,ctl_reg_gp_sel_pla49M1T3_1})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla49M1T3_2 = (pla[49])&(M1&T3);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla49M1T3_2,ctl_reg_gp_hilo_pla49M1T3_2})&(2'b11);
ctl_reg_out_hi = ctl_reg_out_hi | (pla[49])&(M1&T3);
ctl_reg_out_lo = ctl_reg_out_lo | (pla[49])&(M1&T3);
ctl_flags_bus = ctl_flags_bus | (pla[49])&(M1&T3);
ctl_alu_shift_oe = ctl_alu_shift_oe | (pla[49])&(M1&T3)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[49])&(M1&T3);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[49])&(M1&T3);
ctl_flags_sz_we = ctl_flags_sz_we | (pla[49])&(M1&T3);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[49])&(M1&T3);
ctl_flags_hf_we = ctl_flags_hf_we | (pla[49])&(M1&T3);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[49])&(M1&T3);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[49])&(M1&T3);
ctl_flags_cf_we = ctl_flags_cf_we | (pla[49])&(M1&T3);
ctl_state_tbl_we = ctl_state_tbl_we | (pla[49])&(M1&T3);
ctl_state_tbl_cb_set = ctl_state_tbl_cb_set | (pla[49])&(M1&T3);
validPLA = validPLA | (pla[49])&(M1&T4);
nextM = nextM | (pla[49])&(M1&T4);
ctl_mRead = ctl_mRead | (pla[49])&(M1&T4);
fMRead = fMRead | (pla[49])&(M2&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[49])&(M2&T1);
ctl_reg_sys_hilo_pla49M2T1_3 = (pla[49])&(M2&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla49M2T1_3,ctl_reg_sys_hilo_pla49M2T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[49])&(M2&T1);
fMRead = fMRead | (pla[49])&(M2&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[49])&(M2&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[49])&(M2&T2);
ctl_reg_sys_hilo_pla49M2T2_4 = (pla[49])&(M2&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla49M2T2_4,ctl_reg_sys_hilo_pla49M2T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[49])&(M2&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[49])&(M2&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[49])&(M2&T2);
fMRead = fMRead | (pla[49])&(M2&T3);
nextM = nextM | (pla[49])&(M2&T3);
ctl_mRead = ctl_mRead | (pla[49])&(M2&T3);
fMRead = fMRead | (pla[49])&(M3&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[49])&(M3&T1);
ctl_reg_sys_hilo_pla49M3T1_3 = (pla[49])&(M3&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla49M3T1_3,ctl_reg_sys_hilo_pla49M3T1_3})&(2'b11);
ctl_al_we = ctl_al_we | (pla[49])&(M3&T1);
ixy_d = ixy_d | (pla[49])&(M3&T1);
fMRead = fMRead | (pla[49])&(M3&T2);
ctl_reg_sys_we = ctl_reg_sys_we | (pla[49])&(M3&T2);
ctl_reg_sel_pc = ctl_reg_sel_pc | (pla[49])&(M3&T2);
ctl_reg_sys_hilo_pla49M3T2_4 = (pla[49])&(M3&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_pla49M3T2_4,ctl_reg_sys_hilo_pla49M3T2_4})&(2'b11);
pc_inc_hold = pc_inc_hold | (pla[49])&(M3&T2)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (pla[49])&(M3&T2)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (pla[49])&(M3&T2);
ixy_d = ixy_d | (pla[49])&(M3&T2);
fMRead = fMRead | (pla[49])&(M3&T3);
ixy_d = ixy_d | (pla[49])&(M3&T3);
ixy_d = ixy_d | (pla[49])&(M3&T4);
nextM = nextM | (pla[49])&(M3&T5);
ctl_mRead = ctl_mRead | (pla[49])&(M3&T5);
ixy_d = ixy_d | (pla[49])&(M3&T5);
ctl_bus_db_oe = ctl_bus_db_oe | (pla[49])&(M4&T1);
ctl_alu_bs_oe = ctl_alu_bs_oe | (pla[49])&(M4&T1);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (pla[49])&(M4&T1);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (pla[49])&(M4&T1);
ctl_ir_we = ctl_ir_we | (pla[49])&(M4&T1);
ctl_state_ixiy_we = ctl_state_ixiy_we | (pla[3])&(M1&T2);
ctl_state_iy_set = ctl_state_iy_set | (pla[3])&(M1&T2)&(op5);
setIXIY = setIXIY | (pla[3])&(M1&T2);
validPLA = validPLA | (pla[3])&(M1&T4);
setM1 = setM1 | (pla[3])&(M1&T4);
ctl_no_ints = ctl_no_ints | (pla[3])&(M1&T4);
ctl_state_tbl_we = ctl_state_tbl_we | (pla[44])&(M1&T2);
ctl_state_tbl_cb_set = ctl_state_tbl_cb_set | (pla[44])&(M1&T2);
validPLA = validPLA | (pla[44])&(M1&T4);
setM1 = setM1 | (pla[44])&(M1&T4);
ctl_no_ints = ctl_no_ints | (pla[44])&(M1&T4);
ctl_state_tbl_we = ctl_state_tbl_we | (pla[51])&(M1&T2);
ctl_state_tbl_ed_set = ctl_state_tbl_ed_set | (pla[51])&(M1&T2);
validPLA = validPLA | (pla[51])&(M1&T4);
setM1 = setM1 | (pla[51])&(M1&T4);
ctl_no_ints = ctl_no_ints | (pla[51])&(M1&T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[76]);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[76])&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[76])&(~ctl_alu_op_low);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[76]);
ctl_flags_nf_set = ctl_flags_nf_set | (pla[76]);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[76])&(M1&T1);
ctl_pf_sel_pla76M1T1_2 = (pla[76])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla76M1T1_2,ctl_pf_sel_pla76M1T1_2})&(`PFSEL_V);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[78]);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[78])&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[78])&(~ctl_alu_op_low);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[78]);
ctl_flags_nf_set = ctl_flags_nf_set | (pla[78]);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[78])&(M1&T1);
ctl_reg_gp_sel_pla78M1T1_2 = (pla[78])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla78M1T1_2,ctl_reg_gp_sel_pla78M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla78M1T1_3 = (pla[78])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla78M1T1_3,ctl_reg_gp_hilo_pla78M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[78])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[78])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[78])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[78])&(M1&T1);
ctl_pf_sel_pla78M1T1_8 = (pla[78])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla78M1T1_8,ctl_pf_sel_pla78M1T1_8})&(`PFSEL_V);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (pla[79]);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[79])&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[79])&(~ctl_alu_op_low);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[79]);
ctl_flags_nf_set = ctl_flags_nf_set | (pla[79]);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[79])&(M1&T1);
ctl_reg_gp_sel_pla79M1T1_2 = (pla[79])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla79M1T1_2,ctl_reg_gp_sel_pla79M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla79M1T1_3 = (pla[79])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla79M1T1_3,ctl_reg_gp_hilo_pla79M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[79])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[79])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[79])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[79])&(M1&T1);
ctl_pf_sel_pla79M1T1_8 = (pla[79])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla79M1T1_8,ctl_pf_sel_pla79M1T1_8})&(`PFSEL_V);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[80])&(~ctl_alu_op_low);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[80]);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[80]);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[80])&(M1&T1);
ctl_reg_gp_sel_pla80M1T1_2 = (pla[80])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla80M1T1_2,ctl_reg_gp_sel_pla80M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla80M1T1_3 = (pla[80])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla80M1T1_3,ctl_reg_gp_hilo_pla80M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[80])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[80])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[80])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[80])&(M1&T1);
ctl_pf_sel_pla80M1T1_8 = (pla[80])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla80M1T1_8,ctl_pf_sel_pla80M1T1_8})&(`PFSEL_V);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[84])&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[84])&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (pla[84])&(~ctl_alu_op_low);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[84]);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[84]);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[84])&(M1&T1);
ctl_reg_gp_sel_pla84M1T1_2 = (pla[84])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla84M1T1_2,ctl_reg_gp_sel_pla84M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla84M1T1_3 = (pla[84])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla84M1T1_3,ctl_reg_gp_hilo_pla84M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[84])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[84])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[84])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[84])&(M1&T1);
ctl_pf_sel_pla84M1T1_8 = (pla[84])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla84M1T1_8,ctl_pf_sel_pla84M1T1_8})&(`PFSEL_V);
ctl_alu_core_S = ctl_alu_core_S | (pla[85]);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[85]);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[85]);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[85]);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[85])&(M1&T1);
ctl_reg_gp_sel_pla85M1T1_2 = (pla[85])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla85M1T1_2,ctl_reg_gp_sel_pla85M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla85M1T1_3 = (pla[85])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla85M1T1_3,ctl_reg_gp_hilo_pla85M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[85])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[85])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[85])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[85])&(M1&T1);
ctl_pf_sel_pla85M1T1_8 = (pla[85])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla85M1T1_8,ctl_pf_sel_pla85M1T1_8})&(`PFSEL_P);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[85])&(M1&T2);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[85])&(M1&T2);
ctl_alu_core_R = ctl_alu_core_R | (pla[86]);
ctl_alu_core_V = ctl_alu_core_V | (pla[86]);
ctl_alu_core_S = ctl_alu_core_S | (pla[86]);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[86]);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[86]);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[86]);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[86]);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[86])&(M1&T1);
ctl_reg_gp_sel_pla86M1T1_2 = (pla[86])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla86M1T1_2,ctl_reg_gp_sel_pla86M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla86M1T1_3 = (pla[86])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla86M1T1_3,ctl_reg_gp_hilo_pla86M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[86])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[86])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[86])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[86])&(M1&T1);
ctl_pf_sel_pla86M1T1_8 = (pla[86])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla86M1T1_8,ctl_pf_sel_pla86M1T1_8})&(`PFSEL_P);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[86])&(M1&T2);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[86])&(M1&T2);
ctl_alu_core_R = ctl_alu_core_R | (pla[88]);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[88]);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[88]);
ctl_flags_nf_we = ctl_flags_nf_we | (pla[88]);
ctl_flags_nf_clr = ctl_flags_nf_clr | (pla[88]);
ctl_reg_gp_we = ctl_reg_gp_we | (pla[88])&(M1&T1);
ctl_reg_gp_sel_pla88M1T1_2 = (pla[88])&(M1&T1);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_pla88M1T1_2,ctl_reg_gp_sel_pla88M1T1_2})&(`GP_REG_AF);
ctl_reg_gp_hilo_pla88M1T1_3 = (pla[88])&(M1&T1);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_pla88M1T1_3,ctl_reg_gp_hilo_pla88M1T1_3})&(2'b10);
ctl_reg_in_hi = ctl_reg_in_hi | (pla[88])&(M1&T1);
ctl_reg_in_lo = ctl_reg_in_lo | (pla[88])&(M1&T1);
ctl_flags_xy_we = ctl_flags_xy_we | (pla[88])&(M1&T1);
ctl_flags_pf_we = ctl_flags_pf_we | (pla[88])&(M1&T1);
ctl_pf_sel_pla88M1T1_8 = (pla[88])&(M1&T1);
ctl_pf_sel = ctl_pf_sel | ({ctl_pf_sel_pla88M1T1_8,ctl_pf_sel_pla88M1T1_8})&(`PFSEL_P);
ctl_flags_cf_set = ctl_flags_cf_set | (pla[88])&(M1&T2);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (pla[88])&(M1&T2);
ctl_sw_2d = ctl_sw_2d | (ixy_d)&(T1);
ctl_sw_1d = ctl_sw_1d | (ixy_d)&(T1);
ctl_bus_db_oe = ctl_bus_db_oe | (ixy_d)&(T1);
ctl_flags_alu = ctl_flags_alu | (ixy_d)&(T1);
ctl_alu_shift_oe = ctl_alu_shift_oe | (ixy_d)&(T1)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_bus = ctl_alu_op2_sel_bus | (ixy_d)&(T1);
ctl_flags_sz_we = ctl_flags_sz_we | (ixy_d)&(T1);
ctl_reg_gp_sel_ixy_dT2_1 = (ixy_d)&(T2);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_ixy_dT2_1,ctl_reg_gp_sel_ixy_dT2_1})&(`GP_REG_HL);
ctl_reg_gp_hilo_ixy_dT2_2 = (ixy_d)&(T2);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_ixy_dT2_2,ctl_reg_gp_hilo_ixy_dT2_2})&(2'b01);
ctl_reg_out_lo = ctl_reg_out_lo | (ixy_d)&(T2);
ctl_sw_2d = ctl_sw_2d | (ixy_d)&(T2);
ctl_flags_alu = ctl_flags_alu | (ixy_d)&(T2);
ctl_alu_shift_oe = ctl_alu_shift_oe | (ixy_d)&(T2)&(~ctl_alu_bs_oe);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (ixy_d)&(T2);
ctl_alu_op_low = ctl_alu_op_low | (ixy_d)&(T2);
ctl_flags_cf_set = ctl_flags_cf_set | (ixy_d)&(T2)&(ctl_alu_op_low);
ctl_flags_cf_cpl = ctl_flags_cf_cpl | (ixy_d)&(T2)&(ctl_alu_op_low);
ctl_alu_core_hf = ctl_alu_core_hf | (ixy_d)&(T2)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (ixy_d)&(T2);
ctl_reg_sys_we_lo = ctl_reg_sys_we_lo | (ixy_d)&(T3);
ctl_reg_sel_wz = ctl_reg_sel_wz | (ixy_d)&(T3);
ctl_reg_sys_hilo_ixy_dT3_3 = (ixy_d)&(T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_ixy_dT3_3,ctl_reg_sys_hilo_ixy_dT3_3})&({ctl_reg_sys_hilo[1],1'b1});
ctl_reg_in_lo = ctl_reg_in_lo | (ixy_d)&(T3);
ctl_sw_2u = ctl_sw_2u | (ixy_d)&(T3);
ctl_flags_alu = ctl_flags_alu | (ixy_d)&(T3);
ctl_alu_oe = ctl_alu_oe | (ixy_d)&(T3);
ctl_alu_res_oe = ctl_alu_res_oe | (ixy_d)&(T3);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (ixy_d)&(T3);
ctl_alu_core_hf = ctl_alu_core_hf | (ixy_d)&(T3)&(~ctl_alu_op_low);
ctl_flags_cf2_we = ctl_flags_cf2_we | (ixy_d)&(T3);
ctl_reg_gp_sel_ixy_dT4_1 = (ixy_d)&(T4);
ctl_reg_gp_sel = ctl_reg_gp_sel | ({ctl_reg_gp_sel_ixy_dT4_1,ctl_reg_gp_sel_ixy_dT4_1})&(`GP_REG_HL);
ctl_reg_gp_hilo_ixy_dT4_2 = (ixy_d)&(T4);
ctl_reg_gp_hilo = ctl_reg_gp_hilo | ({ctl_reg_gp_hilo_ixy_dT4_2,ctl_reg_gp_hilo_ixy_dT4_2})&(2'b10);
ctl_reg_out_hi = ctl_reg_out_hi | (ixy_d)&(T4);
ctl_reg_out_lo = ctl_reg_out_lo | (ixy_d)&(T4);
ctl_flags_alu = ctl_flags_alu | (ixy_d)&(T4);
ctl_alu_shift_oe = ctl_alu_shift_oe | (ixy_d)&(T4)&(~ctl_alu_bs_oe);
ctl_alu_op2_sel_zero = ctl_alu_op2_sel_zero | (ixy_d)&(T4);
ctl_alu_op1_sel_bus = ctl_alu_op1_sel_bus | (ixy_d)&(T4);
ctl_alu_op_low = ctl_alu_op_low | (ixy_d)&(T4);
ctl_alu_core_hf = ctl_alu_core_hf | (ixy_d)&(T4)&(~ctl_alu_op_low);
ctl_flags_hf_we = ctl_flags_hf_we | (ixy_d)&(T4);
ctl_flags_use_cf2 = ctl_flags_use_cf2 | (ixy_d)&(T4);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (ixy_d)&(T4)&(flags_sf);
ctl_reg_sel_wz = ctl_reg_sel_wz | (ixy_d)&(T5);
ctl_reg_sys_hilo_ixy_dT5_2 = (ixy_d)&(T5);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_ixy_dT5_2,ctl_reg_sys_hilo_ixy_dT5_2})&(2'b11);
ctl_sw_4d = ctl_sw_4d | (ixy_d)&(T5);
ctl_al_we = ctl_al_we | (ixy_d)&(T5);
ctl_reg_sys_we_hi = ctl_reg_sys_we_hi | (ixy_d)&(T5);
ctl_reg_sel_wz = ctl_reg_sel_wz | (ixy_d)&(T5);
ctl_reg_sys_hilo_ixy_dT5_7 = (ixy_d)&(T5);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_ixy_dT5_7,ctl_reg_sys_hilo_ixy_dT5_7})&({1'b1,ctl_reg_sys_hilo[0]});
ctl_reg_in_hi = ctl_reg_in_hi | (ixy_d)&(T5);
ctl_flags_alu = ctl_flags_alu | (ixy_d)&(T5);
ctl_alu_oe = ctl_alu_oe | (ixy_d)&(T5);
ctl_alu_res_oe = ctl_alu_res_oe | (ixy_d)&(T5);
ctl_alu_sel_op2_high = ctl_alu_sel_op2_high | (ixy_d)&(T5);
ctl_alu_core_hf = ctl_alu_core_hf | (ixy_d)&(T5)&(~ctl_alu_op_low);
ctl_flags_xy_we = ctl_flags_xy_we | (ixy_d)&(T5);
ctl_alu_sel_op2_neg = ctl_alu_sel_op2_neg | (ixy_d)&(T5)&(flags_sf);
ctl_state_ixiy_we = ctl_state_ixiy_we | (ixy_d)&(T5);
ctl_state_ixiy_clr = ctl_state_ixiy_clr | (ixy_d)&(T5)&(~setIXIY);
ctl_reg_sys_we = ctl_reg_sys_we | (M1&T1);
ctl_reg_sel_pc = ctl_reg_sel_pc | (M1&T1);
ctl_reg_sys_hilo_1M1T1_3 = (M1&T1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_1M1T1_3,ctl_reg_sys_hilo_1M1T1_3})&(2'b11);
pc_inc_hold = pc_inc_hold | (M1&T1)&((in_halt|in_intr|in_nmi));
ctl_inc_cy = ctl_inc_cy | (M1&T1)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (M1&T1);
ctl_apin_mux2 = ctl_apin_mux2 | (M1&T1);
ctl_reg_sel_ir = ctl_reg_sel_ir | (M1&T2);
ctl_reg_sys_hilo_1M1T2_2 = (M1&T2);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_1M1T2_2,ctl_reg_sys_hilo_1M1T2_2})&(2'b11);
ctl_al_we = ctl_al_we | (M1&T2);
ctl_bus_db_oe = ctl_bus_db_oe | (M1&T2);
ctl_state_ixiy_we = ctl_state_ixiy_we | (M1&T2);
ctl_state_ixiy_clr = ctl_state_ixiy_clr | (M1&T2)&(~setIXIY);
ctl_state_tbl_we = ctl_state_tbl_we | (M1&T2);
ctl_ir_we = ctl_ir_we | (M1&T2);
ctl_bus_zero_oe = ctl_bus_zero_oe | (M1&T2)&(in_halt);
ctl_bus_ff_oe = ctl_bus_ff_oe | (M1&T2)&((in_intr&(im1|im2))|in_nmi);
ctl_reg_sys_we = ctl_reg_sys_we | (M1&T3);
ctl_reg_sel_ir = ctl_reg_sel_ir | (M1&T3);
ctl_reg_sys_hilo_1M1T3_3 = (M1&T3);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_1M1T3_3,ctl_reg_sys_hilo_1M1T3_3})&(2'b11);
ctl_inc_cy = ctl_inc_cy | (M1&T3)&(~pc_inc_hold);
ctl_bus_inc_oe = ctl_bus_inc_oe | (M1&T3);
ctl_apin_mux2 = ctl_apin_mux2 | (M1&T3);
ctl_inc_limit6 = ctl_inc_limit6 | (M1&T3);
ctl_eval_cond = ctl_eval_cond | (M1&T4);
setM1 = setM1 | (~validPLA)&(M1&T4);
ctl_reg_sel_pc = ctl_reg_sel_pc | (setM1);
ctl_reg_sys_hilo_setM1_2 = (setM1);
ctl_reg_sys_hilo = ctl_reg_sys_hilo | ({ctl_reg_sys_hilo_setM1_2,ctl_reg_sys_hilo_setM1_2})&(2'b11);
ctl_al_we = ctl_al_we | (setM1);
